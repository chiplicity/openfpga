magic
tech EFS8A
magscale 1 2
timestamp 1602278301
<< locali >>
rect 24259 41633 24294 41667
rect 26893 41055 26927 41157
rect 31585 41055 31619 41225
rect 23615 41021 23742 41055
rect 29791 40885 29929 40919
rect 14105 40545 14266 40579
rect 23247 40545 23282 40579
rect 28917 40545 29078 40579
rect 34011 40545 34046 40579
rect 38335 40545 38370 40579
rect 14105 40511 14139 40545
rect 28917 40511 28951 40545
rect 24311 39593 24317 39627
rect 24311 39525 24345 39593
rect 34379 39457 34414 39491
rect 40877 38879 40911 39049
rect 25547 38777 25592 38811
rect 11799 38505 11805 38539
rect 38111 38505 38117 38539
rect 11799 38437 11833 38505
rect 38111 38437 38145 38505
rect 28491 38369 28526 38403
rect 39531 38369 39566 38403
rect 32499 37417 32505 37451
rect 32499 37349 32533 37417
rect 25145 36567 25179 36737
rect 26065 36567 26099 36669
rect 16767 36329 16773 36363
rect 36179 36329 36185 36363
rect 16767 36261 16801 36329
rect 36179 36261 36213 36329
rect 14139 36193 14266 36227
rect 15243 36193 15370 36227
rect 34379 36193 34414 36227
rect 39715 36193 39750 36227
rect 24679 35479 24713 35547
rect 24679 35445 24685 35479
rect 24679 35241 24685 35275
rect 24679 35173 24713 35241
rect 19257 34459 19291 34697
rect 19251 34153 19257 34187
rect 21827 34153 21833 34187
rect 19251 34085 19285 34153
rect 21827 34085 21861 34153
rect 11931 34017 11966 34051
rect 30849 33371 30883 33609
rect 40601 33439 40635 33609
rect 43723 33065 43729 33099
rect 43723 32997 43757 33065
rect 34069 32963 34103 32997
rect 25179 32929 25306 32963
rect 34069 32929 34230 32963
rect 22845 32283 22879 32521
rect 25599 32215 25633 32283
rect 25599 32181 25605 32215
rect 32499 31977 32505 32011
rect 32499 31909 32533 31977
rect 26467 31841 26594 31875
rect 42291 31841 42326 31875
rect 45051 31841 45086 31875
rect 29043 30753 29078 30787
rect 14933 30107 14967 30277
rect 23615 30141 23742 30175
rect 25973 30107 26007 30345
rect 17319 29801 17325 29835
rect 22563 29801 22569 29835
rect 43723 29801 43729 29835
rect 17319 29733 17353 29801
rect 22563 29733 22597 29801
rect 43723 29733 43757 29801
rect 9781 29665 9942 29699
rect 26467 29665 26594 29699
rect 35575 29665 35610 29699
rect 45143 29665 45178 29699
rect 9781 29631 9815 29665
rect 22569 29019 22603 29257
rect 21551 28713 21557 28747
rect 30107 28713 30113 28747
rect 33419 28713 33425 28747
rect 21551 28645 21585 28713
rect 30107 28645 30141 28713
rect 33419 28645 33453 28713
rect 14231 28577 14266 28611
rect 19717 28577 19878 28611
rect 43303 28577 43430 28611
rect 19717 28407 19751 28577
rect 26801 27965 26962 27999
rect 26801 27931 26835 27965
rect 18515 27863 18549 27931
rect 18515 27829 18521 27863
rect 38111 27625 38117 27659
rect 41515 27625 41521 27659
rect 38111 27557 38145 27625
rect 41515 27557 41549 27625
rect 9781 27489 9942 27523
rect 9781 27319 9815 27489
rect 12265 27387 12299 27557
rect 24087 26945 24225 26979
rect 10551 26401 10586 26435
rect 13127 26401 13162 26435
rect 23891 26401 23926 26435
rect 30975 26401 31102 26435
rect 34011 26401 34046 26435
rect 36587 26401 36622 26435
rect 44407 26401 44442 26435
rect 28359 25449 28365 25483
rect 28359 25381 28393 25449
rect 12541 24667 12575 24837
rect 44097 24735 44131 24905
rect 38059 24633 38104 24667
rect 24219 24361 24225 24395
rect 24219 24293 24253 24361
rect 41239 23273 41245 23307
rect 41239 23205 41273 23273
rect 14231 23137 14266 23171
rect 36311 23137 36346 23171
rect 21097 22627 21131 22729
rect 23615 22525 23742 22559
rect 29653 22423 29687 22593
rect 31309 22423 31343 22525
rect 38295 22185 38301 22219
rect 18647 22049 18682 22083
rect 19659 22049 19694 22083
rect 23489 21879 23523 22185
rect 38295 22117 38329 22185
rect 36679 22049 36714 22083
rect 28825 21335 28859 21641
rect 32499 21097 32505 21131
rect 32499 21029 32533 21097
rect 14703 20553 14841 20587
rect 32367 20553 32505 20587
rect 40503 20009 40509 20043
rect 40503 19941 40537 20009
rect 18003 19873 18038 19907
rect 29503 19873 29538 19907
rect 35173 19295 35207 19397
rect 32079 18785 32206 18819
rect 18003 18173 18130 18207
rect 18975 17833 18981 17867
rect 21275 17833 21281 17867
rect 18975 17765 19009 17833
rect 21275 17765 21309 17833
rect 36587 17697 36622 17731
rect 18423 16983 18457 17051
rect 18423 16949 18429 16983
rect 10327 16745 10333 16779
rect 10327 16677 10361 16745
rect 21315 16609 21350 16643
rect 21275 15657 21281 15691
rect 28635 15657 28641 15691
rect 21275 15589 21309 15657
rect 28635 15589 28669 15657
rect 9999 15521 10034 15555
rect 43303 15521 43430 15555
rect 32045 14875 32079 15113
rect 34529 14943 34563 15113
rect 39589 14943 39623 15045
rect 10327 14807 10361 14875
rect 10327 14773 10333 14807
rect 10419 14569 10425 14603
rect 32499 14569 32505 14603
rect 10419 14501 10453 14569
rect 32499 14501 32533 14569
rect 35995 13719 36029 13787
rect 35995 13685 36001 13719
rect 28635 13481 28641 13515
rect 28635 13413 28669 13481
rect 15243 13345 15370 13379
rect 23391 12393 23397 12427
rect 39399 12393 39405 12427
rect 10551 12325 10596 12359
rect 23391 12325 23425 12393
rect 39399 12325 39433 12393
rect 23305 11611 23339 11781
rect 14933 10523 14967 10761
rect 23615 10557 23742 10591
rect 30935 10455 30969 10523
rect 30935 10421 30941 10455
rect 22471 10217 22477 10251
rect 22471 10149 22505 10217
rect 8355 9673 8493 9707
rect 21735 9367 21769 9435
rect 21735 9333 21741 9367
rect 27163 9129 27169 9163
rect 27163 9061 27197 9129
rect 13553 7191 13587 7361
rect 16899 7293 17026 7327
rect 20855 7293 20890 7327
rect 22195 7191 22229 7259
rect 27088 7225 27156 7259
rect 22195 7157 22201 7191
rect 32499 6953 32505 6987
rect 32499 6885 32533 6953
rect 36369 6851 36403 6885
rect 36369 6817 36530 6851
rect 10879 5865 10885 5899
rect 10879 5797 10913 5865
rect 37691 5729 37818 5763
rect 28825 4131 28859 4233
rect 16583 3689 16589 3723
rect 16583 3621 16617 3689
rect 30389 3587 30423 3689
rect 26467 3553 26594 3587
rect 12851 2941 12886 2975
rect 16583 2601 16589 2635
rect 16583 2533 16617 2601
<< viali >>
rect 21348 42721 21382 42755
rect 21419 42517 21453 42551
rect 21408 42109 21442 42143
rect 22201 42109 22235 42143
rect 24476 42109 24510 42143
rect 24869 42109 24903 42143
rect 21511 41973 21545 42007
rect 21833 41973 21867 42007
rect 24547 41973 24581 42007
rect 24869 41769 24903 41803
rect 21741 41701 21775 41735
rect 16656 41633 16690 41667
rect 18956 41633 18990 41667
rect 24225 41633 24259 41667
rect 25304 41633 25338 41667
rect 26652 41633 26686 41667
rect 29720 41633 29754 41667
rect 32540 41633 32574 41667
rect 21649 41565 21683 41599
rect 22293 41565 22327 41599
rect 16497 41429 16531 41463
rect 16727 41429 16761 41463
rect 19027 41429 19061 41463
rect 19441 41429 19475 41463
rect 19717 41429 19751 41463
rect 24363 41429 24397 41463
rect 25375 41429 25409 41463
rect 26755 41429 26789 41463
rect 29791 41429 29825 41463
rect 32643 41429 32677 41463
rect 19073 41225 19107 41259
rect 22569 41225 22603 41259
rect 27445 41225 27479 41259
rect 31585 41225 31619 41259
rect 19901 41157 19935 41191
rect 26893 41157 26927 41191
rect 27077 41157 27111 41191
rect 18383 41089 18417 41123
rect 19349 41089 19383 41123
rect 20729 41089 20763 41123
rect 21649 41089 21683 41123
rect 23811 41089 23845 41123
rect 24961 41089 24995 41123
rect 25605 41089 25639 41123
rect 30573 41089 30607 41123
rect 32689 41157 32723 41191
rect 14416 41021 14450 41055
rect 14841 41021 14875 41055
rect 16313 41021 16347 41055
rect 16405 41021 16439 41055
rect 16865 41021 16899 41055
rect 17509 41021 17543 41055
rect 18296 41021 18330 41055
rect 23581 41021 23615 41055
rect 26684 41021 26718 41055
rect 26893 41021 26927 41055
rect 29720 41021 29754 41055
rect 31284 41021 31318 41055
rect 31585 41021 31619 41055
rect 32264 41021 32298 41055
rect 33308 41021 33342 41055
rect 33701 41021 33735 41055
rect 19441 40953 19475 40987
rect 21097 40953 21131 40987
rect 21465 40953 21499 40987
rect 21741 40953 21775 40987
rect 22293 40953 22327 40987
rect 24777 40953 24811 40987
rect 25053 40953 25087 40987
rect 25973 40953 26007 40987
rect 31677 40953 31711 40987
rect 33057 40953 33091 40987
rect 14519 40885 14553 40919
rect 16497 40885 16531 40919
rect 18797 40885 18831 40919
rect 23397 40885 23431 40919
rect 24317 40885 24351 40919
rect 26755 40885 26789 40919
rect 29929 40885 29963 40919
rect 30205 40885 30239 40919
rect 31355 40885 31389 40919
rect 32367 40885 32401 40919
rect 33379 40885 33413 40919
rect 24593 40681 24627 40715
rect 16681 40613 16715 40647
rect 19441 40613 19475 40647
rect 21741 40613 21775 40647
rect 21833 40613 21867 40647
rect 25053 40613 25087 40647
rect 26985 40613 27019 40647
rect 27077 40613 27111 40647
rect 30205 40613 30239 40647
rect 32597 40613 32631 40647
rect 18128 40545 18162 40579
rect 23213 40545 23247 40579
rect 33977 40545 34011 40579
rect 35056 40545 35090 40579
rect 38301 40545 38335 40579
rect 14105 40477 14139 40511
rect 16589 40477 16623 40511
rect 17233 40477 17267 40511
rect 19349 40477 19383 40511
rect 19993 40477 20027 40511
rect 22017 40477 22051 40511
rect 24961 40477 24995 40511
rect 25605 40477 25639 40511
rect 27261 40477 27295 40511
rect 28917 40477 28951 40511
rect 30113 40477 30147 40511
rect 32505 40477 32539 40511
rect 32781 40477 32815 40511
rect 39129 40477 39163 40511
rect 30665 40409 30699 40443
rect 35127 40409 35161 40443
rect 14335 40341 14369 40375
rect 14657 40341 14691 40375
rect 16313 40341 16347 40375
rect 18199 40341 18233 40375
rect 23351 40341 23385 40375
rect 29147 40341 29181 40375
rect 34115 40341 34149 40375
rect 37105 40341 37139 40375
rect 38439 40341 38473 40375
rect 38853 40341 38887 40375
rect 14197 40137 14231 40171
rect 17877 40137 17911 40171
rect 19165 40137 19199 40171
rect 20821 40137 20855 40171
rect 22753 40137 22787 40171
rect 24501 40137 24535 40171
rect 25605 40137 25639 40171
rect 27905 40137 27939 40171
rect 31033 40137 31067 40171
rect 35173 40137 35207 40171
rect 17049 40069 17083 40103
rect 22293 40069 22327 40103
rect 25237 40069 25271 40103
rect 33977 40069 34011 40103
rect 38301 40069 38335 40103
rect 13369 40001 13403 40035
rect 14657 40001 14691 40035
rect 16497 40001 16531 40035
rect 17417 40001 17451 40035
rect 18383 40001 18417 40035
rect 19349 40001 19383 40035
rect 20269 40001 20303 40035
rect 21741 40001 21775 40035
rect 23213 40001 23247 40035
rect 24685 40001 24719 40035
rect 26065 40001 26099 40035
rect 26985 40001 27019 40035
rect 27261 40001 27295 40035
rect 30113 40001 30147 40035
rect 31677 40001 31711 40035
rect 32597 40001 32631 40035
rect 12976 39933 13010 39967
rect 18296 39933 18330 39967
rect 35852 39933 35886 39967
rect 36277 39933 36311 39967
rect 37013 39933 37047 39967
rect 37473 39933 37507 39967
rect 14749 39865 14783 39899
rect 15301 39865 15335 39899
rect 15945 39865 15979 39899
rect 16313 39865 16347 39899
rect 16589 39865 16623 39899
rect 19441 39865 19475 39899
rect 19993 39865 20027 39899
rect 21833 39865 21867 39899
rect 24777 39865 24811 39899
rect 26433 39865 26467 39899
rect 26801 39865 26835 39899
rect 27054 39865 27088 39899
rect 30205 39865 30239 39899
rect 30757 39865 30791 39899
rect 32689 39865 32723 39899
rect 33241 39865 33275 39899
rect 36829 39865 36863 39899
rect 37749 39865 37783 39899
rect 38761 39865 38795 39899
rect 38853 39865 38887 39899
rect 39405 39865 39439 39899
rect 13047 39797 13081 39831
rect 18797 39797 18831 39831
rect 21189 39797 21223 39831
rect 21557 39797 21591 39831
rect 24133 39797 24167 39831
rect 29101 39797 29135 39831
rect 29561 39797 29595 39831
rect 29929 39797 29963 39831
rect 31953 39797 31987 39831
rect 32321 39797 32355 39831
rect 35955 39797 35989 39831
rect 14657 39593 14691 39627
rect 15715 39593 15749 39627
rect 16313 39593 16347 39627
rect 19441 39593 19475 39627
rect 19717 39593 19751 39627
rect 24317 39593 24351 39627
rect 24869 39593 24903 39627
rect 30389 39593 30423 39627
rect 31171 39593 31205 39627
rect 32505 39593 32539 39627
rect 36001 39593 36035 39627
rect 13369 39525 13403 39559
rect 13461 39525 13495 39559
rect 14013 39525 14047 39559
rect 16681 39525 16715 39559
rect 16773 39525 16807 39559
rect 18842 39525 18876 39559
rect 20085 39525 20119 39559
rect 21925 39525 21959 39559
rect 27077 39525 27111 39559
rect 29514 39525 29548 39559
rect 32965 39525 32999 39559
rect 36185 39525 36219 39559
rect 36277 39525 36311 39559
rect 38761 39525 38795 39559
rect 38853 39525 38887 39559
rect 12300 39457 12334 39491
rect 15644 39457 15678 39491
rect 31068 39457 31102 39491
rect 34345 39457 34379 39491
rect 40668 39457 40702 39491
rect 16957 39389 16991 39423
rect 18521 39389 18555 39423
rect 21833 39389 21867 39423
rect 22109 39389 22143 39423
rect 23949 39389 23983 39423
rect 26985 39389 27019 39423
rect 27629 39389 27663 39423
rect 29193 39389 29227 39423
rect 32873 39389 32907 39423
rect 33149 39389 33183 39423
rect 36829 39389 36863 39423
rect 39405 39389 39439 39423
rect 12403 39253 12437 39287
rect 23765 39253 23799 39287
rect 25237 39253 25271 39287
rect 30113 39253 30147 39287
rect 30849 39253 30883 39287
rect 34483 39253 34517 39287
rect 40739 39253 40773 39287
rect 14013 39049 14047 39083
rect 14473 39049 14507 39083
rect 15669 39049 15703 39083
rect 17141 39049 17175 39083
rect 17417 39049 17451 39083
rect 20269 39049 20303 39083
rect 22339 39049 22373 39083
rect 23029 39049 23063 39083
rect 26525 39049 26559 39083
rect 27123 39049 27157 39083
rect 30665 39049 30699 39083
rect 33885 39049 33919 39083
rect 35633 39049 35667 39083
rect 39589 39049 39623 39083
rect 40877 39049 40911 39083
rect 41429 39049 41463 39083
rect 27445 38981 27479 39015
rect 39221 38981 39255 39015
rect 14657 38913 14691 38947
rect 16221 38913 16255 38947
rect 24685 38913 24719 38947
rect 25053 38913 25087 38947
rect 25237 38913 25271 38947
rect 28733 38913 28767 38947
rect 32965 38913 32999 38947
rect 33241 38913 33275 38947
rect 35219 38913 35253 38947
rect 36185 38913 36219 38947
rect 37105 38913 37139 38947
rect 37749 38913 37783 38947
rect 38669 38913 38703 38947
rect 41659 38913 41693 38947
rect 10701 38845 10735 38879
rect 11069 38845 11103 38879
rect 11345 38845 11379 38879
rect 11529 38845 11563 38879
rect 12449 38845 12483 38879
rect 15301 38845 15335 38879
rect 19165 38845 19199 38879
rect 19349 38845 19383 38879
rect 19625 38845 19659 38879
rect 20453 38845 20487 38879
rect 21373 38845 21407 38879
rect 22268 38845 22302 38879
rect 22661 38845 22695 38879
rect 23489 38845 23523 38879
rect 23673 38845 23707 38879
rect 24133 38845 24167 38879
rect 27020 38845 27054 38879
rect 29285 38845 29319 38879
rect 29745 38845 29779 38879
rect 30849 38845 30883 38879
rect 34437 38845 34471 38879
rect 35132 38845 35166 38879
rect 40576 38845 40610 38879
rect 40877 38845 40911 38879
rect 41556 38845 41590 38879
rect 41981 38845 42015 38879
rect 12173 38777 12207 38811
rect 12770 38777 12804 38811
rect 14749 38777 14783 38811
rect 16542 38777 16576 38811
rect 18521 38777 18555 38811
rect 20774 38777 20808 38811
rect 21833 38777 21867 38811
rect 25513 38777 25547 38811
rect 28365 38777 28399 38811
rect 31170 38777 31204 38811
rect 33057 38777 33091 38811
rect 36001 38777 36035 38811
rect 36277 38777 36311 38811
rect 36829 38777 36863 38811
rect 38117 38777 38151 38811
rect 38485 38777 38519 38811
rect 38761 38777 38795 38811
rect 40969 38777 41003 38811
rect 11897 38709 11931 38743
rect 13369 38709 13403 38743
rect 13645 38709 13679 38743
rect 16037 38709 16071 38743
rect 17877 38709 17911 38743
rect 19993 38709 20027 38743
rect 23949 38709 23983 38743
rect 26157 38709 26191 38743
rect 26893 38709 26927 38743
rect 29009 38709 29043 38743
rect 29377 38709 29411 38743
rect 31769 38709 31803 38743
rect 32413 38709 32447 38743
rect 32689 38709 32723 38743
rect 40647 38709 40681 38743
rect 10885 38505 10919 38539
rect 11805 38505 11839 38539
rect 12633 38505 12667 38539
rect 14565 38505 14599 38539
rect 16681 38505 16715 38539
rect 18521 38505 18555 38539
rect 20453 38505 20487 38539
rect 24317 38505 24351 38539
rect 25145 38505 25179 38539
rect 31033 38505 31067 38539
rect 33425 38505 33459 38539
rect 38117 38505 38151 38539
rect 39635 38505 39669 38539
rect 13277 38437 13311 38471
rect 13369 38437 13403 38471
rect 15485 38437 15519 38471
rect 17049 38437 17083 38471
rect 21925 38437 21959 38471
rect 23489 38437 23523 38471
rect 27077 38437 27111 38471
rect 30205 38437 30239 38471
rect 32505 38437 32539 38471
rect 32597 38437 32631 38471
rect 34115 38437 34149 38471
rect 35627 38437 35661 38471
rect 40969 38437 41003 38471
rect 18429 38369 18463 38403
rect 18981 38369 19015 38403
rect 25145 38369 25179 38403
rect 25329 38369 25363 38403
rect 28457 38369 28491 38403
rect 34028 38369 34062 38403
rect 37749 38369 37783 38403
rect 38669 38369 38703 38403
rect 39497 38369 39531 38403
rect 11437 38301 11471 38335
rect 13553 38301 13587 38335
rect 15393 38301 15427 38335
rect 16037 38301 16071 38335
rect 16957 38301 16991 38335
rect 17233 38301 17267 38335
rect 21833 38301 21867 38335
rect 22293 38301 22327 38335
rect 23397 38301 23431 38335
rect 23673 38301 23707 38335
rect 26985 38301 27019 38335
rect 28595 38301 28629 38335
rect 30113 38301 30147 38335
rect 30757 38301 30791 38335
rect 32873 38301 32907 38335
rect 35265 38301 35299 38335
rect 40877 38301 40911 38335
rect 27537 38233 27571 38267
rect 41429 38233 41463 38267
rect 12357 38165 12391 38199
rect 13001 38165 13035 38199
rect 19441 38165 19475 38199
rect 29285 38165 29319 38199
rect 36185 38165 36219 38199
rect 36461 38165 36495 38199
rect 36829 38165 36863 38199
rect 38945 38165 38979 38199
rect 42533 38165 42567 38199
rect 13461 37961 13495 37995
rect 18429 37961 18463 37995
rect 20545 37961 20579 37995
rect 22201 37961 22235 37995
rect 22523 37961 22557 37995
rect 23305 37961 23339 37995
rect 24777 37961 24811 37995
rect 27721 37961 27755 37995
rect 28089 37961 28123 37995
rect 29561 37961 29595 37995
rect 31033 37961 31067 37995
rect 31585 37961 31619 37995
rect 32505 37961 32539 37995
rect 33977 37961 34011 37995
rect 37473 37961 37507 37995
rect 38485 37961 38519 37995
rect 41889 37961 41923 37995
rect 13829 37893 13863 37927
rect 14335 37893 14369 37927
rect 35725 37893 35759 37927
rect 37841 37893 37875 37927
rect 12541 37825 12575 37859
rect 12817 37825 12851 37859
rect 28457 37825 28491 37859
rect 30757 37825 30791 37859
rect 32781 37825 32815 37859
rect 35311 37825 35345 37859
rect 36277 37825 36311 37859
rect 38669 37825 38703 37859
rect 40969 37825 41003 37859
rect 41245 37825 41279 37859
rect 42809 37825 42843 37859
rect 10793 37757 10827 37791
rect 11345 37757 11379 37791
rect 14264 37757 14298 37791
rect 15945 37757 15979 37791
rect 16824 37757 16858 37791
rect 17233 37757 17267 37791
rect 18981 37757 19015 37791
rect 19349 37757 19383 37791
rect 19533 37757 19567 37791
rect 19809 37757 19843 37791
rect 20637 37757 20671 37791
rect 22452 37757 22486 37791
rect 22845 37757 22879 37791
rect 23740 37757 23774 37791
rect 24869 37757 24903 37791
rect 26065 37757 26099 37791
rect 29929 37757 29963 37791
rect 30021 37757 30055 37791
rect 30481 37757 30515 37791
rect 31744 37757 31778 37791
rect 35224 37757 35258 37791
rect 36001 37757 36035 37791
rect 39681 37757 39715 37791
rect 11529 37689 11563 37723
rect 12633 37689 12667 37723
rect 15025 37689 15059 37723
rect 15301 37689 15335 37723
rect 15393 37689 15427 37723
rect 16911 37689 16945 37723
rect 17877 37689 17911 37723
rect 20958 37689 20992 37723
rect 25190 37689 25224 37723
rect 26801 37689 26835 37723
rect 26893 37689 26927 37723
rect 27445 37689 27479 37723
rect 32137 37689 32171 37723
rect 32873 37689 32907 37723
rect 33425 37689 33459 37723
rect 36369 37689 36403 37723
rect 36921 37689 36955 37723
rect 38761 37689 38795 37723
rect 39313 37689 39347 37723
rect 41061 37689 41095 37723
rect 42533 37689 42567 37723
rect 42625 37689 42659 37723
rect 10609 37621 10643 37655
rect 11897 37621 11931 37655
rect 12265 37621 12299 37655
rect 14749 37621 14783 37655
rect 16221 37621 16255 37655
rect 16589 37621 16623 37655
rect 21557 37621 21591 37655
rect 21833 37621 21867 37655
rect 23811 37621 23845 37655
rect 24225 37621 24259 37655
rect 25789 37621 25823 37655
rect 26525 37621 26559 37655
rect 31815 37621 31849 37655
rect 40325 37621 40359 37655
rect 40693 37621 40727 37655
rect 42257 37621 42291 37655
rect 10885 37417 10919 37451
rect 11529 37417 11563 37451
rect 15439 37417 15473 37451
rect 15761 37417 15795 37451
rect 16129 37417 16163 37451
rect 17601 37417 17635 37451
rect 20637 37417 20671 37451
rect 25145 37417 25179 37451
rect 25421 37417 25455 37451
rect 29561 37417 29595 37451
rect 30021 37417 30055 37451
rect 31861 37417 31895 37451
rect 32505 37417 32539 37451
rect 33333 37417 33367 37451
rect 35265 37417 35299 37451
rect 35541 37417 35575 37451
rect 36461 37417 36495 37451
rect 40877 37417 40911 37451
rect 41153 37417 41187 37451
rect 11207 37349 11241 37383
rect 12265 37349 12299 37383
rect 21925 37349 21959 37383
rect 22477 37349 22511 37383
rect 24777 37349 24811 37383
rect 27077 37349 27111 37383
rect 28641 37349 28675 37383
rect 31493 37349 31527 37383
rect 34069 37349 34103 37383
rect 40278 37349 40312 37383
rect 41889 37349 41923 37383
rect 11120 37281 11154 37315
rect 13680 37281 13714 37315
rect 15368 37281 15402 37315
rect 16589 37281 16623 37315
rect 17141 37281 17175 37315
rect 18153 37281 18187 37315
rect 18613 37281 18647 37315
rect 19844 37281 19878 37315
rect 24041 37281 24075 37315
rect 24593 37281 24627 37315
rect 30665 37281 30699 37315
rect 30849 37281 30883 37315
rect 33057 37281 33091 37315
rect 35725 37281 35759 37315
rect 35909 37281 35943 37315
rect 38393 37281 38427 37315
rect 38853 37281 38887 37315
rect 12173 37213 12207 37247
rect 12633 37213 12667 37247
rect 17325 37213 17359 37247
rect 18705 37213 18739 37247
rect 19533 37213 19567 37247
rect 21833 37213 21867 37247
rect 26985 37213 27019 37247
rect 27261 37213 27295 37247
rect 28549 37213 28583 37247
rect 28825 37213 28859 37247
rect 31125 37213 31159 37247
rect 32137 37213 32171 37247
rect 33977 37213 34011 37247
rect 34253 37213 34287 37247
rect 39129 37213 39163 37247
rect 39957 37213 39991 37247
rect 41797 37213 41831 37247
rect 42441 37213 42475 37247
rect 19947 37145 19981 37179
rect 23305 37145 23339 37179
rect 13783 37077 13817 37111
rect 19165 37077 19199 37111
rect 26709 37077 26743 37111
rect 33701 37077 33735 37111
rect 36829 37077 36863 37111
rect 12173 36873 12207 36907
rect 13461 36873 13495 36907
rect 16129 36873 16163 36907
rect 17049 36873 17083 36907
rect 18613 36873 18647 36907
rect 19901 36873 19935 36907
rect 21833 36873 21867 36907
rect 22937 36873 22971 36907
rect 24501 36873 24535 36907
rect 25927 36873 25961 36907
rect 31125 36873 31159 36907
rect 32689 36873 32723 36907
rect 34253 36873 34287 36907
rect 38025 36873 38059 36907
rect 38347 36873 38381 36907
rect 39037 36873 39071 36907
rect 41613 36873 41647 36907
rect 41935 36873 41969 36907
rect 13093 36805 13127 36839
rect 15761 36805 15795 36839
rect 26617 36805 26651 36839
rect 28457 36805 28491 36839
rect 33517 36805 33551 36839
rect 40923 36805 40957 36839
rect 11345 36737 11379 36771
rect 13645 36737 13679 36771
rect 13921 36737 13955 36771
rect 18705 36737 18739 36771
rect 20545 36737 20579 36771
rect 25145 36737 25179 36771
rect 25329 36737 25363 36771
rect 31401 36737 31435 36771
rect 31677 36737 31711 36771
rect 32965 36737 32999 36771
rect 36369 36737 36403 36771
rect 36645 36737 36679 36771
rect 36921 36737 36955 36771
rect 12608 36669 12642 36703
rect 19625 36669 19659 36703
rect 20269 36669 20303 36703
rect 22052 36669 22086 36703
rect 22477 36669 22511 36703
rect 23740 36669 23774 36703
rect 24133 36669 24167 36703
rect 24828 36669 24862 36703
rect 13737 36601 13771 36635
rect 14657 36601 14691 36635
rect 15209 36601 15243 36635
rect 15301 36601 15335 36635
rect 19026 36601 19060 36635
rect 20637 36601 20671 36635
rect 21189 36601 21223 36635
rect 23397 36601 23431 36635
rect 24915 36601 24949 36635
rect 25856 36669 25890 36703
rect 26065 36669 26099 36703
rect 27537 36669 27571 36703
rect 29561 36669 29595 36703
rect 34713 36669 34747 36703
rect 34897 36669 34931 36703
rect 35449 36669 35483 36703
rect 36001 36669 36035 36703
rect 38244 36669 38278 36703
rect 39272 36669 39306 36703
rect 40852 36669 40886 36703
rect 41245 36669 41279 36703
rect 41832 36669 41866 36703
rect 42257 36669 42291 36703
rect 11161 36533 11195 36567
rect 12679 36533 12713 36567
rect 15025 36533 15059 36567
rect 16589 36533 16623 36567
rect 17785 36533 17819 36567
rect 22155 36533 22189 36567
rect 23811 36533 23845 36567
rect 25145 36533 25179 36567
rect 26893 36601 26927 36635
rect 26985 36601 27019 36635
rect 29882 36601 29916 36635
rect 30849 36601 30883 36635
rect 31493 36601 31527 36635
rect 33057 36601 33091 36635
rect 33885 36601 33919 36635
rect 35633 36601 35667 36635
rect 36737 36601 36771 36635
rect 39359 36601 39393 36635
rect 39773 36601 39807 36635
rect 26065 36533 26099 36567
rect 26249 36533 26283 36567
rect 27813 36533 27847 36567
rect 29009 36533 29043 36567
rect 30481 36533 30515 36567
rect 32321 36533 32355 36567
rect 38669 36533 38703 36567
rect 40049 36533 40083 36567
rect 13645 36329 13679 36363
rect 14013 36329 14047 36363
rect 15439 36329 15473 36363
rect 16773 36329 16807 36363
rect 20545 36329 20579 36363
rect 26341 36329 26375 36363
rect 26847 36329 26881 36363
rect 27169 36329 27203 36363
rect 30757 36329 30791 36363
rect 32321 36329 32355 36363
rect 35633 36329 35667 36363
rect 36185 36329 36219 36363
rect 36737 36329 36771 36363
rect 40141 36329 40175 36363
rect 41797 36329 41831 36363
rect 12725 36261 12759 36295
rect 13277 36261 13311 36295
rect 18934 36261 18968 36295
rect 19901 36261 19935 36295
rect 22017 36261 22051 36295
rect 22569 36261 22603 36295
rect 28733 36261 28767 36295
rect 29882 36261 29916 36295
rect 32873 36261 32907 36295
rect 32965 36261 32999 36295
rect 37841 36261 37875 36295
rect 37933 36261 37967 36295
rect 40877 36261 40911 36295
rect 41429 36261 41463 36295
rect 10425 36193 10459 36227
rect 10885 36193 10919 36227
rect 14105 36193 14139 36227
rect 15209 36193 15243 36227
rect 18613 36193 18647 36227
rect 24041 36193 24075 36227
rect 24225 36193 24259 36227
rect 25456 36193 25490 36227
rect 26744 36193 26778 36227
rect 28273 36193 28307 36227
rect 28457 36193 28491 36227
rect 30481 36193 30515 36227
rect 31309 36193 31343 36227
rect 34345 36193 34379 36227
rect 39681 36193 39715 36227
rect 10977 36125 11011 36159
rect 12633 36125 12667 36159
rect 16405 36125 16439 36159
rect 21925 36125 21959 36159
rect 24317 36125 24351 36159
rect 25559 36125 25593 36159
rect 29009 36125 29043 36159
rect 29561 36125 29595 36159
rect 33149 36125 33183 36159
rect 35817 36125 35851 36159
rect 38117 36125 38151 36159
rect 40785 36125 40819 36159
rect 12081 35989 12115 36023
rect 14335 35989 14369 36023
rect 17325 35989 17359 36023
rect 18245 35989 18279 36023
rect 19533 35989 19567 36023
rect 24777 35989 24811 36023
rect 27721 35989 27755 36023
rect 34483 35989 34517 36023
rect 34989 35989 35023 36023
rect 37105 35989 37139 36023
rect 39819 35989 39853 36023
rect 42349 35989 42383 36023
rect 10425 35785 10459 35819
rect 11805 35785 11839 35819
rect 13461 35785 13495 35819
rect 16313 35785 16347 35819
rect 18337 35785 18371 35819
rect 18981 35785 19015 35819
rect 19441 35785 19475 35819
rect 21005 35785 21039 35819
rect 23121 35785 23155 35819
rect 23397 35785 23431 35819
rect 24225 35785 24259 35819
rect 25513 35785 25547 35819
rect 27077 35785 27111 35819
rect 27537 35785 27571 35819
rect 29101 35785 29135 35819
rect 30113 35785 30147 35819
rect 36461 35785 36495 35819
rect 37749 35785 37783 35819
rect 39681 35785 39715 35819
rect 41705 35785 41739 35819
rect 22477 35717 22511 35751
rect 28273 35717 28307 35751
rect 31585 35717 31619 35751
rect 34437 35717 34471 35751
rect 39221 35717 39255 35751
rect 14105 35649 14139 35683
rect 14381 35649 14415 35683
rect 14657 35649 14691 35683
rect 15945 35649 15979 35683
rect 16773 35649 16807 35683
rect 19625 35649 19659 35683
rect 19901 35649 19935 35683
rect 21925 35649 21959 35683
rect 24317 35649 24351 35683
rect 26157 35649 26191 35683
rect 26433 35649 26467 35683
rect 27721 35649 27755 35683
rect 28733 35649 28767 35683
rect 30665 35649 30699 35683
rect 31309 35649 31343 35683
rect 32045 35649 32079 35683
rect 32965 35649 32999 35683
rect 33241 35649 33275 35683
rect 35541 35649 35575 35683
rect 36737 35649 36771 35683
rect 38209 35649 38243 35683
rect 38485 35649 38519 35683
rect 40785 35649 40819 35683
rect 41429 35649 41463 35683
rect 42625 35649 42659 35683
rect 10149 35581 10183 35615
rect 11069 35581 11103 35615
rect 11345 35581 11379 35615
rect 11529 35581 11563 35615
rect 12541 35581 12575 35615
rect 13737 35581 13771 35615
rect 29320 35581 29354 35615
rect 29745 35581 29779 35615
rect 12265 35513 12299 35547
rect 12903 35513 12937 35547
rect 14473 35513 14507 35547
rect 16497 35513 16531 35547
rect 16589 35513 16623 35547
rect 18521 35513 18555 35547
rect 19717 35513 19751 35547
rect 21373 35513 21407 35547
rect 21741 35513 21775 35547
rect 22017 35513 22051 35547
rect 26249 35513 26283 35547
rect 27813 35513 27847 35547
rect 30757 35513 30791 35547
rect 32413 35513 32447 35547
rect 32781 35513 32815 35547
rect 33057 35513 33091 35547
rect 35449 35513 35483 35547
rect 35903 35513 35937 35547
rect 38301 35513 38335 35547
rect 40325 35513 40359 35547
rect 40877 35513 40911 35547
rect 42349 35513 42383 35547
rect 42441 35513 42475 35547
rect 15301 35445 15335 35479
rect 17417 35445 17451 35479
rect 24685 35445 24719 35479
rect 25237 35445 25271 35479
rect 25881 35445 25915 35479
rect 29423 35445 29457 35479
rect 37473 35445 37507 35479
rect 42073 35445 42107 35479
rect 10517 35241 10551 35275
rect 12173 35241 12207 35275
rect 12541 35241 12575 35275
rect 13553 35241 13587 35275
rect 14657 35241 14691 35275
rect 16773 35241 16807 35275
rect 17417 35241 17451 35275
rect 22017 35241 22051 35275
rect 24685 35241 24719 35275
rect 25237 35241 25271 35275
rect 26157 35241 26191 35275
rect 32873 35241 32907 35275
rect 37565 35241 37599 35275
rect 38669 35241 38703 35275
rect 40509 35241 40543 35275
rect 41153 35241 41187 35275
rect 11247 35173 11281 35207
rect 12995 35173 13029 35207
rect 15939 35173 15973 35207
rect 19441 35173 19475 35207
rect 21097 35173 21131 35207
rect 22661 35173 22695 35207
rect 25605 35173 25639 35207
rect 27261 35173 27295 35207
rect 29653 35173 29687 35207
rect 33149 35173 33183 35207
rect 35265 35173 35299 35207
rect 35909 35173 35943 35207
rect 38111 35173 38145 35207
rect 39951 35173 39985 35207
rect 40877 35173 40911 35207
rect 41521 35173 41555 35207
rect 10885 35105 10919 35139
rect 11805 35105 11839 35139
rect 14381 35105 14415 35139
rect 17325 35105 17359 35139
rect 17785 35105 17819 35139
rect 24317 35105 24351 35139
rect 29009 35105 29043 35139
rect 29469 35105 29503 35139
rect 30481 35105 30515 35139
rect 30941 35105 30975 35139
rect 34529 35105 34563 35139
rect 35081 35105 35115 35139
rect 36093 35105 36127 35139
rect 36553 35105 36587 35139
rect 42073 35105 42107 35139
rect 12633 35037 12667 35071
rect 15577 35037 15611 35071
rect 19165 35037 19199 35071
rect 19349 35037 19383 35071
rect 19625 35037 19659 35071
rect 21005 35037 21039 35071
rect 22569 35037 22603 35071
rect 22845 35037 22879 35071
rect 27169 35037 27203 35071
rect 31217 35037 31251 35071
rect 33057 35037 33091 35071
rect 33425 35037 33459 35071
rect 36829 35037 36863 35071
rect 37749 35037 37783 35071
rect 39589 35037 39623 35071
rect 41429 35037 41463 35071
rect 21557 34969 21591 35003
rect 27721 34969 27755 35003
rect 32413 34969 32447 35003
rect 37197 34969 37231 35003
rect 16497 34901 16531 34935
rect 23857 34901 23891 34935
rect 28181 34901 28215 34935
rect 11713 34697 11747 34731
rect 13093 34697 13127 34731
rect 14105 34697 14139 34731
rect 14473 34697 14507 34731
rect 18613 34697 18647 34731
rect 19257 34697 19291 34731
rect 19441 34697 19475 34731
rect 20545 34697 20579 34731
rect 21005 34697 21039 34731
rect 22937 34697 22971 34731
rect 24777 34697 24811 34731
rect 25237 34697 25271 34731
rect 29423 34697 29457 34731
rect 33333 34697 33367 34731
rect 38117 34697 38151 34731
rect 41429 34697 41463 34731
rect 41843 34697 41877 34731
rect 13369 34629 13403 34663
rect 15669 34629 15703 34663
rect 16773 34629 16807 34663
rect 11345 34561 11379 34595
rect 12173 34561 12207 34595
rect 14657 34561 14691 34595
rect 15301 34561 15335 34595
rect 16221 34561 16255 34595
rect 17785 34561 17819 34595
rect 10609 34493 10643 34527
rect 11069 34493 11103 34527
rect 12608 34493 12642 34527
rect 13620 34493 13654 34527
rect 18128 34493 18162 34527
rect 23397 34629 23431 34663
rect 29009 34629 29043 34663
rect 22293 34561 22327 34595
rect 24501 34561 24535 34595
rect 25421 34561 25455 34595
rect 26065 34561 26099 34595
rect 26709 34561 26743 34595
rect 27629 34561 27663 34595
rect 28641 34561 28675 34595
rect 31309 34561 31343 34595
rect 31677 34561 31711 34595
rect 32413 34561 32447 34595
rect 32689 34561 32723 34595
rect 35541 34561 35575 34595
rect 36921 34561 36955 34595
rect 37841 34561 37875 34595
rect 39589 34561 39623 34595
rect 40233 34561 40267 34595
rect 40693 34561 40727 34595
rect 19625 34493 19659 34527
rect 23765 34493 23799 34527
rect 24317 34493 24351 34527
rect 29352 34493 29386 34527
rect 34713 34493 34747 34527
rect 35265 34493 35299 34527
rect 35449 34493 35483 34527
rect 38853 34493 38887 34527
rect 39313 34493 39347 34527
rect 41772 34493 41806 34527
rect 42752 34493 42786 34527
rect 43177 34493 43211 34527
rect 14749 34425 14783 34459
rect 16313 34425 16347 34459
rect 19257 34425 19291 34459
rect 19946 34425 19980 34459
rect 21465 34425 21499 34459
rect 22017 34425 22051 34459
rect 22109 34425 22143 34459
rect 25513 34425 25547 34459
rect 27261 34425 27295 34459
rect 27353 34425 27387 34459
rect 30481 34425 30515 34459
rect 30665 34425 30699 34459
rect 30757 34425 30791 34459
rect 32505 34425 32539 34459
rect 34345 34425 34379 34459
rect 36645 34425 36679 34459
rect 36737 34425 36771 34459
rect 38669 34425 38703 34459
rect 10517 34357 10551 34391
rect 12679 34357 12713 34391
rect 13691 34357 13725 34391
rect 16037 34357 16071 34391
rect 17325 34357 17359 34391
rect 18199 34357 18233 34391
rect 19165 34357 19199 34391
rect 21833 34357 21867 34391
rect 26985 34357 27019 34391
rect 28181 34357 28215 34391
rect 29837 34357 29871 34391
rect 32137 34357 32171 34391
rect 33701 34357 33735 34391
rect 36093 34357 36127 34391
rect 39957 34357 39991 34391
rect 42257 34357 42291 34391
rect 42855 34357 42889 34391
rect 10977 34153 11011 34187
rect 14657 34153 14691 34187
rect 16313 34153 16347 34187
rect 16681 34153 16715 34187
rect 19257 34153 19291 34187
rect 19809 34153 19843 34187
rect 20085 34153 20119 34187
rect 21097 34153 21131 34187
rect 21833 34153 21867 34187
rect 22385 34153 22419 34187
rect 22661 34153 22695 34187
rect 24317 34153 24351 34187
rect 27077 34153 27111 34187
rect 30389 34153 30423 34187
rect 31033 34153 31067 34187
rect 33885 34153 33919 34187
rect 36461 34153 36495 34187
rect 37105 34153 37139 34187
rect 41429 34153 41463 34187
rect 10701 34085 10735 34119
rect 14381 34085 14415 34119
rect 15485 34085 15519 34119
rect 23857 34085 23891 34119
rect 27353 34085 27387 34119
rect 29790 34085 29824 34119
rect 30665 34085 30699 34119
rect 32458 34085 32492 34119
rect 35903 34085 35937 34119
rect 11897 34017 11931 34051
rect 13737 34017 13771 34051
rect 14197 34017 14231 34051
rect 16932 34017 16966 34051
rect 17944 34017 17978 34051
rect 24869 34017 24903 34051
rect 25329 34017 25363 34051
rect 32137 34017 32171 34051
rect 38071 34017 38105 34051
rect 39037 34017 39071 34051
rect 39497 34017 39531 34051
rect 40636 34017 40670 34051
rect 41705 34017 41739 34051
rect 42165 34017 42199 34051
rect 15393 33949 15427 33983
rect 18889 33949 18923 33983
rect 21465 33949 21499 33983
rect 25605 33949 25639 33983
rect 27261 33949 27295 33983
rect 29469 33949 29503 33983
rect 35541 33949 35575 33983
rect 38163 33949 38197 33983
rect 39773 33949 39807 33983
rect 42441 33949 42475 33983
rect 15945 33881 15979 33915
rect 18015 33881 18049 33915
rect 27813 33881 27847 33915
rect 34529 33881 34563 33915
rect 34989 33881 35023 33915
rect 36737 33881 36771 33915
rect 38853 33881 38887 33915
rect 12035 33813 12069 33847
rect 12449 33813 12483 33847
rect 17003 33813 17037 33847
rect 18429 33813 18463 33847
rect 33057 33813 33091 33847
rect 38485 33813 38519 33847
rect 40509 33813 40543 33847
rect 40739 33813 40773 33847
rect 43637 33813 43671 33847
rect 10517 33609 10551 33643
rect 11897 33609 11931 33643
rect 13737 33609 13771 33643
rect 14105 33609 14139 33643
rect 16037 33609 16071 33643
rect 17509 33609 17543 33643
rect 17877 33609 17911 33643
rect 19441 33609 19475 33643
rect 21925 33609 21959 33643
rect 22615 33609 22649 33643
rect 25605 33609 25639 33643
rect 26985 33609 27019 33643
rect 27353 33609 27387 33643
rect 27629 33609 27663 33643
rect 27951 33609 27985 33643
rect 30297 33609 30331 33643
rect 30849 33609 30883 33643
rect 30941 33609 30975 33643
rect 32045 33609 32079 33643
rect 32781 33609 32815 33643
rect 33885 33609 33919 33643
rect 36277 33609 36311 33643
rect 38853 33609 38887 33643
rect 39221 33609 39255 33643
rect 40325 33609 40359 33643
rect 40601 33609 40635 33643
rect 41705 33609 41739 33643
rect 42165 33609 42199 33643
rect 12541 33473 12575 33507
rect 14749 33473 14783 33507
rect 19073 33473 19107 33507
rect 19717 33473 19751 33507
rect 21649 33473 21683 33507
rect 22293 33473 22327 33507
rect 24041 33473 24075 33507
rect 24593 33473 24627 33507
rect 26065 33473 26099 33507
rect 10609 33405 10643 33439
rect 11069 33405 11103 33439
rect 17024 33405 17058 33439
rect 18337 33405 18371 33439
rect 18797 33405 18831 33439
rect 20821 33405 20855 33439
rect 21189 33405 21223 33439
rect 21373 33405 21407 33439
rect 22544 33405 22578 33439
rect 22937 33405 22971 33439
rect 25881 33405 25915 33439
rect 27848 33405 27882 33439
rect 28273 33405 28307 33439
rect 29101 33405 29135 33439
rect 29561 33405 29595 33439
rect 29837 33405 29871 33439
rect 39543 33541 39577 33575
rect 33333 33473 33367 33507
rect 36967 33473 37001 33507
rect 37933 33473 37967 33507
rect 38577 33473 38611 33507
rect 41337 33541 41371 33575
rect 40785 33473 40819 33507
rect 43637 33473 43671 33507
rect 31125 33405 31159 33439
rect 35868 33405 35902 33439
rect 36645 33405 36679 33439
rect 36864 33405 36898 33439
rect 37289 33405 37323 33439
rect 39440 33405 39474 33439
rect 39865 33405 39899 33439
rect 40601 33405 40635 33439
rect 42292 33405 42326 33439
rect 42717 33405 42751 33439
rect 11345 33337 11379 33371
rect 12633 33337 12667 33371
rect 13185 33337 13219 33371
rect 14841 33337 14875 33371
rect 15393 33337 15427 33371
rect 20453 33337 20487 33371
rect 24685 33337 24719 33371
rect 25237 33337 25271 33371
rect 26386 33337 26420 33371
rect 28733 33337 28767 33371
rect 30849 33337 30883 33371
rect 31446 33337 31480 33371
rect 32321 33337 32355 33371
rect 32954 33337 32988 33371
rect 33066 33337 33100 33371
rect 35955 33337 35989 33371
rect 38025 33337 38059 33371
rect 40877 33337 40911 33371
rect 42395 33337 42429 33371
rect 43453 33337 43487 33371
rect 43729 33337 43763 33371
rect 44281 33337 44315 33371
rect 14565 33269 14599 33303
rect 15669 33269 15703 33303
rect 17095 33269 17129 33303
rect 24409 33269 24443 33303
rect 29561 33269 29595 33303
rect 35633 33269 35667 33303
rect 37749 33269 37783 33303
rect 14749 33065 14783 33099
rect 15439 33065 15473 33099
rect 18061 33065 18095 33099
rect 24409 33065 24443 33099
rect 24961 33065 24995 33099
rect 26065 33065 26099 33099
rect 32229 33065 32263 33099
rect 33241 33065 33275 33099
rect 34897 33065 34931 33099
rect 43729 33065 43763 33099
rect 44281 33065 44315 33099
rect 11523 32997 11557 33031
rect 13461 32997 13495 33031
rect 13553 32997 13587 33031
rect 17135 32997 17169 33031
rect 18889 32997 18923 33031
rect 19717 32997 19751 33031
rect 23851 32997 23885 33031
rect 26709 32997 26743 33031
rect 28825 32997 28859 33031
rect 34069 32997 34103 33031
rect 38070 32997 38104 33031
rect 40094 32997 40128 33031
rect 41705 32997 41739 33031
rect 15368 32929 15402 32963
rect 19073 32929 19107 32963
rect 19441 32929 19475 32963
rect 22201 32929 22235 32963
rect 22477 32929 22511 32963
rect 25145 32929 25179 32963
rect 28089 32929 28123 32963
rect 30481 32929 30515 32963
rect 30757 32929 30791 32963
rect 30941 32929 30975 32963
rect 31217 32929 31251 32963
rect 32413 32929 32447 32963
rect 32689 32929 32723 32963
rect 36277 32929 36311 32963
rect 36553 32929 36587 32963
rect 39037 32929 39071 32963
rect 43361 32929 43395 32963
rect 10149 32861 10183 32895
rect 11161 32861 11195 32895
rect 13737 32861 13771 32895
rect 16773 32861 16807 32895
rect 22661 32861 22695 32895
rect 23489 32861 23523 32895
rect 26617 32861 26651 32895
rect 26893 32861 26927 32895
rect 28457 32861 28491 32895
rect 36829 32861 36863 32895
rect 37749 32861 37783 32895
rect 39773 32861 39807 32895
rect 41613 32861 41647 32895
rect 42257 32861 42291 32895
rect 45109 32861 45143 32895
rect 28365 32793 28399 32827
rect 38669 32793 38703 32827
rect 10701 32725 10735 32759
rect 12081 32725 12115 32759
rect 12541 32725 12575 32759
rect 17693 32725 17727 32759
rect 18337 32725 18371 32759
rect 21373 32725 21407 32759
rect 25375 32725 25409 32759
rect 25697 32725 25731 32759
rect 27721 32725 27755 32759
rect 28254 32725 28288 32759
rect 29285 32725 29319 32759
rect 29929 32725 29963 32759
rect 31585 32725 31619 32759
rect 34299 32725 34333 32759
rect 40693 32725 40727 32759
rect 40969 32725 41003 32759
rect 41337 32725 41371 32759
rect 12173 32521 12207 32555
rect 13829 32521 13863 32555
rect 17509 32521 17543 32555
rect 21741 32521 21775 32555
rect 22661 32521 22695 32555
rect 22845 32521 22879 32555
rect 23838 32521 23872 32555
rect 24317 32521 24351 32555
rect 27905 32521 27939 32555
rect 29009 32521 29043 32555
rect 32781 32521 32815 32555
rect 34253 32521 34287 32555
rect 37197 32521 37231 32555
rect 37841 32521 37875 32555
rect 40141 32521 40175 32555
rect 42625 32521 42659 32555
rect 43637 32521 43671 32555
rect 44833 32521 44867 32555
rect 10517 32453 10551 32487
rect 11897 32453 11931 32487
rect 13553 32453 13587 32487
rect 21557 32453 21591 32487
rect 12541 32385 12575 32419
rect 13185 32385 13219 32419
rect 15393 32385 15427 32419
rect 16497 32385 16531 32419
rect 18429 32385 18463 32419
rect 20361 32385 20395 32419
rect 21649 32385 21683 32419
rect 10149 32317 10183 32351
rect 10609 32317 10643 32351
rect 11529 32317 11563 32351
rect 19533 32317 19567 32351
rect 20269 32317 20303 32351
rect 20821 32317 20855 32351
rect 21428 32317 21462 32351
rect 23121 32453 23155 32487
rect 23949 32453 23983 32487
rect 29469 32453 29503 32487
rect 39865 32453 39899 32487
rect 44373 32453 44407 32487
rect 23489 32385 23523 32419
rect 24041 32385 24075 32419
rect 25237 32385 25271 32419
rect 27997 32385 28031 32419
rect 29929 32385 29963 32419
rect 34989 32385 35023 32419
rect 35449 32385 35483 32419
rect 38485 32385 38519 32419
rect 39129 32385 39163 32419
rect 43821 32385 43855 32419
rect 27776 32317 27810 32351
rect 31309 32317 31343 32351
rect 31677 32317 31711 32351
rect 31953 32317 31987 32351
rect 37448 32317 37482 32351
rect 42752 32317 42786 32351
rect 43177 32317 43211 32351
rect 10971 32249 11005 32283
rect 12633 32249 12667 32283
rect 14749 32249 14783 32283
rect 14841 32249 14875 32283
rect 16313 32249 16347 32283
rect 16589 32249 16623 32283
rect 17141 32249 17175 32283
rect 17785 32249 17819 32283
rect 18153 32249 18187 32283
rect 18245 32249 18279 32283
rect 21281 32249 21315 32283
rect 22845 32249 22879 32283
rect 23673 32249 23707 32283
rect 24685 32249 24719 32283
rect 27169 32249 27203 32283
rect 27629 32249 27663 32283
rect 28365 32249 28399 32283
rect 30021 32249 30055 32283
rect 30573 32249 30607 32283
rect 32137 32249 32171 32283
rect 35081 32249 35115 32283
rect 38577 32249 38611 32283
rect 41061 32249 41095 32283
rect 41153 32249 41187 32283
rect 41705 32249 41739 32283
rect 43913 32249 43947 32283
rect 14565 32181 14599 32215
rect 15761 32181 15795 32215
rect 19165 32181 19199 32215
rect 21097 32181 21131 32215
rect 22293 32181 22327 32215
rect 25145 32181 25179 32215
rect 25605 32181 25639 32215
rect 26157 32181 26191 32215
rect 26709 32181 26743 32215
rect 27445 32181 27479 32215
rect 28641 32181 28675 32215
rect 30941 32181 30975 32215
rect 32505 32181 32539 32215
rect 32965 32181 32999 32215
rect 34621 32181 34655 32215
rect 36185 32181 36219 32215
rect 36553 32181 36587 32215
rect 37519 32181 37553 32215
rect 38209 32181 38243 32215
rect 39405 32181 39439 32215
rect 40877 32181 40911 32215
rect 41981 32181 42015 32215
rect 42855 32181 42889 32215
rect 10517 31977 10551 32011
rect 11437 31977 11471 32011
rect 12633 31977 12667 32011
rect 13001 31977 13035 32011
rect 16497 31977 16531 32011
rect 18245 31977 18279 32011
rect 23305 31977 23339 32011
rect 23765 31977 23799 32011
rect 24041 31977 24075 32011
rect 25789 31977 25823 32011
rect 26341 31977 26375 32011
rect 26985 31977 27019 32011
rect 30757 31977 30791 32011
rect 31493 31977 31527 32011
rect 32505 31977 32539 32011
rect 38945 31977 38979 32011
rect 39819 31977 39853 32011
rect 41705 31977 41739 32011
rect 45155 31977 45189 32011
rect 13277 31909 13311 31943
rect 15485 31909 15519 31943
rect 17141 31909 17175 31943
rect 17233 31909 17267 31943
rect 18797 31909 18831 31943
rect 19257 31909 19291 31943
rect 25145 31909 25179 31943
rect 28457 31909 28491 31943
rect 29929 31909 29963 31943
rect 34621 31909 34655 31943
rect 36093 31909 36127 31943
rect 36185 31909 36219 31943
rect 38025 31909 38059 31943
rect 38117 31909 38151 31943
rect 40877 31909 40911 31943
rect 43637 31909 43671 31943
rect 10425 31841 10459 31875
rect 10885 31841 10919 31875
rect 12132 31841 12166 31875
rect 19993 31841 20027 31875
rect 21132 31841 21166 31875
rect 22385 31841 22419 31875
rect 22661 31841 22695 31875
rect 24409 31841 24443 31875
rect 24961 31841 24995 31875
rect 26433 31841 26467 31875
rect 27721 31841 27755 31875
rect 28733 31841 28767 31875
rect 39748 31841 39782 31875
rect 42257 31841 42291 31875
rect 45017 31841 45051 31875
rect 12219 31773 12253 31807
rect 13185 31773 13219 31807
rect 15393 31773 15427 31807
rect 17417 31773 17451 31807
rect 19625 31773 19659 31807
rect 22477 31773 22511 31807
rect 28089 31773 28123 31807
rect 29837 31773 29871 31807
rect 32137 31773 32171 31807
rect 34529 31773 34563 31807
rect 34805 31773 34839 31807
rect 36369 31773 36403 31807
rect 38393 31773 38427 31807
rect 40785 31773 40819 31807
rect 41153 31773 41187 31807
rect 42395 31773 42429 31807
rect 43545 31773 43579 31807
rect 44189 31773 44223 31807
rect 13737 31705 13771 31739
rect 15945 31705 15979 31739
rect 19165 31705 19199 31739
rect 19533 31705 19567 31739
rect 21235 31705 21269 31739
rect 27629 31705 27663 31739
rect 30389 31705 30423 31739
rect 44465 31705 44499 31739
rect 14657 31637 14691 31671
rect 16865 31637 16899 31671
rect 19422 31637 19456 31671
rect 20361 31637 20395 31671
rect 21557 31637 21591 31671
rect 25421 31637 25455 31671
rect 26663 31637 26697 31671
rect 27859 31637 27893 31671
rect 27997 31637 28031 31671
rect 29285 31637 29319 31671
rect 33057 31637 33091 31671
rect 35449 31637 35483 31671
rect 11483 31433 11517 31467
rect 13461 31433 13495 31467
rect 13829 31433 13863 31467
rect 15393 31433 15427 31467
rect 17417 31433 17451 31467
rect 19993 31433 20027 31467
rect 21649 31433 21683 31467
rect 23029 31433 23063 31467
rect 26617 31433 26651 31467
rect 30205 31433 30239 31467
rect 30481 31433 30515 31467
rect 31171 31433 31205 31467
rect 34253 31433 34287 31467
rect 36645 31433 36679 31467
rect 38025 31433 38059 31467
rect 40325 31433 40359 31467
rect 41659 31433 41693 31467
rect 42625 31433 42659 31467
rect 43085 31433 43119 31467
rect 43453 31433 43487 31467
rect 17785 31365 17819 31399
rect 19809 31365 19843 31399
rect 20821 31365 20855 31399
rect 22569 31365 22603 31399
rect 36001 31365 36035 31399
rect 44189 31365 44223 31399
rect 12541 31297 12575 31331
rect 14611 31297 14645 31331
rect 15669 31297 15703 31331
rect 17049 31297 17083 31331
rect 18981 31297 19015 31331
rect 19349 31297 19383 31331
rect 19901 31297 19935 31331
rect 25329 31297 25363 31331
rect 28365 31297 28399 31331
rect 29285 31297 29319 31331
rect 32137 31297 32171 31331
rect 35449 31297 35483 31331
rect 37381 31297 37415 31331
rect 43637 31297 43671 31331
rect 44557 31297 44591 31331
rect 11412 31229 11446 31263
rect 14524 31229 14558 31263
rect 16405 31229 16439 31263
rect 16865 31229 16899 31263
rect 18153 31229 18187 31263
rect 18337 31229 18371 31263
rect 19680 31229 19714 31263
rect 21557 31229 21591 31263
rect 22201 31229 22235 31263
rect 23489 31229 23523 31263
rect 23857 31229 23891 31263
rect 24961 31229 24995 31263
rect 27905 31229 27939 31263
rect 28181 31229 28215 31263
rect 30941 31229 30975 31263
rect 31068 31229 31102 31263
rect 36829 31229 36863 31263
rect 37289 31229 37323 31263
rect 38301 31229 38335 31263
rect 38853 31229 38887 31263
rect 39313 31229 39347 31263
rect 40544 31229 40578 31263
rect 40969 31229 41003 31263
rect 41556 31229 41590 31263
rect 45109 31229 45143 31263
rect 12633 31161 12667 31195
rect 13185 31161 13219 31195
rect 16313 31161 16347 31195
rect 18705 31161 18739 31195
rect 19533 31161 19567 31195
rect 21281 31161 21315 31195
rect 21373 31161 21407 31195
rect 23673 31161 23707 31195
rect 24593 31161 24627 31195
rect 25421 31161 25455 31195
rect 25973 31161 26007 31195
rect 27169 31161 27203 31195
rect 29647 31161 29681 31195
rect 32458 31161 32492 31195
rect 34621 31161 34655 31195
rect 34989 31161 35023 31195
rect 35081 31161 35115 31195
rect 38669 31161 38703 31195
rect 39589 31161 39623 31195
rect 40647 31161 40681 31195
rect 43729 31161 43763 31195
rect 10425 31093 10459 31127
rect 10793 31093 10827 31127
rect 11805 31093 11839 31127
rect 12265 31093 12299 31127
rect 14933 31093 14967 31127
rect 23949 31093 23983 31127
rect 27537 31093 27571 31127
rect 28733 31093 28767 31127
rect 29009 31093 29043 31127
rect 31585 31093 31619 31127
rect 31953 31093 31987 31127
rect 33057 31093 33091 31127
rect 33977 31093 34011 31127
rect 39865 31093 39899 31127
rect 41337 31093 41371 31127
rect 42349 31093 42383 31127
rect 13737 30889 13771 30923
rect 17049 30889 17083 30923
rect 18429 30889 18463 30923
rect 19073 30889 19107 30923
rect 20453 30889 20487 30923
rect 24501 30889 24535 30923
rect 28457 30889 28491 30923
rect 32321 30889 32355 30923
rect 32689 30889 32723 30923
rect 36231 30889 36265 30923
rect 37933 30889 37967 30923
rect 41245 30889 41279 30923
rect 41705 30889 41739 30923
rect 42395 30889 42429 30923
rect 11989 30821 12023 30855
rect 12541 30821 12575 30855
rect 15485 30821 15519 30855
rect 16037 30821 16071 30855
rect 17601 30821 17635 30855
rect 18889 30821 18923 30855
rect 22937 30821 22971 30855
rect 24869 30821 24903 30855
rect 25421 30821 25455 30855
rect 30205 30821 30239 30855
rect 33057 30821 33091 30855
rect 33149 30821 33183 30855
rect 34713 30821 34747 30855
rect 35265 30821 35299 30855
rect 36001 30821 36035 30855
rect 36829 30821 36863 30855
rect 38485 30821 38519 30855
rect 40417 30821 40451 30855
rect 43545 30821 43579 30855
rect 44097 30821 44131 30855
rect 45017 30821 45051 30855
rect 45109 30821 45143 30855
rect 10517 30753 10551 30787
rect 10701 30753 10735 30787
rect 14248 30753 14282 30787
rect 18981 30753 19015 30787
rect 19441 30753 19475 30787
rect 19993 30753 20027 30787
rect 21189 30753 21223 30787
rect 21649 30753 21683 30787
rect 27077 30753 27111 30787
rect 28089 30753 28123 30787
rect 29009 30753 29043 30787
rect 36160 30753 36194 30787
rect 42292 30753 42326 30787
rect 10793 30685 10827 30719
rect 11897 30685 11931 30719
rect 14335 30685 14369 30719
rect 15393 30685 15427 30719
rect 17509 30685 17543 30719
rect 21925 30685 21959 30719
rect 22845 30685 22879 30719
rect 23489 30685 23523 30719
rect 24133 30685 24167 30719
rect 24777 30685 24811 30719
rect 27445 30685 27479 30719
rect 27813 30685 27847 30719
rect 30113 30685 30147 30719
rect 30757 30685 30791 30719
rect 33701 30685 33735 30719
rect 34437 30685 34471 30719
rect 34621 30685 34655 30719
rect 38393 30685 38427 30719
rect 38669 30685 38703 30719
rect 40325 30685 40359 30719
rect 43453 30685 43487 30719
rect 45293 30685 45327 30719
rect 18061 30617 18095 30651
rect 29745 30617 29779 30651
rect 40877 30617 40911 30651
rect 12817 30549 12851 30583
rect 16405 30549 16439 30583
rect 22201 30549 22235 30583
rect 25789 30549 25823 30583
rect 27215 30549 27249 30583
rect 27353 30549 27387 30583
rect 29147 30549 29181 30583
rect 31033 30549 31067 30583
rect 35541 30549 35575 30583
rect 44465 30549 44499 30583
rect 11529 30345 11563 30379
rect 13185 30345 13219 30379
rect 14657 30345 14691 30379
rect 17325 30345 17359 30379
rect 17601 30345 17635 30379
rect 19993 30345 20027 30379
rect 20637 30345 20671 30379
rect 20959 30345 20993 30379
rect 22753 30345 22787 30379
rect 23029 30345 23063 30379
rect 23811 30345 23845 30379
rect 25789 30345 25823 30379
rect 25973 30345 26007 30379
rect 28319 30345 28353 30379
rect 29791 30345 29825 30379
rect 30481 30345 30515 30379
rect 32689 30345 32723 30379
rect 33057 30345 33091 30379
rect 36185 30345 36219 30379
rect 37289 30345 37323 30379
rect 38301 30345 38335 30379
rect 38577 30345 38611 30379
rect 40325 30345 40359 30379
rect 42855 30345 42889 30379
rect 46259 30345 46293 30379
rect 46581 30345 46615 30379
rect 9735 30277 9769 30311
rect 12173 30277 12207 30311
rect 14933 30277 14967 30311
rect 15025 30277 15059 30311
rect 15853 30277 15887 30311
rect 21649 30277 21683 30311
rect 23397 30277 23431 30311
rect 10609 30209 10643 30243
rect 11805 30209 11839 30243
rect 12771 30209 12805 30243
rect 9664 30141 9698 30175
rect 12684 30141 12718 30175
rect 14381 30141 14415 30175
rect 15301 30209 15335 30243
rect 16589 30209 16623 30243
rect 18797 30209 18831 30243
rect 24777 30209 24811 30243
rect 16840 30141 16874 30175
rect 20888 30141 20922 30175
rect 21373 30141 21407 30175
rect 21833 30141 21867 30175
rect 23581 30141 23615 30175
rect 25421 30141 25455 30175
rect 39037 30277 39071 30311
rect 42257 30277 42291 30311
rect 44373 30277 44407 30311
rect 45477 30277 45511 30311
rect 26341 30209 26375 30243
rect 26617 30209 26651 30243
rect 29101 30209 29135 30243
rect 30849 30209 30883 30243
rect 34989 30209 35023 30243
rect 35357 30209 35391 30243
rect 37381 30209 37415 30243
rect 39267 30209 39301 30243
rect 41245 30209 41279 30243
rect 43821 30209 43855 30243
rect 44833 30209 44867 30243
rect 45109 30209 45143 30243
rect 28248 30141 28282 30175
rect 29688 30141 29722 30175
rect 30113 30141 30147 30175
rect 39164 30141 39198 30175
rect 39589 30141 39623 30175
rect 42784 30141 42818 30175
rect 43177 30141 43211 30175
rect 46188 30141 46222 30175
rect 10517 30073 10551 30107
rect 10971 30073 11005 30107
rect 13737 30073 13771 30107
rect 13829 30073 13863 30107
rect 14933 30073 14967 30107
rect 15393 30073 15427 30107
rect 18705 30073 18739 30107
rect 19159 30073 19193 30107
rect 22154 30073 22188 30107
rect 24501 30073 24535 30107
rect 24869 30073 24903 30107
rect 25973 30073 26007 30107
rect 26433 30073 26467 30107
rect 30941 30073 30975 30107
rect 31493 30073 31527 30107
rect 33333 30073 33367 30107
rect 33425 30073 33459 30107
rect 33977 30073 34011 30107
rect 35081 30073 35115 30107
rect 37743 30073 37777 30107
rect 41337 30073 41371 30107
rect 41889 30073 41923 30107
rect 43637 30073 43671 30107
rect 43913 30073 43947 30107
rect 9505 30005 9539 30039
rect 10057 30005 10091 30039
rect 13553 30005 13587 30039
rect 16221 30005 16255 30039
rect 16911 30005 16945 30039
rect 18337 30005 18371 30039
rect 19717 30005 19751 30039
rect 24225 30005 24259 30039
rect 26065 30005 26099 30039
rect 27353 30005 27387 30039
rect 27629 30005 27663 30039
rect 28733 30005 28767 30039
rect 34529 30005 34563 30039
rect 41061 30005 41095 30039
rect 10425 29801 10459 29835
rect 10793 29801 10827 29835
rect 11805 29801 11839 29835
rect 13921 29801 13955 29835
rect 15025 29801 15059 29835
rect 17325 29801 17359 29835
rect 17877 29801 17911 29835
rect 18613 29801 18647 29835
rect 22569 29801 22603 29835
rect 23121 29801 23155 29835
rect 24961 29801 24995 29835
rect 25513 29801 25547 29835
rect 26663 29801 26697 29835
rect 27537 29801 27571 29835
rect 30113 29801 30147 29835
rect 33609 29801 33643 29835
rect 34989 29801 35023 29835
rect 37013 29801 37047 29835
rect 37381 29801 37415 29835
rect 40417 29801 40451 29835
rect 40785 29801 40819 29835
rect 42165 29801 42199 29835
rect 43729 29801 43763 29835
rect 44281 29801 44315 29835
rect 11247 29733 11281 29767
rect 13363 29733 13397 29767
rect 15485 29733 15519 29767
rect 18153 29733 18187 29767
rect 18889 29733 18923 29767
rect 24133 29733 24167 29767
rect 26341 29733 26375 29767
rect 30389 29733 30423 29767
rect 34069 29733 34103 29767
rect 34161 29733 34195 29767
rect 38070 29733 38104 29767
rect 39818 29733 39852 29767
rect 41566 29733 41600 29767
rect 43177 29733 43211 29767
rect 21224 29665 21258 29699
rect 21327 29665 21361 29699
rect 26433 29665 26467 29699
rect 28365 29665 28399 29699
rect 28733 29665 28767 29699
rect 32137 29665 32171 29699
rect 32597 29665 32631 29699
rect 33333 29665 33367 29699
rect 35541 29665 35575 29699
rect 36588 29665 36622 29699
rect 39497 29665 39531 29699
rect 45109 29665 45143 29699
rect 9781 29597 9815 29631
rect 10885 29597 10919 29631
rect 13001 29597 13035 29631
rect 15393 29597 15427 29631
rect 16957 29597 16991 29631
rect 18797 29597 18831 29631
rect 19073 29597 19107 29631
rect 22201 29597 22235 29631
rect 24041 29597 24075 29631
rect 24317 29597 24351 29631
rect 28917 29597 28951 29631
rect 30297 29597 30331 29631
rect 30573 29597 30607 29631
rect 32873 29597 32907 29631
rect 34345 29597 34379 29631
rect 37749 29597 37783 29631
rect 41245 29597 41279 29631
rect 43361 29597 43395 29631
rect 15945 29529 15979 29563
rect 27077 29529 27111 29563
rect 31309 29529 31343 29563
rect 10011 29461 10045 29495
rect 12541 29461 12575 29495
rect 20269 29461 20303 29495
rect 21649 29461 21683 29495
rect 22017 29461 22051 29495
rect 29285 29461 29319 29495
rect 35357 29461 35391 29495
rect 35679 29461 35713 29495
rect 36691 29461 36725 29495
rect 38669 29461 38703 29495
rect 45247 29461 45281 29495
rect 10149 29257 10183 29291
rect 12265 29257 12299 29291
rect 13461 29257 13495 29291
rect 14657 29257 14691 29291
rect 15577 29257 15611 29291
rect 18521 29257 18555 29291
rect 18889 29257 18923 29291
rect 19625 29257 19659 29291
rect 20315 29257 20349 29291
rect 22569 29257 22603 29291
rect 24317 29257 24351 29291
rect 28273 29257 28307 29291
rect 28641 29257 28675 29291
rect 32597 29257 32631 29291
rect 34069 29257 34103 29291
rect 34621 29257 34655 29291
rect 40233 29257 40267 29291
rect 44833 29257 44867 29291
rect 11345 29189 11379 29223
rect 19257 29189 19291 29223
rect 20453 29189 20487 29223
rect 10977 29121 11011 29155
rect 11621 29121 11655 29155
rect 13001 29121 13035 29155
rect 13829 29121 13863 29155
rect 17141 29121 17175 29155
rect 17785 29121 17819 29155
rect 19993 29121 20027 29155
rect 20545 29121 20579 29155
rect 21189 29121 21223 29155
rect 10241 29053 10275 29087
rect 10793 29053 10827 29087
rect 12449 29053 12483 29087
rect 12909 29053 12943 29087
rect 14784 29053 14818 29087
rect 15209 29053 15243 29087
rect 16221 29053 16255 29087
rect 16405 29053 16439 29087
rect 16865 29053 16899 29087
rect 18128 29053 18162 29087
rect 21741 29053 21775 29087
rect 22201 29053 22235 29087
rect 39865 29189 39899 29223
rect 44373 29189 44407 29223
rect 22753 29121 22787 29155
rect 24041 29121 24075 29155
rect 26065 29121 26099 29155
rect 27077 29121 27111 29155
rect 31125 29121 31159 29155
rect 31401 29121 31435 29155
rect 32873 29121 32907 29155
rect 34989 29121 35023 29155
rect 35449 29121 35483 29155
rect 37381 29121 37415 29155
rect 37841 29121 37875 29155
rect 38577 29121 38611 29155
rect 39497 29121 39531 29155
rect 42717 29121 42751 29155
rect 42809 29121 42843 29155
rect 43821 29121 43855 29155
rect 26985 29053 27019 29087
rect 27721 29053 27755 29087
rect 29285 29053 29319 29087
rect 30205 29053 30239 29087
rect 30849 29053 30883 29087
rect 36645 29053 36679 29087
rect 37105 29053 37139 29087
rect 40509 29053 40543 29087
rect 40969 29053 41003 29087
rect 41981 29053 42015 29087
rect 42073 29053 42107 29087
rect 42533 29053 42567 29087
rect 9781 28985 9815 29019
rect 17417 28985 17451 29019
rect 20177 28985 20211 29019
rect 20913 28985 20947 29019
rect 22569 28985 22603 29019
rect 25605 28985 25639 29019
rect 25697 28985 25731 29019
rect 26617 28985 26651 29019
rect 29606 28985 29640 29019
rect 31217 28985 31251 29019
rect 32965 28985 32999 29019
rect 33517 28985 33551 29019
rect 35081 28985 35115 29019
rect 36461 28985 36495 29019
rect 38301 28985 38335 29019
rect 38393 28985 38427 29019
rect 41245 28985 41279 29019
rect 43913 28985 43947 29019
rect 14887 28917 14921 28951
rect 18199 28917 18233 28951
rect 21557 28917 21591 28951
rect 21833 28917 21867 28951
rect 24501 28917 24535 28951
rect 25329 28917 25363 28951
rect 29009 28917 29043 28951
rect 30481 28917 30515 28951
rect 32137 28917 32171 28951
rect 35909 28917 35943 28951
rect 41521 28917 41555 28951
rect 43361 28917 43395 28951
rect 45109 28917 45143 28951
rect 9873 28713 9907 28747
rect 15025 28713 15059 28747
rect 16405 28713 16439 28747
rect 21557 28713 21591 28747
rect 22385 28713 22419 28747
rect 29285 28713 29319 28747
rect 30113 28713 30147 28747
rect 30665 28713 30699 28747
rect 31309 28713 31343 28747
rect 31953 28713 31987 28747
rect 33425 28713 33459 28747
rect 33977 28713 34011 28747
rect 37105 28713 37139 28747
rect 37565 28713 37599 28747
rect 38485 28713 38519 28747
rect 39589 28713 39623 28747
rect 41337 28713 41371 28747
rect 42441 28713 42475 28747
rect 43913 28713 43947 28747
rect 12173 28645 12207 28679
rect 15393 28645 15427 28679
rect 15485 28645 15519 28679
rect 17325 28645 17359 28679
rect 23121 28645 23155 28679
rect 25053 28645 25087 28679
rect 25605 28645 25639 28679
rect 26709 28645 26743 28679
rect 28917 28645 28951 28679
rect 34253 28645 34287 28679
rect 34989 28645 35023 28679
rect 35541 28645 35575 28679
rect 38761 28645 38795 28679
rect 44189 28645 44223 28679
rect 10333 28577 10367 28611
rect 10793 28577 10827 28611
rect 14197 28577 14231 28611
rect 18740 28577 18774 28611
rect 22109 28577 22143 28611
rect 28181 28577 28215 28611
rect 28733 28577 28767 28611
rect 30941 28577 30975 28611
rect 33057 28577 33091 28611
rect 36712 28577 36746 28611
rect 37968 28577 38002 28611
rect 38996 28577 39030 28611
rect 40601 28577 40635 28611
rect 40785 28577 40819 28611
rect 41956 28577 41990 28611
rect 43269 28577 43303 28611
rect 44408 28577 44442 28611
rect 10885 28509 10919 28543
rect 12081 28509 12115 28543
rect 12725 28509 12759 28543
rect 15669 28509 15703 28543
rect 17233 28509 17267 28543
rect 17601 28509 17635 28543
rect 21189 28509 21223 28543
rect 23029 28509 23063 28543
rect 23305 28509 23339 28543
rect 24777 28509 24811 28543
rect 24961 28509 24995 28543
rect 26617 28509 26651 28543
rect 26893 28509 26927 28543
rect 29745 28509 29779 28543
rect 34897 28509 34931 28543
rect 41061 28509 41095 28543
rect 19947 28441 19981 28475
rect 36783 28441 36817 28475
rect 11345 28373 11379 28407
rect 14335 28373 14369 28407
rect 18153 28373 18187 28407
rect 18843 28373 18877 28407
rect 19717 28373 19751 28407
rect 20361 28373 20395 28407
rect 32321 28373 32355 28407
rect 32873 28373 32907 28407
rect 38071 28373 38105 28407
rect 39083 28373 39117 28407
rect 41705 28373 41739 28407
rect 42027 28373 42061 28407
rect 43499 28373 43533 28407
rect 44511 28373 44545 28407
rect 16497 28169 16531 28203
rect 22753 28169 22787 28203
rect 23121 28169 23155 28203
rect 24455 28169 24489 28203
rect 27031 28169 27065 28203
rect 30205 28169 30239 28203
rect 31263 28169 31297 28203
rect 33701 28169 33735 28203
rect 34253 28169 34287 28203
rect 34621 28169 34655 28203
rect 35909 28169 35943 28203
rect 37197 28169 37231 28203
rect 39313 28169 39347 28203
rect 40693 28169 40727 28203
rect 41153 28169 41187 28203
rect 43361 28169 43395 28203
rect 44649 28169 44683 28203
rect 19809 28101 19843 28135
rect 24225 28101 24259 28135
rect 25237 28101 25271 28135
rect 26525 28101 26559 28135
rect 33057 28101 33091 28135
rect 33425 28101 33459 28135
rect 10517 28033 10551 28067
rect 12081 28033 12115 28067
rect 13001 28033 13035 28067
rect 13829 28033 13863 28067
rect 21189 28033 21223 28067
rect 21833 28033 21867 28067
rect 25421 28033 25455 28067
rect 28043 28033 28077 28067
rect 29285 28033 29319 28067
rect 31953 28033 31987 28067
rect 34989 28033 35023 28067
rect 37427 28033 37461 28067
rect 38393 28033 38427 28067
rect 39681 28033 39715 28067
rect 41337 28033 41371 28067
rect 43085 28033 43119 28067
rect 43729 28033 43763 28067
rect 44005 28033 44039 28067
rect 9572 27965 9606 27999
rect 14289 27965 14323 27999
rect 17024 27965 17058 27999
rect 17509 27965 17543 27999
rect 18153 27965 18187 27999
rect 20453 27965 20487 27999
rect 21005 27965 21039 27999
rect 22360 27965 22394 27999
rect 24384 27965 24418 27999
rect 26065 27965 26099 27999
rect 27353 27965 27387 27999
rect 27956 27965 27990 27999
rect 31192 27965 31226 27999
rect 32137 27965 32171 27999
rect 37340 27965 37374 27999
rect 42257 27965 42291 27999
rect 10425 27897 10459 27931
rect 10879 27897 10913 27931
rect 13185 27897 13219 27931
rect 13277 27897 13311 27931
rect 15117 27897 15151 27931
rect 15209 27897 15243 27931
rect 15761 27897 15795 27931
rect 16865 27897 16899 27931
rect 19349 27897 19383 27931
rect 25513 27897 25547 27931
rect 26801 27897 26835 27931
rect 29647 27897 29681 27931
rect 30849 27897 30883 27931
rect 32458 27897 32492 27931
rect 35081 27897 35115 27931
rect 35633 27897 35667 27931
rect 38209 27897 38243 27931
rect 38485 27897 38519 27931
rect 39037 27897 39071 27931
rect 41658 27897 41692 27931
rect 43821 27897 43855 27931
rect 9643 27829 9677 27863
rect 10057 27829 10091 27863
rect 11437 27829 11471 27863
rect 14841 27829 14875 27863
rect 16037 27829 16071 27863
rect 17095 27829 17129 27863
rect 17877 27829 17911 27863
rect 18521 27829 18555 27863
rect 19073 27829 19107 27863
rect 20269 27829 20303 27863
rect 21465 27829 21499 27863
rect 22431 27829 22465 27863
rect 24869 27829 24903 27863
rect 27813 27829 27847 27863
rect 28365 27829 28399 27863
rect 29009 27829 29043 27863
rect 30481 27829 30515 27863
rect 31677 27829 31711 27863
rect 36737 27829 36771 27863
rect 37841 27829 37875 27863
rect 40233 27829 40267 27863
rect 42533 27829 42567 27863
rect 12449 27625 12483 27659
rect 23673 27625 23707 27659
rect 25605 27625 25639 27659
rect 26709 27625 26743 27659
rect 32229 27625 32263 27659
rect 35173 27625 35207 27659
rect 38117 27625 38151 27659
rect 38669 27625 38703 27659
rect 38945 27625 38979 27659
rect 41521 27625 41555 27659
rect 42349 27625 42383 27659
rect 10425 27557 10459 27591
rect 11247 27557 11281 27591
rect 12265 27557 12299 27591
rect 13645 27557 13679 27591
rect 14197 27557 14231 27591
rect 15485 27557 15519 27591
rect 17141 27557 17175 27591
rect 17233 27557 17267 27591
rect 18521 27557 18555 27591
rect 18705 27557 18739 27591
rect 18797 27557 18831 27591
rect 19993 27557 20027 27591
rect 22753 27557 22787 27591
rect 22845 27557 22879 27591
rect 25145 27557 25179 27591
rect 27997 27557 28031 27591
rect 31171 27557 31205 27591
rect 39589 27557 39623 27591
rect 39681 27557 39715 27591
rect 44005 27557 44039 27591
rect 45477 27557 45511 27591
rect 45569 27557 45603 27591
rect 10885 27489 10919 27523
rect 11805 27489 11839 27523
rect 8585 27421 8619 27455
rect 10011 27421 10045 27455
rect 21097 27489 21131 27523
rect 21649 27489 21683 27523
rect 24752 27489 24786 27523
rect 27261 27489 27295 27523
rect 28825 27489 28859 27523
rect 29377 27489 29411 27523
rect 29561 27489 29595 27523
rect 31084 27489 31118 27523
rect 32413 27489 32447 27523
rect 32597 27489 32631 27523
rect 34656 27489 34690 27523
rect 36185 27489 36219 27523
rect 36553 27489 36587 27523
rect 37565 27489 37599 27523
rect 41153 27489 41187 27523
rect 13553 27421 13587 27455
rect 15393 27421 15427 27455
rect 15761 27421 15795 27455
rect 17417 27421 17451 27455
rect 18981 27421 19015 27455
rect 20545 27421 20579 27455
rect 21833 27421 21867 27455
rect 27629 27421 27663 27455
rect 28365 27421 28399 27455
rect 36829 27421 36863 27455
rect 37749 27421 37783 27455
rect 39865 27421 39899 27455
rect 43913 27421 43947 27455
rect 44557 27421 44591 27455
rect 45753 27421 45787 27455
rect 12265 27353 12299 27387
rect 23305 27353 23339 27387
rect 9781 27285 9815 27319
rect 10701 27285 10735 27319
rect 12081 27285 12115 27319
rect 13093 27285 13127 27319
rect 15117 27285 15151 27319
rect 18153 27285 18187 27319
rect 24823 27285 24857 27319
rect 27399 27285 27433 27319
rect 27537 27285 27571 27319
rect 30205 27285 30239 27319
rect 34759 27285 34793 27319
rect 40509 27285 40543 27319
rect 42073 27285 42107 27319
rect 43637 27285 43671 27319
rect 11437 27081 11471 27115
rect 12173 27081 12207 27115
rect 13829 27081 13863 27115
rect 16635 27081 16669 27115
rect 17417 27081 17451 27115
rect 19349 27081 19383 27115
rect 20039 27081 20073 27115
rect 20177 27081 20211 27115
rect 22753 27081 22787 27115
rect 23029 27081 23063 27115
rect 24869 27081 24903 27115
rect 27905 27081 27939 27115
rect 28825 27081 28859 27115
rect 29561 27081 29595 27115
rect 31769 27081 31803 27115
rect 34713 27081 34747 27115
rect 35725 27081 35759 27115
rect 37841 27081 37875 27115
rect 39497 27081 39531 27115
rect 39865 27081 39899 27115
rect 41521 27081 41555 27115
rect 41981 27081 42015 27115
rect 45753 27081 45787 27115
rect 11161 27013 11195 27047
rect 17049 27013 17083 27047
rect 23397 27013 23431 27047
rect 25605 27013 25639 27047
rect 30021 27013 30055 27047
rect 10609 26945 10643 26979
rect 12541 26945 12575 26979
rect 12817 26945 12851 26979
rect 15025 26945 15059 26979
rect 15669 26945 15703 26979
rect 19809 26945 19843 26979
rect 20269 26945 20303 26979
rect 21833 26945 21867 26979
rect 24225 26945 24259 26979
rect 26617 26945 26651 26979
rect 26893 26945 26927 26979
rect 32413 26945 32447 26979
rect 38301 26945 38335 26979
rect 41245 26945 41279 26979
rect 42165 26945 42199 26979
rect 42441 26945 42475 26979
rect 44005 26945 44039 26979
rect 45477 26945 45511 26979
rect 10057 26877 10091 26911
rect 10517 26877 10551 26911
rect 16564 26877 16598 26911
rect 18061 26877 18095 26911
rect 18521 26877 18555 26911
rect 19901 26877 19935 26911
rect 24016 26877 24050 26911
rect 24409 26877 24443 26911
rect 28140 26877 28174 26911
rect 30113 26877 30147 26911
rect 30665 26877 30699 26911
rect 31928 26877 31962 26911
rect 33149 26877 33183 26911
rect 33241 26877 33275 26911
rect 33701 26877 33735 26911
rect 36645 26877 36679 26911
rect 37105 26877 37139 26911
rect 40325 26877 40359 26911
rect 40509 26877 40543 26911
rect 40969 26877 41003 26911
rect 9597 26809 9631 26843
rect 12633 26809 12667 26843
rect 14749 26809 14783 26843
rect 15117 26809 15151 26843
rect 22154 26809 22188 26843
rect 25053 26809 25087 26843
rect 25145 26809 25179 26843
rect 26709 26809 26743 26843
rect 28227 26809 28261 26843
rect 30849 26809 30883 26843
rect 33977 26809 34011 26843
rect 36461 26809 36495 26843
rect 37381 26809 37415 26843
rect 38393 26809 38427 26843
rect 38945 26809 38979 26843
rect 42257 26809 42291 26843
rect 43269 26809 43303 26843
rect 44189 26809 44223 26843
rect 44281 26809 44315 26843
rect 44833 26809 44867 26843
rect 9965 26741 9999 26775
rect 13461 26741 13495 26775
rect 15945 26741 15979 26775
rect 17877 26741 17911 26775
rect 18153 26741 18187 26775
rect 20545 26741 20579 26775
rect 21097 26741 21131 26775
rect 21741 26741 21775 26775
rect 25973 26741 26007 26775
rect 26433 26741 26467 26775
rect 27537 26741 27571 26775
rect 31217 26741 31251 26775
rect 31999 26741 32033 26775
rect 32781 26741 32815 26775
rect 34897 26741 34931 26775
rect 36185 26741 36219 26775
rect 43637 26741 43671 26775
rect 13231 26537 13265 26571
rect 15025 26537 15059 26571
rect 15485 26537 15519 26571
rect 17049 26537 17083 26571
rect 18705 26537 18739 26571
rect 20269 26537 20303 26571
rect 21833 26537 21867 26571
rect 23995 26537 24029 26571
rect 24777 26537 24811 26571
rect 26709 26537 26743 26571
rect 28365 26537 28399 26571
rect 30849 26537 30883 26571
rect 34805 26537 34839 26571
rect 36691 26537 36725 26571
rect 37105 26537 37139 26571
rect 37473 26537 37507 26571
rect 41153 26537 41187 26571
rect 43177 26537 43211 26571
rect 43499 26537 43533 26571
rect 44511 26537 44545 26571
rect 11713 26469 11747 26503
rect 14243 26469 14277 26503
rect 16037 26469 16071 26503
rect 19993 26469 20027 26503
rect 22471 26469 22505 26503
rect 24961 26469 24995 26503
rect 25053 26469 25087 26503
rect 25605 26469 25639 26503
rect 27997 26469 28031 26503
rect 29377 26469 29411 26503
rect 32321 26469 32355 26503
rect 35173 26469 35207 26503
rect 38346 26469 38380 26503
rect 41889 26469 41923 26503
rect 44005 26469 44039 26503
rect 10517 26401 10551 26435
rect 12265 26401 12299 26435
rect 13093 26401 13127 26435
rect 14156 26401 14190 26435
rect 17509 26401 17543 26435
rect 17969 26401 18003 26435
rect 19257 26401 19291 26435
rect 23857 26401 23891 26435
rect 27261 26401 27295 26435
rect 30941 26401 30975 26435
rect 33977 26401 34011 26435
rect 36553 26401 36587 26435
rect 38025 26401 38059 26435
rect 39773 26401 39807 26435
rect 40233 26401 40267 26435
rect 43428 26401 43462 26435
rect 44373 26401 44407 26435
rect 10655 26333 10689 26367
rect 11621 26333 11655 26367
rect 15945 26333 15979 26367
rect 16221 26333 16255 26367
rect 18061 26333 18095 26367
rect 19404 26333 19438 26367
rect 19625 26333 19659 26367
rect 22109 26333 22143 26367
rect 27629 26333 27663 26367
rect 29285 26333 29319 26367
rect 29929 26333 29963 26367
rect 31171 26333 31205 26367
rect 32229 26333 32263 26367
rect 32505 26333 32539 26367
rect 35081 26333 35115 26367
rect 40509 26333 40543 26367
rect 41797 26333 41831 26367
rect 42073 26333 42107 26367
rect 19533 26265 19567 26299
rect 35633 26265 35667 26299
rect 10057 26197 10091 26231
rect 18981 26197 19015 26231
rect 21189 26197 21223 26231
rect 23029 26197 23063 26231
rect 27169 26197 27203 26231
rect 27399 26197 27433 26231
rect 27537 26197 27571 26231
rect 33333 26197 33367 26231
rect 34115 26197 34149 26231
rect 38945 26197 38979 26231
rect 39221 26197 39255 26231
rect 9965 25993 9999 26027
rect 11897 25993 11931 26027
rect 14289 25993 14323 26027
rect 19625 25993 19659 26027
rect 19993 25993 20027 26027
rect 24961 25993 24995 26027
rect 28641 25993 28675 26027
rect 29423 25993 29457 26027
rect 30113 25993 30147 26027
rect 36093 25993 36127 26027
rect 37657 25993 37691 26027
rect 38761 25993 38795 26027
rect 39865 25993 39899 26027
rect 40877 25993 40911 26027
rect 43039 25993 43073 26027
rect 43729 25993 43763 26027
rect 14565 25925 14599 25959
rect 15853 25925 15887 25959
rect 17509 25925 17543 25959
rect 23949 25925 23983 25959
rect 36553 25925 36587 25959
rect 42349 25925 42383 25959
rect 43453 25925 43487 25959
rect 45293 25925 45327 25959
rect 13277 25857 13311 25891
rect 15301 25857 15335 25891
rect 16405 25857 16439 25891
rect 17049 25857 17083 25891
rect 18613 25857 18647 25891
rect 22201 25857 22235 25891
rect 25145 25857 25179 25891
rect 25421 25857 25455 25891
rect 26525 25857 26559 25891
rect 26709 25857 26743 25891
rect 26985 25857 27019 25891
rect 30573 25857 30607 25891
rect 30757 25857 30791 25891
rect 32597 25857 32631 25891
rect 33517 25857 33551 25891
rect 34897 25857 34931 25891
rect 36737 25857 36771 25891
rect 37013 25857 37047 25891
rect 38945 25857 38979 25891
rect 41705 25857 41739 25891
rect 44005 25857 44039 25891
rect 44281 25857 44315 25891
rect 10241 25789 10275 25823
rect 10609 25789 10643 25823
rect 20085 25789 20119 25823
rect 20545 25789 20579 25823
rect 21649 25789 21683 25823
rect 22109 25789 22143 25823
rect 28248 25789 28282 25823
rect 29352 25789 29386 25823
rect 29837 25789 29871 25823
rect 33241 25789 33275 25823
rect 42968 25789 43002 25823
rect 10793 25721 10827 25755
rect 12725 25721 12759 25755
rect 13369 25721 13403 25755
rect 13921 25721 13955 25755
rect 14841 25721 14875 25755
rect 14933 25721 14967 25755
rect 16497 25721 16531 25755
rect 18705 25721 18739 25755
rect 19257 25721 19291 25755
rect 24593 25721 24627 25755
rect 25237 25721 25271 25755
rect 26157 25721 26191 25755
rect 26801 25721 26835 25755
rect 31078 25721 31112 25755
rect 32689 25721 32723 25755
rect 35218 25721 35252 25755
rect 36829 25721 36863 25755
rect 39037 25721 39071 25755
rect 39589 25721 39623 25755
rect 40233 25721 40267 25755
rect 41429 25721 41463 25755
rect 41521 25721 41555 25755
rect 44097 25721 44131 25755
rect 11069 25653 11103 25687
rect 11529 25653 11563 25687
rect 13093 25653 13127 25687
rect 18245 25653 18279 25687
rect 20177 25653 20211 25687
rect 21465 25653 21499 25687
rect 22753 25653 22787 25687
rect 27629 25653 27663 25687
rect 27997 25653 28031 25687
rect 28319 25653 28353 25687
rect 29009 25653 29043 25687
rect 31677 25653 31711 25687
rect 31953 25653 31987 25687
rect 32321 25653 32355 25687
rect 33977 25653 34011 25687
rect 34621 25653 34655 25687
rect 35817 25653 35851 25687
rect 38117 25653 38151 25687
rect 41245 25653 41279 25687
rect 44925 25653 44959 25687
rect 11345 25449 11379 25483
rect 14335 25449 14369 25483
rect 14749 25449 14783 25483
rect 16497 25449 16531 25483
rect 17785 25449 17819 25483
rect 18889 25449 18923 25483
rect 19257 25449 19291 25483
rect 20085 25449 20119 25483
rect 22201 25449 22235 25483
rect 24777 25449 24811 25483
rect 25881 25449 25915 25483
rect 26801 25449 26835 25483
rect 28365 25449 28399 25483
rect 31861 25449 31895 25483
rect 34897 25449 34931 25483
rect 37381 25449 37415 25483
rect 40647 25449 40681 25483
rect 41429 25449 41463 25483
rect 10787 25381 10821 25415
rect 12633 25381 12667 25415
rect 13553 25381 13587 25415
rect 15663 25381 15697 25415
rect 18331 25381 18365 25415
rect 19625 25381 19659 25415
rect 23397 25381 23431 25415
rect 25053 25381 25087 25415
rect 29929 25381 29963 25415
rect 32321 25381 32355 25415
rect 35081 25381 35115 25415
rect 35173 25381 35207 25415
rect 37013 25381 37047 25415
rect 38945 25381 38979 25415
rect 41705 25381 41739 25415
rect 44005 25381 44039 25415
rect 14232 25313 14266 25347
rect 17969 25313 18003 25347
rect 27020 25313 27054 25347
rect 34012 25313 34046 25347
rect 36588 25313 36622 25347
rect 37784 25313 37818 25347
rect 40544 25313 40578 25347
rect 10425 25245 10459 25279
rect 12541 25245 12575 25279
rect 13185 25245 13219 25279
rect 15301 25245 15335 25279
rect 23305 25245 23339 25279
rect 24961 25245 24995 25279
rect 25237 25245 25271 25279
rect 27997 25245 28031 25279
rect 29837 25245 29871 25279
rect 32229 25245 32263 25279
rect 35357 25245 35391 25279
rect 38853 25245 38887 25279
rect 39129 25245 39163 25279
rect 41613 25245 41647 25279
rect 41889 25245 41923 25279
rect 43913 25245 43947 25279
rect 45385 25245 45419 25279
rect 23857 25177 23891 25211
rect 27123 25177 27157 25211
rect 29285 25177 29319 25211
rect 30389 25177 30423 25211
rect 32781 25177 32815 25211
rect 37887 25177 37921 25211
rect 44465 25177 44499 25211
rect 10057 25109 10091 25143
rect 12265 25109 12299 25143
rect 15117 25109 15151 25143
rect 16221 25109 16255 25143
rect 16865 25109 16899 25143
rect 20453 25109 20487 25143
rect 21741 25109 21775 25143
rect 24225 25109 24259 25143
rect 27445 25109 27479 25143
rect 28917 25109 28951 25143
rect 31125 25109 31159 25143
rect 34115 25109 34149 25143
rect 34437 25109 34471 25143
rect 36691 25109 36725 25143
rect 38209 25109 38243 25143
rect 10333 24905 10367 24939
rect 11529 24905 11563 24939
rect 13553 24905 13587 24939
rect 15485 24905 15519 24939
rect 17141 24905 17175 24939
rect 23029 24905 23063 24939
rect 24869 24905 24903 24939
rect 25145 24905 25179 24939
rect 26617 24905 26651 24939
rect 27077 24905 27111 24939
rect 34621 24905 34655 24939
rect 35909 24905 35943 24939
rect 36369 24905 36403 24939
rect 37289 24905 37323 24939
rect 38945 24905 38979 24939
rect 40693 24905 40727 24939
rect 41705 24905 41739 24939
rect 43637 24905 43671 24939
rect 43867 24905 43901 24939
rect 44097 24905 44131 24939
rect 44281 24905 44315 24939
rect 44649 24905 44683 24939
rect 12173 24837 12207 24871
rect 12541 24837 12575 24871
rect 33149 24837 33183 24871
rect 39313 24837 39347 24871
rect 42533 24837 42567 24871
rect 9965 24769 9999 24803
rect 10425 24701 10459 24735
rect 10977 24701 11011 24735
rect 11897 24701 11931 24735
rect 16037 24769 16071 24803
rect 17785 24769 17819 24803
rect 20177 24769 20211 24803
rect 22753 24769 22787 24803
rect 23949 24769 23983 24803
rect 29377 24769 29411 24803
rect 30021 24769 30055 24803
rect 34989 24769 35023 24803
rect 35265 24769 35299 24803
rect 37749 24769 37783 24803
rect 42901 24769 42935 24803
rect 12633 24701 12667 24735
rect 14381 24701 14415 24735
rect 14841 24701 14875 24735
rect 17509 24701 17543 24735
rect 18061 24701 18095 24735
rect 18613 24701 18647 24735
rect 21925 24701 21959 24735
rect 22293 24701 22327 24735
rect 22569 24701 22603 24735
rect 25697 24701 25731 24735
rect 27445 24701 27479 24735
rect 27997 24701 28031 24735
rect 33276 24701 33310 24735
rect 36496 24701 36530 24735
rect 40912 24701 40946 24735
rect 41337 24701 41371 24735
rect 43796 24701 43830 24735
rect 44097 24701 44131 24735
rect 11161 24633 11195 24667
rect 12541 24633 12575 24667
rect 12955 24633 12989 24667
rect 13829 24633 13863 24667
rect 15117 24633 15151 24667
rect 16129 24633 16163 24667
rect 16681 24633 16715 24667
rect 20539 24633 20573 24667
rect 23397 24633 23431 24667
rect 24270 24633 24304 24667
rect 25513 24633 25547 24667
rect 26018 24633 26052 24667
rect 28181 24633 28215 24667
rect 29101 24633 29135 24667
rect 29469 24633 29503 24667
rect 31769 24633 31803 24667
rect 31861 24633 31895 24667
rect 32413 24633 32447 24667
rect 33379 24633 33413 24667
rect 35081 24633 35115 24667
rect 37657 24633 37691 24667
rect 38025 24633 38059 24667
rect 41015 24633 41049 24667
rect 41981 24633 42015 24667
rect 42073 24633 42107 24667
rect 14197 24565 14231 24599
rect 15853 24565 15887 24599
rect 18153 24565 18187 24599
rect 19165 24565 19199 24599
rect 20085 24565 20119 24599
rect 21097 24565 21131 24599
rect 28457 24565 28491 24599
rect 30297 24565 30331 24599
rect 31585 24565 31619 24599
rect 32689 24565 32723 24599
rect 33977 24565 34011 24599
rect 36599 24565 36633 24599
rect 38669 24565 38703 24599
rect 10425 24361 10459 24395
rect 10793 24361 10827 24395
rect 12081 24361 12115 24395
rect 13001 24361 13035 24395
rect 14381 24361 14415 24395
rect 15485 24361 15519 24395
rect 15807 24361 15841 24395
rect 20177 24361 20211 24395
rect 21189 24361 21223 24395
rect 23305 24361 23339 24395
rect 24225 24361 24259 24395
rect 24777 24361 24811 24395
rect 25145 24361 25179 24395
rect 27905 24361 27939 24395
rect 28181 24361 28215 24395
rect 28825 24361 28859 24395
rect 30113 24361 30147 24395
rect 31769 24361 31803 24395
rect 32275 24361 32309 24395
rect 32597 24361 32631 24395
rect 35081 24361 35115 24395
rect 36461 24361 36495 24395
rect 38853 24361 38887 24395
rect 41429 24361 41463 24395
rect 42073 24361 42107 24395
rect 42395 24361 42429 24395
rect 11482 24293 11516 24327
rect 16129 24293 16163 24327
rect 18331 24293 18365 24327
rect 22109 24293 22143 24327
rect 30481 24293 30515 24327
rect 35357 24293 35391 24327
rect 35909 24293 35943 24327
rect 38254 24293 38288 24327
rect 40830 24293 40864 24327
rect 41705 24293 41739 24327
rect 43545 24293 43579 24327
rect 12909 24225 12943 24259
rect 13461 24225 13495 24259
rect 15736 24225 15770 24259
rect 16732 24225 16766 24259
rect 17969 24225 18003 24259
rect 19784 24225 19818 24259
rect 21189 24225 21223 24259
rect 21373 24225 21407 24259
rect 22544 24225 22578 24259
rect 26560 24225 26594 24259
rect 28733 24225 28767 24259
rect 29193 24225 29227 24259
rect 32172 24225 32206 24259
rect 33793 24225 33827 24259
rect 34069 24225 34103 24259
rect 40509 24225 40543 24259
rect 42324 24225 42358 24259
rect 11161 24157 11195 24191
rect 16819 24157 16853 24191
rect 23857 24157 23891 24191
rect 27445 24157 27479 24191
rect 30389 24157 30423 24191
rect 31033 24157 31067 24191
rect 34345 24157 34379 24191
rect 34713 24157 34747 24191
rect 35265 24157 35299 24191
rect 37933 24157 37967 24191
rect 43453 24157 43487 24191
rect 44097 24157 44131 24191
rect 19855 24089 19889 24123
rect 22615 24089 22649 24123
rect 12449 24021 12483 24055
rect 18889 24021 18923 24055
rect 19165 24021 19199 24055
rect 23765 24021 23799 24055
rect 25697 24021 25731 24055
rect 26663 24021 26697 24055
rect 29745 24021 29779 24055
rect 11529 23817 11563 23851
rect 12265 23817 12299 23851
rect 13461 23817 13495 23851
rect 17417 23817 17451 23851
rect 17877 23817 17911 23851
rect 18337 23817 18371 23851
rect 18705 23817 18739 23851
rect 19901 23817 19935 23851
rect 20545 23817 20579 23851
rect 22201 23817 22235 23851
rect 22937 23817 22971 23851
rect 24685 23817 24719 23851
rect 26433 23817 26467 23851
rect 27261 23817 27295 23851
rect 28733 23817 28767 23851
rect 29469 23817 29503 23851
rect 30757 23817 30791 23851
rect 33701 23817 33735 23851
rect 36553 23817 36587 23851
rect 36921 23817 36955 23851
rect 38577 23817 38611 23851
rect 40325 23817 40359 23851
rect 41245 23817 41279 23851
rect 43729 23817 43763 23851
rect 11253 23749 11287 23783
rect 14933 23749 14967 23783
rect 19441 23749 19475 23783
rect 30389 23749 30423 23783
rect 32965 23749 32999 23783
rect 35817 23749 35851 23783
rect 40923 23749 40957 23783
rect 43361 23749 43395 23783
rect 13001 23681 13035 23715
rect 18889 23681 18923 23715
rect 21005 23681 21039 23715
rect 22569 23681 22603 23715
rect 24409 23681 24443 23715
rect 26893 23681 26927 23715
rect 29837 23681 29871 23715
rect 31493 23681 31527 23715
rect 32413 23681 32447 23715
rect 35265 23681 35299 23715
rect 37749 23681 37783 23715
rect 38761 23681 38795 23715
rect 41889 23681 41923 23715
rect 12449 23613 12483 23647
rect 12909 23613 12943 23647
rect 14064 23613 14098 23647
rect 14473 23613 14507 23647
rect 16656 23613 16690 23647
rect 17049 23613 17083 23647
rect 23489 23613 23523 23647
rect 23949 23613 23983 23647
rect 24133 23613 24167 23647
rect 27629 23613 27663 23647
rect 27905 23613 27939 23647
rect 37105 23613 37139 23647
rect 37565 23613 37599 23647
rect 40820 23613 40854 23647
rect 41613 23613 41647 23647
rect 14151 23545 14185 23579
rect 15117 23545 15151 23579
rect 15218 23545 15252 23579
rect 15761 23545 15795 23579
rect 16037 23545 16071 23579
rect 18981 23545 19015 23579
rect 21326 23545 21360 23579
rect 28089 23545 28123 23579
rect 29929 23545 29963 23579
rect 31861 23545 31895 23579
rect 32505 23545 32539 23579
rect 33977 23545 34011 23579
rect 34713 23545 34747 23579
rect 35350 23545 35384 23579
rect 36185 23545 36219 23579
rect 38853 23545 38887 23579
rect 39405 23545 39439 23579
rect 41981 23545 42015 23579
rect 42533 23545 42567 23579
rect 16727 23477 16761 23511
rect 20821 23477 20855 23511
rect 21925 23477 21959 23511
rect 32137 23477 32171 23511
rect 38117 23477 38151 23511
rect 42809 23477 42843 23511
rect 13001 23273 13035 23307
rect 14335 23273 14369 23307
rect 15117 23273 15151 23307
rect 18797 23273 18831 23307
rect 23949 23273 23983 23307
rect 27445 23273 27479 23307
rect 29377 23273 29411 23307
rect 30389 23273 30423 23307
rect 33057 23273 33091 23307
rect 37105 23273 37139 23307
rect 38025 23273 38059 23307
rect 38761 23273 38795 23307
rect 39221 23273 39255 23307
rect 41245 23273 41279 23307
rect 41797 23273 41831 23307
rect 42073 23273 42107 23307
rect 42441 23273 42475 23307
rect 15485 23205 15519 23239
rect 17141 23205 17175 23239
rect 19073 23205 19107 23239
rect 21097 23205 21131 23239
rect 23673 23205 23707 23239
rect 28083 23205 28117 23239
rect 29790 23205 29824 23239
rect 32499 23205 32533 23239
rect 34850 23205 34884 23239
rect 11897 23137 11931 23171
rect 12357 23137 12391 23171
rect 14197 23137 14231 23171
rect 22937 23137 22971 23171
rect 23489 23137 23523 23171
rect 24501 23137 24535 23171
rect 25237 23137 25271 23171
rect 26525 23137 26559 23171
rect 30665 23137 30699 23171
rect 36277 23137 36311 23171
rect 37933 23137 37967 23171
rect 38301 23137 38335 23171
rect 39313 23137 39347 23171
rect 39773 23137 39807 23171
rect 12449 23069 12483 23103
rect 15393 23069 15427 23103
rect 17049 23069 17083 23103
rect 17325 23069 17359 23103
rect 18981 23069 19015 23103
rect 19625 23069 19659 23103
rect 21005 23069 21039 23103
rect 24869 23069 24903 23103
rect 27077 23069 27111 23103
rect 27721 23069 27755 23103
rect 29469 23069 29503 23103
rect 32137 23069 32171 23103
rect 34529 23069 34563 23103
rect 40049 23069 40083 23103
rect 40877 23069 40911 23103
rect 15945 23001 15979 23035
rect 21557 23001 21591 23035
rect 26709 22933 26743 22967
rect 28641 22933 28675 22967
rect 35449 22933 35483 22967
rect 35725 22933 35759 22967
rect 36415 22933 36449 22967
rect 13369 22729 13403 22763
rect 14289 22729 14323 22763
rect 16589 22729 16623 22763
rect 16819 22729 16853 22763
rect 17233 22729 17267 22763
rect 20177 22729 20211 22763
rect 21005 22729 21039 22763
rect 21097 22729 21131 22763
rect 22937 22729 22971 22763
rect 23397 22729 23431 22763
rect 24501 22729 24535 22763
rect 28365 22729 28399 22763
rect 29009 22729 29043 22763
rect 36277 22729 36311 22763
rect 38393 22729 38427 22763
rect 39773 22729 39807 22763
rect 41061 22729 41095 22763
rect 41705 22729 41739 22763
rect 15669 22661 15703 22695
rect 22201 22661 22235 22695
rect 39313 22661 39347 22695
rect 42487 22661 42521 22695
rect 12449 22593 12483 22627
rect 15117 22593 15151 22627
rect 18797 22593 18831 22627
rect 19073 22593 19107 22627
rect 21097 22593 21131 22627
rect 21281 22593 21315 22627
rect 21557 22593 21591 22627
rect 27905 22593 27939 22627
rect 29653 22593 29687 22627
rect 29837 22593 29871 22627
rect 30481 22593 30515 22627
rect 32321 22593 32355 22627
rect 32965 22593 32999 22627
rect 35541 22593 35575 22627
rect 41337 22593 41371 22627
rect 16748 22525 16782 22559
rect 23581 22525 23615 22559
rect 24225 22525 24259 22559
rect 25329 22525 25363 22559
rect 26157 22525 26191 22559
rect 26249 22525 26283 22559
rect 27261 22525 27295 22559
rect 27537 22525 27571 22559
rect 27813 22525 27847 22559
rect 11805 22457 11839 22491
rect 12265 22457 12299 22491
rect 12770 22457 12804 22491
rect 15209 22457 15243 22491
rect 17509 22457 17543 22491
rect 18613 22457 18647 22491
rect 18889 22457 18923 22491
rect 21373 22457 21407 22491
rect 24685 22457 24719 22491
rect 26709 22457 26743 22491
rect 31309 22525 31343 22559
rect 31585 22525 31619 22559
rect 32045 22525 32079 22559
rect 33701 22525 33735 22559
rect 33828 22525 33862 22559
rect 36921 22525 36955 22559
rect 37381 22525 37415 22559
rect 38536 22525 38570 22559
rect 38945 22525 38979 22559
rect 40544 22525 40578 22559
rect 42384 22525 42418 22559
rect 42809 22525 42843 22559
rect 43428 22525 43462 22559
rect 43821 22525 43855 22559
rect 29929 22457 29963 22491
rect 11437 22389 11471 22423
rect 14933 22389 14967 22423
rect 16037 22389 16071 22423
rect 19717 22389 19751 22423
rect 20637 22389 20671 22423
rect 23811 22389 23845 22423
rect 25789 22389 25823 22423
rect 26433 22389 26467 22423
rect 29469 22389 29503 22423
rect 29653 22389 29687 22423
rect 33931 22457 33965 22491
rect 35265 22457 35299 22491
rect 35357 22457 35391 22491
rect 37657 22457 37691 22491
rect 31309 22389 31343 22423
rect 31401 22389 31435 22423
rect 32597 22389 32631 22423
rect 34529 22389 34563 22423
rect 36737 22389 36771 22423
rect 37933 22389 37967 22423
rect 38623 22389 38657 22423
rect 40647 22389 40681 22423
rect 43499 22389 43533 22423
rect 12449 22185 12483 22219
rect 14749 22185 14783 22219
rect 19441 22185 19475 22219
rect 19763 22185 19797 22219
rect 23489 22185 23523 22219
rect 23673 22185 23707 22219
rect 29009 22185 29043 22219
rect 29837 22185 29871 22219
rect 30113 22185 30147 22219
rect 31677 22185 31711 22219
rect 34529 22185 34563 22219
rect 34897 22185 34931 22219
rect 38301 22185 38335 22219
rect 13322 22117 13356 22151
rect 15117 22117 15151 22151
rect 15485 22117 15519 22151
rect 16037 22117 16071 22151
rect 17233 22117 17267 22151
rect 17785 22117 17819 22151
rect 18751 22117 18785 22151
rect 21281 22117 21315 22151
rect 11713 22049 11747 22083
rect 11989 22049 12023 22083
rect 13001 22049 13035 22083
rect 18613 22049 18647 22083
rect 19625 22049 19659 22083
rect 23305 22049 23339 22083
rect 12173 21981 12207 22015
rect 15393 21981 15427 22015
rect 17141 21981 17175 22015
rect 21189 21981 21223 22015
rect 21557 21981 21591 22015
rect 28410 22117 28444 22151
rect 33425 22117 33459 22151
rect 35173 22117 35207 22151
rect 35265 22117 35299 22151
rect 40049 22117 40083 22151
rect 43545 22117 43579 22151
rect 24501 22049 24535 22083
rect 24685 22049 24719 22083
rect 26985 22049 27019 22083
rect 31068 22049 31102 22083
rect 32264 22049 32298 22083
rect 36645 22049 36679 22083
rect 37933 22049 37967 22083
rect 41429 22049 41463 22083
rect 41889 22049 41923 22083
rect 27261 21981 27295 22015
rect 28089 21981 28123 22015
rect 31171 21981 31205 22015
rect 33333 21981 33367 22015
rect 33701 21981 33735 22015
rect 35817 21981 35851 22015
rect 39957 21981 39991 22015
rect 40601 21981 40635 22015
rect 42165 21981 42199 22015
rect 42441 21981 42475 22015
rect 43453 21981 43487 22015
rect 43729 21981 43763 22015
rect 27629 21913 27663 21947
rect 13921 21845 13955 21879
rect 19073 21845 19107 21879
rect 23121 21845 23155 21879
rect 23489 21845 23523 21879
rect 24777 21845 24811 21879
rect 32367 21845 32401 21879
rect 33057 21845 33091 21879
rect 36783 21845 36817 21879
rect 37105 21845 37139 21879
rect 38853 21845 38887 21879
rect 11253 21641 11287 21675
rect 11897 21641 11931 21675
rect 12817 21641 12851 21675
rect 14105 21641 14139 21675
rect 16589 21641 16623 21675
rect 16911 21641 16945 21675
rect 17601 21641 17635 21675
rect 18613 21641 18647 21675
rect 20453 21641 20487 21675
rect 21833 21641 21867 21675
rect 22753 21641 22787 21675
rect 24501 21641 24535 21675
rect 24869 21641 24903 21675
rect 27169 21641 27203 21675
rect 27767 21641 27801 21675
rect 28641 21641 28675 21675
rect 28825 21641 28859 21675
rect 30849 21641 30883 21675
rect 31401 21641 31435 21675
rect 31861 21641 31895 21675
rect 33977 21641 34011 21675
rect 35909 21641 35943 21675
rect 38301 21641 38335 21675
rect 40233 21641 40267 21675
rect 40647 21641 40681 21675
rect 41429 21641 41463 21675
rect 44925 21641 44959 21675
rect 17325 21573 17359 21607
rect 24225 21573 24259 21607
rect 27905 21573 27939 21607
rect 11483 21505 11517 21539
rect 15301 21505 15335 21539
rect 16221 21505 16255 21539
rect 27997 21505 28031 21539
rect 28365 21505 28399 21539
rect 11396 21437 11430 21471
rect 12909 21437 12943 21471
rect 16840 21437 16874 21471
rect 18797 21437 18831 21471
rect 19257 21437 19291 21471
rect 20913 21437 20947 21471
rect 22109 21437 22143 21471
rect 23740 21437 23774 21471
rect 25421 21437 25455 21471
rect 26157 21437 26191 21471
rect 27629 21437 27663 21471
rect 13230 21369 13264 21403
rect 14749 21369 14783 21403
rect 15117 21369 15151 21403
rect 15393 21369 15427 21403
rect 15945 21369 15979 21403
rect 19717 21369 19751 21403
rect 21234 21369 21268 21403
rect 26249 21369 26283 21403
rect 32091 21573 32125 21607
rect 41981 21573 42015 21607
rect 32413 21505 32447 21539
rect 33057 21505 33091 21539
rect 33701 21505 33735 21539
rect 34989 21505 35023 21539
rect 35265 21505 35299 21539
rect 36921 21505 36955 21539
rect 37289 21505 37323 21539
rect 39957 21505 39991 21539
rect 42165 21505 42199 21539
rect 44005 21505 44039 21539
rect 44281 21505 44315 21539
rect 29101 21437 29135 21471
rect 29561 21437 29595 21471
rect 29745 21437 29779 21471
rect 31008 21437 31042 21471
rect 31988 21437 32022 21471
rect 32873 21437 32907 21471
rect 40544 21437 40578 21471
rect 40969 21437 41003 21471
rect 30021 21369 30055 21403
rect 33149 21369 33183 21403
rect 35081 21369 35115 21403
rect 37013 21369 37047 21403
rect 38945 21369 38979 21403
rect 39037 21369 39071 21403
rect 39589 21369 39623 21403
rect 42486 21369 42520 21403
rect 44097 21369 44131 21403
rect 12173 21301 12207 21335
rect 13829 21301 13863 21335
rect 18981 21301 19015 21335
rect 20729 21301 20763 21335
rect 23811 21301 23845 21335
rect 26617 21301 26651 21335
rect 27537 21301 27571 21335
rect 28825 21301 28859 21335
rect 31079 21301 31113 21335
rect 34713 21301 34747 21335
rect 36369 21301 36403 21335
rect 36645 21301 36679 21335
rect 37933 21301 37967 21335
rect 38761 21301 38795 21335
rect 43085 21301 43119 21335
rect 43453 21301 43487 21335
rect 43729 21301 43763 21335
rect 13737 21097 13771 21131
rect 17141 21097 17175 21131
rect 19993 21097 20027 21131
rect 21925 21097 21959 21131
rect 26663 21097 26697 21131
rect 27261 21097 27295 21131
rect 28825 21097 28859 21131
rect 32505 21097 32539 21131
rect 33333 21097 33367 21131
rect 34989 21097 35023 21131
rect 35357 21097 35391 21131
rect 38439 21097 38473 21131
rect 38945 21097 38979 21131
rect 42257 21097 42291 21131
rect 44373 21097 44407 21131
rect 13001 21029 13035 21063
rect 15669 21029 15703 21063
rect 17601 21029 17635 21063
rect 19394 21029 19428 21063
rect 21097 21029 21131 21063
rect 24777 21029 24811 21063
rect 28549 21029 28583 21063
rect 29285 21029 29319 21063
rect 34069 21029 34103 21063
rect 34621 21029 34655 21063
rect 36461 21029 36495 21063
rect 39497 21029 39531 21063
rect 41429 21029 41463 21063
rect 43545 21029 43579 21063
rect 10609 20961 10643 20995
rect 12316 20961 12350 20995
rect 13312 20961 13346 20995
rect 19073 20961 19107 20995
rect 23581 20961 23615 20995
rect 26560 20961 26594 20995
rect 27813 20961 27847 20995
rect 27960 20961 27994 20995
rect 29536 20961 29570 20995
rect 30481 20961 30515 20995
rect 30941 20961 30975 20995
rect 33057 20961 33091 20995
rect 35725 20961 35759 20995
rect 36185 20961 36219 20995
rect 38368 20961 38402 20995
rect 12403 20893 12437 20927
rect 15577 20893 15611 20927
rect 17509 20893 17543 20927
rect 18153 20893 18187 20927
rect 21005 20893 21039 20927
rect 24685 20893 24719 20927
rect 25329 20893 25363 20927
rect 28181 20893 28215 20927
rect 31217 20893 31251 20927
rect 32137 20893 32171 20927
rect 33977 20893 34011 20927
rect 39405 20893 39439 20927
rect 40049 20893 40083 20927
rect 41337 20893 41371 20927
rect 41613 20893 41647 20927
rect 43453 20893 43487 20927
rect 43729 20893 43763 20927
rect 13415 20825 13449 20859
rect 16129 20825 16163 20859
rect 21557 20825 21591 20859
rect 10977 20757 11011 20791
rect 18705 20757 18739 20791
rect 23397 20757 23431 20791
rect 23949 20757 23983 20791
rect 27721 20757 27755 20791
rect 28089 20757 28123 20791
rect 29607 20757 29641 20791
rect 33701 20757 33735 20791
rect 36921 20757 36955 20791
rect 37197 20757 37231 20791
rect 10149 20553 10183 20587
rect 12633 20553 12667 20587
rect 14013 20553 14047 20587
rect 14841 20553 14875 20587
rect 16957 20553 16991 20587
rect 17509 20553 17543 20587
rect 17785 20553 17819 20587
rect 19441 20553 19475 20587
rect 21557 20553 21591 20587
rect 21925 20553 21959 20587
rect 22247 20553 22281 20587
rect 23397 20553 23431 20587
rect 24777 20553 24811 20587
rect 25697 20553 25731 20587
rect 27794 20553 27828 20587
rect 28641 20553 28675 20587
rect 29101 20553 29135 20587
rect 31493 20553 31527 20587
rect 32045 20553 32079 20587
rect 32505 20553 32539 20587
rect 33057 20553 33091 20587
rect 34253 20553 34287 20587
rect 34621 20553 34655 20587
rect 35035 20553 35069 20587
rect 35449 20553 35483 20587
rect 37381 20553 37415 20587
rect 38945 20553 38979 20587
rect 39313 20553 39347 20587
rect 39681 20553 39715 20587
rect 42717 20553 42751 20587
rect 42947 20553 42981 20587
rect 44281 20553 44315 20587
rect 16221 20485 16255 20519
rect 19165 20485 19199 20519
rect 23029 20485 23063 20519
rect 27905 20485 27939 20519
rect 31125 20485 31159 20519
rect 16589 20417 16623 20451
rect 18153 20417 18187 20451
rect 21281 20417 21315 20451
rect 24041 20417 24075 20451
rect 27997 20417 28031 20451
rect 29929 20417 29963 20451
rect 33333 20417 33367 20451
rect 33793 20417 33827 20451
rect 36001 20417 36035 20451
rect 36185 20417 36219 20451
rect 38025 20417 38059 20451
rect 41613 20417 41647 20451
rect 9724 20349 9758 20383
rect 9827 20349 9861 20383
rect 10609 20349 10643 20383
rect 10793 20349 10827 20383
rect 12265 20349 12299 20383
rect 13093 20349 13127 20383
rect 14632 20349 14666 20383
rect 15025 20349 15059 20383
rect 20545 20349 20579 20383
rect 21005 20349 21039 20383
rect 22144 20349 22178 20383
rect 22569 20349 22603 20383
rect 25329 20349 25363 20383
rect 26065 20349 26099 20383
rect 26801 20349 26835 20383
rect 27629 20349 27663 20383
rect 32296 20349 32330 20383
rect 34964 20349 34998 20383
rect 42876 20349 42910 20383
rect 43269 20349 43303 20383
rect 43872 20349 43906 20383
rect 10701 20281 10735 20315
rect 13737 20281 13771 20315
rect 15669 20281 15703 20315
rect 15761 20281 15795 20315
rect 18245 20281 18279 20315
rect 18797 20281 18831 20315
rect 23765 20281 23799 20315
rect 23857 20281 23891 20315
rect 28365 20281 28399 20315
rect 30291 20281 30325 20315
rect 33425 20281 33459 20315
rect 36506 20281 36540 20315
rect 37749 20281 37783 20315
rect 38117 20281 38151 20315
rect 38669 20281 38703 20315
rect 41337 20281 41371 20315
rect 41429 20281 41463 20315
rect 43959 20281 43993 20315
rect 15393 20213 15427 20247
rect 19901 20213 19935 20247
rect 20361 20213 20395 20247
rect 27077 20213 27111 20247
rect 27445 20213 27479 20247
rect 29837 20213 29871 20247
rect 30849 20213 30883 20247
rect 32689 20213 32723 20247
rect 37105 20213 37139 20247
rect 40785 20213 40819 20247
rect 41061 20213 41095 20247
rect 42257 20213 42291 20247
rect 43637 20213 43671 20247
rect 10057 20009 10091 20043
rect 10609 20009 10643 20043
rect 16313 20009 16347 20043
rect 17509 20009 17543 20043
rect 20545 20009 20579 20043
rect 26341 20009 26375 20043
rect 28549 20009 28583 20043
rect 30021 20009 30055 20043
rect 32735 20009 32769 20043
rect 40509 20009 40543 20043
rect 11069 19941 11103 19975
rect 13277 19941 13311 19975
rect 15393 19941 15427 19975
rect 15485 19941 15519 19975
rect 16037 19941 16071 19975
rect 18107 19941 18141 19975
rect 19165 19941 19199 19975
rect 20913 19941 20947 19975
rect 23397 19941 23431 19975
rect 25053 19941 25087 19975
rect 26709 19941 26743 19975
rect 30665 19941 30699 19975
rect 33241 19941 33275 19975
rect 33793 19941 33827 19975
rect 36185 19941 36219 19975
rect 36277 19941 36311 19975
rect 38577 19941 38611 19975
rect 43453 19941 43487 19975
rect 43545 19941 43579 19975
rect 9873 19873 9907 19907
rect 16992 19873 17026 19907
rect 17969 19873 18003 19907
rect 19257 19873 19291 19907
rect 28089 19873 28123 19907
rect 29469 19873 29503 19907
rect 32664 19873 32698 19907
rect 41061 19873 41095 19907
rect 41924 19873 41958 19907
rect 44960 19873 44994 19907
rect 10977 19805 11011 19839
rect 13185 19805 13219 19839
rect 13461 19805 13495 19839
rect 18797 19805 18831 19839
rect 19625 19805 19659 19839
rect 21281 19805 21315 19839
rect 23121 19805 23155 19839
rect 23305 19805 23339 19839
rect 23581 19805 23615 19839
rect 24961 19805 24995 19839
rect 25605 19805 25639 19839
rect 26617 19805 26651 19839
rect 26893 19805 26927 19839
rect 29607 19805 29641 19839
rect 30573 19805 30607 19839
rect 33701 19805 33735 19839
rect 33977 19805 34011 19839
rect 36829 19805 36863 19839
rect 38485 19805 38519 19839
rect 39129 19805 39163 19839
rect 40141 19805 40175 19839
rect 43729 19805 43763 19839
rect 11529 19737 11563 19771
rect 19717 19737 19751 19771
rect 21373 19737 21407 19771
rect 31125 19737 31159 19771
rect 35725 19737 35759 19771
rect 42027 19737 42061 19771
rect 14105 19669 14139 19703
rect 17095 19669 17129 19703
rect 19395 19669 19429 19703
rect 19533 19669 19567 19703
rect 21051 19669 21085 19703
rect 21189 19669 21223 19703
rect 24225 19669 24259 19703
rect 24593 19669 24627 19703
rect 27629 19669 27663 19703
rect 28273 19669 28307 19703
rect 38025 19669 38059 19703
rect 41337 19669 41371 19703
rect 41797 19669 41831 19703
rect 45063 19669 45097 19703
rect 9965 19465 9999 19499
rect 10701 19465 10735 19499
rect 12173 19465 12207 19499
rect 12633 19465 12667 19499
rect 15209 19465 15243 19499
rect 15853 19465 15887 19499
rect 17417 19465 17451 19499
rect 18199 19465 18233 19499
rect 19717 19465 19751 19499
rect 20959 19465 20993 19499
rect 22477 19465 22511 19499
rect 23121 19465 23155 19499
rect 24961 19465 24995 19499
rect 26525 19465 26559 19499
rect 28273 19465 28307 19499
rect 28641 19465 28675 19499
rect 29101 19465 29135 19499
rect 31401 19465 31435 19499
rect 32781 19465 32815 19499
rect 34621 19465 34655 19499
rect 35817 19465 35851 19499
rect 36185 19465 36219 19499
rect 40233 19465 40267 19499
rect 40831 19465 40865 19499
rect 42717 19465 42751 19499
rect 43177 19465 43211 19499
rect 44097 19465 44131 19499
rect 44925 19465 44959 19499
rect 14289 19397 14323 19431
rect 19395 19397 19429 19431
rect 20729 19397 20763 19431
rect 31125 19397 31159 19431
rect 33149 19397 33183 19431
rect 34253 19397 34287 19431
rect 35173 19397 35207 19431
rect 35449 19397 35483 19431
rect 37289 19397 37323 19431
rect 38761 19397 38795 19431
rect 42349 19397 42383 19431
rect 10333 19329 10367 19363
rect 10885 19329 10919 19363
rect 11529 19329 11563 19363
rect 15393 19329 15427 19363
rect 19165 19329 19199 19363
rect 19625 19329 19659 19363
rect 21741 19329 21775 19363
rect 23765 19329 23799 19363
rect 25697 19329 25731 19363
rect 33609 19329 33643 19363
rect 41153 19329 41187 19363
rect 41797 19329 41831 19363
rect 12449 19261 12483 19295
rect 16313 19261 16347 19295
rect 16957 19261 16991 19295
rect 18096 19261 18130 19295
rect 19487 19261 19521 19295
rect 20856 19261 20890 19295
rect 22017 19261 22051 19295
rect 27169 19261 27203 19295
rect 27905 19261 27939 19295
rect 29837 19261 29871 19295
rect 32264 19261 32298 19295
rect 34964 19261 34998 19295
rect 35173 19261 35207 19295
rect 38853 19261 38887 19295
rect 39313 19261 39347 19295
rect 39589 19261 39623 19295
rect 40728 19261 40762 19295
rect 43320 19261 43354 19295
rect 10977 19193 11011 19227
rect 13737 19193 13771 19227
rect 13829 19193 13863 19227
rect 17141 19193 17175 19227
rect 19257 19193 19291 19227
rect 20269 19193 20303 19227
rect 21281 19193 21315 19227
rect 23857 19193 23891 19227
rect 24409 19193 24443 19227
rect 25421 19193 25455 19227
rect 25513 19193 25547 19227
rect 30159 19193 30193 19227
rect 32367 19193 32401 19227
rect 33333 19193 33367 19227
rect 33425 19193 33459 19227
rect 36737 19193 36771 19227
rect 36829 19193 36863 19227
rect 38301 19193 38335 19227
rect 41889 19193 41923 19227
rect 43407 19193 43441 19227
rect 13093 19125 13127 19159
rect 13461 19125 13495 19159
rect 17785 19125 17819 19159
rect 18797 19125 18831 19159
rect 22201 19125 22235 19159
rect 23397 19125 23431 19159
rect 27537 19125 27571 19159
rect 29745 19125 29779 19159
rect 30757 19125 30791 19159
rect 35035 19125 35069 19159
rect 36553 19125 36587 19159
rect 37933 19125 37967 19159
rect 41613 19125 41647 19159
rect 43729 19125 43763 19159
rect 10977 18921 11011 18955
rect 11253 18921 11287 18955
rect 13185 18921 13219 18955
rect 19165 18921 19199 18955
rect 20729 18921 20763 18955
rect 21097 18921 21131 18955
rect 22017 18921 22051 18955
rect 23673 18921 23707 18955
rect 25697 18921 25731 18955
rect 32873 18921 32907 18955
rect 39129 18921 39163 18955
rect 40141 18921 40175 18955
rect 40555 18921 40589 18955
rect 12725 18853 12759 18887
rect 13737 18853 13771 18887
rect 14289 18853 14323 18887
rect 18797 18853 18831 18887
rect 19257 18853 19291 18887
rect 23121 18853 23155 18887
rect 29653 18853 29687 18887
rect 29929 18853 29963 18887
rect 30665 18853 30699 18887
rect 31217 18853 31251 18887
rect 33333 18853 33367 18887
rect 33701 18853 33735 18887
rect 34253 18853 34287 18887
rect 35173 18853 35207 18887
rect 35265 18853 35299 18887
rect 35817 18853 35851 18887
rect 38301 18853 38335 18887
rect 41521 18853 41555 18887
rect 41613 18853 41647 18887
rect 10492 18785 10526 18819
rect 12633 18785 12667 18819
rect 15644 18785 15678 18819
rect 17233 18785 17267 18819
rect 18153 18785 18187 18819
rect 21419 18785 21453 18819
rect 21511 18785 21545 18819
rect 22477 18785 22511 18819
rect 24593 18785 24627 18819
rect 25421 18785 25455 18819
rect 27077 18785 27111 18819
rect 29193 18785 29227 18819
rect 29469 18785 29503 18819
rect 32045 18785 32079 18819
rect 36696 18785 36730 18819
rect 40452 18785 40486 18819
rect 43428 18785 43462 18819
rect 13645 18717 13679 18751
rect 16589 18717 16623 18751
rect 19404 18717 19438 18751
rect 19625 18717 19659 18751
rect 19993 18717 20027 18751
rect 24685 18717 24719 18751
rect 27721 18717 27755 18751
rect 30389 18717 30423 18751
rect 30573 18717 30607 18751
rect 32275 18717 32309 18751
rect 33609 18717 33643 18751
rect 36783 18717 36817 18751
rect 38209 18717 38243 18751
rect 41797 18717 41831 18751
rect 17969 18649 18003 18683
rect 38761 18649 38795 18683
rect 10563 18581 10597 18615
rect 15715 18581 15749 18615
rect 18337 18581 18371 18615
rect 19533 18581 19567 18615
rect 25053 18581 25087 18615
rect 26709 18581 26743 18615
rect 37105 18581 37139 18615
rect 43085 18581 43119 18615
rect 43499 18581 43533 18615
rect 10885 18377 10919 18411
rect 12081 18377 12115 18411
rect 17509 18377 17543 18411
rect 18613 18377 18647 18411
rect 18981 18377 19015 18411
rect 19349 18377 19383 18411
rect 21373 18377 21407 18411
rect 23029 18377 23063 18411
rect 23489 18377 23523 18411
rect 24685 18377 24719 18411
rect 27077 18377 27111 18411
rect 29009 18377 29043 18411
rect 29745 18377 29779 18411
rect 33057 18377 33091 18411
rect 34069 18377 34103 18411
rect 35725 18377 35759 18411
rect 36461 18377 36495 18411
rect 37657 18377 37691 18411
rect 39865 18377 39899 18411
rect 41889 18377 41923 18411
rect 44005 18377 44039 18411
rect 12817 18309 12851 18343
rect 17785 18309 17819 18343
rect 25513 18309 25547 18343
rect 40233 18309 40267 18343
rect 41613 18309 41647 18343
rect 13369 18241 13403 18275
rect 16497 18241 16531 18275
rect 20453 18241 20487 18275
rect 23765 18241 23799 18275
rect 24225 18241 24259 18275
rect 25973 18241 26007 18275
rect 27997 18241 28031 18275
rect 36645 18241 36679 18275
rect 38485 18241 38519 18275
rect 40601 18241 40635 18275
rect 43085 18241 43119 18275
rect 43729 18241 43763 18275
rect 9689 18173 9723 18207
rect 10057 18173 10091 18207
rect 10333 18173 10367 18207
rect 11380 18173 11414 18207
rect 14632 18173 14666 18207
rect 15117 18173 15151 18207
rect 17969 18173 18003 18207
rect 19625 18173 19659 18207
rect 19993 18173 20027 18207
rect 20361 18173 20395 18207
rect 29320 18173 29354 18207
rect 30113 18173 30147 18207
rect 30665 18173 30699 18207
rect 33184 18173 33218 18207
rect 33287 18173 33321 18207
rect 34948 18173 34982 18207
rect 35357 18173 35391 18207
rect 10517 18105 10551 18139
rect 13001 18105 13035 18139
rect 13093 18105 13127 18139
rect 14381 18105 14415 18139
rect 16313 18105 16347 18139
rect 16589 18105 16623 18139
rect 17141 18105 17175 18139
rect 22109 18105 22143 18139
rect 22201 18105 22235 18139
rect 22753 18105 22787 18139
rect 23857 18105 23891 18139
rect 25145 18105 25179 18139
rect 25697 18105 25731 18139
rect 25789 18105 25823 18139
rect 27721 18105 27755 18139
rect 27813 18105 27847 18139
rect 30986 18105 31020 18139
rect 32229 18105 32263 18139
rect 35035 18105 35069 18139
rect 36737 18105 36771 18139
rect 37289 18105 37323 18139
rect 38209 18105 38243 18139
rect 38301 18105 38335 18139
rect 40693 18105 40727 18139
rect 41245 18105 41279 18139
rect 42901 18105 42935 18139
rect 43177 18105 43211 18139
rect 9229 18037 9263 18071
rect 11161 18037 11195 18071
rect 11483 18037 11517 18071
rect 13921 18037 13955 18071
rect 14703 18037 14737 18071
rect 15669 18037 15703 18071
rect 18199 18037 18233 18071
rect 21925 18037 21959 18071
rect 27445 18037 27479 18071
rect 29423 18037 29457 18071
rect 30573 18037 30607 18071
rect 31585 18037 31619 18071
rect 33701 18037 33735 18071
rect 34621 18037 34655 18071
rect 37933 18037 37967 18071
rect 39129 18037 39163 18071
rect 9873 17833 9907 17867
rect 10793 17833 10827 17867
rect 13001 17833 13035 17867
rect 16497 17833 16531 17867
rect 18981 17833 19015 17867
rect 19993 17833 20027 17867
rect 21281 17833 21315 17867
rect 27123 17833 27157 17867
rect 31125 17833 31159 17867
rect 36691 17833 36725 17867
rect 37381 17833 37415 17867
rect 38853 17833 38887 17867
rect 45063 17833 45097 17867
rect 11713 17765 11747 17799
rect 13185 17765 13219 17799
rect 13277 17765 13311 17799
rect 15485 17765 15519 17799
rect 17049 17765 17083 17799
rect 23305 17765 23339 17799
rect 23857 17765 23891 17799
rect 24869 17765 24903 17799
rect 28181 17765 28215 17799
rect 28733 17765 28767 17799
rect 30757 17765 30791 17799
rect 31401 17765 31435 17799
rect 33333 17765 33367 17799
rect 33517 17765 33551 17799
rect 33609 17765 33643 17799
rect 35173 17765 35207 17799
rect 37105 17765 37139 17799
rect 39726 17765 39760 17799
rect 41474 17765 41508 17799
rect 43177 17765 43211 17799
rect 43453 17765 43487 17799
rect 43545 17765 43579 17799
rect 10057 17697 10091 17731
rect 10333 17697 10367 17731
rect 18153 17697 18187 17731
rect 19533 17697 19567 17731
rect 27052 17697 27086 17731
rect 30297 17697 30331 17731
rect 30481 17697 30515 17731
rect 36553 17697 36587 17731
rect 37841 17697 37875 17731
rect 38393 17697 38427 17731
rect 40693 17697 40727 17731
rect 42073 17697 42107 17731
rect 44992 17697 45026 17731
rect 11621 17629 11655 17663
rect 13461 17629 13495 17663
rect 15393 17629 15427 17663
rect 16037 17629 16071 17663
rect 16957 17629 16991 17663
rect 18613 17629 18647 17663
rect 20913 17629 20947 17663
rect 23213 17629 23247 17663
rect 24777 17629 24811 17663
rect 25053 17629 25087 17663
rect 28089 17629 28123 17663
rect 32137 17629 32171 17663
rect 33793 17629 33827 17663
rect 35081 17629 35115 17663
rect 38577 17629 38611 17663
rect 39405 17629 39439 17663
rect 41153 17629 41187 17663
rect 43729 17629 43763 17663
rect 12173 17561 12207 17595
rect 12633 17561 12667 17595
rect 17509 17561 17543 17595
rect 21833 17561 21867 17595
rect 35633 17561 35667 17595
rect 18429 17493 18463 17527
rect 20269 17493 20303 17527
rect 22109 17493 22143 17527
rect 25697 17493 25731 17527
rect 27721 17493 27755 17527
rect 40325 17493 40359 17527
rect 9689 17289 9723 17323
rect 13829 17289 13863 17323
rect 15761 17289 15795 17323
rect 17417 17289 17451 17323
rect 19257 17289 19291 17323
rect 21373 17289 21407 17323
rect 23121 17289 23155 17323
rect 24777 17289 24811 17323
rect 25329 17289 25363 17323
rect 29009 17289 29043 17323
rect 29423 17289 29457 17323
rect 30481 17289 30515 17323
rect 34345 17289 34379 17323
rect 39497 17289 39531 17323
rect 39865 17289 39899 17323
rect 40325 17289 40359 17323
rect 41521 17289 41555 17323
rect 42257 17289 42291 17323
rect 43361 17289 43395 17323
rect 43637 17289 43671 17323
rect 45201 17289 45235 17323
rect 13461 17221 13495 17255
rect 18981 17221 19015 17255
rect 22523 17221 22557 17255
rect 32689 17221 32723 17255
rect 36553 17221 36587 17255
rect 37289 17221 37323 17255
rect 37841 17221 37875 17255
rect 38393 17221 38427 17255
rect 41153 17221 41187 17255
rect 10149 17153 10183 17187
rect 12541 17153 12575 17187
rect 13001 17153 13035 17187
rect 20453 17153 20487 17187
rect 22293 17153 22327 17187
rect 24409 17153 24443 17187
rect 25881 17153 25915 17187
rect 27077 17153 27111 17187
rect 31033 17153 31067 17187
rect 31217 17153 31251 17187
rect 31493 17153 31527 17187
rect 33701 17153 33735 17187
rect 36737 17153 36771 17187
rect 39221 17153 39255 17187
rect 41889 17153 41923 17187
rect 44557 17153 44591 17187
rect 14289 17085 14323 17119
rect 14473 17085 14507 17119
rect 16037 17085 16071 17119
rect 18061 17085 18095 17119
rect 22452 17085 22486 17119
rect 27537 17085 27571 17119
rect 27997 17085 28031 17119
rect 29320 17085 29354 17119
rect 34713 17085 34747 17119
rect 35081 17085 35115 17119
rect 35541 17085 35575 17119
rect 38485 17085 38519 17119
rect 38945 17085 38979 17119
rect 42441 17085 42475 17119
rect 10057 17017 10091 17051
rect 10470 17017 10504 17051
rect 12265 17017 12299 17051
rect 12633 17017 12667 17051
rect 15117 17017 15151 17051
rect 15945 17017 15979 17051
rect 20269 17017 20303 17051
rect 20774 17017 20808 17051
rect 21649 17017 21683 17051
rect 23765 17017 23799 17051
rect 23857 17017 23891 17051
rect 25605 17017 25639 17051
rect 25697 17017 25731 17051
rect 30113 17017 30147 17051
rect 31309 17017 31343 17051
rect 33333 17017 33367 17051
rect 33425 17017 33459 17051
rect 35817 17017 35851 17051
rect 36185 17017 36219 17051
rect 36829 17017 36863 17051
rect 40601 17017 40635 17051
rect 40693 17017 40727 17051
rect 42763 17017 42797 17051
rect 44281 17017 44315 17051
rect 44373 17017 44407 17051
rect 9229 16949 9263 16983
rect 11069 16949 11103 16983
rect 11621 16949 11655 16983
rect 15393 16949 15427 16983
rect 17049 16949 17083 16983
rect 17877 16949 17911 16983
rect 18429 16949 18463 16983
rect 23489 16949 23523 16983
rect 27353 16949 27387 16983
rect 27813 16949 27847 16983
rect 28641 16949 28675 16983
rect 33149 16949 33183 16983
rect 44005 16949 44039 16983
rect 10333 16745 10367 16779
rect 10885 16745 10919 16779
rect 14381 16745 14415 16779
rect 15117 16745 15151 16779
rect 18613 16745 18647 16779
rect 18889 16745 18923 16779
rect 20453 16745 20487 16779
rect 23305 16745 23339 16779
rect 23765 16745 23799 16779
rect 24777 16745 24811 16779
rect 28825 16745 28859 16779
rect 31217 16745 31251 16779
rect 32643 16745 32677 16779
rect 33333 16745 33367 16779
rect 35081 16745 35115 16779
rect 35449 16745 35483 16779
rect 36829 16745 36863 16779
rect 37887 16745 37921 16779
rect 38209 16745 38243 16779
rect 38577 16745 38611 16779
rect 40877 16745 40911 16779
rect 42441 16745 42475 16779
rect 12725 16677 12759 16711
rect 15485 16677 15519 16711
rect 16037 16677 16071 16711
rect 17049 16677 17083 16711
rect 22477 16677 22511 16711
rect 23029 16677 23063 16711
rect 25053 16677 25087 16711
rect 28267 16677 28301 16711
rect 33609 16677 33643 16711
rect 33701 16677 33735 16711
rect 36230 16677 36264 16711
rect 41245 16677 41279 16711
rect 43177 16677 43211 16711
rect 43522 16677 43556 16711
rect 9965 16609 9999 16643
rect 14197 16609 14231 16643
rect 18981 16609 19015 16643
rect 19257 16609 19291 16643
rect 21281 16609 21315 16643
rect 23892 16609 23926 16643
rect 26560 16609 26594 16643
rect 27905 16609 27939 16643
rect 29653 16609 29687 16643
rect 30113 16609 30147 16643
rect 32572 16609 32606 16643
rect 37784 16609 37818 16643
rect 39405 16609 39439 16643
rect 39865 16609 39899 16643
rect 12633 16541 12667 16575
rect 13001 16541 13035 16575
rect 15393 16541 15427 16575
rect 16957 16541 16991 16575
rect 17233 16541 17267 16575
rect 22385 16541 22419 16575
rect 24961 16541 24995 16575
rect 25605 16541 25639 16575
rect 30205 16541 30239 16575
rect 33885 16541 33919 16575
rect 35909 16541 35943 16575
rect 40141 16541 40175 16575
rect 40509 16541 40543 16575
rect 41153 16541 41187 16575
rect 41429 16541 41463 16575
rect 43453 16541 43487 16575
rect 43729 16541 43763 16575
rect 21419 16473 21453 16507
rect 23995 16473 24029 16507
rect 26663 16473 26697 16507
rect 11529 16405 11563 16439
rect 18153 16405 18187 16439
rect 19901 16405 19935 16439
rect 21097 16405 21131 16439
rect 22109 16405 22143 16439
rect 24317 16405 24351 16439
rect 27537 16405 27571 16439
rect 29285 16405 29319 16439
rect 37105 16405 37139 16439
rect 39037 16405 39071 16439
rect 9321 16201 9355 16235
rect 9689 16201 9723 16235
rect 12265 16201 12299 16235
rect 12725 16201 12759 16235
rect 13001 16201 13035 16235
rect 14289 16201 14323 16235
rect 14933 16201 14967 16235
rect 15853 16201 15887 16235
rect 17417 16201 17451 16235
rect 19809 16201 19843 16235
rect 24133 16201 24167 16235
rect 25329 16201 25363 16235
rect 29653 16201 29687 16235
rect 33333 16201 33367 16235
rect 33563 16201 33597 16235
rect 35219 16201 35253 16235
rect 37749 16201 37783 16235
rect 40233 16201 40267 16235
rect 41429 16201 41463 16235
rect 41705 16201 41739 16235
rect 43453 16201 43487 16235
rect 9919 16133 9953 16167
rect 11437 16133 11471 16167
rect 15301 16133 15335 16167
rect 35541 16133 35575 16167
rect 36001 16133 36035 16167
rect 39865 16133 39899 16167
rect 42073 16133 42107 16167
rect 13553 16065 13587 16099
rect 15531 16065 15565 16099
rect 17141 16065 17175 16099
rect 20637 16065 20671 16099
rect 22109 16065 22143 16099
rect 22753 16065 22787 16099
rect 26157 16065 26191 16099
rect 30113 16065 30147 16099
rect 31953 16065 31987 16099
rect 32597 16065 32631 16099
rect 37289 16065 37323 16099
rect 38209 16065 38243 16099
rect 40509 16065 40543 16099
rect 43821 16065 43855 16099
rect 9848 15997 9882 16031
rect 15439 15997 15473 16031
rect 17877 15997 17911 16031
rect 18061 15997 18095 16031
rect 18613 15997 18647 16031
rect 19993 15997 20027 16031
rect 20361 15997 20395 16031
rect 27629 15997 27663 16031
rect 28089 15997 28123 16031
rect 33492 15997 33526 16031
rect 33977 15997 34011 16031
rect 34713 15997 34747 16031
rect 35116 15997 35150 16031
rect 36093 15997 36127 16031
rect 42257 15997 42291 16031
rect 42717 15997 42751 16031
rect 10885 15929 10919 15963
rect 10977 15929 11011 15963
rect 13277 15929 13311 15963
rect 13369 15929 13403 15963
rect 16497 15929 16531 15963
rect 16589 15929 16623 15963
rect 21925 15929 21959 15963
rect 22201 15929 22235 15963
rect 24317 15929 24351 15963
rect 24409 15929 24443 15963
rect 24961 15929 24995 15963
rect 25881 15929 25915 15963
rect 25973 15929 26007 15963
rect 28365 15929 28399 15963
rect 30434 15929 30468 15963
rect 32045 15929 32079 15963
rect 36414 15929 36448 15963
rect 38301 15929 38335 15963
rect 38853 15929 38887 15963
rect 40830 15929 40864 15963
rect 44281 15929 44315 15963
rect 10333 15861 10367 15895
rect 10701 15861 10735 15895
rect 16313 15861 16347 15895
rect 18153 15861 18187 15895
rect 19165 15861 19199 15895
rect 21373 15861 21407 15895
rect 23029 15861 23063 15895
rect 23397 15861 23431 15895
rect 25697 15861 25731 15895
rect 26801 15861 26835 15895
rect 27445 15861 27479 15895
rect 28641 15861 28675 15895
rect 29929 15861 29963 15895
rect 31033 15861 31067 15895
rect 31677 15861 31711 15895
rect 32965 15861 32999 15895
rect 34253 15861 34287 15895
rect 37013 15861 37047 15895
rect 39405 15861 39439 15895
rect 42349 15861 42383 15895
rect 13553 15657 13587 15691
rect 17325 15657 17359 15691
rect 18797 15657 18831 15691
rect 21281 15657 21315 15691
rect 21833 15657 21867 15691
rect 22293 15657 22327 15691
rect 25421 15657 25455 15691
rect 27997 15657 28031 15691
rect 28641 15657 28675 15691
rect 29193 15657 29227 15691
rect 29745 15657 29779 15691
rect 30205 15657 30239 15691
rect 31953 15657 31987 15691
rect 33333 15657 33367 15691
rect 36001 15657 36035 15691
rect 38209 15657 38243 15691
rect 40417 15657 40451 15691
rect 43499 15657 43533 15691
rect 11161 15589 11195 15623
rect 11713 15589 11747 15623
rect 12725 15589 12759 15623
rect 15485 15589 15519 15623
rect 18239 15589 18273 15623
rect 24454 15589 24488 15623
rect 26709 15589 26743 15623
rect 32734 15589 32768 15623
rect 33977 15589 34011 15623
rect 34345 15589 34379 15623
rect 36737 15589 36771 15623
rect 38485 15589 38519 15623
rect 9965 15521 9999 15555
rect 16932 15521 16966 15555
rect 19692 15521 19726 15555
rect 22696 15521 22730 15555
rect 25053 15521 25087 15555
rect 30757 15521 30791 15555
rect 30941 15521 30975 15555
rect 36001 15521 36035 15555
rect 36185 15521 36219 15555
rect 40509 15521 40543 15555
rect 40969 15521 41003 15555
rect 42257 15521 42291 15555
rect 43269 15521 43303 15555
rect 10103 15453 10137 15487
rect 11069 15453 11103 15487
rect 12633 15453 12667 15487
rect 15393 15453 15427 15487
rect 17877 15453 17911 15487
rect 20913 15453 20947 15487
rect 24133 15453 24167 15487
rect 26617 15453 26651 15487
rect 27629 15453 27663 15487
rect 28273 15453 28307 15487
rect 31217 15453 31251 15487
rect 32413 15453 32447 15487
rect 34253 15453 34287 15487
rect 34529 15453 34563 15487
rect 38393 15453 38427 15487
rect 38853 15453 38887 15487
rect 41153 15453 41187 15487
rect 13185 15385 13219 15419
rect 15945 15385 15979 15419
rect 16497 15385 16531 15419
rect 19763 15385 19797 15419
rect 27169 15385 27203 15419
rect 10885 15317 10919 15351
rect 17003 15317 17037 15351
rect 19073 15317 19107 15351
rect 22799 15317 22833 15351
rect 25881 15317 25915 15351
rect 37197 15317 37231 15351
rect 41889 15317 41923 15351
rect 9505 15113 9539 15147
rect 10885 15113 10919 15147
rect 11529 15113 11563 15147
rect 12633 15113 12667 15147
rect 14565 15113 14599 15147
rect 15669 15113 15703 15147
rect 16037 15113 16071 15147
rect 17877 15113 17911 15147
rect 18337 15113 18371 15147
rect 19349 15113 19383 15147
rect 19717 15113 19751 15147
rect 21925 15113 21959 15147
rect 24685 15113 24719 15147
rect 25421 15113 25455 15147
rect 27169 15113 27203 15147
rect 27491 15113 27525 15147
rect 28641 15113 28675 15147
rect 29837 15113 29871 15147
rect 30297 15113 30331 15147
rect 31769 15113 31803 15147
rect 32045 15113 32079 15147
rect 32137 15113 32171 15147
rect 33885 15113 33919 15147
rect 34529 15113 34563 15147
rect 34621 15113 34655 15147
rect 36001 15113 36035 15147
rect 36277 15113 36311 15147
rect 38439 15113 38473 15147
rect 39451 15113 39485 15147
rect 40233 15113 40267 15147
rect 41429 15113 41463 15147
rect 43361 15113 43395 15147
rect 26801 15045 26835 15079
rect 15025 14977 15059 15011
rect 18429 14977 18463 15011
rect 22201 14977 22235 15011
rect 24225 14977 24259 15011
rect 28273 14977 28307 15011
rect 9137 14909 9171 14943
rect 9965 14909 9999 14943
rect 13436 14909 13470 14943
rect 16256 14909 16290 14943
rect 16681 14909 16715 14943
rect 20177 14909 20211 14943
rect 21005 14909 21039 14943
rect 23397 14909 23431 14943
rect 23673 14909 23707 14943
rect 24133 14909 24167 14943
rect 25145 14909 25179 14943
rect 25605 14909 25639 14943
rect 26525 14909 26559 14943
rect 27388 14909 27422 14943
rect 27813 14909 27847 14943
rect 29101 14909 29135 14943
rect 29320 14909 29354 14943
rect 30665 14909 30699 14943
rect 31033 14909 31067 14943
rect 31217 14909 31251 14943
rect 31493 14909 31527 14943
rect 39129 15045 39163 15079
rect 39589 15045 39623 15079
rect 39773 15045 39807 15079
rect 40969 15045 41003 15079
rect 42441 15045 42475 15079
rect 42901 15045 42935 15079
rect 36829 14977 36863 15011
rect 38209 14977 38243 15011
rect 40647 14977 40681 15011
rect 41889 14977 41923 15011
rect 32321 14909 32355 14943
rect 33517 14909 33551 14943
rect 34529 14909 34563 14943
rect 34897 14909 34931 14943
rect 35357 14909 35391 14943
rect 38336 14909 38370 14943
rect 38761 14909 38795 14943
rect 39380 14909 39414 14943
rect 39589 14909 39623 14943
rect 40560 14909 40594 14943
rect 13001 14841 13035 14875
rect 14749 14841 14783 14875
rect 14841 14841 14875 14875
rect 18750 14841 18784 14875
rect 20453 14841 20487 14875
rect 20821 14841 20855 14875
rect 21326 14841 21360 14875
rect 25926 14841 25960 14875
rect 32045 14841 32079 14875
rect 32642 14841 32676 14875
rect 35633 14841 35667 14875
rect 36921 14841 36955 14875
rect 37473 14841 37507 14875
rect 41981 14841 42015 14875
rect 9873 14773 9907 14807
rect 10333 14773 10367 14807
rect 11253 14773 11287 14807
rect 13507 14773 13541 14807
rect 13921 14773 13955 14807
rect 16359 14773 16393 14807
rect 17141 14773 17175 14807
rect 17509 14773 17543 14807
rect 22661 14773 22695 14807
rect 29423 14773 29457 14807
rect 33241 14773 33275 14807
rect 34253 14773 34287 14807
rect 10425 14569 10459 14603
rect 18429 14569 18463 14603
rect 21005 14569 21039 14603
rect 23765 14569 23799 14603
rect 24225 14569 24259 14603
rect 25145 14569 25179 14603
rect 30389 14569 30423 14603
rect 32505 14569 32539 14603
rect 33057 14569 33091 14603
rect 34989 14569 35023 14603
rect 42073 14569 42107 14603
rect 11989 14501 12023 14535
rect 13461 14501 13495 14535
rect 13553 14501 13587 14535
rect 15669 14501 15703 14535
rect 15761 14501 15795 14535
rect 22661 14501 22695 14535
rect 23213 14501 23247 14535
rect 26709 14501 26743 14535
rect 27261 14501 27295 14535
rect 28365 14501 28399 14535
rect 28457 14501 28491 14535
rect 34069 14501 34103 14535
rect 36277 14501 36311 14535
rect 37197 14501 37231 14535
rect 38577 14501 38611 14535
rect 41474 14501 41508 14535
rect 17392 14433 17426 14467
rect 18337 14433 18371 14467
rect 18797 14433 18831 14467
rect 20913 14433 20947 14467
rect 21465 14433 21499 14467
rect 24869 14433 24903 14467
rect 25329 14433 25363 14467
rect 30757 14433 30791 14467
rect 30941 14433 30975 14467
rect 36829 14433 36863 14467
rect 41153 14433 41187 14467
rect 10057 14365 10091 14399
rect 11897 14365 11931 14399
rect 12173 14365 12207 14399
rect 13737 14365 13771 14399
rect 15945 14365 15979 14399
rect 22569 14365 22603 14399
rect 26617 14365 26651 14399
rect 29009 14365 29043 14399
rect 31217 14365 31251 14399
rect 32137 14365 32171 14399
rect 33977 14365 34011 14399
rect 36185 14365 36219 14399
rect 38485 14365 38519 14399
rect 39129 14365 39163 14399
rect 14749 14297 14783 14331
rect 34529 14297 34563 14331
rect 9873 14229 9907 14263
rect 10977 14229 11011 14263
rect 13277 14229 13311 14263
rect 16589 14229 16623 14263
rect 17463 14229 17497 14263
rect 18245 14229 18279 14263
rect 29377 14229 29411 14263
rect 11483 14025 11517 14059
rect 12725 14025 12759 14059
rect 14289 14025 14323 14059
rect 15761 14025 15795 14059
rect 16129 14025 16163 14059
rect 20177 14025 20211 14059
rect 24961 14025 24995 14059
rect 25651 14025 25685 14059
rect 27537 14025 27571 14059
rect 27997 14025 28031 14059
rect 30941 14025 30975 14059
rect 31677 14025 31711 14059
rect 32413 14025 32447 14059
rect 33609 14025 33643 14059
rect 34161 14025 34195 14059
rect 34529 14025 34563 14059
rect 35541 14025 35575 14059
rect 37197 14025 37231 14059
rect 41521 14025 41555 14059
rect 11897 13957 11931 13991
rect 15393 13957 15427 13991
rect 21373 13957 21407 13991
rect 25329 13957 25363 13991
rect 26433 13957 26467 13991
rect 30573 13957 30607 13991
rect 40325 13957 40359 13991
rect 9321 13889 9355 13923
rect 12173 13889 12207 13923
rect 13093 13889 13127 13923
rect 13553 13889 13587 13923
rect 14841 13889 14875 13923
rect 16681 13889 16715 13923
rect 20913 13889 20947 13923
rect 24685 13889 24719 13923
rect 26065 13889 26099 13923
rect 27261 13889 27295 13923
rect 29653 13889 29687 13923
rect 32689 13889 32723 13923
rect 35633 13889 35667 13923
rect 38853 13889 38887 13923
rect 41153 13889 41187 13923
rect 10057 13821 10091 13855
rect 10241 13821 10275 13855
rect 11380 13821 11414 13855
rect 18889 13821 18923 13855
rect 19073 13821 19107 13855
rect 20361 13821 20395 13855
rect 20821 13821 20855 13855
rect 22636 13821 22670 13855
rect 25548 13821 25582 13855
rect 28156 13821 28190 13855
rect 29101 13821 29135 13855
rect 31896 13821 31930 13855
rect 33768 13821 33802 13855
rect 40576 13821 40610 13855
rect 10885 13753 10919 13787
rect 13277 13753 13311 13787
rect 13369 13753 13403 13787
rect 14565 13753 14599 13787
rect 14933 13753 14967 13787
rect 16405 13753 16439 13787
rect 16497 13753 16531 13787
rect 23489 13753 23523 13787
rect 24041 13753 24075 13787
rect 24133 13753 24167 13787
rect 26617 13753 26651 13787
rect 26709 13753 26743 13787
rect 28549 13753 28583 13787
rect 29377 13753 29411 13787
rect 29469 13753 29503 13787
rect 37381 13753 37415 13787
rect 38209 13753 38243 13787
rect 38485 13753 38519 13787
rect 38577 13753 38611 13787
rect 9597 13685 9631 13719
rect 9873 13685 9907 13719
rect 11161 13685 11195 13719
rect 17417 13685 17451 13719
rect 17785 13685 17819 13719
rect 18337 13685 18371 13719
rect 18705 13685 18739 13719
rect 21741 13685 21775 13719
rect 22385 13685 22419 13719
rect 22707 13685 22741 13719
rect 23121 13685 23155 13719
rect 28227 13685 28261 13719
rect 31999 13685 32033 13719
rect 33839 13685 33873 13719
rect 36001 13685 36035 13719
rect 36553 13685 36587 13719
rect 36921 13685 36955 13719
rect 37933 13685 37967 13719
rect 39405 13685 39439 13719
rect 40647 13685 40681 13719
rect 9873 13481 9907 13515
rect 14105 13481 14139 13515
rect 14841 13481 14875 13515
rect 15761 13481 15795 13515
rect 18705 13481 18739 13515
rect 19165 13481 19199 13515
rect 21005 13481 21039 13515
rect 24041 13481 24075 13515
rect 26341 13481 26375 13515
rect 27445 13481 27479 13515
rect 28181 13481 28215 13515
rect 28641 13481 28675 13515
rect 30159 13481 30193 13515
rect 35633 13481 35667 13515
rect 38761 13481 38795 13515
rect 11621 13413 11655 13447
rect 12173 13413 12207 13447
rect 13547 13413 13581 13447
rect 15439 13413 15473 13447
rect 16957 13413 16991 13447
rect 22753 13413 22787 13447
rect 22845 13413 22879 13447
rect 24409 13413 24443 13447
rect 26887 13413 26921 13447
rect 35357 13413 35391 13447
rect 36179 13413 36213 13447
rect 37933 13413 37967 13447
rect 39497 13413 39531 13447
rect 10057 13345 10091 13379
rect 10241 13345 10275 13379
rect 15209 13345 15243 13379
rect 18889 13345 18923 13379
rect 19073 13345 19107 13379
rect 20913 13345 20947 13379
rect 21373 13345 21407 13379
rect 29193 13345 29227 13379
rect 30056 13345 30090 13379
rect 32204 13345 32238 13379
rect 33149 13345 33183 13379
rect 34840 13345 34874 13379
rect 11529 13277 11563 13311
rect 13185 13277 13219 13311
rect 16865 13277 16899 13311
rect 17141 13277 17175 13311
rect 23121 13277 23155 13311
rect 24317 13277 24351 13311
rect 24777 13277 24811 13311
rect 26525 13277 26559 13311
rect 28273 13277 28307 13311
rect 35817 13277 35851 13311
rect 37841 13277 37875 13311
rect 39405 13277 39439 13311
rect 34943 13209 34977 13243
rect 38393 13209 38427 13243
rect 39957 13209 39991 13243
rect 10793 13141 10827 13175
rect 16589 13141 16623 13175
rect 17877 13141 17911 13175
rect 20453 13141 20487 13175
rect 22569 13141 22603 13175
rect 25605 13141 25639 13175
rect 27813 13141 27847 13175
rect 29469 13141 29503 13175
rect 31033 13141 31067 13175
rect 32275 13141 32309 13175
rect 33333 13141 33367 13175
rect 36737 13141 36771 13175
rect 9275 12937 9309 12971
rect 11529 12937 11563 12971
rect 13093 12937 13127 12971
rect 16129 12937 16163 12971
rect 16405 12937 16439 12971
rect 19349 12937 19383 12971
rect 23029 12937 23063 12971
rect 23811 12937 23845 12971
rect 24593 12937 24627 12971
rect 26525 12937 26559 12971
rect 30205 12937 30239 12971
rect 30481 12937 30515 12971
rect 32597 12937 32631 12971
rect 36783 12937 36817 12971
rect 37657 12937 37691 12971
rect 38301 12937 38335 12971
rect 39865 12937 39899 12971
rect 40233 12937 40267 12971
rect 8263 12869 8297 12903
rect 12173 12869 12207 12903
rect 18337 12869 18371 12903
rect 22753 12869 22787 12903
rect 24225 12869 24259 12903
rect 25513 12869 25547 12903
rect 26893 12869 26927 12903
rect 32321 12869 32355 12903
rect 33885 12869 33919 12903
rect 37979 12869 38013 12903
rect 9873 12801 9907 12835
rect 13921 12801 13955 12835
rect 17141 12801 17175 12835
rect 20085 12801 20119 12835
rect 20913 12801 20947 12835
rect 28365 12801 28399 12835
rect 29285 12801 29319 12835
rect 35817 12801 35851 12835
rect 36461 12801 36495 12835
rect 39221 12801 39255 12835
rect 8192 12733 8226 12767
rect 9045 12733 9079 12767
rect 9172 12733 9206 12767
rect 10149 12733 10183 12767
rect 10609 12733 10643 12767
rect 11805 12733 11839 12767
rect 12725 12733 12759 12767
rect 13185 12733 13219 12767
rect 13645 12733 13679 12767
rect 14197 12733 14231 12767
rect 14841 12733 14875 12767
rect 14933 12733 14967 12767
rect 15393 12733 15427 12767
rect 16773 12733 16807 12767
rect 17877 12733 17911 12767
rect 18429 12733 18463 12767
rect 23489 12733 23523 12767
rect 23708 12733 23742 12767
rect 25145 12733 25179 12767
rect 25605 12733 25639 12767
rect 27629 12733 27663 12767
rect 28181 12733 28215 12767
rect 31033 12733 31067 12767
rect 32873 12733 32907 12767
rect 35357 12733 35391 12767
rect 35541 12733 35575 12767
rect 36680 12733 36714 12767
rect 37908 12733 37942 12767
rect 16589 12665 16623 12699
rect 18750 12665 18784 12699
rect 20729 12665 20763 12699
rect 21234 12665 21268 12699
rect 25926 12665 25960 12699
rect 28641 12665 28675 12699
rect 29101 12665 29135 12699
rect 29647 12665 29681 12699
rect 30941 12665 30975 12699
rect 31395 12665 31429 12699
rect 32781 12665 32815 12699
rect 37105 12665 37139 12699
rect 38945 12665 38979 12699
rect 39037 12665 39071 12699
rect 8677 12597 8711 12631
rect 10241 12597 10275 12631
rect 15025 12597 15059 12631
rect 17509 12597 17543 12631
rect 19625 12597 19659 12631
rect 20453 12597 20487 12631
rect 21833 12597 21867 12631
rect 27445 12597 27479 12631
rect 31953 12597 31987 12631
rect 34713 12597 34747 12631
rect 36185 12597 36219 12631
rect 38761 12597 38795 12631
rect 11161 12393 11195 12427
rect 13829 12393 13863 12427
rect 14933 12393 14967 12427
rect 18705 12393 18739 12427
rect 19947 12393 19981 12427
rect 22201 12393 22235 12427
rect 23397 12393 23431 12427
rect 23949 12393 23983 12427
rect 25145 12393 25179 12427
rect 31217 12393 31251 12427
rect 35173 12393 35207 12427
rect 37933 12393 37967 12427
rect 38945 12393 38979 12427
rect 39405 12393 39439 12427
rect 39957 12393 39991 12427
rect 41705 12393 41739 12427
rect 9965 12325 9999 12359
rect 10517 12325 10551 12359
rect 12903 12325 12937 12359
rect 16399 12325 16433 12359
rect 18147 12325 18181 12359
rect 21602 12325 21636 12359
rect 27905 12325 27939 12359
rect 28273 12325 28307 12359
rect 29469 12325 29503 12359
rect 30659 12325 30693 12359
rect 33057 12325 33091 12359
rect 34069 12325 34103 12359
rect 41147 12325 41181 12359
rect 10241 12257 10275 12291
rect 13461 12257 13495 12291
rect 15485 12257 15519 12291
rect 19876 12257 19910 12291
rect 24869 12257 24903 12291
rect 25329 12257 25363 12291
rect 27169 12257 27203 12291
rect 27721 12257 27755 12291
rect 28733 12257 28767 12291
rect 29285 12257 29319 12291
rect 32413 12257 32447 12291
rect 35484 12257 35518 12291
rect 36461 12257 36495 12291
rect 12541 12189 12575 12223
rect 16037 12189 16071 12223
rect 17785 12189 17819 12223
rect 20729 12189 20763 12223
rect 21281 12189 21315 12223
rect 23029 12189 23063 12223
rect 30297 12189 30331 12223
rect 33977 12189 34011 12223
rect 34253 12189 34287 12223
rect 38485 12189 38519 12223
rect 39037 12189 39071 12223
rect 40785 12189 40819 12223
rect 18981 12121 19015 12155
rect 16957 12053 16991 12087
rect 21097 12053 21131 12087
rect 24225 12053 24259 12087
rect 26709 12053 26743 12087
rect 29929 12053 29963 12087
rect 35587 12053 35621 12087
rect 36645 12053 36679 12087
rect 36921 12053 36955 12087
rect 9505 11849 9539 11883
rect 15853 11849 15887 11883
rect 16497 11849 16531 11883
rect 17141 11849 17175 11883
rect 17877 11849 17911 11883
rect 19901 11849 19935 11883
rect 21465 11849 21499 11883
rect 24593 11849 24627 11883
rect 30941 11849 30975 11883
rect 31493 11849 31527 11883
rect 32137 11849 32171 11883
rect 34253 11849 34287 11883
rect 36185 11849 36219 11883
rect 38301 11849 38335 11883
rect 39589 11849 39623 11883
rect 40877 11849 40911 11883
rect 11253 11781 11287 11815
rect 12265 11781 12299 11815
rect 14841 11781 14875 11815
rect 16221 11781 16255 11815
rect 16819 11781 16853 11815
rect 23029 11781 23063 11815
rect 23305 11781 23339 11815
rect 23397 11781 23431 11815
rect 31723 11781 31757 11815
rect 33885 11781 33919 11815
rect 13185 11713 13219 11747
rect 13829 11713 13863 11747
rect 14933 11713 14967 11747
rect 21005 11713 21039 11747
rect 21925 11713 21959 11747
rect 10333 11645 10367 11679
rect 11897 11645 11931 11679
rect 12725 11645 12759 11679
rect 12909 11645 12943 11679
rect 13461 11645 13495 11679
rect 16748 11645 16782 11679
rect 18521 11645 18555 11679
rect 18889 11645 18923 11679
rect 19073 11645 19107 11679
rect 20361 11645 20395 11679
rect 20729 11645 20763 11679
rect 20913 11645 20947 11679
rect 22293 11645 22327 11679
rect 22477 11645 22511 11679
rect 23673 11713 23707 11747
rect 26525 11713 26559 11747
rect 27445 11713 27479 11747
rect 32689 11713 32723 11747
rect 33333 11713 33367 11747
rect 36737 11713 36771 11747
rect 39221 11713 39255 11747
rect 39865 11713 39899 11747
rect 24869 11645 24903 11679
rect 25605 11645 25639 11679
rect 25789 11645 25823 11679
rect 26249 11645 26283 11679
rect 30113 11645 30147 11679
rect 30297 11645 30331 11679
rect 31652 11645 31686 11679
rect 34713 11645 34747 11679
rect 35541 11645 35575 11679
rect 38485 11645 38519 11679
rect 38945 11645 38979 11679
rect 9873 11577 9907 11611
rect 10241 11577 10275 11611
rect 10695 11577 10729 11611
rect 15254 11577 15288 11611
rect 22753 11577 22787 11611
rect 23305 11577 23339 11611
rect 24035 11577 24069 11611
rect 26801 11577 26835 11611
rect 27261 11577 27295 11611
rect 27537 11577 27571 11611
rect 28089 11577 28123 11611
rect 29745 11577 29779 11611
rect 30573 11577 30607 11611
rect 32505 11577 32539 11611
rect 32781 11577 32815 11611
rect 34897 11577 34931 11611
rect 36553 11577 36587 11611
rect 37099 11577 37133 11611
rect 18705 11509 18739 11543
rect 25237 11509 25271 11543
rect 28365 11509 28399 11543
rect 28733 11509 28767 11543
rect 37657 11509 37691 11543
rect 41153 11509 41187 11543
rect 9965 11305 9999 11339
rect 10333 11305 10367 11339
rect 11069 11305 11103 11339
rect 13185 11305 13219 11339
rect 15025 11305 15059 11339
rect 16037 11305 16071 11339
rect 17785 11305 17819 11339
rect 17969 11305 18003 11339
rect 19717 11305 19751 11339
rect 23857 11305 23891 11339
rect 24685 11305 24719 11339
rect 26617 11305 26651 11339
rect 27629 11305 27663 11339
rect 30573 11305 30607 11339
rect 32689 11305 32723 11339
rect 35633 11305 35667 11339
rect 12357 11237 12391 11271
rect 19441 11237 19475 11271
rect 20913 11237 20947 11271
rect 23581 11237 23615 11271
rect 24225 11237 24259 11271
rect 36829 11237 36863 11271
rect 37933 11237 37967 11271
rect 40049 11237 40083 11271
rect 10241 11169 10275 11203
rect 10517 11169 10551 11203
rect 12541 11169 12575 11203
rect 12909 11169 12943 11203
rect 13737 11169 13771 11203
rect 13921 11169 13955 11203
rect 16221 11169 16255 11203
rect 16405 11169 16439 11203
rect 18153 11169 18187 11203
rect 18337 11169 18371 11203
rect 18889 11169 18923 11203
rect 19625 11169 19659 11203
rect 21097 11169 21131 11203
rect 21465 11169 21499 11203
rect 23029 11169 23063 11203
rect 23305 11169 23339 11203
rect 24409 11169 24443 11203
rect 24869 11169 24903 11203
rect 26525 11169 26559 11203
rect 26985 11169 27019 11203
rect 28156 11169 28190 11203
rect 29561 11169 29595 11203
rect 30021 11169 30055 11203
rect 32172 11169 32206 11203
rect 35173 11169 35207 11203
rect 36277 11169 36311 11203
rect 36553 11169 36587 11203
rect 39589 11169 39623 11203
rect 39773 11169 39807 11203
rect 14289 11101 14323 11135
rect 25789 11101 25823 11135
rect 30297 11101 30331 11135
rect 30941 11101 30975 11135
rect 37841 11101 37875 11135
rect 38301 11101 38335 11135
rect 22017 11033 22051 11067
rect 28227 11033 28261 11067
rect 20545 10965 20579 10999
rect 22661 10965 22695 10999
rect 27997 10965 28031 10999
rect 29285 10965 29319 10999
rect 32275 10965 32309 10999
rect 34805 10965 34839 10999
rect 10793 10761 10827 10795
rect 11897 10761 11931 10795
rect 12725 10761 12759 10795
rect 14565 10761 14599 10795
rect 14933 10761 14967 10795
rect 18613 10761 18647 10795
rect 19073 10761 19107 10795
rect 21833 10761 21867 10795
rect 23029 10761 23063 10795
rect 24317 10761 24351 10795
rect 27537 10761 27571 10795
rect 28181 10761 28215 10795
rect 29423 10761 29457 10795
rect 29745 10761 29779 10795
rect 30481 10761 30515 10795
rect 34345 10761 34379 10795
rect 36185 10761 36219 10795
rect 36553 10761 36587 10795
rect 37289 10761 37323 10795
rect 38301 10761 38335 10795
rect 39405 10761 39439 10795
rect 9689 10625 9723 10659
rect 9321 10557 9355 10591
rect 10057 10557 10091 10591
rect 10701 10557 10735 10591
rect 12449 10557 12483 10591
rect 12633 10557 12667 10591
rect 13369 10557 13403 10591
rect 14473 10557 14507 10591
rect 17141 10693 17175 10727
rect 17417 10693 17451 10727
rect 17785 10693 17819 10727
rect 29009 10693 29043 10727
rect 34713 10693 34747 10727
rect 37933 10693 37967 10727
rect 39681 10693 39715 10727
rect 15577 10625 15611 10659
rect 16129 10625 16163 10659
rect 16773 10625 16807 10659
rect 22293 10625 22327 10659
rect 26617 10625 26651 10659
rect 30573 10625 30607 10659
rect 32505 10625 32539 10659
rect 16037 10557 16071 10591
rect 16313 10557 16347 10591
rect 18797 10557 18831 10591
rect 18981 10557 19015 10591
rect 20821 10557 20855 10591
rect 21373 10557 21407 10591
rect 22636 10557 22670 10591
rect 23581 10557 23615 10591
rect 24869 10557 24903 10591
rect 25789 10557 25823 10591
rect 29320 10557 29354 10591
rect 37540 10557 37574 10591
rect 9045 10489 9079 10523
rect 9137 10489 9171 10523
rect 10425 10489 10459 10523
rect 10517 10489 10551 10523
rect 11437 10489 11471 10523
rect 12265 10489 12299 10523
rect 14105 10489 14139 10523
rect 14289 10489 14323 10523
rect 14933 10489 14967 10523
rect 15945 10489 15979 10523
rect 19993 10489 20027 10523
rect 20637 10489 20671 10523
rect 21557 10489 21591 10523
rect 23811 10489 23845 10523
rect 24777 10489 24811 10523
rect 25231 10489 25265 10523
rect 26525 10489 26559 10523
rect 26979 10489 27013 10523
rect 32321 10489 32355 10523
rect 32597 10489 32631 10523
rect 33149 10489 33183 10523
rect 34989 10489 35023 10523
rect 35081 10489 35115 10523
rect 35633 10489 35667 10523
rect 13829 10421 13863 10455
rect 15209 10421 15243 10455
rect 18337 10421 18371 10455
rect 19625 10421 19659 10455
rect 22707 10421 22741 10455
rect 23397 10421 23431 10455
rect 26065 10421 26099 10455
rect 30941 10421 30975 10455
rect 31493 10421 31527 10455
rect 31861 10421 31895 10455
rect 33517 10421 33551 10455
rect 37611 10421 37645 10455
rect 10149 10217 10183 10251
rect 10793 10217 10827 10251
rect 12173 10217 12207 10251
rect 13737 10217 13771 10251
rect 14289 10217 14323 10251
rect 19349 10217 19383 10251
rect 21235 10217 21269 10251
rect 22477 10217 22511 10251
rect 23029 10217 23063 10251
rect 23673 10217 23707 10251
rect 26341 10217 26375 10251
rect 31217 10217 31251 10251
rect 35541 10217 35575 10251
rect 10517 10149 10551 10183
rect 18061 10149 18095 10183
rect 18613 10149 18647 10183
rect 25053 10149 25087 10183
rect 25329 10149 25363 10183
rect 27261 10149 27295 10183
rect 27353 10149 27387 10183
rect 27905 10149 27939 10183
rect 30659 10149 30693 10183
rect 32505 10149 32539 10183
rect 32597 10149 32631 10183
rect 33149 10149 33183 10183
rect 34069 10149 34103 10183
rect 34345 10149 34379 10183
rect 35173 10149 35207 10183
rect 36277 10149 36311 10183
rect 37749 10149 37783 10183
rect 10701 10081 10735 10115
rect 11897 10081 11931 10115
rect 12082 10081 12116 10115
rect 13277 10081 13311 10115
rect 13507 10081 13541 10115
rect 16865 10081 16899 10115
rect 18245 10081 18279 10115
rect 19441 10081 19475 10115
rect 19625 10081 19659 10115
rect 21164 10081 21198 10115
rect 24317 10081 24351 10115
rect 24777 10081 24811 10115
rect 28825 10081 28859 10115
rect 29193 10081 29227 10115
rect 37841 10081 37875 10115
rect 15761 10013 15795 10047
rect 16221 10013 16255 10047
rect 20269 10013 20303 10047
rect 22109 10013 22143 10047
rect 29469 10013 29503 10047
rect 30297 10013 30331 10047
rect 34253 10013 34287 10047
rect 34897 10013 34931 10047
rect 36185 10013 36219 10047
rect 36829 10013 36863 10047
rect 13185 9945 13219 9979
rect 13369 9945 13403 9979
rect 21557 9945 21591 9979
rect 24133 9945 24167 9979
rect 11345 9877 11379 9911
rect 12725 9877 12759 9911
rect 16037 9877 16071 9911
rect 19717 9877 19751 9911
rect 21925 9877 21959 9911
rect 26709 9877 26743 9911
rect 8493 9673 8527 9707
rect 10517 9673 10551 9707
rect 14841 9673 14875 9707
rect 17049 9673 17083 9707
rect 17509 9673 17543 9707
rect 18337 9673 18371 9707
rect 20913 9673 20947 9707
rect 21281 9673 21315 9707
rect 22569 9673 22603 9707
rect 25145 9673 25179 9707
rect 27261 9673 27295 9707
rect 28733 9673 28767 9707
rect 29561 9673 29595 9707
rect 30941 9673 30975 9707
rect 31217 9673 31251 9707
rect 33931 9673 33965 9707
rect 34345 9673 34379 9707
rect 34621 9673 34655 9707
rect 36461 9673 36495 9707
rect 38301 9673 38335 9707
rect 13645 9605 13679 9639
rect 15807 9605 15841 9639
rect 15945 9605 15979 9639
rect 16129 9605 16163 9639
rect 33609 9605 33643 9639
rect 39037 9605 39071 9639
rect 8769 9537 8803 9571
rect 13737 9537 13771 9571
rect 16037 9537 16071 9571
rect 20545 9537 20579 9571
rect 21373 9537 21407 9571
rect 24225 9537 24259 9571
rect 28365 9537 28399 9571
rect 34989 9537 35023 9571
rect 36185 9537 36219 9571
rect 8284 9469 8318 9503
rect 9413 9469 9447 9503
rect 10057 9469 10091 9503
rect 13516 9469 13550 9503
rect 14105 9469 14139 9503
rect 18061 9469 18095 9503
rect 18245 9469 18279 9503
rect 19809 9469 19843 9503
rect 20361 9469 20395 9503
rect 25973 9469 26007 9503
rect 26157 9469 26191 9503
rect 26617 9469 26651 9503
rect 27756 9469 27790 9503
rect 29653 9469 29687 9503
rect 33828 9469 33862 9503
rect 37197 9469 37231 9503
rect 37933 9469 37967 9503
rect 38853 9469 38887 9503
rect 39313 9469 39347 9503
rect 9137 9401 9171 9435
rect 9229 9401 9263 9435
rect 9781 9401 9815 9435
rect 10701 9401 10735 9435
rect 10793 9401 10827 9435
rect 11345 9401 11379 9435
rect 13369 9401 13403 9435
rect 15669 9401 15703 9435
rect 19533 9401 19567 9435
rect 22937 9401 22971 9435
rect 24317 9401 24351 9435
rect 24869 9401 24903 9435
rect 26893 9401 26927 9435
rect 30015 9401 30049 9435
rect 31769 9401 31803 9435
rect 32321 9401 32355 9435
rect 32413 9401 32447 9435
rect 32965 9401 32999 9435
rect 35081 9401 35115 9435
rect 35633 9401 35667 9435
rect 11897 9333 11931 9367
rect 12909 9333 12943 9367
rect 13277 9333 13311 9367
rect 14381 9333 14415 9367
rect 15117 9333 15151 9367
rect 15485 9333 15519 9367
rect 16681 9333 16715 9367
rect 17785 9333 17819 9367
rect 18889 9333 18923 9367
rect 21741 9333 21775 9367
rect 22293 9333 22327 9367
rect 23489 9333 23523 9367
rect 24041 9333 24075 9367
rect 27629 9333 27663 9367
rect 27859 9333 27893 9367
rect 30573 9333 30607 9367
rect 32045 9333 32079 9367
rect 33241 9333 33275 9367
rect 37749 9333 37783 9367
rect 8723 9129 8757 9163
rect 9965 9129 9999 9163
rect 10977 9129 11011 9163
rect 11253 9129 11287 9163
rect 18889 9129 18923 9163
rect 20269 9129 20303 9163
rect 21465 9129 21499 9163
rect 21833 9129 21867 9163
rect 22845 9129 22879 9163
rect 27169 9129 27203 9163
rect 27997 9129 28031 9163
rect 33793 9129 33827 9163
rect 10378 9061 10412 9095
rect 14013 9061 14047 9095
rect 18061 9061 18095 9095
rect 19993 9061 20027 9095
rect 22287 9061 22321 9095
rect 24317 9061 24351 9095
rect 29377 9061 29411 9095
rect 29653 9061 29687 9095
rect 32321 9061 32355 9095
rect 32873 9061 32907 9095
rect 34161 9061 34195 9095
rect 35725 9061 35759 9095
rect 37933 9061 37967 9095
rect 8652 8993 8686 9027
rect 11897 8993 11931 9027
rect 12081 8993 12115 9027
rect 13277 8993 13311 9027
rect 13553 8993 13587 9027
rect 15669 8993 15703 9027
rect 15899 8993 15933 9027
rect 18245 8993 18279 9027
rect 19441 8993 19475 9027
rect 19625 8993 19659 9027
rect 20980 8993 21014 9027
rect 26801 8993 26835 9027
rect 28641 8993 28675 9027
rect 29101 8993 29135 9027
rect 30205 8993 30239 9027
rect 30665 8993 30699 9027
rect 34713 8993 34747 9027
rect 10057 8925 10091 8959
rect 13369 8925 13403 8959
rect 16129 8925 16163 8959
rect 21925 8925 21959 8959
rect 24225 8925 24259 8959
rect 24869 8925 24903 8959
rect 30941 8925 30975 8959
rect 32229 8925 32263 8959
rect 34069 8925 34103 8959
rect 35633 8925 35667 8959
rect 35909 8925 35943 8959
rect 37841 8925 37875 8959
rect 38117 8925 38151 8959
rect 12725 8857 12759 8891
rect 15761 8857 15795 8891
rect 21051 8857 21085 8891
rect 12173 8789 12207 8823
rect 13185 8789 13219 8823
rect 15485 8789 15519 8823
rect 18337 8789 18371 8823
rect 26157 8789 26191 8823
rect 27721 8789 27755 8823
rect 34989 8789 35023 8823
rect 36553 8789 36587 8823
rect 8677 8585 8711 8619
rect 11621 8585 11655 8619
rect 14289 8585 14323 8619
rect 17877 8585 17911 8619
rect 19993 8585 20027 8619
rect 20729 8585 20763 8619
rect 22293 8585 22327 8619
rect 22569 8585 22603 8619
rect 25145 8585 25179 8619
rect 25605 8585 25639 8619
rect 27445 8585 27479 8619
rect 28641 8585 28675 8619
rect 29929 8585 29963 8619
rect 30297 8585 30331 8619
rect 31769 8585 31803 8619
rect 32689 8585 32723 8619
rect 34253 8585 34287 8619
rect 34713 8585 34747 8619
rect 35909 8585 35943 8619
rect 36277 8585 36311 8619
rect 38853 8585 38887 8619
rect 16037 8517 16071 8551
rect 16957 8517 16991 8551
rect 17325 8517 17359 8551
rect 23489 8517 23523 8551
rect 26893 8517 26927 8551
rect 33885 8517 33919 8551
rect 9597 8449 9631 8483
rect 12817 8449 12851 8483
rect 13277 8449 13311 8483
rect 15025 8449 15059 8483
rect 15393 8449 15427 8483
rect 16681 8449 16715 8483
rect 21925 8449 21959 8483
rect 24225 8449 24259 8483
rect 28365 8449 28399 8483
rect 32367 8449 32401 8483
rect 33333 8449 33367 8483
rect 34989 8449 35023 8483
rect 35265 8449 35299 8483
rect 36553 8449 36587 8483
rect 37197 8449 37231 8483
rect 10333 8381 10367 8415
rect 10517 8381 10551 8415
rect 13921 8381 13955 8415
rect 15945 8381 15979 8415
rect 16221 8381 16255 8415
rect 18797 8381 18831 8415
rect 18981 8381 19015 8415
rect 21005 8381 21039 8415
rect 21189 8381 21223 8415
rect 21649 8381 21683 8415
rect 30481 8381 30515 8415
rect 31401 8381 31435 8415
rect 32045 8381 32079 8415
rect 32264 8381 32298 8415
rect 38025 8381 38059 8415
rect 38485 8381 38519 8415
rect 9229 8313 9263 8347
rect 11989 8313 12023 8347
rect 18337 8313 18371 8347
rect 18705 8313 18739 8347
rect 19717 8313 19751 8347
rect 24041 8313 24075 8347
rect 24317 8313 24351 8347
rect 24869 8313 24903 8347
rect 25789 8313 25823 8347
rect 25881 8313 25915 8347
rect 26433 8313 26467 8347
rect 27721 8313 27755 8347
rect 27813 8313 27847 8347
rect 30802 8313 30836 8347
rect 33149 8313 33183 8347
rect 33425 8313 33459 8347
rect 35081 8313 35115 8347
rect 36645 8313 36679 8347
rect 9873 8245 9907 8279
rect 10149 8245 10183 8279
rect 13185 8245 13219 8279
rect 15853 8245 15887 8279
rect 19073 8245 19107 8279
rect 29009 8245 29043 8279
rect 29561 8245 29595 8279
rect 37749 8245 37783 8279
rect 38209 8245 38243 8279
rect 13369 8041 13403 8075
rect 17509 8041 17543 8075
rect 18797 8041 18831 8075
rect 24041 8041 24075 8075
rect 26341 8041 26375 8075
rect 27721 8041 27755 8075
rect 28227 8041 28261 8075
rect 29561 8041 29595 8075
rect 31079 8041 31113 8075
rect 32229 8041 32263 8075
rect 34069 8041 34103 8075
rect 35541 8041 35575 8075
rect 36001 8041 36035 8075
rect 10609 7973 10643 8007
rect 12173 7973 12207 8007
rect 13645 7973 13679 8007
rect 16589 7973 16623 8007
rect 19441 7973 19475 8007
rect 19993 7973 20027 8007
rect 24409 7973 24443 8007
rect 24961 7973 24995 8007
rect 26709 7973 26743 8007
rect 33241 7973 33275 8007
rect 34345 7973 34379 8007
rect 34897 7973 34931 8007
rect 36277 7973 36311 8007
rect 36829 7973 36863 8007
rect 37933 7973 37967 8007
rect 13737 7905 13771 7939
rect 15853 7905 15887 7939
rect 17417 7905 17451 7939
rect 17969 7905 18003 7939
rect 19625 7905 19659 7939
rect 21097 7905 21131 7939
rect 21373 7905 21407 7939
rect 22937 7905 22971 7939
rect 23121 7905 23155 7939
rect 28124 7905 28158 7939
rect 29285 7905 29319 7939
rect 29745 7905 29779 7939
rect 30976 7905 31010 7939
rect 31401 7905 31435 7939
rect 32137 7905 32171 7939
rect 32597 7905 32631 7939
rect 39348 7905 39382 7939
rect 8585 7837 8619 7871
rect 10517 7837 10551 7871
rect 12081 7837 12115 7871
rect 12357 7837 12391 7871
rect 16221 7837 16255 7871
rect 21649 7837 21683 7871
rect 21925 7837 21959 7871
rect 23397 7837 23431 7871
rect 24317 7837 24351 7871
rect 26617 7837 26651 7871
rect 27261 7837 27295 7871
rect 34253 7837 34287 7871
rect 36185 7837 36219 7871
rect 37841 7837 37875 7871
rect 38117 7837 38151 7871
rect 11069 7769 11103 7803
rect 15991 7769 16025 7803
rect 30297 7769 30331 7803
rect 30665 7769 30699 7803
rect 10149 7701 10183 7735
rect 15577 7701 15611 7735
rect 16129 7701 16163 7735
rect 16957 7701 16991 7735
rect 23673 7701 23707 7735
rect 25697 7701 25731 7735
rect 39451 7701 39485 7735
rect 9873 7497 9907 7531
rect 10885 7497 10919 7531
rect 11161 7497 11195 7531
rect 14381 7497 14415 7531
rect 15466 7497 15500 7531
rect 15761 7497 15795 7531
rect 17095 7497 17129 7531
rect 20729 7497 20763 7531
rect 21741 7497 21775 7531
rect 23029 7497 23063 7531
rect 24869 7497 24903 7531
rect 26341 7497 26375 7531
rect 26709 7497 26743 7531
rect 27721 7497 27755 7531
rect 28365 7497 28399 7531
rect 29469 7497 29503 7531
rect 31309 7497 31343 7531
rect 33149 7497 33183 7531
rect 33517 7497 33551 7531
rect 34253 7497 34287 7531
rect 36093 7497 36127 7531
rect 38761 7497 38795 7531
rect 39313 7497 39347 7531
rect 9505 7429 9539 7463
rect 11897 7429 11931 7463
rect 13369 7429 13403 7463
rect 15577 7429 15611 7463
rect 17417 7429 17451 7463
rect 17877 7429 17911 7463
rect 20959 7429 20993 7463
rect 23489 7429 23523 7463
rect 25559 7429 25593 7463
rect 27997 7429 28031 7463
rect 29929 7429 29963 7463
rect 31677 7429 31711 7463
rect 32781 7429 32815 7463
rect 36829 7429 36863 7463
rect 9137 7361 9171 7395
rect 13553 7361 13587 7395
rect 15117 7361 15151 7395
rect 15669 7361 15703 7395
rect 18889 7361 18923 7395
rect 21373 7361 21407 7395
rect 21833 7361 21867 7395
rect 23673 7361 23707 7395
rect 36277 7361 36311 7395
rect 37657 7361 37691 7395
rect 37749 7361 37783 7395
rect 8493 7293 8527 7327
rect 8585 7293 8619 7327
rect 8769 7293 8803 7327
rect 9965 7293 9999 7327
rect 12449 7293 12483 7327
rect 10286 7225 10320 7259
rect 12173 7225 12207 7259
rect 12770 7225 12804 7259
rect 14013 7293 14047 7327
rect 14841 7293 14875 7327
rect 15301 7293 15335 7327
rect 16865 7293 16899 7327
rect 19533 7293 19567 7327
rect 20821 7293 20855 7327
rect 22753 7293 22787 7327
rect 24593 7293 24627 7327
rect 25456 7293 25490 7327
rect 25881 7293 25915 7327
rect 26801 7293 26835 7327
rect 30113 7293 30147 7327
rect 30573 7293 30607 7327
rect 31861 7293 31895 7327
rect 33609 7293 33643 7327
rect 34932 7293 34966 7327
rect 35357 7293 35391 7327
rect 37289 7293 37323 7327
rect 38209 7293 38243 7327
rect 16313 7225 16347 7259
rect 20085 7225 20119 7259
rect 24035 7225 24069 7259
rect 27054 7225 27088 7259
rect 30849 7225 30883 7259
rect 32182 7225 32216 7259
rect 36369 7225 36403 7259
rect 13553 7157 13587 7191
rect 13645 7157 13679 7191
rect 16773 7157 16807 7191
rect 19441 7157 19475 7191
rect 22201 7157 22235 7191
rect 29009 7157 29043 7191
rect 33793 7157 33827 7191
rect 34529 7157 34563 7191
rect 35035 7157 35069 7191
rect 9505 6953 9539 6987
rect 10057 6953 10091 6987
rect 10977 6953 11011 6987
rect 12541 6953 12575 6987
rect 14151 6953 14185 6987
rect 16037 6953 16071 6987
rect 16405 6953 16439 6987
rect 17509 6953 17543 6987
rect 19441 6953 19475 6987
rect 22937 6953 22971 6987
rect 23765 6953 23799 6987
rect 24501 6953 24535 6987
rect 25191 6953 25225 6987
rect 26341 6953 26375 6987
rect 26617 6953 26651 6987
rect 27721 6953 27755 6987
rect 30297 6953 30331 6987
rect 31309 6953 31343 6987
rect 32505 6953 32539 6987
rect 33057 6953 33091 6987
rect 37013 6953 37047 6987
rect 16910 6885 16944 6919
rect 18061 6885 18095 6919
rect 18521 6885 18555 6919
rect 22103 6885 22137 6919
rect 28825 6885 28859 6919
rect 34069 6885 34103 6919
rect 36369 6885 36403 6919
rect 10241 6817 10275 6851
rect 10517 6817 10551 6851
rect 12725 6817 12759 6851
rect 12909 6817 12943 6851
rect 14048 6817 14082 6851
rect 15577 6817 15611 6851
rect 21189 6817 21223 6851
rect 22661 6817 22695 6851
rect 23489 6817 23523 6851
rect 23949 6817 23983 6851
rect 25088 6817 25122 6851
rect 26525 6817 26559 6851
rect 26985 6817 27019 6851
rect 30205 6817 30239 6851
rect 30665 6817 30699 6851
rect 32137 6817 32171 6851
rect 35484 6817 35518 6851
rect 38393 6817 38427 6851
rect 16589 6749 16623 6783
rect 18429 6749 18463 6783
rect 21741 6749 21775 6783
rect 28733 6749 28767 6783
rect 29377 6749 29411 6783
rect 33793 6749 33827 6783
rect 33977 6749 34011 6783
rect 35587 6749 35621 6783
rect 36277 6749 36311 6783
rect 37749 6749 37783 6783
rect 18981 6681 19015 6715
rect 34529 6681 34563 6715
rect 36599 6681 36633 6715
rect 11989 6613 12023 6647
rect 21557 6613 21591 6647
rect 29653 6613 29687 6647
rect 31953 6613 31987 6647
rect 9321 6409 9355 6443
rect 12265 6409 12299 6443
rect 14749 6409 14783 6443
rect 19073 6409 19107 6443
rect 21833 6409 21867 6443
rect 23857 6409 23891 6443
rect 25513 6409 25547 6443
rect 25973 6409 26007 6443
rect 27537 6409 27571 6443
rect 30297 6409 30331 6443
rect 30849 6409 30883 6443
rect 32137 6409 32171 6443
rect 34621 6409 34655 6443
rect 35909 6409 35943 6443
rect 36921 6409 36955 6443
rect 37289 6409 37323 6443
rect 38025 6409 38059 6443
rect 10057 6341 10091 6375
rect 15853 6341 15887 6375
rect 20453 6341 20487 6375
rect 24317 6341 24351 6375
rect 27077 6341 27111 6375
rect 12541 6273 12575 6307
rect 16773 6273 16807 6307
rect 17417 6273 17451 6307
rect 21373 6273 21407 6307
rect 23489 6273 23523 6307
rect 27721 6273 27755 6307
rect 28365 6273 28399 6307
rect 29377 6273 29411 6307
rect 30941 6273 30975 6307
rect 32781 6273 32815 6307
rect 33333 6273 33367 6307
rect 10425 6205 10459 6239
rect 10609 6205 10643 6239
rect 14565 6205 14599 6239
rect 16037 6205 16071 6239
rect 16497 6205 16531 6239
rect 18061 6205 18095 6239
rect 18521 6205 18555 6239
rect 19676 6205 19710 6239
rect 20177 6205 20211 6239
rect 20637 6205 20671 6239
rect 21189 6205 21223 6239
rect 22385 6205 22419 6239
rect 23029 6205 23063 6239
rect 24501 6205 24535 6239
rect 25053 6205 25087 6239
rect 26065 6205 26099 6239
rect 26525 6205 26559 6239
rect 26801 6205 26835 6239
rect 34989 6205 35023 6239
rect 36528 6205 36562 6239
rect 37540 6205 37574 6239
rect 38301 6205 38335 6239
rect 9689 6137 9723 6171
rect 10885 6137 10919 6171
rect 12633 6137 12667 6171
rect 13185 6137 13219 6171
rect 13921 6137 13955 6171
rect 15577 6137 15611 6171
rect 19763 6137 19797 6171
rect 22201 6137 22235 6171
rect 25237 6137 25271 6171
rect 27813 6137 27847 6171
rect 29469 6137 29503 6171
rect 30021 6137 30055 6171
rect 31303 6137 31337 6171
rect 33425 6137 33459 6171
rect 33977 6137 34011 6171
rect 34897 6137 34931 6171
rect 11805 6069 11839 6103
rect 14381 6069 14415 6103
rect 17049 6069 17083 6103
rect 17877 6069 17911 6103
rect 18153 6069 18187 6103
rect 22477 6069 22511 6103
rect 28733 6069 28767 6103
rect 29101 6069 29135 6103
rect 31861 6069 31895 6103
rect 33149 6069 33183 6103
rect 34345 6069 34379 6103
rect 36599 6069 36633 6103
rect 37611 6069 37645 6103
rect 10241 5865 10275 5899
rect 10885 5865 10919 5899
rect 12541 5865 12575 5899
rect 13093 5865 13127 5899
rect 18153 5865 18187 5899
rect 18521 5865 18555 5899
rect 21005 5865 21039 5899
rect 22201 5865 22235 5899
rect 26709 5865 26743 5899
rect 31033 5865 31067 5899
rect 31953 5865 31987 5899
rect 32229 5865 32263 5899
rect 33241 5865 33275 5899
rect 17325 5797 17359 5831
rect 18889 5797 18923 5831
rect 20729 5797 20763 5831
rect 24593 5797 24627 5831
rect 24869 5797 24903 5831
rect 27398 5797 27432 5831
rect 29831 5797 29865 5831
rect 30757 5797 30791 5831
rect 33793 5797 33827 5831
rect 35817 5797 35851 5831
rect 36369 5797 36403 5831
rect 13001 5729 13035 5763
rect 13461 5729 13495 5763
rect 15853 5729 15887 5763
rect 16129 5729 16163 5763
rect 20913 5729 20947 5763
rect 21465 5729 21499 5763
rect 22753 5729 22787 5763
rect 22937 5729 22971 5763
rect 27077 5729 27111 5763
rect 29469 5729 29503 5763
rect 32137 5729 32171 5763
rect 32597 5729 32631 5763
rect 34437 5729 34471 5763
rect 37657 5729 37691 5763
rect 10517 5661 10551 5695
rect 16221 5661 16255 5695
rect 17233 5661 17267 5695
rect 17509 5661 17543 5695
rect 18797 5661 18831 5695
rect 19073 5661 19107 5695
rect 23121 5661 23155 5695
rect 24777 5661 24811 5695
rect 25421 5661 25455 5695
rect 28733 5661 28767 5695
rect 35725 5661 35759 5695
rect 11437 5525 11471 5559
rect 12817 5525 12851 5559
rect 26065 5525 26099 5559
rect 27997 5525 28031 5559
rect 29377 5525 29411 5559
rect 30389 5525 30423 5559
rect 37887 5525 37921 5559
rect 10149 5321 10183 5355
rect 10517 5321 10551 5355
rect 11529 5321 11563 5355
rect 12725 5321 12759 5355
rect 15393 5321 15427 5355
rect 16865 5321 16899 5355
rect 17233 5321 17267 5355
rect 18981 5321 19015 5355
rect 19257 5321 19291 5355
rect 20177 5321 20211 5355
rect 21281 5321 21315 5355
rect 22845 5321 22879 5355
rect 23213 5321 23247 5355
rect 24133 5321 24167 5355
rect 27905 5321 27939 5355
rect 30297 5321 30331 5355
rect 30849 5321 30883 5355
rect 32137 5321 32171 5355
rect 34161 5321 34195 5355
rect 36921 5321 36955 5355
rect 37933 5321 37967 5355
rect 38301 5321 38335 5355
rect 13001 5253 13035 5287
rect 25789 5253 25823 5287
rect 26249 5253 26283 5287
rect 27537 5253 27571 5287
rect 31861 5253 31895 5287
rect 34621 5253 34655 5287
rect 13185 5185 13219 5219
rect 14381 5185 14415 5219
rect 17785 5185 17819 5219
rect 18061 5185 18095 5219
rect 26341 5185 26375 5219
rect 29837 5185 29871 5219
rect 30941 5185 30975 5219
rect 10609 5117 10643 5151
rect 11805 5117 11839 5151
rect 15577 5117 15611 5151
rect 16129 5117 16163 5151
rect 20269 5117 20303 5151
rect 20821 5117 20855 5151
rect 21741 5117 21775 5151
rect 21833 5117 21867 5151
rect 22385 5117 22419 5151
rect 24593 5117 24627 5151
rect 28124 5117 28158 5151
rect 28549 5117 28583 5151
rect 32597 5117 32631 5151
rect 32689 5117 32723 5151
rect 33241 5117 33275 5151
rect 33701 5117 33735 5151
rect 34932 5117 34966 5151
rect 36553 5117 36587 5151
rect 37473 5117 37507 5151
rect 10930 5049 10964 5083
rect 13506 5049 13540 5083
rect 15117 5049 15151 5083
rect 18382 5049 18416 5083
rect 21005 5049 21039 5083
rect 22569 5049 22603 5083
rect 24501 5049 24535 5083
rect 24955 5049 24989 5083
rect 26703 5049 26737 5083
rect 29377 5049 29411 5083
rect 29469 5049 29503 5083
rect 31262 5049 31296 5083
rect 36645 5049 36679 5083
rect 9597 4981 9631 5015
rect 14105 4981 14139 5015
rect 15669 4981 15703 5015
rect 25513 4981 25547 5015
rect 27261 4981 27295 5015
rect 28227 4981 28261 5015
rect 29101 4981 29135 5015
rect 32781 4981 32815 5015
rect 35035 4981 35069 5015
rect 35725 4981 35759 5015
rect 37657 4981 37691 5015
rect 10609 4777 10643 4811
rect 11345 4777 11379 4811
rect 12035 4777 12069 4811
rect 15669 4777 15703 4811
rect 16037 4777 16071 4811
rect 17049 4777 17083 4811
rect 18889 4777 18923 4811
rect 20361 4777 20395 4811
rect 21097 4777 21131 4811
rect 22569 4777 22603 4811
rect 24409 4777 24443 4811
rect 27537 4777 27571 4811
rect 30297 4777 30331 4811
rect 36001 4777 36035 4811
rect 12449 4709 12483 4743
rect 13461 4709 13495 4743
rect 14657 4709 14691 4743
rect 16450 4709 16484 4743
rect 23483 4709 23517 4743
rect 24777 4709 24811 4743
rect 25053 4709 25087 4743
rect 26709 4709 26743 4743
rect 29463 4709 29497 4743
rect 32597 4709 32631 4743
rect 34161 4709 34195 4743
rect 36093 4709 36127 4743
rect 10517 4641 10551 4675
rect 10793 4641 10827 4675
rect 11964 4641 11998 4675
rect 16129 4641 16163 4675
rect 17877 4641 17911 4675
rect 18429 4641 18463 4675
rect 19441 4641 19475 4675
rect 19625 4641 19659 4675
rect 21465 4641 21499 4675
rect 22017 4641 22051 4675
rect 23121 4641 23155 4675
rect 28156 4641 28190 4675
rect 31100 4641 31134 4675
rect 36737 4641 36771 4675
rect 13001 4573 13035 4607
rect 13369 4573 13403 4607
rect 13645 4573 13679 4607
rect 18521 4573 18555 4607
rect 22201 4573 22235 4607
rect 24961 4573 24995 4607
rect 26617 4573 26651 4607
rect 27261 4573 27295 4607
rect 29009 4573 29043 4607
rect 29101 4573 29135 4607
rect 32505 4573 32539 4607
rect 34069 4573 34103 4607
rect 25513 4505 25547 4539
rect 33057 4505 33091 4539
rect 34621 4505 34655 4539
rect 14289 4437 14323 4471
rect 15117 4437 15151 4471
rect 17785 4437 17819 4471
rect 19717 4437 19751 4471
rect 22937 4437 22971 4471
rect 24041 4437 24075 4471
rect 28227 4437 28261 4471
rect 30021 4437 30055 4471
rect 30941 4437 30975 4471
rect 31171 4437 31205 4471
rect 34989 4437 35023 4471
rect 38025 4437 38059 4471
rect 10057 4233 10091 4267
rect 12265 4233 12299 4267
rect 16497 4233 16531 4267
rect 17095 4233 17129 4267
rect 17509 4233 17543 4267
rect 17877 4233 17911 4267
rect 19533 4233 19567 4267
rect 20177 4233 20211 4267
rect 22017 4233 22051 4267
rect 22477 4233 22511 4267
rect 28641 4233 28675 4267
rect 28825 4233 28859 4267
rect 30389 4233 30423 4267
rect 30757 4233 30791 4267
rect 33517 4233 33551 4267
rect 36001 4233 36035 4267
rect 37841 4233 37875 4267
rect 10425 4165 10459 4199
rect 11437 4165 11471 4199
rect 26709 4165 26743 4199
rect 28181 4165 28215 4199
rect 29101 4165 29135 4199
rect 32229 4165 32263 4199
rect 33057 4165 33091 4199
rect 10885 4097 10919 4131
rect 11805 4097 11839 4131
rect 12909 4097 12943 4131
rect 14197 4097 14231 4131
rect 18429 4097 18463 4131
rect 19763 4097 19797 4131
rect 20821 4097 20855 4131
rect 26801 4097 26835 4131
rect 28825 4097 28859 4131
rect 29377 4097 29411 4131
rect 30021 4097 30055 4131
rect 32505 4097 32539 4131
rect 34989 4097 35023 4131
rect 35633 4097 35667 4131
rect 36553 4097 36587 4131
rect 36829 4097 36863 4131
rect 38117 4097 38151 4131
rect 38393 4097 38427 4131
rect 12449 4029 12483 4063
rect 12633 4029 12667 4063
rect 13277 4029 13311 4063
rect 13829 4029 13863 4063
rect 15669 4029 15703 4063
rect 16992 4029 17026 4063
rect 19660 4029 19694 4063
rect 22636 4029 22670 4063
rect 23673 4029 23707 4063
rect 25640 4029 25674 4063
rect 10977 3961 11011 3995
rect 18153 3961 18187 3995
rect 18245 3961 18279 3995
rect 20729 3961 20763 3995
rect 21142 3961 21176 3995
rect 23213 3961 23247 3995
rect 24035 3961 24069 3995
rect 27163 3961 27197 3995
rect 29469 3961 29503 3995
rect 30941 3961 30975 3995
rect 31033 3961 31067 3995
rect 31585 3961 31619 3995
rect 32597 3961 32631 3995
rect 34713 3961 34747 3995
rect 35081 3961 35115 3995
rect 36645 3961 36679 3995
rect 38209 3961 38243 3995
rect 13645 3893 13679 3927
rect 16129 3893 16163 3927
rect 16773 3893 16807 3927
rect 19073 3893 19107 3927
rect 21741 3893 21775 3927
rect 22707 3893 22741 3927
rect 24593 3893 24627 3927
rect 24961 3893 24995 3927
rect 25237 3893 25271 3927
rect 25743 3893 25777 3927
rect 26341 3893 26375 3927
rect 27721 3893 27755 3927
rect 31953 3893 31987 3927
rect 33977 3893 34011 3927
rect 36369 3893 36403 3927
rect 11023 3689 11057 3723
rect 11437 3689 11471 3723
rect 14565 3689 14599 3723
rect 16037 3689 16071 3723
rect 16589 3689 16623 3723
rect 17141 3689 17175 3723
rect 17877 3689 17911 3723
rect 20729 3689 20763 3723
rect 24133 3689 24167 3723
rect 25881 3689 25915 3723
rect 26663 3689 26697 3723
rect 26985 3689 27019 3723
rect 29745 3689 29779 3723
rect 30389 3689 30423 3723
rect 33149 3689 33183 3723
rect 34713 3689 34747 3723
rect 36553 3689 36587 3723
rect 18153 3621 18187 3655
rect 22931 3621 22965 3655
rect 23857 3621 23891 3655
rect 25053 3621 25087 3655
rect 25605 3621 25639 3655
rect 28181 3621 28215 3655
rect 28733 3621 28767 3655
rect 30573 3621 30607 3655
rect 30665 3621 30699 3655
rect 32321 3621 32355 3655
rect 33885 3621 33919 3655
rect 35541 3621 35575 3655
rect 10952 3553 10986 3587
rect 13737 3553 13771 3587
rect 19568 3553 19602 3587
rect 20913 3553 20947 3587
rect 21373 3553 21407 3587
rect 22569 3553 22603 3587
rect 26433 3553 26467 3587
rect 29377 3553 29411 3587
rect 30389 3553 30423 3587
rect 35633 3553 35667 3587
rect 37749 3553 37783 3587
rect 11897 3485 11931 3519
rect 12265 3485 12299 3519
rect 16221 3485 16255 3519
rect 18061 3485 18095 3519
rect 18337 3485 18371 3519
rect 21465 3485 21499 3519
rect 24961 3485 24995 3519
rect 28089 3485 28123 3519
rect 31217 3485 31251 3519
rect 32229 3485 32263 3519
rect 32505 3485 32539 3519
rect 33793 3485 33827 3519
rect 37105 3485 37139 3519
rect 14841 3417 14875 3451
rect 21925 3417 21959 3451
rect 34345 3417 34379 3451
rect 9229 3349 9263 3383
rect 11713 3349 11747 3383
rect 14197 3349 14231 3383
rect 19073 3349 19107 3383
rect 19671 3349 19705 3383
rect 23489 3349 23523 3383
rect 24777 3349 24811 3383
rect 27721 3349 27755 3383
rect 37933 3349 37967 3383
rect 8677 3145 8711 3179
rect 11529 3145 11563 3179
rect 12955 3145 12989 3179
rect 16129 3145 16163 3179
rect 16773 3145 16807 3179
rect 17095 3145 17129 3179
rect 17877 3145 17911 3179
rect 19901 3145 19935 3179
rect 20729 3145 20763 3179
rect 22937 3145 22971 3179
rect 23305 3145 23339 3179
rect 23811 3145 23845 3179
rect 26065 3145 26099 3179
rect 26525 3145 26559 3179
rect 26755 3145 26789 3179
rect 27169 3145 27203 3179
rect 29009 3145 29043 3179
rect 30389 3145 30423 3179
rect 32045 3145 32079 3179
rect 33241 3145 33275 3179
rect 34253 3145 34287 3179
rect 38209 3145 38243 3179
rect 16497 3077 16531 3111
rect 20361 3077 20395 3111
rect 22661 3077 22695 3111
rect 9597 3009 9631 3043
rect 13645 3009 13679 3043
rect 13829 3009 13863 3043
rect 18981 3009 19015 3043
rect 19257 3009 19291 3043
rect 21189 3009 21223 3043
rect 25421 3009 25455 3043
rect 27721 3009 27755 3043
rect 28365 3009 28399 3043
rect 31217 3009 31251 3043
rect 32229 3009 32263 3043
rect 36277 3009 36311 3043
rect 36921 3009 36955 3043
rect 37197 3009 37231 3043
rect 37841 3009 37875 3043
rect 9229 2941 9263 2975
rect 11069 2941 11103 2975
rect 12633 2941 12667 2975
rect 12817 2941 12851 2975
rect 14197 2941 14231 2975
rect 15669 2941 15703 2975
rect 16992 2941 17026 2975
rect 17417 2941 17451 2975
rect 23708 2941 23742 2975
rect 24133 2941 24167 2975
rect 26684 2941 26718 2975
rect 29520 2941 29554 2975
rect 31769 2941 31803 2975
rect 32321 2941 32355 2975
rect 33828 2941 33862 2975
rect 34713 2941 34747 2975
rect 36185 2941 36219 2975
rect 13277 2873 13311 2907
rect 18797 2873 18831 2907
rect 19073 2873 19107 2907
rect 21097 2873 21131 2907
rect 21551 2873 21585 2907
rect 24777 2873 24811 2907
rect 24869 2873 24903 2907
rect 27537 2873 27571 2907
rect 27813 2873 27847 2907
rect 29607 2873 29641 2907
rect 30573 2873 30607 2907
rect 30665 2873 30699 2907
rect 37289 2873 37323 2907
rect 9045 2805 9079 2839
rect 11897 2805 11931 2839
rect 18245 2805 18279 2839
rect 22109 2805 22143 2839
rect 24593 2805 24627 2839
rect 25789 2805 25823 2839
rect 28733 2805 28767 2839
rect 30021 2805 30055 2839
rect 33609 2805 33643 2839
rect 33931 2805 33965 2839
rect 35449 2805 35483 2839
rect 11989 2601 12023 2635
rect 12449 2601 12483 2635
rect 12909 2601 12943 2635
rect 14289 2601 14323 2635
rect 15669 2601 15703 2635
rect 16129 2601 16163 2635
rect 16589 2601 16623 2635
rect 17141 2601 17175 2635
rect 19441 2601 19475 2635
rect 21005 2601 21039 2635
rect 22293 2601 22327 2635
rect 24409 2601 24443 2635
rect 28595 2601 28629 2635
rect 31125 2601 31159 2635
rect 31631 2601 31665 2635
rect 34345 2601 34379 2635
rect 35265 2601 35299 2635
rect 37151 2601 37185 2635
rect 37565 2601 37599 2635
rect 10655 2533 10689 2567
rect 18061 2533 18095 2567
rect 18842 2533 18876 2567
rect 21694 2533 21728 2567
rect 25053 2533 25087 2567
rect 25145 2533 25179 2567
rect 26709 2533 26743 2567
rect 27077 2533 27111 2567
rect 28273 2533 28307 2567
rect 29561 2533 29595 2567
rect 29929 2533 29963 2567
rect 30757 2533 30791 2567
rect 33793 2533 33827 2567
rect 35633 2533 35667 2567
rect 36185 2533 36219 2567
rect 10568 2465 10602 2499
rect 11564 2465 11598 2499
rect 13829 2465 13863 2499
rect 14432 2465 14466 2499
rect 14841 2465 14875 2499
rect 16221 2465 16255 2499
rect 17785 2465 17819 2499
rect 18521 2465 18555 2499
rect 20637 2465 20671 2499
rect 21373 2465 21407 2499
rect 28492 2465 28526 2499
rect 31560 2465 31594 2499
rect 31953 2465 31987 2499
rect 32413 2465 32447 2499
rect 33241 2465 33275 2499
rect 34161 2465 34195 2499
rect 34621 2465 34655 2499
rect 37080 2465 37114 2499
rect 13369 2397 13403 2431
rect 14519 2397 14553 2431
rect 24869 2397 24903 2431
rect 25421 2397 25455 2431
rect 26985 2397 27019 2431
rect 27261 2397 27295 2431
rect 29837 2397 29871 2431
rect 30113 2397 30147 2431
rect 33333 2397 33367 2431
rect 35541 2397 35575 2431
rect 36461 2397 36495 2431
rect 29101 2329 29135 2363
rect 9229 2261 9263 2295
rect 11069 2261 11103 2295
rect 11437 2261 11471 2295
rect 11667 2261 11701 2295
rect 26249 2261 26283 2295
<< metal1 >>
rect 13814 49512 13820 49564
rect 13872 49552 13878 49564
rect 16114 49552 16120 49564
rect 13872 49524 16120 49552
rect 13872 49512 13878 49524
rect 16114 49512 16120 49524
rect 16172 49512 16178 49564
rect 19426 49512 19432 49564
rect 19484 49552 19490 49564
rect 20254 49552 20260 49564
rect 19484 49524 20260 49552
rect 19484 49512 19490 49524
rect 20254 49512 20260 49524
rect 20312 49512 20318 49564
rect 24210 49512 24216 49564
rect 24268 49552 24274 49564
rect 24946 49552 24952 49564
rect 24268 49524 24952 49552
rect 24268 49512 24274 49524
rect 24946 49512 24952 49524
rect 25004 49512 25010 49564
rect 1104 47354 48852 47376
rect 1104 47302 19606 47354
rect 19658 47302 19670 47354
rect 19722 47302 19734 47354
rect 19786 47302 19798 47354
rect 19850 47302 48852 47354
rect 1104 47280 48852 47302
rect 1104 46810 48852 46832
rect 1104 46758 4246 46810
rect 4298 46758 4310 46810
rect 4362 46758 4374 46810
rect 4426 46758 4438 46810
rect 4490 46758 34966 46810
rect 35018 46758 35030 46810
rect 35082 46758 35094 46810
rect 35146 46758 35158 46810
rect 35210 46758 48852 46810
rect 1104 46736 48852 46758
rect 1104 46266 48852 46288
rect 1104 46214 19606 46266
rect 19658 46214 19670 46266
rect 19722 46214 19734 46266
rect 19786 46214 19798 46266
rect 19850 46214 48852 46266
rect 1104 46192 48852 46214
rect 1104 45722 48852 45744
rect 1104 45670 4246 45722
rect 4298 45670 4310 45722
rect 4362 45670 4374 45722
rect 4426 45670 4438 45722
rect 4490 45670 34966 45722
rect 35018 45670 35030 45722
rect 35082 45670 35094 45722
rect 35146 45670 35158 45722
rect 35210 45670 48852 45722
rect 1104 45648 48852 45670
rect 1104 45178 48852 45200
rect 1104 45126 19606 45178
rect 19658 45126 19670 45178
rect 19722 45126 19734 45178
rect 19786 45126 19798 45178
rect 19850 45126 48852 45178
rect 1104 45104 48852 45126
rect 1104 44634 48852 44656
rect 1104 44582 4246 44634
rect 4298 44582 4310 44634
rect 4362 44582 4374 44634
rect 4426 44582 4438 44634
rect 4490 44582 34966 44634
rect 35018 44582 35030 44634
rect 35082 44582 35094 44634
rect 35146 44582 35158 44634
rect 35210 44582 48852 44634
rect 1104 44560 48852 44582
rect 1104 44090 48852 44112
rect 1104 44038 19606 44090
rect 19658 44038 19670 44090
rect 19722 44038 19734 44090
rect 19786 44038 19798 44090
rect 19850 44038 48852 44090
rect 1104 44016 48852 44038
rect 1104 43546 48852 43568
rect 1104 43494 4246 43546
rect 4298 43494 4310 43546
rect 4362 43494 4374 43546
rect 4426 43494 4438 43546
rect 4490 43494 34966 43546
rect 35018 43494 35030 43546
rect 35082 43494 35094 43546
rect 35146 43494 35158 43546
rect 35210 43494 48852 43546
rect 1104 43472 48852 43494
rect 1104 43002 48852 43024
rect 1104 42950 19606 43002
rect 19658 42950 19670 43002
rect 19722 42950 19734 43002
rect 19786 42950 19798 43002
rect 19850 42950 48852 43002
rect 1104 42928 48852 42950
rect 21336 42755 21394 42761
rect 21336 42721 21348 42755
rect 21382 42752 21394 42755
rect 21818 42752 21824 42764
rect 21382 42724 21824 42752
rect 21382 42721 21394 42724
rect 21336 42715 21394 42721
rect 21818 42712 21824 42724
rect 21876 42712 21882 42764
rect 21407 42551 21465 42557
rect 21407 42517 21419 42551
rect 21453 42548 21465 42551
rect 21634 42548 21640 42560
rect 21453 42520 21640 42548
rect 21453 42517 21465 42520
rect 21407 42511 21465 42517
rect 21634 42508 21640 42520
rect 21692 42508 21698 42560
rect 1104 42458 48852 42480
rect 1104 42406 4246 42458
rect 4298 42406 4310 42458
rect 4362 42406 4374 42458
rect 4426 42406 4438 42458
rect 4490 42406 34966 42458
rect 35018 42406 35030 42458
rect 35082 42406 35094 42458
rect 35146 42406 35158 42458
rect 35210 42406 48852 42458
rect 1104 42384 48852 42406
rect 14182 42100 14188 42152
rect 14240 42140 14246 42152
rect 21396 42143 21454 42149
rect 21396 42140 21408 42143
rect 14240 42112 21408 42140
rect 14240 42100 14246 42112
rect 21396 42109 21408 42112
rect 21442 42140 21454 42143
rect 22189 42143 22247 42149
rect 22189 42140 22201 42143
rect 21442 42112 22201 42140
rect 21442 42109 21454 42112
rect 21396 42103 21454 42109
rect 22189 42109 22201 42112
rect 22235 42140 22247 42143
rect 24302 42140 24308 42152
rect 22235 42112 24308 42140
rect 22235 42109 22247 42112
rect 22189 42103 22247 42109
rect 24302 42100 24308 42112
rect 24360 42100 24366 42152
rect 24464 42143 24522 42149
rect 24464 42109 24476 42143
rect 24510 42140 24522 42143
rect 24854 42140 24860 42152
rect 24510 42112 24860 42140
rect 24510 42109 24522 42112
rect 24464 42103 24522 42109
rect 24854 42100 24860 42112
rect 24912 42100 24918 42152
rect 21499 42007 21557 42013
rect 21499 41973 21511 42007
rect 21545 42004 21557 42007
rect 21726 42004 21732 42016
rect 21545 41976 21732 42004
rect 21545 41973 21557 41976
rect 21499 41967 21557 41973
rect 21726 41964 21732 41976
rect 21784 41964 21790 42016
rect 21818 41964 21824 42016
rect 21876 42004 21882 42016
rect 24535 42007 24593 42013
rect 21876 41976 21921 42004
rect 21876 41964 21882 41976
rect 24535 41973 24547 42007
rect 24581 42004 24593 42007
rect 24762 42004 24768 42016
rect 24581 41976 24768 42004
rect 24581 41973 24593 41976
rect 24535 41967 24593 41973
rect 24762 41964 24768 41976
rect 24820 41964 24826 42016
rect 24854 41964 24860 42016
rect 24912 42004 24918 42016
rect 30374 42004 30380 42016
rect 24912 41976 30380 42004
rect 24912 41964 24918 41976
rect 30374 41964 30380 41976
rect 30432 41964 30438 42016
rect 1104 41914 48852 41936
rect 1104 41862 19606 41914
rect 19658 41862 19670 41914
rect 19722 41862 19734 41914
rect 19786 41862 19798 41914
rect 19850 41862 48852 41914
rect 1104 41840 48852 41862
rect 24762 41760 24768 41812
rect 24820 41800 24826 41812
rect 24857 41803 24915 41809
rect 24857 41800 24869 41803
rect 24820 41772 24869 41800
rect 24820 41760 24826 41772
rect 24857 41769 24869 41772
rect 24903 41769 24915 41803
rect 24857 41763 24915 41769
rect 21729 41735 21787 41741
rect 21729 41701 21741 41735
rect 21775 41732 21787 41735
rect 21910 41732 21916 41744
rect 21775 41704 21916 41732
rect 21775 41701 21787 41704
rect 21729 41695 21787 41701
rect 21910 41692 21916 41704
rect 21968 41692 21974 41744
rect 16644 41667 16702 41673
rect 16644 41633 16656 41667
rect 16690 41664 16702 41667
rect 17494 41664 17500 41676
rect 16690 41636 17500 41664
rect 16690 41633 16702 41636
rect 16644 41627 16702 41633
rect 17494 41624 17500 41636
rect 17552 41624 17558 41676
rect 18944 41667 19002 41673
rect 18944 41633 18956 41667
rect 18990 41664 19002 41667
rect 19058 41664 19064 41676
rect 18990 41636 19064 41664
rect 18990 41633 19002 41636
rect 18944 41627 19002 41633
rect 19058 41624 19064 41636
rect 19116 41624 19122 41676
rect 24210 41664 24216 41676
rect 24171 41636 24216 41664
rect 24210 41624 24216 41636
rect 24268 41624 24274 41676
rect 25292 41667 25350 41673
rect 25292 41633 25304 41667
rect 25338 41664 25350 41667
rect 25958 41664 25964 41676
rect 25338 41636 25964 41664
rect 25338 41633 25350 41636
rect 25292 41627 25350 41633
rect 25958 41624 25964 41636
rect 26016 41624 26022 41676
rect 26640 41667 26698 41673
rect 26640 41664 26652 41667
rect 26620 41633 26652 41664
rect 26686 41633 26698 41667
rect 26620 41627 26698 41633
rect 29708 41667 29766 41673
rect 29708 41633 29720 41667
rect 29754 41664 29766 41667
rect 30190 41664 30196 41676
rect 29754 41636 30196 41664
rect 29754 41633 29766 41636
rect 29708 41627 29766 41633
rect 21634 41596 21640 41608
rect 21595 41568 21640 41596
rect 21634 41556 21640 41568
rect 21692 41556 21698 41608
rect 22278 41596 22284 41608
rect 22239 41568 22284 41596
rect 22278 41556 22284 41568
rect 22336 41556 22342 41608
rect 26620 41596 26648 41627
rect 30190 41624 30196 41636
rect 30248 41624 30254 41676
rect 32122 41624 32128 41676
rect 32180 41664 32186 41676
rect 32528 41667 32586 41673
rect 32528 41664 32540 41667
rect 32180 41636 32540 41664
rect 32180 41624 32186 41636
rect 32528 41633 32540 41636
rect 32574 41633 32586 41667
rect 32528 41627 32586 41633
rect 27430 41596 27436 41608
rect 23446 41568 27436 41596
rect 23198 41488 23204 41540
rect 23256 41528 23262 41540
rect 23446 41528 23474 41568
rect 27430 41556 27436 41568
rect 27488 41556 27494 41608
rect 23256 41500 23474 41528
rect 23256 41488 23262 41500
rect 16482 41460 16488 41472
rect 16443 41432 16488 41460
rect 16482 41420 16488 41432
rect 16540 41420 16546 41472
rect 16574 41420 16580 41472
rect 16632 41460 16638 41472
rect 16715 41463 16773 41469
rect 16715 41460 16727 41463
rect 16632 41432 16727 41460
rect 16632 41420 16638 41432
rect 16715 41429 16727 41432
rect 16761 41429 16773 41463
rect 16715 41423 16773 41429
rect 19015 41463 19073 41469
rect 19015 41429 19027 41463
rect 19061 41460 19073 41463
rect 19150 41460 19156 41472
rect 19061 41432 19156 41460
rect 19061 41429 19073 41432
rect 19015 41423 19073 41429
rect 19150 41420 19156 41432
rect 19208 41420 19214 41472
rect 19426 41460 19432 41472
rect 19387 41432 19432 41460
rect 19426 41420 19432 41432
rect 19484 41420 19490 41472
rect 19702 41460 19708 41472
rect 19663 41432 19708 41460
rect 19702 41420 19708 41432
rect 19760 41420 19766 41472
rect 24351 41463 24409 41469
rect 24351 41429 24363 41463
rect 24397 41460 24409 41463
rect 24578 41460 24584 41472
rect 24397 41432 24584 41460
rect 24397 41429 24409 41432
rect 24351 41423 24409 41429
rect 24578 41420 24584 41432
rect 24636 41420 24642 41472
rect 24946 41420 24952 41472
rect 25004 41460 25010 41472
rect 25363 41463 25421 41469
rect 25363 41460 25375 41463
rect 25004 41432 25375 41460
rect 25004 41420 25010 41432
rect 25363 41429 25375 41432
rect 25409 41429 25421 41463
rect 25363 41423 25421 41429
rect 26743 41463 26801 41469
rect 26743 41429 26755 41463
rect 26789 41460 26801 41463
rect 26878 41460 26884 41472
rect 26789 41432 26884 41460
rect 26789 41429 26801 41432
rect 26743 41423 26801 41429
rect 26878 41420 26884 41432
rect 26936 41420 26942 41472
rect 29779 41463 29837 41469
rect 29779 41429 29791 41463
rect 29825 41460 29837 41463
rect 30098 41460 30104 41472
rect 29825 41432 30104 41460
rect 29825 41429 29837 41432
rect 29779 41423 29837 41429
rect 30098 41420 30104 41432
rect 30156 41420 30162 41472
rect 32631 41463 32689 41469
rect 32631 41429 32643 41463
rect 32677 41460 32689 41463
rect 32766 41460 32772 41472
rect 32677 41432 32772 41460
rect 32677 41429 32689 41432
rect 32631 41423 32689 41429
rect 32766 41420 32772 41432
rect 32824 41420 32830 41472
rect 1104 41370 48852 41392
rect 1104 41318 4246 41370
rect 4298 41318 4310 41370
rect 4362 41318 4374 41370
rect 4426 41318 4438 41370
rect 4490 41318 34966 41370
rect 35018 41318 35030 41370
rect 35082 41318 35094 41370
rect 35146 41318 35158 41370
rect 35210 41318 48852 41370
rect 1104 41296 48852 41318
rect 19058 41256 19064 41268
rect 19019 41228 19064 41256
rect 19058 41216 19064 41228
rect 19116 41216 19122 41268
rect 21634 41216 21640 41268
rect 21692 41256 21698 41268
rect 22557 41259 22615 41265
rect 22557 41256 22569 41259
rect 21692 41228 22569 41256
rect 21692 41216 21698 41228
rect 22557 41225 22569 41228
rect 22603 41225 22615 41259
rect 27430 41256 27436 41268
rect 27391 41228 27436 41256
rect 22557 41219 22615 41225
rect 27430 41216 27436 41228
rect 27488 41256 27494 41268
rect 31573 41259 31631 41265
rect 31573 41256 31585 41259
rect 27488 41228 31585 41256
rect 27488 41216 27494 41228
rect 31573 41225 31585 41228
rect 31619 41225 31631 41259
rect 31573 41219 31631 41225
rect 19886 41188 19892 41200
rect 19799 41160 19892 41188
rect 19886 41148 19892 41160
rect 19944 41188 19950 41200
rect 22278 41188 22284 41200
rect 19944 41160 22284 41188
rect 19944 41148 19950 41160
rect 22278 41148 22284 41160
rect 22336 41148 22342 41200
rect 24302 41148 24308 41200
rect 24360 41188 24366 41200
rect 26881 41191 26939 41197
rect 26881 41188 26893 41191
rect 24360 41160 26893 41188
rect 24360 41148 24366 41160
rect 26881 41157 26893 41160
rect 26927 41188 26939 41191
rect 27065 41191 27123 41197
rect 27065 41188 27077 41191
rect 26927 41160 27077 41188
rect 26927 41157 26939 41160
rect 26881 41151 26939 41157
rect 27065 41157 27077 41160
rect 27111 41188 27123 41191
rect 30926 41188 30932 41200
rect 27111 41160 30932 41188
rect 27111 41157 27123 41160
rect 27065 41151 27123 41157
rect 30926 41148 30932 41160
rect 30984 41148 30990 41200
rect 32122 41148 32128 41200
rect 32180 41188 32186 41200
rect 32677 41191 32735 41197
rect 32677 41188 32689 41191
rect 32180 41160 32689 41188
rect 32180 41148 32186 41160
rect 32677 41157 32689 41160
rect 32723 41157 32735 41191
rect 32677 41151 32735 41157
rect 14550 41080 14556 41132
rect 14608 41120 14614 41132
rect 16482 41120 16488 41132
rect 14608 41092 16488 41120
rect 14608 41080 14614 41092
rect 16482 41080 16488 41092
rect 16540 41120 16546 41132
rect 18371 41123 18429 41129
rect 16540 41092 16896 41120
rect 16540 41080 16546 41092
rect 14274 41012 14280 41064
rect 14332 41052 14338 41064
rect 16868 41061 16896 41092
rect 18371 41089 18383 41123
rect 18417 41120 18429 41123
rect 19337 41123 19395 41129
rect 19337 41120 19349 41123
rect 18417 41092 19349 41120
rect 18417 41089 18429 41092
rect 18371 41083 18429 41089
rect 19337 41089 19349 41092
rect 19383 41120 19395 41123
rect 19702 41120 19708 41132
rect 19383 41092 19708 41120
rect 19383 41089 19395 41092
rect 19337 41083 19395 41089
rect 19702 41080 19708 41092
rect 19760 41080 19766 41132
rect 20717 41123 20775 41129
rect 20717 41089 20729 41123
rect 20763 41120 20775 41123
rect 21637 41123 21695 41129
rect 21637 41120 21649 41123
rect 20763 41092 21649 41120
rect 20763 41089 20775 41092
rect 20717 41083 20775 41089
rect 21637 41089 21649 41092
rect 21683 41120 21695 41123
rect 23799 41123 23857 41129
rect 23799 41120 23811 41123
rect 21683 41092 23811 41120
rect 21683 41089 21695 41092
rect 21637 41083 21695 41089
rect 23799 41089 23811 41092
rect 23845 41089 23857 41123
rect 23799 41083 23857 41089
rect 24762 41080 24768 41132
rect 24820 41120 24826 41132
rect 24949 41123 25007 41129
rect 24949 41120 24961 41123
rect 24820 41092 24961 41120
rect 24820 41080 24826 41092
rect 24949 41089 24961 41092
rect 24995 41089 25007 41123
rect 24949 41083 25007 41089
rect 25593 41123 25651 41129
rect 25593 41089 25605 41123
rect 25639 41120 25651 41123
rect 27246 41120 27252 41132
rect 25639 41092 27252 41120
rect 25639 41089 25651 41092
rect 25593 41083 25651 41089
rect 27246 41080 27252 41092
rect 27304 41080 27310 41132
rect 30561 41123 30619 41129
rect 30561 41089 30573 41123
rect 30607 41120 30619 41123
rect 35526 41120 35532 41132
rect 30607 41092 35532 41120
rect 30607 41089 30619 41092
rect 30561 41083 30619 41089
rect 14404 41055 14462 41061
rect 14404 41052 14416 41055
rect 14332 41024 14416 41052
rect 14332 41012 14338 41024
rect 14404 41021 14416 41024
rect 14450 41052 14462 41055
rect 14829 41055 14887 41061
rect 14829 41052 14841 41055
rect 14450 41024 14841 41052
rect 14450 41021 14462 41024
rect 14404 41015 14462 41021
rect 14829 41021 14841 41024
rect 14875 41021 14887 41055
rect 14829 41015 14887 41021
rect 16301 41055 16359 41061
rect 16301 41021 16313 41055
rect 16347 41052 16359 41055
rect 16393 41055 16451 41061
rect 16393 41052 16405 41055
rect 16347 41024 16405 41052
rect 16347 41021 16359 41024
rect 16301 41015 16359 41021
rect 16393 41021 16405 41024
rect 16439 41021 16451 41055
rect 16393 41015 16451 41021
rect 16853 41055 16911 41061
rect 16853 41021 16865 41055
rect 16899 41021 16911 41055
rect 17494 41052 17500 41064
rect 17407 41024 17500 41052
rect 16853 41015 16911 41021
rect 16408 40984 16436 41015
rect 17494 41012 17500 41024
rect 17552 41052 17558 41064
rect 18284 41055 18342 41061
rect 18284 41052 18296 41055
rect 17552 41024 18296 41052
rect 17552 41012 17558 41024
rect 18284 41021 18296 41024
rect 18330 41052 18342 41055
rect 18598 41052 18604 41064
rect 18330 41024 18604 41052
rect 18330 41021 18342 41024
rect 18284 41015 18342 41021
rect 18598 41012 18604 41024
rect 18656 41052 18662 41064
rect 18782 41052 18788 41064
rect 18656 41024 18788 41052
rect 18656 41012 18662 41024
rect 18782 41012 18788 41024
rect 18840 41012 18846 41064
rect 23569 41055 23627 41061
rect 23569 41021 23581 41055
rect 23615 41021 23627 41055
rect 23569 41015 23627 41021
rect 26672 41055 26730 41061
rect 26672 41021 26684 41055
rect 26718 41052 26730 41055
rect 26881 41055 26939 41061
rect 26881 41052 26893 41055
rect 26718 41024 26893 41052
rect 26718 41021 26730 41024
rect 26672 41015 26730 41021
rect 26881 41021 26893 41024
rect 26927 41021 26939 41055
rect 26881 41015 26939 41021
rect 29708 41055 29766 41061
rect 29708 41021 29720 41055
rect 29754 41052 29766 41055
rect 30374 41052 30380 41064
rect 29754 41024 30380 41052
rect 29754 41021 29766 41024
rect 29708 41015 29766 41021
rect 18414 40984 18420 40996
rect 16408 40956 18420 40984
rect 18414 40944 18420 40956
rect 18472 40944 18478 40996
rect 19426 40984 19432 40996
rect 19387 40956 19432 40984
rect 19426 40944 19432 40956
rect 19484 40944 19490 40996
rect 21085 40987 21143 40993
rect 21085 40953 21097 40987
rect 21131 40984 21143 40987
rect 21453 40987 21511 40993
rect 21453 40984 21465 40987
rect 21131 40956 21465 40984
rect 21131 40953 21143 40956
rect 21085 40947 21143 40953
rect 21453 40953 21465 40956
rect 21499 40984 21511 40987
rect 21729 40987 21787 40993
rect 21729 40984 21741 40987
rect 21499 40956 21741 40984
rect 21499 40953 21511 40956
rect 21453 40947 21511 40953
rect 21729 40953 21741 40956
rect 21775 40984 21787 40987
rect 21910 40984 21916 40996
rect 21775 40956 21916 40984
rect 21775 40953 21787 40956
rect 21729 40947 21787 40953
rect 21910 40944 21916 40956
rect 21968 40944 21974 40996
rect 22094 40944 22100 40996
rect 22152 40984 22158 40996
rect 22281 40987 22339 40993
rect 22281 40984 22293 40987
rect 22152 40956 22293 40984
rect 22152 40944 22158 40956
rect 22281 40953 22293 40956
rect 22327 40953 22339 40987
rect 22281 40947 22339 40953
rect 14366 40876 14372 40928
rect 14424 40916 14430 40928
rect 14507 40919 14565 40925
rect 14507 40916 14519 40919
rect 14424 40888 14519 40916
rect 14424 40876 14430 40888
rect 14507 40885 14519 40888
rect 14553 40885 14565 40919
rect 16482 40916 16488 40928
rect 16443 40888 16488 40916
rect 14507 40879 14565 40885
rect 16482 40876 16488 40888
rect 16540 40876 16546 40928
rect 18782 40916 18788 40928
rect 18743 40888 18788 40916
rect 18782 40876 18788 40888
rect 18840 40876 18846 40928
rect 23014 40876 23020 40928
rect 23072 40916 23078 40928
rect 23385 40919 23443 40925
rect 23385 40916 23397 40919
rect 23072 40888 23397 40916
rect 23072 40876 23078 40888
rect 23385 40885 23397 40888
rect 23431 40916 23443 40919
rect 23584 40916 23612 41015
rect 30374 41012 30380 41024
rect 30432 41052 30438 41064
rect 30576 41052 30604 41083
rect 35526 41080 35532 41092
rect 35584 41080 35590 41132
rect 30432 41024 30604 41052
rect 31272 41055 31330 41061
rect 30432 41012 30438 41024
rect 31272 41021 31284 41055
rect 31318 41021 31330 41055
rect 31272 41015 31330 41021
rect 31573 41055 31631 41061
rect 31573 41021 31585 41055
rect 31619 41052 31631 41055
rect 32252 41055 32310 41061
rect 32252 41052 32264 41055
rect 31619 41024 32264 41052
rect 31619 41021 31631 41024
rect 31573 41015 31631 41021
rect 32252 41021 32264 41024
rect 32298 41052 32310 41055
rect 32298 41021 32327 41052
rect 32252 41015 32327 41021
rect 24765 40987 24823 40993
rect 24765 40953 24777 40987
rect 24811 40984 24823 40987
rect 25038 40984 25044 40996
rect 24811 40956 25044 40984
rect 24811 40953 24823 40956
rect 24765 40947 24823 40953
rect 25038 40944 25044 40956
rect 25096 40944 25102 40996
rect 25958 40984 25964 40996
rect 25871 40956 25964 40984
rect 25958 40944 25964 40956
rect 26016 40984 26022 40996
rect 31287 40984 31315 41015
rect 31662 40984 31668 40996
rect 26016 40956 30236 40984
rect 31287 40956 31668 40984
rect 26016 40944 26022 40956
rect 30208 40928 30236 40956
rect 31662 40944 31668 40956
rect 31720 40944 31726 40996
rect 32299 40984 32327 41015
rect 32858 41012 32864 41064
rect 32916 41052 32922 41064
rect 33296 41055 33354 41061
rect 33296 41052 33308 41055
rect 32916 41024 33308 41052
rect 32916 41012 32922 41024
rect 33296 41021 33308 41024
rect 33342 41052 33354 41055
rect 33689 41055 33747 41061
rect 33689 41052 33701 41055
rect 33342 41024 33701 41052
rect 33342 41021 33354 41024
rect 33296 41015 33354 41021
rect 33689 41021 33701 41024
rect 33735 41021 33747 41055
rect 33689 41015 33747 41021
rect 33042 40984 33048 40996
rect 32299 40956 33048 40984
rect 33042 40944 33048 40956
rect 33100 40944 33106 40996
rect 24302 40916 24308 40928
rect 23431 40888 23612 40916
rect 24263 40888 24308 40916
rect 23431 40885 23443 40888
rect 23385 40879 23443 40885
rect 24302 40876 24308 40888
rect 24360 40876 24366 40928
rect 26743 40919 26801 40925
rect 26743 40885 26755 40919
rect 26789 40916 26801 40919
rect 26970 40916 26976 40928
rect 26789 40888 26976 40916
rect 26789 40885 26801 40888
rect 26743 40879 26801 40885
rect 26970 40876 26976 40888
rect 27028 40876 27034 40928
rect 29914 40916 29920 40928
rect 29875 40888 29920 40916
rect 29914 40876 29920 40888
rect 29972 40876 29978 40928
rect 30190 40916 30196 40928
rect 30151 40888 30196 40916
rect 30190 40876 30196 40888
rect 30248 40876 30254 40928
rect 31343 40919 31401 40925
rect 31343 40885 31355 40919
rect 31389 40916 31401 40919
rect 31478 40916 31484 40928
rect 31389 40888 31484 40916
rect 31389 40885 31401 40888
rect 31343 40879 31401 40885
rect 31478 40876 31484 40888
rect 31536 40876 31542 40928
rect 32355 40919 32413 40925
rect 32355 40885 32367 40919
rect 32401 40916 32413 40919
rect 32582 40916 32588 40928
rect 32401 40888 32588 40916
rect 32401 40885 32413 40888
rect 32355 40879 32413 40885
rect 32582 40876 32588 40888
rect 32640 40876 32646 40928
rect 33367 40919 33425 40925
rect 33367 40885 33379 40919
rect 33413 40916 33425 40919
rect 33778 40916 33784 40928
rect 33413 40888 33784 40916
rect 33413 40885 33425 40888
rect 33367 40879 33425 40885
rect 33778 40876 33784 40888
rect 33836 40876 33842 40928
rect 1104 40826 48852 40848
rect 1104 40774 19606 40826
rect 19658 40774 19670 40826
rect 19722 40774 19734 40826
rect 19786 40774 19798 40826
rect 19850 40774 48852 40826
rect 1104 40752 48852 40774
rect 24578 40712 24584 40724
rect 24539 40684 24584 40712
rect 24578 40672 24584 40684
rect 24636 40672 24642 40724
rect 26878 40672 26884 40724
rect 26936 40712 26942 40724
rect 26936 40684 27016 40712
rect 26936 40672 26942 40684
rect 16669 40647 16727 40653
rect 16669 40613 16681 40647
rect 16715 40644 16727 40647
rect 16758 40644 16764 40656
rect 16715 40616 16764 40644
rect 16715 40613 16727 40616
rect 16669 40607 16727 40613
rect 16758 40604 16764 40616
rect 16816 40604 16822 40656
rect 19426 40644 19432 40656
rect 19387 40616 19432 40644
rect 19426 40604 19432 40616
rect 19484 40604 19490 40656
rect 21726 40644 21732 40656
rect 21687 40616 21732 40644
rect 21726 40604 21732 40616
rect 21784 40604 21790 40656
rect 21821 40647 21879 40653
rect 21821 40613 21833 40647
rect 21867 40644 21879 40647
rect 22002 40644 22008 40656
rect 21867 40616 22008 40644
rect 21867 40613 21879 40616
rect 21821 40607 21879 40613
rect 22002 40604 22008 40616
rect 22060 40604 22066 40656
rect 25038 40644 25044 40656
rect 24999 40616 25044 40644
rect 25038 40604 25044 40616
rect 25096 40604 25102 40656
rect 26988 40653 27016 40684
rect 26973 40647 27031 40653
rect 26973 40613 26985 40647
rect 27019 40613 27031 40647
rect 26973 40607 27031 40613
rect 27062 40604 27068 40656
rect 27120 40644 27126 40656
rect 30190 40644 30196 40656
rect 27120 40616 27165 40644
rect 30151 40616 30196 40644
rect 27120 40604 27126 40616
rect 30190 40604 30196 40616
rect 30248 40604 30254 40656
rect 32585 40647 32643 40653
rect 32585 40613 32597 40647
rect 32631 40644 32643 40647
rect 32674 40644 32680 40656
rect 32631 40616 32680 40644
rect 32631 40613 32643 40616
rect 32585 40607 32643 40613
rect 32674 40604 32680 40616
rect 32732 40604 32738 40656
rect 17862 40536 17868 40588
rect 17920 40576 17926 40588
rect 18116 40579 18174 40585
rect 18116 40576 18128 40579
rect 17920 40548 18128 40576
rect 17920 40536 17926 40548
rect 18116 40545 18128 40548
rect 18162 40576 18174 40579
rect 19058 40576 19064 40588
rect 18162 40548 19064 40576
rect 18162 40545 18174 40548
rect 18116 40539 18174 40545
rect 19058 40536 19064 40548
rect 19116 40536 19122 40588
rect 23198 40576 23204 40588
rect 23159 40548 23204 40576
rect 23198 40536 23204 40548
rect 23256 40536 23262 40588
rect 33962 40576 33968 40588
rect 33923 40548 33968 40576
rect 33962 40536 33968 40548
rect 34020 40536 34026 40588
rect 35044 40579 35102 40585
rect 35044 40545 35056 40579
rect 35090 40576 35102 40579
rect 35250 40576 35256 40588
rect 35090 40548 35256 40576
rect 35090 40545 35102 40548
rect 35044 40539 35102 40545
rect 35250 40536 35256 40548
rect 35308 40536 35314 40588
rect 38286 40576 38292 40588
rect 38247 40548 38292 40576
rect 38286 40536 38292 40548
rect 38344 40536 38350 40588
rect 14093 40511 14151 40517
rect 14093 40477 14105 40511
rect 14139 40508 14151 40511
rect 14182 40508 14188 40520
rect 14139 40480 14188 40508
rect 14139 40477 14151 40480
rect 14093 40471 14151 40477
rect 14182 40468 14188 40480
rect 14240 40468 14246 40520
rect 16577 40511 16635 40517
rect 16577 40508 16589 40511
rect 16316 40480 16589 40508
rect 14323 40375 14381 40381
rect 14323 40341 14335 40375
rect 14369 40372 14381 40375
rect 14642 40372 14648 40384
rect 14369 40344 14648 40372
rect 14369 40341 14381 40344
rect 14323 40335 14381 40341
rect 14642 40332 14648 40344
rect 14700 40332 14706 40384
rect 16206 40332 16212 40384
rect 16264 40372 16270 40384
rect 16316 40381 16344 40480
rect 16577 40477 16589 40480
rect 16623 40477 16635 40511
rect 17218 40508 17224 40520
rect 17179 40480 17224 40508
rect 16577 40471 16635 40477
rect 17218 40468 17224 40480
rect 17276 40468 17282 40520
rect 19150 40468 19156 40520
rect 19208 40508 19214 40520
rect 19337 40511 19395 40517
rect 19337 40508 19349 40511
rect 19208 40480 19349 40508
rect 19208 40468 19214 40480
rect 19337 40477 19349 40480
rect 19383 40477 19395 40511
rect 19337 40471 19395 40477
rect 19981 40511 20039 40517
rect 19981 40477 19993 40511
rect 20027 40508 20039 40511
rect 20530 40508 20536 40520
rect 20027 40480 20536 40508
rect 20027 40477 20039 40480
rect 19981 40471 20039 40477
rect 20530 40468 20536 40480
rect 20588 40508 20594 40520
rect 22005 40511 22063 40517
rect 22005 40508 22017 40511
rect 20588 40480 22017 40508
rect 20588 40468 20594 40480
rect 22005 40477 22017 40480
rect 22051 40508 22063 40511
rect 22094 40508 22100 40520
rect 22051 40480 22100 40508
rect 22051 40477 22063 40480
rect 22005 40471 22063 40477
rect 22094 40468 22100 40480
rect 22152 40468 22158 40520
rect 24946 40508 24952 40520
rect 24907 40480 24952 40508
rect 24946 40468 24952 40480
rect 25004 40468 25010 40520
rect 25593 40511 25651 40517
rect 25593 40477 25605 40511
rect 25639 40508 25651 40511
rect 26142 40508 26148 40520
rect 25639 40480 26148 40508
rect 25639 40477 25651 40480
rect 25593 40471 25651 40477
rect 26142 40468 26148 40480
rect 26200 40508 26206 40520
rect 27249 40511 27307 40517
rect 27249 40508 27261 40511
rect 26200 40480 27261 40508
rect 26200 40468 26206 40480
rect 27249 40477 27261 40480
rect 27295 40477 27307 40511
rect 27249 40471 27307 40477
rect 28905 40511 28963 40517
rect 28905 40477 28917 40511
rect 28951 40508 28963 40511
rect 29086 40508 29092 40520
rect 28951 40480 29092 40508
rect 28951 40477 28963 40480
rect 28905 40471 28963 40477
rect 24302 40400 24308 40452
rect 24360 40440 24366 40452
rect 28920 40440 28948 40471
rect 29086 40468 29092 40480
rect 29144 40468 29150 40520
rect 29914 40468 29920 40520
rect 29972 40508 29978 40520
rect 30101 40511 30159 40517
rect 30101 40508 30113 40511
rect 29972 40480 30113 40508
rect 29972 40468 29978 40480
rect 30101 40477 30113 40480
rect 30147 40508 30159 40511
rect 31018 40508 31024 40520
rect 30147 40480 31024 40508
rect 30147 40477 30159 40480
rect 30101 40471 30159 40477
rect 31018 40468 31024 40480
rect 31076 40468 31082 40520
rect 32490 40508 32496 40520
rect 32451 40480 32496 40508
rect 32490 40468 32496 40480
rect 32548 40468 32554 40520
rect 32769 40511 32827 40517
rect 32769 40477 32781 40511
rect 32815 40477 32827 40511
rect 32769 40471 32827 40477
rect 24360 40412 28948 40440
rect 30653 40443 30711 40449
rect 24360 40400 24366 40412
rect 30653 40409 30665 40443
rect 30699 40440 30711 40443
rect 32398 40440 32404 40452
rect 30699 40412 32404 40440
rect 30699 40409 30711 40412
rect 30653 40403 30711 40409
rect 32398 40400 32404 40412
rect 32456 40440 32462 40452
rect 32784 40440 32812 40471
rect 38746 40468 38752 40520
rect 38804 40508 38810 40520
rect 39117 40511 39175 40517
rect 39117 40508 39129 40511
rect 38804 40480 39129 40508
rect 38804 40468 38810 40480
rect 39117 40477 39129 40480
rect 39163 40477 39175 40511
rect 39117 40471 39175 40477
rect 32456 40412 32812 40440
rect 32456 40400 32462 40412
rect 33226 40400 33232 40452
rect 33284 40440 33290 40452
rect 35115 40443 35173 40449
rect 35115 40440 35127 40443
rect 33284 40412 35127 40440
rect 33284 40400 33290 40412
rect 35115 40409 35127 40412
rect 35161 40409 35173 40443
rect 35115 40403 35173 40409
rect 16301 40375 16359 40381
rect 16301 40372 16313 40375
rect 16264 40344 16313 40372
rect 16264 40332 16270 40344
rect 16301 40341 16313 40344
rect 16347 40341 16359 40375
rect 16301 40335 16359 40341
rect 16666 40332 16672 40384
rect 16724 40372 16730 40384
rect 18187 40375 18245 40381
rect 18187 40372 18199 40375
rect 16724 40344 18199 40372
rect 16724 40332 16730 40344
rect 18187 40341 18199 40344
rect 18233 40341 18245 40375
rect 18187 40335 18245 40341
rect 22738 40332 22744 40384
rect 22796 40372 22802 40384
rect 23339 40375 23397 40381
rect 23339 40372 23351 40375
rect 22796 40344 23351 40372
rect 22796 40332 22802 40344
rect 23339 40341 23351 40344
rect 23385 40341 23397 40375
rect 23339 40335 23397 40341
rect 29135 40375 29193 40381
rect 29135 40341 29147 40375
rect 29181 40372 29193 40375
rect 29914 40372 29920 40384
rect 29181 40344 29920 40372
rect 29181 40341 29193 40344
rect 29135 40335 29193 40341
rect 29914 40332 29920 40344
rect 29972 40332 29978 40384
rect 32950 40332 32956 40384
rect 33008 40372 33014 40384
rect 34103 40375 34161 40381
rect 34103 40372 34115 40375
rect 33008 40344 34115 40372
rect 33008 40332 33014 40344
rect 34103 40341 34115 40344
rect 34149 40341 34161 40375
rect 34103 40335 34161 40341
rect 37093 40375 37151 40381
rect 37093 40341 37105 40375
rect 37139 40372 37151 40375
rect 37458 40372 37464 40384
rect 37139 40344 37464 40372
rect 37139 40341 37151 40344
rect 37093 40335 37151 40341
rect 37458 40332 37464 40344
rect 37516 40332 37522 40384
rect 38427 40375 38485 40381
rect 38427 40341 38439 40375
rect 38473 40372 38485 40375
rect 38562 40372 38568 40384
rect 38473 40344 38568 40372
rect 38473 40341 38485 40344
rect 38427 40335 38485 40341
rect 38562 40332 38568 40344
rect 38620 40332 38626 40384
rect 38838 40372 38844 40384
rect 38799 40344 38844 40372
rect 38838 40332 38844 40344
rect 38896 40332 38902 40384
rect 1104 40282 48852 40304
rect 1104 40230 4246 40282
rect 4298 40230 4310 40282
rect 4362 40230 4374 40282
rect 4426 40230 4438 40282
rect 4490 40230 34966 40282
rect 35018 40230 35030 40282
rect 35082 40230 35094 40282
rect 35146 40230 35158 40282
rect 35210 40230 48852 40282
rect 1104 40208 48852 40230
rect 14182 40168 14188 40180
rect 14143 40140 14188 40168
rect 14182 40128 14188 40140
rect 14240 40128 14246 40180
rect 17862 40168 17868 40180
rect 17823 40140 17868 40168
rect 17862 40128 17868 40140
rect 17920 40128 17926 40180
rect 19153 40171 19211 40177
rect 19153 40137 19165 40171
rect 19199 40168 19211 40171
rect 19426 40168 19432 40180
rect 19199 40140 19432 40168
rect 19199 40137 19211 40140
rect 19153 40131 19211 40137
rect 19426 40128 19432 40140
rect 19484 40128 19490 40180
rect 20809 40171 20867 40177
rect 20809 40137 20821 40171
rect 20855 40168 20867 40171
rect 21726 40168 21732 40180
rect 20855 40140 21732 40168
rect 20855 40137 20867 40140
rect 20809 40131 20867 40137
rect 21726 40128 21732 40140
rect 21784 40128 21790 40180
rect 22738 40168 22744 40180
rect 22699 40140 22744 40168
rect 22738 40128 22744 40140
rect 22796 40128 22802 40180
rect 24489 40171 24547 40177
rect 24489 40137 24501 40171
rect 24535 40168 24547 40171
rect 25038 40168 25044 40180
rect 24535 40140 25044 40168
rect 24535 40137 24547 40140
rect 24489 40131 24547 40137
rect 25038 40128 25044 40140
rect 25096 40168 25102 40180
rect 25593 40171 25651 40177
rect 25593 40168 25605 40171
rect 25096 40140 25605 40168
rect 25096 40128 25102 40140
rect 25593 40137 25605 40140
rect 25639 40137 25651 40171
rect 25593 40131 25651 40137
rect 26878 40128 26884 40180
rect 26936 40168 26942 40180
rect 27893 40171 27951 40177
rect 27893 40168 27905 40171
rect 26936 40140 27905 40168
rect 26936 40128 26942 40140
rect 27893 40137 27905 40140
rect 27939 40137 27951 40171
rect 31018 40168 31024 40180
rect 30979 40140 31024 40168
rect 27893 40131 27951 40137
rect 31018 40128 31024 40140
rect 31076 40128 31082 40180
rect 33042 40128 33048 40180
rect 33100 40168 33106 40180
rect 35161 40171 35219 40177
rect 33100 40140 35112 40168
rect 33100 40128 33106 40140
rect 16022 40060 16028 40112
rect 16080 40100 16086 40112
rect 17037 40103 17095 40109
rect 17037 40100 17049 40103
rect 16080 40072 17049 40100
rect 16080 40060 16086 40072
rect 17037 40069 17049 40072
rect 17083 40069 17095 40103
rect 22278 40100 22284 40112
rect 22239 40072 22284 40100
rect 17037 40063 17095 40069
rect 22278 40060 22284 40072
rect 22336 40060 22342 40112
rect 13354 40032 13360 40044
rect 13315 40004 13360 40032
rect 13354 39992 13360 40004
rect 13412 39992 13418 40044
rect 14642 40032 14648 40044
rect 14603 40004 14648 40032
rect 14642 39992 14648 40004
rect 14700 39992 14706 40044
rect 16485 40035 16543 40041
rect 16485 40001 16497 40035
rect 16531 40032 16543 40035
rect 16574 40032 16580 40044
rect 16531 40004 16580 40032
rect 16531 40001 16543 40004
rect 16485 39995 16543 40001
rect 16574 39992 16580 40004
rect 16632 40032 16638 40044
rect 17405 40035 17463 40041
rect 17405 40032 17417 40035
rect 16632 40004 17417 40032
rect 16632 39992 16638 40004
rect 17405 40001 17417 40004
rect 17451 40001 17463 40035
rect 17405 39995 17463 40001
rect 18371 40035 18429 40041
rect 18371 40001 18383 40035
rect 18417 40032 18429 40035
rect 19337 40035 19395 40041
rect 19337 40032 19349 40035
rect 18417 40004 19349 40032
rect 18417 40001 18429 40004
rect 18371 39995 18429 40001
rect 19337 40001 19349 40004
rect 19383 40032 19395 40035
rect 20257 40035 20315 40041
rect 20257 40032 20269 40035
rect 19383 40004 20269 40032
rect 19383 40001 19395 40004
rect 19337 39995 19395 40001
rect 20257 40001 20269 40004
rect 20303 40001 20315 40035
rect 20257 39995 20315 40001
rect 21729 40035 21787 40041
rect 21729 40001 21741 40035
rect 21775 40032 21787 40035
rect 22756 40032 22784 40128
rect 24578 40060 24584 40112
rect 24636 40100 24642 40112
rect 25225 40103 25283 40109
rect 24636 40072 24716 40100
rect 24636 40060 24642 40072
rect 23198 40032 23204 40044
rect 21775 40004 22784 40032
rect 23159 40004 23204 40032
rect 21775 40001 21787 40004
rect 21729 39995 21787 40001
rect 23198 39992 23204 40004
rect 23256 39992 23262 40044
rect 24688 40041 24716 40072
rect 25225 40069 25237 40103
rect 25271 40100 25283 40103
rect 27798 40100 27804 40112
rect 25271 40072 27804 40100
rect 25271 40069 25283 40072
rect 25225 40063 25283 40069
rect 27798 40060 27804 40072
rect 27856 40060 27862 40112
rect 32214 40060 32220 40112
rect 32272 40100 32278 40112
rect 33962 40100 33968 40112
rect 32272 40072 33968 40100
rect 32272 40060 32278 40072
rect 33962 40060 33968 40072
rect 34020 40060 34026 40112
rect 35084 40100 35112 40140
rect 35161 40137 35173 40171
rect 35207 40168 35219 40171
rect 35250 40168 35256 40180
rect 35207 40140 35256 40168
rect 35207 40137 35219 40140
rect 35161 40131 35219 40137
rect 35250 40128 35256 40140
rect 35308 40168 35314 40180
rect 39666 40168 39672 40180
rect 35308 40140 39672 40168
rect 35308 40128 35314 40140
rect 39666 40128 39672 40140
rect 39724 40128 39730 40180
rect 38286 40100 38292 40112
rect 35084 40072 38292 40100
rect 38286 40060 38292 40072
rect 38344 40100 38350 40112
rect 39206 40100 39212 40112
rect 38344 40072 39212 40100
rect 38344 40060 38350 40072
rect 39206 40060 39212 40072
rect 39264 40060 39270 40112
rect 24673 40035 24731 40041
rect 24673 40001 24685 40035
rect 24719 40001 24731 40035
rect 24673 39995 24731 40001
rect 26053 40035 26111 40041
rect 26053 40001 26065 40035
rect 26099 40032 26111 40035
rect 26970 40032 26976 40044
rect 26099 40004 26976 40032
rect 26099 40001 26111 40004
rect 26053 39995 26111 40001
rect 26970 39992 26976 40004
rect 27028 39992 27034 40044
rect 27246 40032 27252 40044
rect 27207 40004 27252 40032
rect 27246 39992 27252 40004
rect 27304 39992 27310 40044
rect 30098 40032 30104 40044
rect 30059 40004 30104 40032
rect 30098 39992 30104 40004
rect 30156 39992 30162 40044
rect 31665 40035 31723 40041
rect 31665 40001 31677 40035
rect 31711 40032 31723 40035
rect 32582 40032 32588 40044
rect 31711 40004 32588 40032
rect 31711 40001 31723 40004
rect 31665 39995 31723 40001
rect 32582 39992 32588 40004
rect 32640 39992 32646 40044
rect 12986 39973 12992 39976
rect 12964 39967 12992 39973
rect 12964 39964 12976 39967
rect 12899 39936 12976 39964
rect 12964 39933 12976 39936
rect 13044 39964 13050 39976
rect 13372 39964 13400 39992
rect 13044 39936 13400 39964
rect 18284 39967 18342 39973
rect 12964 39927 12992 39933
rect 12986 39924 12992 39927
rect 13044 39924 13050 39936
rect 18284 39933 18296 39967
rect 18330 39964 18342 39967
rect 18330 39936 18828 39964
rect 18330 39933 18342 39936
rect 18284 39927 18342 39933
rect 14734 39896 14740 39908
rect 14695 39868 14740 39896
rect 14734 39856 14740 39868
rect 14792 39856 14798 39908
rect 15286 39896 15292 39908
rect 15247 39868 15292 39896
rect 15286 39856 15292 39868
rect 15344 39856 15350 39908
rect 15933 39899 15991 39905
rect 15933 39865 15945 39899
rect 15979 39896 15991 39899
rect 16301 39899 16359 39905
rect 16301 39896 16313 39899
rect 15979 39868 16313 39896
rect 15979 39865 15991 39868
rect 15933 39859 15991 39865
rect 16301 39865 16313 39868
rect 16347 39896 16359 39899
rect 16577 39899 16635 39905
rect 16577 39896 16589 39899
rect 16347 39868 16589 39896
rect 16347 39865 16359 39868
rect 16301 39859 16359 39865
rect 16577 39865 16589 39868
rect 16623 39896 16635 39899
rect 16758 39896 16764 39908
rect 16623 39868 16764 39896
rect 16623 39865 16635 39868
rect 16577 39859 16635 39865
rect 16758 39856 16764 39868
rect 16816 39856 16822 39908
rect 17494 39896 17500 39908
rect 16868 39868 17500 39896
rect 13035 39831 13093 39837
rect 13035 39797 13047 39831
rect 13081 39828 13093 39831
rect 13170 39828 13176 39840
rect 13081 39800 13176 39828
rect 13081 39797 13093 39800
rect 13035 39791 13093 39797
rect 13170 39788 13176 39800
rect 13228 39788 13234 39840
rect 16390 39788 16396 39840
rect 16448 39828 16454 39840
rect 16868 39828 16896 39868
rect 17494 39856 17500 39868
rect 17552 39896 17558 39908
rect 18299 39896 18327 39927
rect 17552 39868 18327 39896
rect 17552 39856 17558 39868
rect 18800 39840 18828 39936
rect 35526 39924 35532 39976
rect 35584 39964 35590 39976
rect 35840 39967 35898 39973
rect 35840 39964 35852 39967
rect 35584 39936 35852 39964
rect 35584 39924 35590 39936
rect 35840 39933 35852 39936
rect 35886 39964 35898 39967
rect 36265 39967 36323 39973
rect 36265 39964 36277 39967
rect 35886 39936 36277 39964
rect 35886 39933 35898 39936
rect 35840 39927 35898 39933
rect 36265 39933 36277 39936
rect 36311 39933 36323 39967
rect 36265 39927 36323 39933
rect 37001 39967 37059 39973
rect 37001 39933 37013 39967
rect 37047 39933 37059 39967
rect 37458 39964 37464 39976
rect 37419 39936 37464 39964
rect 37001 39927 37059 39933
rect 19426 39896 19432 39908
rect 19387 39868 19432 39896
rect 19426 39856 19432 39868
rect 19484 39856 19490 39908
rect 19978 39896 19984 39908
rect 19939 39868 19984 39896
rect 19978 39856 19984 39868
rect 20036 39856 20042 39908
rect 21821 39899 21879 39905
rect 21821 39865 21833 39899
rect 21867 39865 21879 39899
rect 21821 39859 21879 39865
rect 24765 39899 24823 39905
rect 24765 39865 24777 39899
rect 24811 39896 24823 39899
rect 25038 39896 25044 39908
rect 24811 39868 25044 39896
rect 24811 39865 24823 39868
rect 24765 39859 24823 39865
rect 18782 39828 18788 39840
rect 16448 39800 16896 39828
rect 18743 39800 18788 39828
rect 16448 39788 16454 39800
rect 18782 39788 18788 39800
rect 18840 39788 18846 39840
rect 21177 39831 21235 39837
rect 21177 39797 21189 39831
rect 21223 39828 21235 39831
rect 21545 39831 21603 39837
rect 21545 39828 21557 39831
rect 21223 39800 21557 39828
rect 21223 39797 21235 39800
rect 21177 39791 21235 39797
rect 21545 39797 21557 39800
rect 21591 39828 21603 39831
rect 21836 39828 21864 39859
rect 25038 39856 25044 39868
rect 25096 39856 25102 39908
rect 27062 39905 27068 39908
rect 26421 39899 26479 39905
rect 26421 39865 26433 39899
rect 26467 39896 26479 39899
rect 26789 39899 26847 39905
rect 26789 39896 26801 39899
rect 26467 39868 26801 39896
rect 26467 39865 26479 39868
rect 26421 39859 26479 39865
rect 26789 39865 26801 39868
rect 26835 39896 26847 39899
rect 27042 39899 27068 39905
rect 27042 39896 27054 39899
rect 26835 39868 27054 39896
rect 26835 39865 26847 39868
rect 26789 39859 26847 39865
rect 27042 39865 27054 39868
rect 27042 39859 27068 39865
rect 27062 39856 27068 39859
rect 27120 39856 27126 39908
rect 30190 39896 30196 39908
rect 30024 39868 30196 39896
rect 30024 39840 30052 39868
rect 30190 39856 30196 39868
rect 30248 39856 30254 39908
rect 30745 39899 30803 39905
rect 30745 39865 30757 39899
rect 30791 39896 30803 39899
rect 30791 39868 32489 39896
rect 30791 39865 30803 39868
rect 30745 39859 30803 39865
rect 22002 39828 22008 39840
rect 21591 39800 22008 39828
rect 21591 39797 21603 39800
rect 21545 39791 21603 39797
rect 22002 39788 22008 39800
rect 22060 39788 22066 39840
rect 24121 39831 24179 39837
rect 24121 39797 24133 39831
rect 24167 39828 24179 39831
rect 24946 39828 24952 39840
rect 24167 39800 24952 39828
rect 24167 39797 24179 39800
rect 24121 39791 24179 39797
rect 24946 39788 24952 39800
rect 25004 39788 25010 39840
rect 29086 39828 29092 39840
rect 29047 39800 29092 39828
rect 29086 39788 29092 39800
rect 29144 39788 29150 39840
rect 29549 39831 29607 39837
rect 29549 39797 29561 39831
rect 29595 39828 29607 39831
rect 29917 39831 29975 39837
rect 29917 39828 29929 39831
rect 29595 39800 29929 39828
rect 29595 39797 29607 39800
rect 29549 39791 29607 39797
rect 29917 39797 29929 39800
rect 29963 39828 29975 39831
rect 30006 39828 30012 39840
rect 29963 39800 30012 39828
rect 29963 39797 29975 39800
rect 29917 39791 29975 39797
rect 30006 39788 30012 39800
rect 30064 39788 30070 39840
rect 31754 39788 31760 39840
rect 31812 39828 31818 39840
rect 31941 39831 31999 39837
rect 31941 39828 31953 39831
rect 31812 39800 31953 39828
rect 31812 39788 31818 39800
rect 31941 39797 31953 39800
rect 31987 39828 31999 39831
rect 32309 39831 32367 39837
rect 32309 39828 32321 39831
rect 31987 39800 32321 39828
rect 31987 39797 31999 39800
rect 31941 39791 31999 39797
rect 32309 39797 32321 39800
rect 32355 39797 32367 39831
rect 32461 39828 32489 39868
rect 32582 39856 32588 39908
rect 32640 39896 32646 39908
rect 32677 39899 32735 39905
rect 32677 39896 32689 39899
rect 32640 39868 32689 39896
rect 32640 39856 32646 39868
rect 32677 39865 32689 39868
rect 32723 39865 32735 39899
rect 33229 39899 33287 39905
rect 33229 39896 33241 39899
rect 32677 39859 32735 39865
rect 33152 39868 33241 39896
rect 33152 39840 33180 39868
rect 33229 39865 33241 39868
rect 33275 39865 33287 39899
rect 33229 39859 33287 39865
rect 35710 39856 35716 39908
rect 35768 39896 35774 39908
rect 36817 39899 36875 39905
rect 36817 39896 36829 39899
rect 35768 39868 36829 39896
rect 35768 39856 35774 39868
rect 36817 39865 36829 39868
rect 36863 39896 36875 39899
rect 37016 39896 37044 39927
rect 37458 39924 37464 39936
rect 37516 39924 37522 39976
rect 37734 39896 37740 39908
rect 36863 39868 37044 39896
rect 37695 39868 37740 39896
rect 36863 39865 36875 39868
rect 36817 39859 36875 39865
rect 37734 39856 37740 39868
rect 37792 39856 37798 39908
rect 38746 39896 38752 39908
rect 38707 39868 38752 39896
rect 38746 39856 38752 39868
rect 38804 39856 38810 39908
rect 38838 39856 38844 39908
rect 38896 39896 38902 39908
rect 39393 39899 39451 39905
rect 38896 39868 38941 39896
rect 38896 39856 38902 39868
rect 39393 39865 39405 39899
rect 39439 39896 39451 39899
rect 42150 39896 42156 39908
rect 39439 39868 42156 39896
rect 39439 39865 39451 39868
rect 39393 39859 39451 39865
rect 42150 39856 42156 39868
rect 42208 39856 42214 39908
rect 33134 39828 33140 39840
rect 32461 39800 33140 39828
rect 32309 39791 32367 39797
rect 33134 39788 33140 39800
rect 33192 39788 33198 39840
rect 35943 39831 36001 39837
rect 35943 39797 35955 39831
rect 35989 39828 36001 39831
rect 36078 39828 36084 39840
rect 35989 39800 36084 39828
rect 35989 39797 36001 39800
rect 35943 39791 36001 39797
rect 36078 39788 36084 39800
rect 36136 39788 36142 39840
rect 1104 39738 48852 39760
rect 1104 39686 19606 39738
rect 19658 39686 19670 39738
rect 19722 39686 19734 39738
rect 19786 39686 19798 39738
rect 19850 39686 48852 39738
rect 1104 39664 48852 39686
rect 14645 39627 14703 39633
rect 14645 39624 14657 39627
rect 13786 39596 14657 39624
rect 13170 39516 13176 39568
rect 13228 39556 13234 39568
rect 13357 39559 13415 39565
rect 13357 39556 13369 39559
rect 13228 39528 13369 39556
rect 13228 39516 13234 39528
rect 13357 39525 13369 39528
rect 13403 39525 13415 39559
rect 13357 39519 13415 39525
rect 13449 39559 13507 39565
rect 13449 39525 13461 39559
rect 13495 39556 13507 39559
rect 13786 39556 13814 39596
rect 14645 39593 14657 39596
rect 14691 39624 14703 39627
rect 14734 39624 14740 39636
rect 14691 39596 14740 39624
rect 14691 39593 14703 39596
rect 14645 39587 14703 39593
rect 14734 39584 14740 39596
rect 14792 39584 14798 39636
rect 15703 39627 15761 39633
rect 15703 39593 15715 39627
rect 15749 39624 15761 39627
rect 16206 39624 16212 39636
rect 15749 39596 16212 39624
rect 15749 39593 15761 39596
rect 15703 39587 15761 39593
rect 16206 39584 16212 39596
rect 16264 39584 16270 39636
rect 16301 39627 16359 39633
rect 16301 39593 16313 39627
rect 16347 39624 16359 39627
rect 16482 39624 16488 39636
rect 16347 39596 16488 39624
rect 16347 39593 16359 39596
rect 16301 39587 16359 39593
rect 16482 39584 16488 39596
rect 16540 39584 16546 39636
rect 19426 39624 19432 39636
rect 19387 39596 19432 39624
rect 19426 39584 19432 39596
rect 19484 39624 19490 39636
rect 19705 39627 19763 39633
rect 19705 39624 19717 39627
rect 19484 39596 19717 39624
rect 19484 39584 19490 39596
rect 19705 39593 19717 39596
rect 19751 39593 19763 39627
rect 24302 39624 24308 39636
rect 24263 39596 24308 39624
rect 19705 39587 19763 39593
rect 24302 39584 24308 39596
rect 24360 39584 24366 39636
rect 24857 39627 24915 39633
rect 24857 39593 24869 39627
rect 24903 39624 24915 39627
rect 25038 39624 25044 39636
rect 24903 39596 25044 39624
rect 24903 39593 24915 39596
rect 24857 39587 24915 39593
rect 25038 39584 25044 39596
rect 25096 39584 25102 39636
rect 30098 39584 30104 39636
rect 30156 39624 30162 39636
rect 30377 39627 30435 39633
rect 30377 39624 30389 39627
rect 30156 39596 30389 39624
rect 30156 39584 30162 39596
rect 30377 39593 30389 39596
rect 30423 39593 30435 39627
rect 30377 39587 30435 39593
rect 31159 39627 31217 39633
rect 31159 39593 31171 39627
rect 31205 39624 31217 39627
rect 32490 39624 32496 39636
rect 31205 39596 32496 39624
rect 31205 39593 31217 39596
rect 31159 39587 31217 39593
rect 32490 39584 32496 39596
rect 32548 39584 32554 39636
rect 35989 39627 36047 39633
rect 35989 39593 36001 39627
rect 36035 39624 36047 39627
rect 36078 39624 36084 39636
rect 36035 39596 36084 39624
rect 36035 39593 36047 39596
rect 35989 39587 36047 39593
rect 36078 39584 36084 39596
rect 36136 39624 36142 39636
rect 36136 39596 36216 39624
rect 36136 39584 36142 39596
rect 13998 39556 14004 39568
rect 13495 39528 13814 39556
rect 13911 39528 14004 39556
rect 13495 39525 13507 39528
rect 13449 39519 13507 39525
rect 13998 39516 14004 39528
rect 14056 39556 14062 39568
rect 16022 39556 16028 39568
rect 14056 39528 16028 39556
rect 14056 39516 14062 39528
rect 16022 39516 16028 39528
rect 16080 39516 16086 39568
rect 16390 39516 16396 39568
rect 16448 39516 16454 39568
rect 16666 39556 16672 39568
rect 16627 39528 16672 39556
rect 16666 39516 16672 39528
rect 16724 39516 16730 39568
rect 16758 39516 16764 39568
rect 16816 39556 16822 39568
rect 16816 39528 16861 39556
rect 16816 39516 16822 39528
rect 18690 39516 18696 39568
rect 18748 39556 18754 39568
rect 18830 39559 18888 39565
rect 18830 39556 18842 39559
rect 18748 39528 18842 39556
rect 18748 39516 18754 39528
rect 18830 39525 18842 39528
rect 18876 39525 18888 39559
rect 18830 39519 18888 39525
rect 19150 39516 19156 39568
rect 19208 39556 19214 39568
rect 20073 39559 20131 39565
rect 20073 39556 20085 39559
rect 19208 39528 20085 39556
rect 19208 39516 19214 39528
rect 20073 39525 20085 39528
rect 20119 39525 20131 39559
rect 20073 39519 20131 39525
rect 21913 39559 21971 39565
rect 21913 39525 21925 39559
rect 21959 39556 21971 39559
rect 22002 39556 22008 39568
rect 21959 39528 22008 39556
rect 21959 39525 21971 39528
rect 21913 39519 21971 39525
rect 22002 39516 22008 39528
rect 22060 39516 22066 39568
rect 27062 39556 27068 39568
rect 27023 39528 27068 39556
rect 27062 39516 27068 39528
rect 27120 39516 27126 39568
rect 28994 39516 29000 39568
rect 29052 39556 29058 39568
rect 29502 39559 29560 39565
rect 29502 39556 29514 39559
rect 29052 39528 29514 39556
rect 29052 39516 29058 39528
rect 29502 39525 29514 39528
rect 29548 39525 29560 39559
rect 29502 39519 29560 39525
rect 32674 39516 32680 39568
rect 32732 39556 32738 39568
rect 36188 39565 36216 39596
rect 32953 39559 33011 39565
rect 32953 39556 32965 39559
rect 32732 39528 32965 39556
rect 32732 39516 32738 39528
rect 32953 39525 32965 39528
rect 32999 39525 33011 39559
rect 32953 39519 33011 39525
rect 36173 39559 36231 39565
rect 36173 39525 36185 39559
rect 36219 39525 36231 39559
rect 36173 39519 36231 39525
rect 36265 39559 36323 39565
rect 36265 39525 36277 39559
rect 36311 39556 36323 39559
rect 36446 39556 36452 39568
rect 36311 39528 36452 39556
rect 36311 39525 36323 39528
rect 36265 39519 36323 39525
rect 36446 39516 36452 39528
rect 36504 39516 36510 39568
rect 38562 39516 38568 39568
rect 38620 39556 38626 39568
rect 38749 39559 38807 39565
rect 38749 39556 38761 39559
rect 38620 39528 38761 39556
rect 38620 39516 38626 39528
rect 38749 39525 38761 39528
rect 38795 39525 38807 39559
rect 38749 39519 38807 39525
rect 38838 39516 38844 39568
rect 38896 39556 38902 39568
rect 38896 39528 38941 39556
rect 38896 39516 38902 39528
rect 11882 39448 11888 39500
rect 11940 39488 11946 39500
rect 15654 39497 15660 39500
rect 12288 39491 12346 39497
rect 12288 39488 12300 39491
rect 11940 39460 12300 39488
rect 11940 39448 11946 39460
rect 12288 39457 12300 39460
rect 12334 39457 12346 39491
rect 15632 39491 15660 39497
rect 15632 39488 15644 39491
rect 15567 39460 15644 39488
rect 12288 39451 12346 39457
rect 15632 39457 15644 39460
rect 15712 39488 15718 39500
rect 16408 39488 16436 39516
rect 15712 39460 16436 39488
rect 15632 39451 15660 39457
rect 15654 39448 15660 39451
rect 15712 39448 15718 39460
rect 30926 39448 30932 39500
rect 30984 39488 30990 39500
rect 31056 39491 31114 39497
rect 31056 39488 31068 39491
rect 30984 39460 31068 39488
rect 30984 39448 30990 39460
rect 31056 39457 31068 39460
rect 31102 39457 31114 39491
rect 31056 39451 31114 39457
rect 34333 39491 34391 39497
rect 34333 39457 34345 39491
rect 34379 39488 34391 39491
rect 34422 39488 34428 39500
rect 34379 39460 34428 39488
rect 34379 39457 34391 39460
rect 34333 39451 34391 39457
rect 34422 39448 34428 39460
rect 34480 39448 34486 39500
rect 40656 39491 40714 39497
rect 40656 39457 40668 39491
rect 40702 39488 40714 39491
rect 40770 39488 40776 39500
rect 40702 39460 40776 39488
rect 40702 39457 40714 39460
rect 40656 39451 40714 39457
rect 40770 39448 40776 39460
rect 40828 39448 40834 39500
rect 15286 39380 15292 39432
rect 15344 39420 15350 39432
rect 15930 39420 15936 39432
rect 15344 39392 15936 39420
rect 15344 39380 15350 39392
rect 15930 39380 15936 39392
rect 15988 39420 15994 39432
rect 16945 39423 17003 39429
rect 16945 39420 16957 39423
rect 15988 39392 16957 39420
rect 15988 39380 15994 39392
rect 16945 39389 16957 39392
rect 16991 39389 17003 39423
rect 18506 39420 18512 39432
rect 18467 39392 18512 39420
rect 16945 39383 17003 39389
rect 18506 39380 18512 39392
rect 18564 39380 18570 39432
rect 21818 39420 21824 39432
rect 21779 39392 21824 39420
rect 21818 39380 21824 39392
rect 21876 39380 21882 39432
rect 22097 39423 22155 39429
rect 22097 39389 22109 39423
rect 22143 39389 22155 39423
rect 23934 39420 23940 39432
rect 23895 39392 23940 39420
rect 22097 39383 22155 39389
rect 19426 39312 19432 39364
rect 19484 39352 19490 39364
rect 19978 39352 19984 39364
rect 19484 39324 19984 39352
rect 19484 39312 19490 39324
rect 19978 39312 19984 39324
rect 20036 39352 20042 39364
rect 22112 39352 22140 39383
rect 23934 39380 23940 39392
rect 23992 39380 23998 39432
rect 26970 39420 26976 39432
rect 26931 39392 26976 39420
rect 26970 39380 26976 39392
rect 27028 39380 27034 39432
rect 27617 39423 27675 39429
rect 27617 39389 27629 39423
rect 27663 39420 27675 39423
rect 27798 39420 27804 39432
rect 27663 39392 27804 39420
rect 27663 39389 27675 39392
rect 27617 39383 27675 39389
rect 27798 39380 27804 39392
rect 27856 39380 27862 39432
rect 29178 39420 29184 39432
rect 29139 39392 29184 39420
rect 29178 39380 29184 39392
rect 29236 39380 29242 39432
rect 32858 39420 32864 39432
rect 32819 39392 32864 39420
rect 32858 39380 32864 39392
rect 32916 39380 32922 39432
rect 33137 39423 33195 39429
rect 33137 39389 33149 39423
rect 33183 39389 33195 39423
rect 36814 39420 36820 39432
rect 36775 39392 36820 39420
rect 33137 39383 33195 39389
rect 22278 39352 22284 39364
rect 20036 39324 22284 39352
rect 20036 39312 20042 39324
rect 22278 39312 22284 39324
rect 22336 39312 22342 39364
rect 32398 39312 32404 39364
rect 32456 39352 32462 39364
rect 33152 39352 33180 39383
rect 36814 39380 36820 39392
rect 36872 39380 36878 39432
rect 39393 39423 39451 39429
rect 39393 39389 39405 39423
rect 39439 39420 39451 39423
rect 41414 39420 41420 39432
rect 39439 39392 41420 39420
rect 39439 39389 39451 39392
rect 39393 39383 39451 39389
rect 41414 39380 41420 39392
rect 41472 39380 41478 39432
rect 32456 39324 33180 39352
rect 32456 39312 32462 39324
rect 12391 39287 12449 39293
rect 12391 39253 12403 39287
rect 12437 39284 12449 39287
rect 13262 39284 13268 39296
rect 12437 39256 13268 39284
rect 12437 39253 12449 39256
rect 12391 39247 12449 39253
rect 13262 39244 13268 39256
rect 13320 39244 13326 39296
rect 23750 39284 23756 39296
rect 23711 39256 23756 39284
rect 23750 39244 23756 39256
rect 23808 39244 23814 39296
rect 25222 39284 25228 39296
rect 25183 39256 25228 39284
rect 25222 39244 25228 39256
rect 25280 39244 25286 39296
rect 30098 39284 30104 39296
rect 30059 39256 30104 39284
rect 30098 39244 30104 39256
rect 30156 39244 30162 39296
rect 30742 39244 30748 39296
rect 30800 39284 30806 39296
rect 30837 39287 30895 39293
rect 30837 39284 30849 39287
rect 30800 39256 30849 39284
rect 30800 39244 30806 39256
rect 30837 39253 30849 39256
rect 30883 39253 30895 39287
rect 30837 39247 30895 39253
rect 33042 39244 33048 39296
rect 33100 39284 33106 39296
rect 34471 39287 34529 39293
rect 34471 39284 34483 39287
rect 33100 39256 34483 39284
rect 33100 39244 33106 39256
rect 34471 39253 34483 39256
rect 34517 39253 34529 39287
rect 34471 39247 34529 39253
rect 40727 39287 40785 39293
rect 40727 39253 40739 39287
rect 40773 39284 40785 39287
rect 40954 39284 40960 39296
rect 40773 39256 40960 39284
rect 40773 39253 40785 39256
rect 40727 39247 40785 39253
rect 40954 39244 40960 39256
rect 41012 39244 41018 39296
rect 1104 39194 48852 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 34966 39194
rect 35018 39142 35030 39194
rect 35082 39142 35094 39194
rect 35146 39142 35158 39194
rect 35210 39142 48852 39194
rect 1104 39120 48852 39142
rect 13170 39040 13176 39092
rect 13228 39080 13234 39092
rect 14001 39083 14059 39089
rect 14001 39080 14013 39083
rect 13228 39052 14013 39080
rect 13228 39040 13234 39052
rect 14001 39049 14013 39052
rect 14047 39049 14059 39083
rect 14001 39043 14059 39049
rect 14461 39083 14519 39089
rect 14461 39049 14473 39083
rect 14507 39080 14519 39083
rect 14734 39080 14740 39092
rect 14507 39052 14740 39080
rect 14507 39049 14519 39052
rect 14461 39043 14519 39049
rect 14734 39040 14740 39052
rect 14792 39040 14798 39092
rect 15654 39080 15660 39092
rect 15615 39052 15660 39080
rect 15654 39040 15660 39052
rect 15712 39040 15718 39092
rect 16758 39040 16764 39092
rect 16816 39080 16822 39092
rect 17129 39083 17187 39089
rect 17129 39080 17141 39083
rect 16816 39052 17141 39080
rect 16816 39040 16822 39052
rect 17129 39049 17141 39052
rect 17175 39080 17187 39083
rect 17405 39083 17463 39089
rect 17405 39080 17417 39083
rect 17175 39052 17417 39080
rect 17175 39049 17187 39052
rect 17129 39043 17187 39049
rect 17405 39049 17417 39052
rect 17451 39049 17463 39083
rect 17405 39043 17463 39049
rect 18690 39040 18696 39092
rect 18748 39080 18754 39092
rect 20257 39083 20315 39089
rect 20257 39080 20269 39083
rect 18748 39052 20269 39080
rect 18748 39040 18754 39052
rect 20257 39049 20269 39052
rect 20303 39049 20315 39083
rect 20257 39043 20315 39049
rect 13556 38984 19196 39012
rect 13556 38944 13584 38984
rect 11072 38916 13584 38944
rect 10502 38836 10508 38888
rect 10560 38876 10566 38888
rect 11072 38885 11100 38916
rect 13722 38904 13728 38956
rect 13780 38944 13786 38956
rect 14366 38944 14372 38956
rect 13780 38916 14372 38944
rect 13780 38904 13786 38916
rect 14366 38904 14372 38916
rect 14424 38944 14430 38956
rect 14645 38947 14703 38953
rect 14645 38944 14657 38947
rect 14424 38916 14657 38944
rect 14424 38904 14430 38916
rect 14645 38913 14657 38916
rect 14691 38913 14703 38947
rect 14645 38907 14703 38913
rect 16209 38947 16267 38953
rect 16209 38913 16221 38947
rect 16255 38944 16267 38947
rect 16482 38944 16488 38956
rect 16255 38916 16488 38944
rect 16255 38913 16267 38916
rect 16209 38907 16267 38913
rect 16482 38904 16488 38916
rect 16540 38904 16546 38956
rect 10689 38879 10747 38885
rect 10689 38876 10701 38879
rect 10560 38848 10701 38876
rect 10560 38836 10566 38848
rect 10689 38845 10701 38848
rect 10735 38876 10747 38879
rect 11057 38879 11115 38885
rect 11057 38876 11069 38879
rect 10735 38848 11069 38876
rect 10735 38845 10747 38848
rect 10689 38839 10747 38845
rect 11057 38845 11069 38848
rect 11103 38845 11115 38879
rect 11330 38876 11336 38888
rect 11291 38848 11336 38876
rect 11057 38839 11115 38845
rect 11330 38836 11336 38848
rect 11388 38836 11394 38888
rect 11517 38879 11575 38885
rect 11517 38845 11529 38879
rect 11563 38876 11575 38879
rect 12437 38879 12495 38885
rect 12437 38876 12449 38879
rect 11563 38848 12449 38876
rect 11563 38845 11575 38848
rect 11517 38839 11575 38845
rect 12437 38845 12449 38848
rect 12483 38876 12495 38879
rect 12618 38876 12624 38888
rect 12483 38848 12624 38876
rect 12483 38845 12495 38848
rect 12437 38839 12495 38845
rect 12618 38836 12624 38848
rect 12676 38836 12682 38888
rect 15289 38879 15347 38885
rect 15289 38845 15301 38879
rect 15335 38876 15347 38879
rect 15378 38876 15384 38888
rect 15335 38848 15384 38876
rect 15335 38845 15347 38848
rect 15289 38839 15347 38845
rect 15378 38836 15384 38848
rect 15436 38876 15442 38888
rect 17218 38876 17224 38888
rect 15436 38848 17224 38876
rect 15436 38836 15442 38848
rect 17218 38836 17224 38848
rect 17276 38836 17282 38888
rect 19168 38885 19196 38984
rect 20272 38944 20300 39043
rect 21818 39040 21824 39092
rect 21876 39080 21882 39092
rect 22327 39083 22385 39089
rect 22327 39080 22339 39083
rect 21876 39052 22339 39080
rect 21876 39040 21882 39052
rect 22327 39049 22339 39052
rect 22373 39080 22385 39083
rect 23017 39083 23075 39089
rect 23017 39080 23029 39083
rect 22373 39052 23029 39080
rect 22373 39049 22385 39052
rect 22327 39043 22385 39049
rect 23017 39049 23029 39052
rect 23063 39049 23075 39083
rect 23017 39043 23075 39049
rect 26513 39083 26571 39089
rect 26513 39049 26525 39083
rect 26559 39080 26571 39083
rect 26970 39080 26976 39092
rect 26559 39052 26976 39080
rect 26559 39049 26571 39052
rect 26513 39043 26571 39049
rect 26970 39040 26976 39052
rect 27028 39080 27034 39092
rect 27111 39083 27169 39089
rect 27111 39080 27123 39083
rect 27028 39052 27123 39080
rect 27028 39040 27034 39052
rect 27111 39049 27123 39052
rect 27157 39049 27169 39083
rect 27111 39043 27169 39049
rect 28994 39040 29000 39092
rect 29052 39080 29058 39092
rect 30650 39080 30656 39092
rect 29052 39052 30656 39080
rect 29052 39040 29058 39052
rect 30650 39040 30656 39052
rect 30708 39040 30714 39092
rect 32858 39040 32864 39092
rect 32916 39080 32922 39092
rect 33873 39083 33931 39089
rect 33873 39080 33885 39083
rect 32916 39052 33885 39080
rect 32916 39040 32922 39052
rect 33873 39049 33885 39052
rect 33919 39049 33931 39083
rect 35618 39080 35624 39092
rect 35579 39052 35624 39080
rect 33873 39043 33931 39049
rect 35618 39040 35624 39052
rect 35676 39040 35682 39092
rect 38562 39040 38568 39092
rect 38620 39080 38626 39092
rect 39577 39083 39635 39089
rect 39577 39080 39589 39083
rect 38620 39052 39589 39080
rect 38620 39040 38626 39052
rect 39577 39049 39589 39052
rect 39623 39049 39635 39083
rect 39577 39043 39635 39049
rect 40865 39083 40923 39089
rect 40865 39049 40877 39083
rect 40911 39080 40923 39083
rect 41417 39083 41475 39089
rect 41417 39080 41429 39083
rect 40911 39052 41429 39080
rect 40911 39049 40923 39052
rect 40865 39043 40923 39049
rect 41417 39049 41429 39052
rect 41463 39080 41475 39083
rect 41506 39080 41512 39092
rect 41463 39052 41512 39080
rect 41463 39049 41475 39052
rect 41417 39043 41475 39049
rect 41506 39040 41512 39052
rect 41564 39040 41570 39092
rect 27433 39015 27491 39021
rect 27433 39012 27445 39015
rect 23446 38984 27445 39012
rect 23446 38944 23474 38984
rect 24302 38944 24308 38956
rect 20272 38916 20576 38944
rect 19153 38879 19211 38885
rect 19153 38845 19165 38879
rect 19199 38845 19211 38879
rect 19153 38839 19211 38845
rect 11698 38768 11704 38820
rect 11756 38808 11762 38820
rect 12161 38811 12219 38817
rect 12161 38808 12173 38811
rect 11756 38780 12173 38808
rect 11756 38768 11762 38780
rect 12161 38777 12173 38780
rect 12207 38808 12219 38811
rect 12758 38811 12816 38817
rect 12758 38808 12770 38811
rect 12207 38780 12770 38808
rect 12207 38777 12219 38780
rect 12161 38771 12219 38777
rect 12758 38777 12770 38780
rect 12804 38777 12816 38811
rect 12758 38771 12816 38777
rect 13648 38780 13814 38808
rect 11882 38740 11888 38752
rect 11843 38712 11888 38740
rect 11882 38700 11888 38712
rect 11940 38700 11946 38752
rect 13357 38743 13415 38749
rect 13357 38709 13369 38743
rect 13403 38740 13415 38743
rect 13446 38740 13452 38752
rect 13403 38712 13452 38740
rect 13403 38709 13415 38712
rect 13357 38703 13415 38709
rect 13446 38700 13452 38712
rect 13504 38740 13510 38752
rect 13648 38749 13676 38780
rect 13633 38743 13691 38749
rect 13633 38740 13645 38743
rect 13504 38712 13645 38740
rect 13504 38700 13510 38712
rect 13633 38709 13645 38712
rect 13679 38709 13691 38743
rect 13786 38740 13814 38780
rect 14734 38768 14740 38820
rect 14792 38808 14798 38820
rect 16530 38811 16588 38817
rect 16530 38808 16542 38811
rect 14792 38780 14837 38808
rect 16040 38780 16542 38808
rect 14792 38768 14798 38780
rect 14752 38740 14780 38768
rect 16040 38749 16068 38780
rect 16530 38777 16542 38780
rect 16576 38808 16588 38811
rect 18509 38811 18567 38817
rect 18509 38808 18521 38811
rect 16576 38780 18521 38808
rect 16576 38777 16588 38780
rect 16530 38771 16588 38777
rect 18509 38777 18521 38780
rect 18555 38808 18567 38811
rect 18690 38808 18696 38820
rect 18555 38780 18696 38808
rect 18555 38777 18567 38780
rect 18509 38771 18567 38777
rect 18690 38768 18696 38780
rect 18748 38768 18754 38820
rect 13786 38712 14780 38740
rect 16025 38743 16083 38749
rect 13633 38703 13691 38709
rect 16025 38709 16037 38743
rect 16071 38709 16083 38743
rect 17862 38740 17868 38752
rect 17823 38712 17868 38740
rect 16025 38703 16083 38709
rect 17862 38700 17868 38712
rect 17920 38700 17926 38752
rect 19168 38740 19196 38839
rect 19242 38836 19248 38888
rect 19300 38876 19306 38888
rect 19337 38879 19395 38885
rect 19337 38876 19349 38879
rect 19300 38848 19349 38876
rect 19300 38836 19306 38848
rect 19337 38845 19349 38848
rect 19383 38845 19395 38879
rect 19337 38839 19395 38845
rect 19613 38879 19671 38885
rect 19613 38845 19625 38879
rect 19659 38876 19671 38879
rect 20438 38876 20444 38888
rect 19659 38848 20444 38876
rect 19659 38845 19671 38848
rect 19613 38839 19671 38845
rect 20438 38836 20444 38848
rect 20496 38836 20502 38888
rect 20548 38808 20576 38916
rect 22664 38916 23474 38944
rect 24215 38916 24308 38944
rect 22664 38888 22692 38916
rect 24302 38904 24308 38916
rect 24360 38944 24366 38956
rect 24673 38947 24731 38953
rect 24673 38944 24685 38947
rect 24360 38916 24685 38944
rect 24360 38904 24366 38916
rect 24673 38913 24685 38916
rect 24719 38944 24731 38947
rect 24762 38944 24768 38956
rect 24719 38916 24768 38944
rect 24719 38913 24731 38916
rect 24673 38907 24731 38913
rect 24762 38904 24768 38916
rect 24820 38944 24826 38956
rect 25041 38947 25099 38953
rect 25041 38944 25053 38947
rect 24820 38916 25053 38944
rect 24820 38904 24826 38916
rect 25041 38913 25053 38916
rect 25087 38913 25099 38947
rect 25222 38944 25228 38956
rect 25183 38916 25228 38944
rect 25041 38907 25099 38913
rect 25222 38904 25228 38916
rect 25280 38904 25286 38956
rect 21361 38879 21419 38885
rect 21361 38845 21373 38879
rect 21407 38876 21419 38879
rect 22256 38879 22314 38885
rect 21407 38848 21864 38876
rect 21407 38845 21419 38848
rect 21361 38839 21419 38845
rect 20622 38808 20628 38820
rect 20535 38780 20628 38808
rect 20622 38768 20628 38780
rect 20680 38808 20686 38820
rect 21836 38817 21864 38848
rect 22256 38845 22268 38879
rect 22302 38876 22314 38879
rect 22646 38876 22652 38888
rect 22302 38848 22652 38876
rect 22302 38845 22314 38848
rect 22256 38839 22314 38845
rect 22646 38836 22652 38848
rect 22704 38836 22710 38888
rect 23474 38836 23480 38888
rect 23532 38876 23538 38888
rect 23661 38879 23719 38885
rect 23661 38876 23673 38879
rect 23532 38848 23673 38876
rect 23532 38836 23538 38848
rect 23661 38845 23673 38848
rect 23707 38845 23719 38879
rect 23661 38839 23719 38845
rect 20762 38811 20820 38817
rect 20762 38808 20774 38811
rect 20680 38780 20774 38808
rect 20680 38768 20686 38780
rect 20762 38777 20774 38780
rect 20808 38777 20820 38811
rect 20762 38771 20820 38777
rect 21821 38811 21879 38817
rect 21821 38777 21833 38811
rect 21867 38808 21879 38811
rect 22002 38808 22008 38820
rect 21867 38780 22008 38808
rect 21867 38777 21879 38780
rect 21821 38771 21879 38777
rect 22002 38768 22008 38780
rect 22060 38808 22066 38820
rect 23198 38808 23204 38820
rect 22060 38780 23204 38808
rect 22060 38768 22066 38780
rect 23198 38768 23204 38780
rect 23256 38768 23262 38820
rect 23676 38808 23704 38839
rect 23750 38836 23756 38888
rect 23808 38876 23814 38888
rect 24121 38879 24179 38885
rect 24121 38876 24133 38879
rect 23808 38848 24133 38876
rect 23808 38836 23814 38848
rect 24121 38845 24133 38848
rect 24167 38876 24179 38879
rect 25314 38876 25320 38888
rect 24167 38848 25320 38876
rect 24167 38845 24179 38848
rect 24121 38839 24179 38845
rect 25314 38836 25320 38848
rect 25372 38836 25378 38888
rect 27023 38885 27051 38984
rect 27433 38981 27445 38984
rect 27479 39012 27491 39015
rect 31662 39012 31668 39024
rect 27479 38984 31668 39012
rect 27479 38981 27491 38984
rect 27433 38975 27491 38981
rect 31662 38972 31668 38984
rect 31720 38972 31726 39024
rect 32398 38972 32404 39024
rect 32456 39012 32462 39024
rect 33134 39012 33140 39024
rect 32456 38984 33140 39012
rect 32456 38972 32462 38984
rect 33134 38972 33140 38984
rect 33192 39012 33198 39024
rect 33192 38984 33285 39012
rect 33192 38972 33198 38984
rect 36814 38972 36820 39024
rect 36872 39012 36878 39024
rect 37826 39012 37832 39024
rect 36872 38984 37832 39012
rect 36872 38972 36878 38984
rect 37826 38972 37832 38984
rect 37884 39012 37890 39024
rect 39209 39015 39267 39021
rect 39209 39012 39221 39015
rect 37884 38984 39221 39012
rect 37884 38972 37890 38984
rect 39209 38981 39221 38984
rect 39255 38981 39267 39015
rect 39209 38975 39267 38981
rect 28721 38947 28779 38953
rect 28721 38913 28733 38947
rect 28767 38944 28779 38947
rect 32953 38947 33011 38953
rect 28767 38916 29776 38944
rect 28767 38913 28779 38916
rect 28721 38907 28779 38913
rect 27008 38879 27066 38885
rect 27008 38845 27020 38879
rect 27054 38845 27066 38879
rect 29270 38876 29276 38888
rect 27008 38839 27066 38845
rect 27126 38848 29276 38876
rect 25498 38808 25504 38820
rect 23676 38780 25176 38808
rect 25459 38780 25504 38808
rect 19978 38740 19984 38752
rect 19168 38712 19984 38740
rect 19978 38700 19984 38712
rect 20036 38700 20042 38752
rect 23382 38700 23388 38752
rect 23440 38740 23446 38752
rect 23934 38740 23940 38752
rect 23440 38712 23940 38740
rect 23440 38700 23446 38712
rect 23934 38700 23940 38712
rect 23992 38700 23998 38752
rect 25148 38740 25176 38780
rect 25498 38768 25504 38780
rect 25556 38768 25562 38820
rect 27126 38808 27154 38848
rect 29270 38836 29276 38848
rect 29328 38836 29334 38888
rect 29748 38885 29776 38916
rect 32953 38913 32965 38947
rect 32999 38944 33011 38947
rect 33042 38944 33048 38956
rect 32999 38916 33048 38944
rect 32999 38913 33011 38916
rect 32953 38907 33011 38913
rect 33042 38904 33048 38916
rect 33100 38904 33106 38956
rect 33152 38944 33180 38972
rect 33229 38947 33287 38953
rect 33229 38944 33241 38947
rect 33152 38916 33241 38944
rect 33229 38913 33241 38916
rect 33275 38913 33287 38947
rect 33229 38907 33287 38913
rect 35207 38947 35265 38953
rect 35207 38913 35219 38947
rect 35253 38944 35265 38947
rect 36173 38947 36231 38953
rect 36173 38944 36185 38947
rect 35253 38916 36185 38944
rect 35253 38913 35265 38916
rect 35207 38907 35265 38913
rect 36173 38913 36185 38916
rect 36219 38944 36231 38947
rect 37093 38947 37151 38953
rect 37093 38944 37105 38947
rect 36219 38916 37105 38944
rect 36219 38913 36231 38916
rect 36173 38907 36231 38913
rect 37093 38913 37105 38916
rect 37139 38913 37151 38947
rect 37093 38907 37151 38913
rect 37737 38947 37795 38953
rect 37737 38913 37749 38947
rect 37783 38944 37795 38947
rect 38657 38947 38715 38953
rect 38657 38944 38669 38947
rect 37783 38916 38669 38944
rect 37783 38913 37795 38916
rect 37737 38907 37795 38913
rect 38657 38913 38669 38916
rect 38703 38944 38715 38947
rect 41647 38947 41705 38953
rect 41647 38944 41659 38947
rect 38703 38916 41659 38944
rect 38703 38913 38715 38916
rect 38657 38907 38715 38913
rect 41647 38913 41659 38916
rect 41693 38913 41705 38947
rect 41647 38907 41705 38913
rect 29733 38879 29791 38885
rect 29733 38845 29745 38879
rect 29779 38876 29791 38879
rect 30006 38876 30012 38888
rect 29779 38848 30012 38876
rect 29779 38845 29791 38848
rect 29733 38839 29791 38845
rect 30006 38836 30012 38848
rect 30064 38836 30070 38888
rect 30742 38836 30748 38888
rect 30800 38876 30806 38888
rect 30837 38879 30895 38885
rect 30837 38876 30849 38879
rect 30800 38848 30849 38876
rect 30800 38836 30806 38848
rect 30837 38845 30849 38848
rect 30883 38845 30895 38879
rect 34422 38876 34428 38888
rect 34383 38848 34428 38876
rect 30837 38839 30895 38845
rect 34422 38836 34428 38848
rect 34480 38836 34486 38888
rect 35120 38879 35178 38885
rect 35120 38845 35132 38879
rect 35166 38876 35178 38879
rect 35618 38876 35624 38888
rect 35166 38848 35624 38876
rect 35166 38845 35178 38848
rect 35120 38839 35178 38845
rect 35618 38836 35624 38848
rect 35676 38836 35682 38888
rect 39298 38836 39304 38888
rect 39356 38876 39362 38888
rect 39942 38876 39948 38888
rect 39356 38848 39948 38876
rect 39356 38836 39362 38848
rect 39942 38836 39948 38848
rect 40000 38876 40006 38888
rect 40564 38879 40622 38885
rect 40564 38876 40576 38879
rect 40000 38848 40576 38876
rect 40000 38836 40006 38848
rect 40564 38845 40576 38848
rect 40610 38876 40622 38879
rect 40865 38879 40923 38885
rect 40865 38876 40877 38879
rect 40610 38848 40877 38876
rect 40610 38845 40622 38848
rect 40564 38839 40622 38845
rect 40865 38845 40877 38848
rect 40911 38845 40923 38879
rect 40865 38839 40923 38845
rect 41322 38836 41328 38888
rect 41380 38876 41386 38888
rect 41544 38879 41602 38885
rect 41544 38876 41556 38879
rect 41380 38848 41556 38876
rect 41380 38836 41386 38848
rect 41544 38845 41556 38848
rect 41590 38876 41602 38879
rect 41969 38879 42027 38885
rect 41969 38876 41981 38879
rect 41590 38848 41981 38876
rect 41590 38845 41602 38848
rect 41544 38839 41602 38845
rect 41969 38845 41981 38848
rect 42015 38876 42027 38879
rect 46934 38876 46940 38888
rect 42015 38848 46940 38876
rect 42015 38845 42027 38848
rect 41969 38839 42027 38845
rect 46934 38836 46940 38848
rect 46992 38836 46998 38888
rect 25700 38780 27154 38808
rect 28353 38811 28411 38817
rect 25700 38740 25728 38780
rect 28353 38777 28365 38811
rect 28399 38808 28411 38811
rect 28399 38780 29224 38808
rect 28399 38777 28411 38780
rect 28353 38771 28411 38777
rect 29196 38752 29224 38780
rect 30650 38768 30656 38820
rect 30708 38808 30714 38820
rect 31158 38811 31216 38817
rect 31158 38808 31170 38811
rect 30708 38780 31170 38808
rect 30708 38768 30714 38780
rect 31158 38777 31170 38780
rect 31204 38777 31216 38811
rect 31158 38771 31216 38777
rect 33045 38811 33103 38817
rect 33045 38777 33057 38811
rect 33091 38777 33103 38811
rect 33045 38771 33103 38777
rect 35989 38811 36047 38817
rect 35989 38777 36001 38811
rect 36035 38808 36047 38811
rect 36265 38811 36323 38817
rect 36265 38808 36277 38811
rect 36035 38780 36277 38808
rect 36035 38777 36047 38780
rect 35989 38771 36047 38777
rect 36265 38777 36277 38780
rect 36311 38808 36323 38811
rect 36446 38808 36452 38820
rect 36311 38780 36452 38808
rect 36311 38777 36323 38780
rect 36265 38771 36323 38777
rect 25148 38712 25728 38740
rect 26145 38743 26203 38749
rect 26145 38709 26157 38743
rect 26191 38740 26203 38743
rect 26881 38743 26939 38749
rect 26881 38740 26893 38743
rect 26191 38712 26893 38740
rect 26191 38709 26203 38712
rect 26145 38703 26203 38709
rect 26881 38709 26893 38712
rect 26927 38740 26939 38743
rect 27062 38740 27068 38752
rect 26927 38712 27068 38740
rect 26927 38709 26939 38712
rect 26881 38703 26939 38709
rect 27062 38700 27068 38712
rect 27120 38700 27126 38752
rect 28994 38740 29000 38752
rect 28955 38712 29000 38740
rect 28994 38700 29000 38712
rect 29052 38700 29058 38752
rect 29178 38700 29184 38752
rect 29236 38740 29242 38752
rect 29365 38743 29423 38749
rect 29365 38740 29377 38743
rect 29236 38712 29377 38740
rect 29236 38700 29242 38712
rect 29365 38709 29377 38712
rect 29411 38709 29423 38743
rect 31754 38740 31760 38752
rect 31715 38712 31760 38740
rect 29365 38703 29423 38709
rect 31754 38700 31760 38712
rect 31812 38700 31818 38752
rect 32401 38743 32459 38749
rect 32401 38709 32413 38743
rect 32447 38740 32459 38743
rect 32674 38740 32680 38752
rect 32447 38712 32680 38740
rect 32447 38709 32459 38712
rect 32401 38703 32459 38709
rect 32674 38700 32680 38712
rect 32732 38740 32738 38752
rect 33060 38740 33088 38771
rect 36446 38768 36452 38780
rect 36504 38768 36510 38820
rect 36817 38811 36875 38817
rect 36817 38777 36829 38811
rect 36863 38808 36875 38811
rect 36998 38808 37004 38820
rect 36863 38780 37004 38808
rect 36863 38777 36875 38780
rect 36817 38771 36875 38777
rect 36998 38768 37004 38780
rect 37056 38768 37062 38820
rect 38105 38811 38163 38817
rect 38105 38777 38117 38811
rect 38151 38808 38163 38811
rect 38473 38811 38531 38817
rect 38473 38808 38485 38811
rect 38151 38780 38485 38808
rect 38151 38777 38163 38780
rect 38105 38771 38163 38777
rect 38473 38777 38485 38780
rect 38519 38808 38531 38811
rect 38749 38811 38807 38817
rect 38749 38808 38761 38811
rect 38519 38780 38761 38808
rect 38519 38777 38531 38780
rect 38473 38771 38531 38777
rect 38749 38777 38761 38780
rect 38795 38808 38807 38811
rect 38838 38808 38844 38820
rect 38795 38780 38844 38808
rect 38795 38777 38807 38780
rect 38749 38771 38807 38777
rect 38838 38768 38844 38780
rect 38896 38768 38902 38820
rect 40770 38808 40776 38820
rect 40281 38780 40776 38808
rect 32732 38712 33088 38740
rect 32732 38700 32738 38712
rect 35894 38700 35900 38752
rect 35952 38740 35958 38752
rect 38562 38740 38568 38752
rect 35952 38712 38568 38740
rect 35952 38700 35958 38712
rect 38562 38700 38568 38712
rect 38620 38740 38626 38752
rect 40281 38740 40309 38780
rect 40770 38768 40776 38780
rect 40828 38808 40834 38820
rect 40957 38811 41015 38817
rect 40957 38808 40969 38811
rect 40828 38780 40969 38808
rect 40828 38768 40834 38780
rect 40957 38777 40969 38780
rect 41003 38777 41015 38811
rect 40957 38771 41015 38777
rect 38620 38712 40309 38740
rect 40635 38743 40693 38749
rect 38620 38700 38626 38712
rect 40635 38709 40647 38743
rect 40681 38740 40693 38743
rect 40862 38740 40868 38752
rect 40681 38712 40868 38740
rect 40681 38709 40693 38712
rect 40635 38703 40693 38709
rect 40862 38700 40868 38712
rect 40920 38700 40926 38752
rect 1104 38650 48852 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 48852 38650
rect 1104 38576 48852 38598
rect 10873 38539 10931 38545
rect 10873 38505 10885 38539
rect 10919 38536 10931 38539
rect 11330 38536 11336 38548
rect 10919 38508 11336 38536
rect 10919 38505 10931 38508
rect 10873 38499 10931 38505
rect 11330 38496 11336 38508
rect 11388 38496 11394 38548
rect 11698 38496 11704 38548
rect 11756 38536 11762 38548
rect 11793 38539 11851 38545
rect 11793 38536 11805 38539
rect 11756 38508 11805 38536
rect 11756 38496 11762 38508
rect 11793 38505 11805 38508
rect 11839 38505 11851 38539
rect 12618 38536 12624 38548
rect 12579 38508 12624 38536
rect 11793 38499 11851 38505
rect 12618 38496 12624 38508
rect 12676 38496 12682 38548
rect 13722 38496 13728 38548
rect 13780 38536 13786 38548
rect 14553 38539 14611 38545
rect 14553 38536 14565 38539
rect 13780 38508 14565 38536
rect 13780 38496 13786 38508
rect 14553 38505 14565 38508
rect 14599 38505 14611 38539
rect 16666 38536 16672 38548
rect 16627 38508 16672 38536
rect 14553 38499 14611 38505
rect 16666 38496 16672 38508
rect 16724 38496 16730 38548
rect 17862 38496 17868 38548
rect 17920 38536 17926 38548
rect 18506 38536 18512 38548
rect 17920 38508 18512 38536
rect 17920 38496 17926 38508
rect 18506 38496 18512 38508
rect 18564 38496 18570 38548
rect 20438 38536 20444 38548
rect 20399 38508 20444 38536
rect 20438 38496 20444 38508
rect 20496 38496 20502 38548
rect 23382 38496 23388 38548
rect 23440 38536 23446 38548
rect 24305 38539 24363 38545
rect 24305 38536 24317 38539
rect 23440 38508 24317 38536
rect 23440 38496 23446 38508
rect 24305 38505 24317 38508
rect 24351 38505 24363 38539
rect 24305 38499 24363 38505
rect 25133 38539 25191 38545
rect 25133 38505 25145 38539
rect 25179 38536 25191 38539
rect 25222 38536 25228 38548
rect 25179 38508 25228 38536
rect 25179 38505 25191 38508
rect 25133 38499 25191 38505
rect 25222 38496 25228 38508
rect 25280 38496 25286 38548
rect 25498 38496 25504 38548
rect 25556 38536 25562 38548
rect 28994 38536 29000 38548
rect 25556 38508 29000 38536
rect 25556 38496 25562 38508
rect 28994 38496 29000 38508
rect 29052 38496 29058 38548
rect 30282 38496 30288 38548
rect 30340 38536 30346 38548
rect 30926 38536 30932 38548
rect 30340 38508 30932 38536
rect 30340 38496 30346 38508
rect 30926 38496 30932 38508
rect 30984 38536 30990 38548
rect 31021 38539 31079 38545
rect 31021 38536 31033 38539
rect 30984 38508 31033 38536
rect 30984 38496 30990 38508
rect 31021 38505 31033 38508
rect 31067 38505 31079 38539
rect 31021 38499 31079 38505
rect 33042 38496 33048 38548
rect 33100 38536 33106 38548
rect 33413 38539 33471 38545
rect 33413 38536 33425 38539
rect 33100 38508 33425 38536
rect 33100 38496 33106 38508
rect 33413 38505 33425 38508
rect 33459 38505 33471 38539
rect 38102 38536 38108 38548
rect 38063 38508 38108 38536
rect 33413 38499 33471 38505
rect 38102 38496 38108 38508
rect 38160 38496 38166 38548
rect 38746 38496 38752 38548
rect 38804 38536 38810 38548
rect 39623 38539 39681 38545
rect 39623 38536 39635 38539
rect 38804 38508 39635 38536
rect 38804 38496 38810 38508
rect 39623 38505 39635 38508
rect 39669 38505 39681 38539
rect 39623 38499 39681 38505
rect 13262 38468 13268 38480
rect 13223 38440 13268 38468
rect 13262 38428 13268 38440
rect 13320 38428 13326 38480
rect 13357 38471 13415 38477
rect 13357 38437 13369 38471
rect 13403 38468 13415 38471
rect 13446 38468 13452 38480
rect 13403 38440 13452 38468
rect 13403 38437 13415 38440
rect 13357 38431 13415 38437
rect 13446 38428 13452 38440
rect 13504 38428 13510 38480
rect 15470 38468 15476 38480
rect 15431 38440 15476 38468
rect 15470 38428 15476 38440
rect 15528 38468 15534 38480
rect 17037 38471 17095 38477
rect 17037 38468 17049 38471
rect 15528 38440 17049 38468
rect 15528 38428 15534 38440
rect 17037 38437 17049 38440
rect 17083 38437 17095 38471
rect 17037 38431 17095 38437
rect 21818 38428 21824 38480
rect 21876 38468 21882 38480
rect 21913 38471 21971 38477
rect 21913 38468 21925 38471
rect 21876 38440 21925 38468
rect 21876 38428 21882 38440
rect 21913 38437 21925 38440
rect 21959 38437 21971 38471
rect 21913 38431 21971 38437
rect 23198 38428 23204 38480
rect 23256 38468 23262 38480
rect 23477 38471 23535 38477
rect 23477 38468 23489 38471
rect 23256 38440 23489 38468
rect 23256 38428 23262 38440
rect 23477 38437 23489 38440
rect 23523 38437 23535 38471
rect 27062 38468 27068 38480
rect 26975 38440 27068 38468
rect 23477 38431 23535 38437
rect 27062 38428 27068 38440
rect 27120 38468 27126 38480
rect 27706 38468 27712 38480
rect 27120 38440 27712 38468
rect 27120 38428 27126 38440
rect 27706 38428 27712 38440
rect 27764 38428 27770 38480
rect 29546 38428 29552 38480
rect 29604 38468 29610 38480
rect 30098 38468 30104 38480
rect 29604 38440 30104 38468
rect 29604 38428 29610 38440
rect 30098 38428 30104 38440
rect 30156 38468 30162 38480
rect 30193 38471 30251 38477
rect 30193 38468 30205 38471
rect 30156 38440 30205 38468
rect 30156 38428 30162 38440
rect 30193 38437 30205 38440
rect 30239 38437 30251 38471
rect 30193 38431 30251 38437
rect 31570 38428 31576 38480
rect 31628 38468 31634 38480
rect 32493 38471 32551 38477
rect 32493 38468 32505 38471
rect 31628 38440 32505 38468
rect 31628 38428 31634 38440
rect 32493 38437 32505 38440
rect 32539 38437 32551 38471
rect 32493 38431 32551 38437
rect 32582 38428 32588 38480
rect 32640 38468 32646 38480
rect 32640 38440 32685 38468
rect 32640 38428 32646 38440
rect 32858 38428 32864 38480
rect 32916 38468 32922 38480
rect 34103 38471 34161 38477
rect 34103 38468 34115 38471
rect 32916 38440 34115 38468
rect 32916 38428 32922 38440
rect 34103 38437 34115 38440
rect 34149 38437 34161 38471
rect 34103 38431 34161 38437
rect 35615 38471 35673 38477
rect 35615 38437 35627 38471
rect 35661 38468 35673 38471
rect 35802 38468 35808 38480
rect 35661 38440 35808 38468
rect 35661 38437 35673 38440
rect 35615 38431 35673 38437
rect 35802 38428 35808 38440
rect 35860 38428 35866 38480
rect 40957 38471 41015 38477
rect 40957 38437 40969 38471
rect 41003 38468 41015 38471
rect 41046 38468 41052 38480
rect 41003 38440 41052 38468
rect 41003 38437 41015 38440
rect 40957 38431 41015 38437
rect 41046 38428 41052 38440
rect 41104 38428 41110 38480
rect 18414 38400 18420 38412
rect 18375 38372 18420 38400
rect 18414 38360 18420 38372
rect 18472 38360 18478 38412
rect 18969 38403 19027 38409
rect 18969 38369 18981 38403
rect 19015 38400 19027 38403
rect 19150 38400 19156 38412
rect 19015 38372 19156 38400
rect 19015 38369 19027 38372
rect 18969 38363 19027 38369
rect 19150 38360 19156 38372
rect 19208 38360 19214 38412
rect 25130 38400 25136 38412
rect 25091 38372 25136 38400
rect 25130 38360 25136 38372
rect 25188 38360 25194 38412
rect 25314 38400 25320 38412
rect 25275 38372 25320 38400
rect 25314 38360 25320 38372
rect 25372 38360 25378 38412
rect 28442 38400 28448 38412
rect 28403 38372 28448 38400
rect 28442 38360 28448 38372
rect 28500 38360 28506 38412
rect 33962 38400 33968 38412
rect 33926 38372 33968 38400
rect 33962 38360 33968 38372
rect 34020 38409 34026 38412
rect 34020 38403 34074 38409
rect 34020 38369 34028 38403
rect 34062 38400 34074 38403
rect 35894 38400 35900 38412
rect 34062 38372 35900 38400
rect 34062 38369 34074 38372
rect 34020 38363 34074 38369
rect 34020 38360 34026 38363
rect 35894 38360 35900 38372
rect 35952 38360 35958 38412
rect 37734 38400 37740 38412
rect 37695 38372 37740 38400
rect 37734 38360 37740 38372
rect 37792 38360 37798 38412
rect 38657 38403 38715 38409
rect 38657 38369 38669 38403
rect 38703 38400 38715 38403
rect 38838 38400 38844 38412
rect 38703 38372 38844 38400
rect 38703 38369 38715 38372
rect 38657 38363 38715 38369
rect 38838 38360 38844 38372
rect 38896 38360 38902 38412
rect 39485 38403 39543 38409
rect 39485 38369 39497 38403
rect 39531 38400 39543 38403
rect 39574 38400 39580 38412
rect 39531 38372 39580 38400
rect 39531 38369 39543 38372
rect 39485 38363 39543 38369
rect 39574 38360 39580 38372
rect 39632 38360 39638 38412
rect 11425 38335 11483 38341
rect 11425 38301 11437 38335
rect 11471 38332 11483 38335
rect 11514 38332 11520 38344
rect 11471 38304 11520 38332
rect 11471 38301 11483 38304
rect 11425 38295 11483 38301
rect 11514 38292 11520 38304
rect 11572 38292 11578 38344
rect 12618 38292 12624 38344
rect 12676 38332 12682 38344
rect 13541 38335 13599 38341
rect 13541 38332 13553 38335
rect 12676 38304 13553 38332
rect 12676 38292 12682 38304
rect 13541 38301 13553 38304
rect 13587 38301 13599 38335
rect 13541 38295 13599 38301
rect 15381 38335 15439 38341
rect 15381 38301 15393 38335
rect 15427 38332 15439 38335
rect 15838 38332 15844 38344
rect 15427 38304 15844 38332
rect 15427 38301 15439 38304
rect 15381 38295 15439 38301
rect 15838 38292 15844 38304
rect 15896 38292 15902 38344
rect 16022 38332 16028 38344
rect 15983 38304 16028 38332
rect 16022 38292 16028 38304
rect 16080 38292 16086 38344
rect 16942 38332 16948 38344
rect 16903 38304 16948 38332
rect 16942 38292 16948 38304
rect 17000 38292 17006 38344
rect 17218 38332 17224 38344
rect 17179 38304 17224 38332
rect 17218 38292 17224 38304
rect 17276 38292 17282 38344
rect 21821 38335 21879 38341
rect 21821 38301 21833 38335
rect 21867 38332 21879 38335
rect 22186 38332 22192 38344
rect 21867 38304 22192 38332
rect 21867 38301 21879 38304
rect 21821 38295 21879 38301
rect 22186 38292 22192 38304
rect 22244 38292 22250 38344
rect 22278 38292 22284 38344
rect 22336 38332 22342 38344
rect 22336 38304 22381 38332
rect 22336 38292 22342 38304
rect 23198 38292 23204 38344
rect 23256 38332 23262 38344
rect 23385 38335 23443 38341
rect 23385 38332 23397 38335
rect 23256 38304 23397 38332
rect 23256 38292 23262 38304
rect 23385 38301 23397 38304
rect 23431 38301 23443 38335
rect 23658 38332 23664 38344
rect 23619 38304 23664 38332
rect 23385 38295 23443 38301
rect 23658 38292 23664 38304
rect 23716 38292 23722 38344
rect 26973 38335 27031 38341
rect 26973 38301 26985 38335
rect 27019 38332 27031 38335
rect 28074 38332 28080 38344
rect 27019 38304 28080 38332
rect 27019 38301 27031 38304
rect 26973 38295 27031 38301
rect 28074 38292 28080 38304
rect 28132 38332 28138 38344
rect 28583 38335 28641 38341
rect 28583 38332 28595 38335
rect 28132 38304 28595 38332
rect 28132 38292 28138 38304
rect 28583 38301 28595 38304
rect 28629 38301 28641 38335
rect 28583 38295 28641 38301
rect 29914 38292 29920 38344
rect 29972 38332 29978 38344
rect 30101 38335 30159 38341
rect 30101 38332 30113 38335
rect 29972 38304 30113 38332
rect 29972 38292 29978 38304
rect 30101 38301 30113 38304
rect 30147 38301 30159 38335
rect 30101 38295 30159 38301
rect 30745 38335 30803 38341
rect 30745 38301 30757 38335
rect 30791 38332 30803 38335
rect 31846 38332 31852 38344
rect 30791 38304 31852 38332
rect 30791 38301 30803 38304
rect 30745 38295 30803 38301
rect 31846 38292 31852 38304
rect 31904 38332 31910 38344
rect 32030 38332 32036 38344
rect 31904 38304 32036 38332
rect 31904 38292 31910 38304
rect 32030 38292 32036 38304
rect 32088 38292 32094 38344
rect 32858 38292 32864 38344
rect 32916 38332 32922 38344
rect 34238 38332 34244 38344
rect 32916 38304 34244 38332
rect 32916 38292 32922 38304
rect 34238 38292 34244 38304
rect 34296 38292 34302 38344
rect 35250 38332 35256 38344
rect 35211 38304 35256 38332
rect 35250 38292 35256 38304
rect 35308 38292 35314 38344
rect 40862 38332 40868 38344
rect 40823 38304 40868 38332
rect 40862 38292 40868 38304
rect 40920 38292 40926 38344
rect 27522 38264 27528 38276
rect 27483 38236 27528 38264
rect 27522 38224 27528 38236
rect 27580 38224 27586 38276
rect 41414 38264 41420 38276
rect 41375 38236 41420 38264
rect 41414 38224 41420 38236
rect 41472 38224 41478 38276
rect 12342 38196 12348 38208
rect 12303 38168 12348 38196
rect 12342 38156 12348 38168
rect 12400 38156 12406 38208
rect 12526 38156 12532 38208
rect 12584 38196 12590 38208
rect 12989 38199 13047 38205
rect 12989 38196 13001 38199
rect 12584 38168 13001 38196
rect 12584 38156 12590 38168
rect 12989 38165 13001 38168
rect 13035 38165 13047 38199
rect 12989 38159 13047 38165
rect 19150 38156 19156 38208
rect 19208 38196 19214 38208
rect 19429 38199 19487 38205
rect 19429 38196 19441 38199
rect 19208 38168 19441 38196
rect 19208 38156 19214 38168
rect 19429 38165 19441 38168
rect 19475 38165 19487 38199
rect 19429 38159 19487 38165
rect 19978 38156 19984 38208
rect 20036 38196 20042 38208
rect 25130 38196 25136 38208
rect 20036 38168 25136 38196
rect 20036 38156 20042 38168
rect 25130 38156 25136 38168
rect 25188 38156 25194 38208
rect 29270 38196 29276 38208
rect 29183 38168 29276 38196
rect 29270 38156 29276 38168
rect 29328 38156 29334 38208
rect 31938 38156 31944 38208
rect 31996 38196 32002 38208
rect 35710 38196 35716 38208
rect 31996 38168 35716 38196
rect 31996 38156 32002 38168
rect 35710 38156 35716 38168
rect 35768 38156 35774 38208
rect 36173 38199 36231 38205
rect 36173 38165 36185 38199
rect 36219 38196 36231 38199
rect 36446 38196 36452 38208
rect 36219 38168 36452 38196
rect 36219 38165 36231 38168
rect 36173 38159 36231 38165
rect 36446 38156 36452 38168
rect 36504 38156 36510 38208
rect 36538 38156 36544 38208
rect 36596 38196 36602 38208
rect 36817 38199 36875 38205
rect 36817 38196 36829 38199
rect 36596 38168 36829 38196
rect 36596 38156 36602 38168
rect 36817 38165 36829 38168
rect 36863 38165 36875 38199
rect 38930 38196 38936 38208
rect 38891 38168 38936 38196
rect 36817 38159 36875 38165
rect 38930 38156 38936 38168
rect 38988 38156 38994 38208
rect 42518 38196 42524 38208
rect 42479 38168 42524 38196
rect 42518 38156 42524 38168
rect 42576 38156 42582 38208
rect 1104 38106 48852 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 48852 38106
rect 1104 38032 48852 38054
rect 13446 37992 13452 38004
rect 13407 37964 13452 37992
rect 13446 37952 13452 37964
rect 13504 37952 13510 38004
rect 17678 37952 17684 38004
rect 17736 37992 17742 38004
rect 18414 37992 18420 38004
rect 17736 37964 18420 37992
rect 17736 37952 17742 37964
rect 18414 37952 18420 37964
rect 18472 37952 18478 38004
rect 20533 37995 20591 38001
rect 20533 37961 20545 37995
rect 20579 37992 20591 37995
rect 20622 37992 20628 38004
rect 20579 37964 20628 37992
rect 20579 37961 20591 37964
rect 20533 37955 20591 37961
rect 20622 37952 20628 37964
rect 20680 37952 20686 38004
rect 22186 37992 22192 38004
rect 22147 37964 22192 37992
rect 22186 37952 22192 37964
rect 22244 37992 22250 38004
rect 22511 37995 22569 38001
rect 22511 37992 22523 37995
rect 22244 37964 22523 37992
rect 22244 37952 22250 37964
rect 22511 37961 22523 37964
rect 22557 37961 22569 37995
rect 23290 37992 23296 38004
rect 23251 37964 23296 37992
rect 22511 37955 22569 37961
rect 23290 37952 23296 37964
rect 23348 37952 23354 38004
rect 24762 37992 24768 38004
rect 24723 37964 24768 37992
rect 24762 37952 24768 37964
rect 24820 37952 24826 38004
rect 27706 37992 27712 38004
rect 27667 37964 27712 37992
rect 27706 37952 27712 37964
rect 27764 37952 27770 38004
rect 28074 37992 28080 38004
rect 28035 37964 28080 37992
rect 28074 37952 28080 37964
rect 28132 37952 28138 38004
rect 29546 37992 29552 38004
rect 29507 37964 29552 37992
rect 29546 37952 29552 37964
rect 29604 37952 29610 38004
rect 29914 37952 29920 38004
rect 29972 37992 29978 38004
rect 31021 37995 31079 38001
rect 31021 37992 31033 37995
rect 29972 37964 31033 37992
rect 29972 37952 29978 37964
rect 31021 37961 31033 37964
rect 31067 37961 31079 37995
rect 31021 37955 31079 37961
rect 31573 37995 31631 38001
rect 31573 37961 31585 37995
rect 31619 37992 31631 37995
rect 31754 37992 31760 38004
rect 31619 37964 31760 37992
rect 31619 37961 31631 37964
rect 31573 37955 31631 37961
rect 31754 37952 31760 37964
rect 31812 37992 31818 38004
rect 32493 37995 32551 38001
rect 32493 37992 32505 37995
rect 31812 37964 32505 37992
rect 31812 37952 31818 37964
rect 32493 37961 32505 37964
rect 32539 37992 32551 37995
rect 32582 37992 32588 38004
rect 32539 37964 32588 37992
rect 32539 37961 32551 37964
rect 32493 37955 32551 37961
rect 32582 37952 32588 37964
rect 32640 37992 32646 38004
rect 32858 37992 32864 38004
rect 32640 37964 32864 37992
rect 32640 37952 32646 37964
rect 32858 37952 32864 37964
rect 32916 37952 32922 38004
rect 33962 37992 33968 38004
rect 33923 37964 33968 37992
rect 33962 37952 33968 37964
rect 34020 37952 34026 38004
rect 37461 37995 37519 38001
rect 37461 37961 37473 37995
rect 37507 37992 37519 37995
rect 37734 37992 37740 38004
rect 37507 37964 37740 37992
rect 37507 37961 37519 37964
rect 37461 37955 37519 37961
rect 37734 37952 37740 37964
rect 37792 37952 37798 38004
rect 38473 37995 38531 38001
rect 38473 37961 38485 37995
rect 38519 37992 38531 37995
rect 38838 37992 38844 38004
rect 38519 37964 38844 37992
rect 38519 37961 38531 37964
rect 38473 37955 38531 37961
rect 38838 37952 38844 37964
rect 38896 37952 38902 38004
rect 40862 37952 40868 38004
rect 40920 37992 40926 38004
rect 41877 37995 41935 38001
rect 41877 37992 41889 37995
rect 40920 37964 41889 37992
rect 40920 37952 40926 37964
rect 41877 37961 41889 37964
rect 41923 37961 41935 37995
rect 41877 37955 41935 37961
rect 10796 37896 12940 37924
rect 10796 37797 10824 37896
rect 12526 37856 12532 37868
rect 12487 37828 12532 37856
rect 12526 37816 12532 37828
rect 12584 37816 12590 37868
rect 12618 37816 12624 37868
rect 12676 37856 12682 37868
rect 12805 37859 12863 37865
rect 12805 37856 12817 37859
rect 12676 37828 12817 37856
rect 12676 37816 12682 37828
rect 12805 37825 12817 37828
rect 12851 37825 12863 37859
rect 12912 37856 12940 37896
rect 13262 37884 13268 37936
rect 13320 37924 13326 37936
rect 13817 37927 13875 37933
rect 13817 37924 13829 37927
rect 13320 37896 13829 37924
rect 13320 37884 13326 37896
rect 13817 37893 13829 37896
rect 13863 37893 13875 37927
rect 13817 37887 13875 37893
rect 14323 37927 14381 37933
rect 14323 37893 14335 37927
rect 14369 37924 14381 37927
rect 15838 37924 15844 37936
rect 14369 37896 15844 37924
rect 14369 37893 14381 37896
rect 14323 37887 14381 37893
rect 15838 37884 15844 37896
rect 15896 37884 15902 37936
rect 17218 37884 17224 37936
rect 17276 37924 17282 37936
rect 17276 37896 22462 37924
rect 17276 37884 17282 37896
rect 12912 37828 19012 37856
rect 12805 37819 12863 37825
rect 10781 37791 10839 37797
rect 10781 37788 10793 37791
rect 10612 37760 10793 37788
rect 10226 37612 10232 37664
rect 10284 37652 10290 37664
rect 10612 37661 10640 37760
rect 10781 37757 10793 37760
rect 10827 37757 10839 37791
rect 11330 37788 11336 37800
rect 11291 37760 11336 37788
rect 10781 37751 10839 37757
rect 11330 37748 11336 37760
rect 11388 37748 11394 37800
rect 14252 37791 14310 37797
rect 14252 37757 14264 37791
rect 14298 37788 14310 37791
rect 14734 37788 14740 37800
rect 14298 37760 14740 37788
rect 14298 37757 14310 37760
rect 14252 37751 14310 37757
rect 14734 37748 14740 37760
rect 14792 37748 14798 37800
rect 15930 37748 15936 37800
rect 15988 37788 15994 37800
rect 16812 37791 16870 37797
rect 15988 37760 16033 37788
rect 15988 37748 15994 37760
rect 16812 37757 16824 37791
rect 16858 37788 16870 37791
rect 17218 37788 17224 37800
rect 16858 37760 17224 37788
rect 16858 37757 16870 37760
rect 16812 37751 16870 37757
rect 17218 37748 17224 37760
rect 17276 37748 17282 37800
rect 18984 37797 19012 37828
rect 18969 37791 19027 37797
rect 18969 37757 18981 37791
rect 19015 37788 19027 37791
rect 19334 37788 19340 37800
rect 19015 37760 19340 37788
rect 19015 37757 19027 37760
rect 18969 37751 19027 37757
rect 19334 37748 19340 37760
rect 19392 37748 19398 37800
rect 19521 37791 19579 37797
rect 19521 37757 19533 37791
rect 19567 37757 19579 37791
rect 19521 37751 19579 37757
rect 19797 37791 19855 37797
rect 19797 37757 19809 37791
rect 19843 37788 19855 37791
rect 20622 37788 20628 37800
rect 19843 37760 20628 37788
rect 19843 37757 19855 37760
rect 19797 37751 19855 37757
rect 11514 37720 11520 37732
rect 11475 37692 11520 37720
rect 11514 37680 11520 37692
rect 11572 37680 11578 37732
rect 12621 37723 12679 37729
rect 12621 37689 12633 37723
rect 12667 37689 12679 37723
rect 15013 37723 15071 37729
rect 15013 37720 15025 37723
rect 12621 37683 12679 37689
rect 13280 37692 15025 37720
rect 10597 37655 10655 37661
rect 10597 37652 10609 37655
rect 10284 37624 10609 37652
rect 10284 37612 10290 37624
rect 10597 37621 10609 37624
rect 10643 37621 10655 37655
rect 10597 37615 10655 37621
rect 11698 37612 11704 37664
rect 11756 37652 11762 37664
rect 11885 37655 11943 37661
rect 11885 37652 11897 37655
rect 11756 37624 11897 37652
rect 11756 37612 11762 37624
rect 11885 37621 11897 37624
rect 11931 37652 11943 37655
rect 11974 37652 11980 37664
rect 11931 37624 11980 37652
rect 11931 37621 11943 37624
rect 11885 37615 11943 37621
rect 11974 37612 11980 37624
rect 12032 37612 12038 37664
rect 12253 37655 12311 37661
rect 12253 37621 12265 37655
rect 12299 37652 12311 37655
rect 12342 37652 12348 37664
rect 12299 37624 12348 37652
rect 12299 37621 12311 37624
rect 12253 37615 12311 37621
rect 12342 37612 12348 37624
rect 12400 37652 12406 37664
rect 12636 37652 12664 37683
rect 13280 37652 13308 37692
rect 15013 37689 15025 37692
rect 15059 37689 15071 37723
rect 15286 37720 15292 37732
rect 15247 37692 15292 37720
rect 15013 37683 15071 37689
rect 14734 37652 14740 37664
rect 12400 37624 13308 37652
rect 14695 37624 14740 37652
rect 12400 37612 12406 37624
rect 14734 37612 14740 37624
rect 14792 37612 14798 37664
rect 15028 37652 15056 37683
rect 15286 37680 15292 37692
rect 15344 37680 15350 37732
rect 15381 37723 15439 37729
rect 15381 37689 15393 37723
rect 15427 37720 15439 37723
rect 15470 37720 15476 37732
rect 15427 37692 15476 37720
rect 15427 37689 15439 37692
rect 15381 37683 15439 37689
rect 15396 37652 15424 37683
rect 15470 37680 15476 37692
rect 15528 37680 15534 37732
rect 16942 37729 16948 37732
rect 16899 37723 16948 37729
rect 16899 37720 16911 37723
rect 16855 37692 16911 37720
rect 16899 37689 16911 37692
rect 16945 37689 16948 37723
rect 16899 37683 16948 37689
rect 16942 37680 16948 37683
rect 17000 37720 17006 37732
rect 17586 37720 17592 37732
rect 17000 37692 17592 37720
rect 17000 37680 17006 37692
rect 17586 37680 17592 37692
rect 17644 37680 17650 37732
rect 17865 37723 17923 37729
rect 17865 37689 17877 37723
rect 17911 37720 17923 37723
rect 19150 37720 19156 37732
rect 17911 37692 19156 37720
rect 17911 37689 17923 37692
rect 17865 37683 17923 37689
rect 19150 37680 19156 37692
rect 19208 37720 19214 37732
rect 19536 37720 19564 37751
rect 20622 37748 20628 37760
rect 20680 37748 20686 37800
rect 22434 37797 22462 37896
rect 24780 37856 24808 37952
rect 25130 37884 25136 37936
rect 25188 37924 25194 37936
rect 25188 37896 31202 37924
rect 25188 37884 25194 37896
rect 24688 37828 24808 37856
rect 22434 37791 22498 37797
rect 22434 37760 22452 37791
rect 22440 37757 22452 37760
rect 22486 37788 22498 37791
rect 22554 37788 22560 37800
rect 22486 37760 22560 37788
rect 22486 37757 22498 37760
rect 22440 37751 22498 37757
rect 22554 37748 22560 37760
rect 22612 37788 22618 37800
rect 22833 37791 22891 37797
rect 22833 37788 22845 37791
rect 22612 37760 22845 37788
rect 22612 37748 22618 37760
rect 22833 37757 22845 37760
rect 22879 37757 22891 37791
rect 22833 37751 22891 37757
rect 23728 37791 23786 37797
rect 23728 37757 23740 37791
rect 23774 37788 23786 37791
rect 23774 37760 24256 37788
rect 23774 37757 23786 37760
rect 23728 37751 23786 37757
rect 19208 37692 19564 37720
rect 19208 37680 19214 37692
rect 20714 37680 20720 37732
rect 20772 37720 20778 37732
rect 20946 37723 21004 37729
rect 20946 37720 20958 37723
rect 20772 37692 20958 37720
rect 20772 37680 20778 37692
rect 20946 37689 20958 37692
rect 20992 37689 21004 37723
rect 20946 37683 21004 37689
rect 16209 37655 16267 37661
rect 16209 37652 16221 37655
rect 15028 37624 16221 37652
rect 16209 37621 16221 37624
rect 16255 37652 16267 37655
rect 16577 37655 16635 37661
rect 16577 37652 16589 37655
rect 16255 37624 16589 37652
rect 16255 37621 16267 37624
rect 16209 37615 16267 37621
rect 16577 37621 16589 37624
rect 16623 37621 16635 37655
rect 16577 37615 16635 37621
rect 21545 37655 21603 37661
rect 21545 37621 21557 37655
rect 21591 37652 21603 37655
rect 21818 37652 21824 37664
rect 21591 37624 21824 37652
rect 21591 37621 21603 37624
rect 21545 37615 21603 37621
rect 21818 37612 21824 37624
rect 21876 37612 21882 37664
rect 23382 37612 23388 37664
rect 23440 37652 23446 37664
rect 24228 37661 24256 37760
rect 24688 37732 24716 37828
rect 26510 37816 26516 37868
rect 26568 37856 26574 37868
rect 28442 37856 28448 37868
rect 26568 37828 28448 37856
rect 26568 37816 26574 37828
rect 28442 37816 28448 37828
rect 28500 37816 28506 37868
rect 24762 37748 24768 37800
rect 24820 37788 24826 37800
rect 30024 37797 30052 37896
rect 30742 37856 30748 37868
rect 30703 37828 30748 37856
rect 30742 37816 30748 37828
rect 30800 37816 30806 37868
rect 31174 37856 31202 37896
rect 31662 37884 31668 37936
rect 31720 37924 31726 37936
rect 35713 37927 35771 37933
rect 31720 37896 35163 37924
rect 31720 37884 31726 37896
rect 31938 37856 31944 37868
rect 31174 37828 31944 37856
rect 31938 37816 31944 37828
rect 31996 37816 32002 37868
rect 32766 37856 32772 37868
rect 32727 37828 32772 37856
rect 32766 37816 32772 37828
rect 32824 37856 32830 37868
rect 33226 37856 33232 37868
rect 32824 37828 33232 37856
rect 32824 37816 32830 37828
rect 33226 37816 33232 37828
rect 33284 37816 33290 37868
rect 24857 37791 24915 37797
rect 24857 37788 24869 37791
rect 24820 37760 24869 37788
rect 24820 37748 24826 37760
rect 24857 37757 24869 37760
rect 24903 37788 24915 37791
rect 26053 37791 26111 37797
rect 26053 37788 26065 37791
rect 24903 37760 26065 37788
rect 24903 37757 24915 37760
rect 24857 37751 24915 37757
rect 26053 37757 26065 37760
rect 26099 37757 26111 37791
rect 26053 37751 26111 37757
rect 29917 37791 29975 37797
rect 29917 37757 29929 37791
rect 29963 37788 29975 37791
rect 30009 37791 30067 37797
rect 30009 37788 30021 37791
rect 29963 37760 30021 37788
rect 29963 37757 29975 37760
rect 29917 37751 29975 37757
rect 30009 37757 30021 37760
rect 30055 37757 30067 37791
rect 30009 37751 30067 37757
rect 30098 37748 30104 37800
rect 30156 37788 30162 37800
rect 30469 37791 30527 37797
rect 30469 37788 30481 37791
rect 30156 37760 30481 37788
rect 30156 37748 30162 37760
rect 30469 37757 30481 37760
rect 30515 37757 30527 37791
rect 30469 37751 30527 37757
rect 31732 37791 31790 37797
rect 31732 37757 31744 37791
rect 31778 37757 31790 37791
rect 31732 37751 31790 37757
rect 24670 37720 24676 37732
rect 24583 37692 24676 37720
rect 24670 37680 24676 37692
rect 24728 37720 24734 37732
rect 25178 37723 25236 37729
rect 25178 37720 25190 37723
rect 24728 37692 25190 37720
rect 24728 37680 24734 37692
rect 25178 37689 25190 37692
rect 25224 37720 25236 37723
rect 25498 37720 25504 37732
rect 25224 37692 25504 37720
rect 25224 37689 25236 37692
rect 25178 37683 25236 37689
rect 25498 37680 25504 37692
rect 25556 37680 25562 37732
rect 26789 37723 26847 37729
rect 26789 37689 26801 37723
rect 26835 37689 26847 37723
rect 26789 37683 26847 37689
rect 23799 37655 23857 37661
rect 23799 37652 23811 37655
rect 23440 37624 23811 37652
rect 23440 37612 23446 37624
rect 23799 37621 23811 37624
rect 23845 37621 23857 37655
rect 23799 37615 23857 37621
rect 24213 37655 24271 37661
rect 24213 37621 24225 37655
rect 24259 37652 24271 37655
rect 24302 37652 24308 37664
rect 24259 37624 24308 37652
rect 24259 37621 24271 37624
rect 24213 37615 24271 37621
rect 24302 37612 24308 37624
rect 24360 37612 24366 37664
rect 25777 37655 25835 37661
rect 25777 37621 25789 37655
rect 25823 37652 25835 37655
rect 26513 37655 26571 37661
rect 26513 37652 26525 37655
rect 25823 37624 26525 37652
rect 25823 37621 25835 37624
rect 25777 37615 25835 37621
rect 26513 37621 26525 37624
rect 26559 37652 26571 37655
rect 26602 37652 26608 37664
rect 26559 37624 26608 37652
rect 26559 37621 26571 37624
rect 26513 37615 26571 37621
rect 26602 37612 26608 37624
rect 26660 37612 26666 37664
rect 26694 37612 26700 37664
rect 26752 37652 26758 37664
rect 26804 37652 26832 37683
rect 26878 37680 26884 37732
rect 26936 37720 26942 37732
rect 27433 37723 27491 37729
rect 26936 37692 26981 37720
rect 26936 37680 26942 37692
rect 27433 37689 27445 37723
rect 27479 37720 27491 37723
rect 27798 37720 27804 37732
rect 27479 37692 27804 37720
rect 27479 37689 27491 37692
rect 27433 37683 27491 37689
rect 27798 37680 27804 37692
rect 27856 37680 27862 37732
rect 29730 37680 29736 37732
rect 29788 37720 29794 37732
rect 31747 37720 31775 37751
rect 32125 37723 32183 37729
rect 32125 37720 32137 37723
rect 29788 37692 32137 37720
rect 29788 37680 29794 37692
rect 32125 37689 32137 37692
rect 32171 37689 32183 37723
rect 32125 37683 32183 37689
rect 32858 37680 32864 37732
rect 32916 37720 32922 37732
rect 33410 37720 33416 37732
rect 32916 37692 32961 37720
rect 33371 37692 33416 37720
rect 32916 37680 32922 37692
rect 33410 37680 33416 37692
rect 33468 37680 33474 37732
rect 26752 37624 26832 37652
rect 31803 37655 31861 37661
rect 26752 37612 26758 37624
rect 31803 37621 31815 37655
rect 31849 37652 31861 37655
rect 32030 37652 32036 37664
rect 31849 37624 32036 37652
rect 31849 37621 31861 37624
rect 31803 37615 31861 37621
rect 32030 37612 32036 37624
rect 32088 37612 32094 37664
rect 35135 37652 35163 37896
rect 35713 37893 35725 37927
rect 35759 37924 35771 37927
rect 35802 37924 35808 37936
rect 35759 37896 35808 37924
rect 35759 37893 35771 37896
rect 35713 37887 35771 37893
rect 35802 37884 35808 37896
rect 35860 37924 35866 37936
rect 37829 37927 37887 37933
rect 37829 37924 37841 37927
rect 35860 37896 37841 37924
rect 35860 37884 35866 37896
rect 37829 37893 37841 37896
rect 37875 37924 37887 37927
rect 38102 37924 38108 37936
rect 37875 37896 38108 37924
rect 37875 37893 37887 37896
rect 37829 37887 37887 37893
rect 38102 37884 38108 37896
rect 38160 37924 38166 37936
rect 40034 37924 40040 37936
rect 38160 37896 40040 37924
rect 38160 37884 38166 37896
rect 40034 37884 40040 37896
rect 40092 37884 40098 37936
rect 42150 37884 42156 37936
rect 42208 37924 42214 37936
rect 42208 37896 42840 37924
rect 42208 37884 42214 37896
rect 35299 37859 35357 37865
rect 35299 37825 35311 37859
rect 35345 37856 35357 37859
rect 36265 37859 36323 37865
rect 36265 37856 36277 37859
rect 35345 37828 36277 37856
rect 35345 37825 35357 37828
rect 35299 37819 35357 37825
rect 36265 37825 36277 37828
rect 36311 37856 36323 37859
rect 36538 37856 36544 37868
rect 36311 37828 36544 37856
rect 36311 37825 36323 37828
rect 36265 37819 36323 37825
rect 36538 37816 36544 37828
rect 36596 37816 36602 37868
rect 38657 37859 38715 37865
rect 38657 37825 38669 37859
rect 38703 37856 38715 37859
rect 38930 37856 38936 37868
rect 38703 37828 38936 37856
rect 38703 37825 38715 37828
rect 38657 37819 38715 37825
rect 38930 37816 38936 37828
rect 38988 37816 38994 37868
rect 40954 37856 40960 37868
rect 40915 37828 40960 37856
rect 40954 37816 40960 37828
rect 41012 37816 41018 37868
rect 41230 37856 41236 37868
rect 41191 37828 41236 37856
rect 41230 37816 41236 37828
rect 41288 37816 41294 37868
rect 42812 37865 42840 37896
rect 42797 37859 42855 37865
rect 42797 37825 42809 37859
rect 42843 37825 42855 37859
rect 42797 37819 42855 37825
rect 35212 37791 35270 37797
rect 35212 37757 35224 37791
rect 35258 37788 35270 37791
rect 35986 37788 35992 37800
rect 35258 37760 35992 37788
rect 35258 37757 35270 37760
rect 35212 37751 35270 37757
rect 35986 37748 35992 37760
rect 36044 37748 36050 37800
rect 39574 37748 39580 37800
rect 39632 37788 39638 37800
rect 39669 37791 39727 37797
rect 39669 37788 39681 37791
rect 39632 37760 39681 37788
rect 39632 37748 39638 37760
rect 39669 37757 39681 37760
rect 39715 37788 39727 37791
rect 40678 37788 40684 37800
rect 39715 37760 40684 37788
rect 39715 37757 39727 37760
rect 39669 37751 39727 37757
rect 40678 37748 40684 37760
rect 40736 37748 40742 37800
rect 36357 37723 36415 37729
rect 36357 37689 36369 37723
rect 36403 37720 36415 37723
rect 36446 37720 36452 37732
rect 36403 37692 36452 37720
rect 36403 37689 36415 37692
rect 36357 37683 36415 37689
rect 36446 37680 36452 37692
rect 36504 37680 36510 37732
rect 36909 37723 36967 37729
rect 36909 37689 36921 37723
rect 36955 37720 36967 37723
rect 37182 37720 37188 37732
rect 36955 37692 37188 37720
rect 36955 37689 36967 37692
rect 36909 37683 36967 37689
rect 37182 37680 37188 37692
rect 37240 37680 37246 37732
rect 38749 37723 38807 37729
rect 38749 37689 38761 37723
rect 38795 37720 38807 37723
rect 38838 37720 38844 37732
rect 38795 37692 38844 37720
rect 38795 37689 38807 37692
rect 38749 37683 38807 37689
rect 38838 37680 38844 37692
rect 38896 37680 38902 37732
rect 39298 37720 39304 37732
rect 39259 37692 39304 37720
rect 39298 37680 39304 37692
rect 39356 37680 39362 37732
rect 39592 37652 39620 37748
rect 41046 37720 41052 37732
rect 40959 37692 41052 37720
rect 41046 37680 41052 37692
rect 41104 37680 41110 37732
rect 42518 37720 42524 37732
rect 42479 37692 42524 37720
rect 42518 37680 42524 37692
rect 42576 37680 42582 37732
rect 42613 37723 42671 37729
rect 42613 37689 42625 37723
rect 42659 37689 42671 37723
rect 42613 37683 42671 37689
rect 35135 37624 39620 37652
rect 40313 37655 40371 37661
rect 40313 37621 40325 37655
rect 40359 37652 40371 37655
rect 40681 37655 40739 37661
rect 40681 37652 40693 37655
rect 40359 37624 40693 37652
rect 40359 37621 40371 37624
rect 40313 37615 40371 37621
rect 40681 37621 40693 37624
rect 40727 37652 40739 37655
rect 40862 37652 40868 37664
rect 40727 37624 40868 37652
rect 40727 37621 40739 37624
rect 40681 37615 40739 37621
rect 40862 37612 40868 37624
rect 40920 37652 40926 37664
rect 41064 37652 41092 37680
rect 42245 37655 42303 37661
rect 42245 37652 42257 37655
rect 40920 37624 42257 37652
rect 40920 37612 40926 37624
rect 42245 37621 42257 37624
rect 42291 37652 42303 37655
rect 42628 37652 42656 37683
rect 42291 37624 42656 37652
rect 42291 37621 42303 37624
rect 42245 37615 42303 37621
rect 1104 37562 48852 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 48852 37562
rect 1104 37488 48852 37510
rect 10870 37448 10876 37460
rect 10783 37420 10876 37448
rect 10870 37408 10876 37420
rect 10928 37448 10934 37460
rect 11330 37448 11336 37460
rect 10928 37420 11336 37448
rect 10928 37408 10934 37420
rect 11330 37408 11336 37420
rect 11388 37408 11394 37460
rect 11514 37448 11520 37460
rect 11475 37420 11520 37448
rect 11514 37408 11520 37420
rect 11572 37408 11578 37460
rect 12526 37448 12532 37460
rect 11808 37420 12532 37448
rect 11195 37383 11253 37389
rect 11195 37349 11207 37383
rect 11241 37380 11253 37383
rect 11808 37380 11836 37420
rect 12526 37408 12532 37420
rect 12584 37408 12590 37460
rect 15286 37408 15292 37460
rect 15344 37448 15350 37460
rect 15427 37451 15485 37457
rect 15427 37448 15439 37451
rect 15344 37420 15439 37448
rect 15344 37408 15350 37420
rect 15427 37417 15439 37420
rect 15473 37448 15485 37451
rect 15749 37451 15807 37457
rect 15749 37448 15761 37451
rect 15473 37420 15761 37448
rect 15473 37417 15485 37420
rect 15427 37411 15485 37417
rect 15749 37417 15761 37420
rect 15795 37417 15807 37451
rect 15749 37411 15807 37417
rect 15838 37408 15844 37460
rect 15896 37448 15902 37460
rect 16117 37451 16175 37457
rect 16117 37448 16129 37451
rect 15896 37420 16129 37448
rect 15896 37408 15902 37420
rect 16117 37417 16129 37420
rect 16163 37417 16175 37451
rect 17586 37448 17592 37460
rect 17547 37420 17592 37448
rect 16117 37411 16175 37417
rect 17586 37408 17592 37420
rect 17644 37408 17650 37460
rect 20622 37448 20628 37460
rect 20583 37420 20628 37448
rect 20622 37408 20628 37420
rect 20680 37408 20686 37460
rect 25130 37448 25136 37460
rect 25091 37420 25136 37448
rect 25130 37408 25136 37420
rect 25188 37408 25194 37460
rect 25314 37408 25320 37460
rect 25372 37448 25378 37460
rect 25409 37451 25467 37457
rect 25409 37448 25421 37451
rect 25372 37420 25421 37448
rect 25372 37408 25378 37420
rect 25409 37417 25421 37420
rect 25455 37417 25467 37451
rect 25409 37411 25467 37417
rect 28994 37408 29000 37460
rect 29052 37448 29058 37460
rect 29549 37451 29607 37457
rect 29549 37448 29561 37451
rect 29052 37420 29561 37448
rect 29052 37408 29058 37420
rect 29549 37417 29561 37420
rect 29595 37448 29607 37451
rect 29638 37448 29644 37460
rect 29595 37420 29644 37448
rect 29595 37417 29607 37420
rect 29549 37411 29607 37417
rect 29638 37408 29644 37420
rect 29696 37408 29702 37460
rect 30006 37448 30012 37460
rect 29967 37420 30012 37448
rect 30006 37408 30012 37420
rect 30064 37408 30070 37460
rect 31570 37408 31576 37460
rect 31628 37448 31634 37460
rect 31849 37451 31907 37457
rect 31849 37448 31861 37451
rect 31628 37420 31861 37448
rect 31628 37408 31634 37420
rect 31849 37417 31861 37420
rect 31895 37417 31907 37451
rect 32490 37448 32496 37460
rect 32451 37420 32496 37448
rect 31849 37411 31907 37417
rect 32490 37408 32496 37420
rect 32548 37408 32554 37460
rect 33226 37408 33232 37460
rect 33284 37448 33290 37460
rect 33321 37451 33379 37457
rect 33321 37448 33333 37451
rect 33284 37420 33333 37448
rect 33284 37408 33290 37420
rect 33321 37417 33333 37420
rect 33367 37417 33379 37451
rect 35250 37448 35256 37460
rect 35211 37420 35256 37448
rect 33321 37411 33379 37417
rect 35250 37408 35256 37420
rect 35308 37448 35314 37460
rect 35529 37451 35587 37457
rect 35529 37448 35541 37451
rect 35308 37420 35541 37448
rect 35308 37408 35314 37420
rect 35529 37417 35541 37420
rect 35575 37417 35587 37451
rect 36446 37448 36452 37460
rect 36407 37420 36452 37448
rect 35529 37411 35587 37417
rect 36446 37408 36452 37420
rect 36504 37408 36510 37460
rect 40862 37448 40868 37460
rect 40823 37420 40868 37448
rect 40862 37408 40868 37420
rect 40920 37408 40926 37460
rect 40954 37408 40960 37460
rect 41012 37448 41018 37460
rect 41141 37451 41199 37457
rect 41141 37448 41153 37451
rect 41012 37420 41153 37448
rect 41012 37408 41018 37420
rect 41141 37417 41153 37420
rect 41187 37417 41199 37451
rect 41141 37411 41199 37417
rect 11241 37352 11836 37380
rect 11241 37349 11253 37352
rect 11195 37343 11253 37349
rect 12158 37340 12164 37392
rect 12216 37380 12222 37392
rect 12253 37383 12311 37389
rect 12253 37380 12265 37383
rect 12216 37352 12265 37380
rect 12216 37340 12222 37352
rect 12253 37349 12265 37352
rect 12299 37349 12311 37383
rect 12253 37343 12311 37349
rect 14274 37340 14280 37392
rect 14332 37380 14338 37392
rect 17218 37380 17224 37392
rect 14332 37352 17224 37380
rect 14332 37340 14338 37352
rect 17218 37340 17224 37352
rect 17276 37340 17282 37392
rect 21818 37340 21824 37392
rect 21876 37380 21882 37392
rect 21913 37383 21971 37389
rect 21913 37380 21925 37383
rect 21876 37352 21925 37380
rect 21876 37340 21882 37352
rect 21913 37349 21925 37352
rect 21959 37349 21971 37383
rect 21913 37343 21971 37349
rect 22465 37383 22523 37389
rect 22465 37349 22477 37383
rect 22511 37380 22523 37383
rect 23658 37380 23664 37392
rect 22511 37352 23664 37380
rect 22511 37349 22523 37352
rect 22465 37343 22523 37349
rect 23658 37340 23664 37352
rect 23716 37340 23722 37392
rect 24762 37380 24768 37392
rect 24723 37352 24768 37380
rect 24762 37340 24768 37352
rect 24820 37340 24826 37392
rect 11108 37315 11166 37321
rect 11108 37281 11120 37315
rect 11154 37281 11166 37315
rect 11108 37275 11166 37281
rect 11123 37244 11151 37275
rect 13446 37272 13452 37324
rect 13504 37312 13510 37324
rect 13668 37315 13726 37321
rect 13668 37312 13680 37315
rect 13504 37284 13680 37312
rect 13504 37272 13510 37284
rect 13668 37281 13680 37284
rect 13714 37281 13726 37315
rect 13668 37275 13726 37281
rect 15356 37315 15414 37321
rect 15356 37281 15368 37315
rect 15402 37312 15414 37315
rect 16022 37312 16028 37324
rect 15402 37284 16028 37312
rect 15402 37281 15414 37284
rect 15356 37275 15414 37281
rect 16022 37272 16028 37284
rect 16080 37272 16086 37324
rect 16482 37272 16488 37324
rect 16540 37312 16546 37324
rect 16577 37315 16635 37321
rect 16577 37312 16589 37315
rect 16540 37284 16589 37312
rect 16540 37272 16546 37284
rect 16577 37281 16589 37284
rect 16623 37281 16635 37315
rect 16577 37275 16635 37281
rect 17034 37272 17040 37324
rect 17092 37312 17098 37324
rect 17129 37315 17187 37321
rect 17129 37312 17141 37315
rect 17092 37284 17141 37312
rect 17092 37272 17098 37284
rect 17129 37281 17141 37284
rect 17175 37312 17187 37315
rect 17175 37284 18092 37312
rect 17175 37281 17187 37284
rect 17129 37275 17187 37281
rect 11238 37244 11244 37256
rect 11123 37216 11244 37244
rect 11238 37204 11244 37216
rect 11296 37204 11302 37256
rect 12158 37244 12164 37256
rect 12119 37216 12164 37244
rect 12158 37204 12164 37216
rect 12216 37204 12222 37256
rect 12618 37244 12624 37256
rect 12579 37216 12624 37244
rect 12618 37204 12624 37216
rect 12676 37204 12682 37256
rect 17310 37244 17316 37256
rect 17271 37216 17316 37244
rect 17310 37204 17316 37216
rect 17368 37204 17374 37256
rect 18064 37244 18092 37284
rect 18138 37272 18144 37324
rect 18196 37312 18202 37324
rect 18601 37315 18659 37321
rect 18601 37312 18613 37315
rect 18196 37284 18241 37312
rect 18524 37284 18613 37312
rect 18196 37272 18202 37284
rect 18524 37244 18552 37284
rect 18601 37281 18613 37284
rect 18647 37281 18659 37315
rect 19832 37315 19890 37321
rect 19832 37312 19844 37315
rect 18601 37275 18659 37281
rect 19720 37284 19844 37312
rect 19720 37256 19748 37284
rect 19832 37281 19844 37284
rect 19878 37281 19890 37315
rect 24026 37312 24032 37324
rect 23987 37284 24032 37312
rect 19832 37275 19890 37281
rect 24026 37272 24032 37284
rect 24084 37272 24090 37324
rect 24578 37312 24584 37324
rect 24491 37284 24584 37312
rect 24578 37272 24584 37284
rect 24636 37312 24642 37324
rect 25332 37312 25360 37408
rect 26786 37340 26792 37392
rect 26844 37380 26850 37392
rect 27065 37383 27123 37389
rect 27065 37380 27077 37383
rect 26844 37352 27077 37380
rect 26844 37340 26850 37352
rect 27065 37349 27077 37352
rect 27111 37349 27123 37383
rect 28626 37380 28632 37392
rect 28587 37352 28632 37380
rect 27065 37343 27123 37349
rect 28626 37340 28632 37352
rect 28684 37340 28690 37392
rect 30024 37380 30052 37408
rect 30024 37352 30880 37380
rect 30852 37324 30880 37352
rect 31386 37340 31392 37392
rect 31444 37380 31450 37392
rect 31481 37383 31539 37389
rect 31481 37380 31493 37383
rect 31444 37352 31493 37380
rect 31444 37340 31450 37352
rect 31481 37349 31493 37352
rect 31527 37380 31539 37383
rect 32306 37380 32312 37392
rect 31527 37352 32312 37380
rect 31527 37349 31539 37352
rect 31481 37343 31539 37349
rect 32306 37340 32312 37352
rect 32364 37340 32370 37392
rect 34057 37383 34115 37389
rect 34057 37380 34069 37383
rect 33612 37352 34069 37380
rect 24636 37284 25360 37312
rect 30653 37315 30711 37321
rect 24636 37272 24642 37284
rect 30653 37281 30665 37315
rect 30699 37312 30711 37315
rect 30742 37312 30748 37324
rect 30699 37284 30748 37312
rect 30699 37281 30711 37284
rect 30653 37275 30711 37281
rect 30742 37272 30748 37284
rect 30800 37272 30806 37324
rect 30834 37272 30840 37324
rect 30892 37312 30898 37324
rect 30892 37284 30985 37312
rect 30892 37272 30898 37284
rect 32674 37272 32680 37324
rect 32732 37312 32738 37324
rect 33045 37315 33103 37321
rect 33045 37312 33057 37315
rect 32732 37284 33057 37312
rect 32732 37272 32738 37284
rect 33045 37281 33057 37284
rect 33091 37312 33103 37315
rect 33612 37312 33640 37352
rect 34057 37349 34069 37352
rect 34103 37349 34115 37383
rect 34057 37343 34115 37349
rect 40034 37340 40040 37392
rect 40092 37380 40098 37392
rect 40266 37383 40324 37389
rect 40266 37380 40278 37383
rect 40092 37352 40278 37380
rect 40092 37340 40098 37352
rect 40266 37349 40278 37352
rect 40312 37349 40324 37383
rect 40880 37380 40908 37408
rect 41598 37380 41604 37392
rect 40880 37352 41604 37380
rect 40266 37343 40324 37349
rect 41598 37340 41604 37352
rect 41656 37380 41662 37392
rect 41877 37383 41935 37389
rect 41877 37380 41889 37383
rect 41656 37352 41889 37380
rect 41656 37340 41662 37352
rect 41877 37349 41889 37352
rect 41923 37349 41935 37383
rect 41877 37343 41935 37349
rect 35710 37312 35716 37324
rect 33091 37284 33640 37312
rect 35671 37284 35716 37312
rect 33091 37281 33103 37284
rect 33045 37275 33103 37281
rect 35710 37272 35716 37284
rect 35768 37272 35774 37324
rect 35894 37312 35900 37324
rect 35855 37284 35900 37312
rect 35894 37272 35900 37284
rect 35952 37272 35958 37324
rect 38381 37315 38439 37321
rect 38381 37281 38393 37315
rect 38427 37281 38439 37315
rect 38838 37312 38844 37324
rect 38799 37284 38844 37312
rect 38381 37275 38439 37281
rect 18690 37244 18696 37256
rect 18064 37216 18552 37244
rect 18651 37216 18696 37244
rect 13771 37111 13829 37117
rect 13771 37077 13783 37111
rect 13817 37108 13829 37111
rect 14366 37108 14372 37120
rect 13817 37080 14372 37108
rect 13817 37077 13829 37080
rect 13771 37071 13829 37077
rect 14366 37068 14372 37080
rect 14424 37068 14430 37120
rect 18414 37068 18420 37120
rect 18472 37108 18478 37120
rect 18524 37108 18552 37216
rect 18690 37204 18696 37216
rect 18748 37244 18754 37256
rect 19521 37247 19579 37253
rect 19521 37244 19533 37247
rect 18748 37216 19533 37244
rect 18748 37204 18754 37216
rect 19521 37213 19533 37216
rect 19567 37213 19579 37247
rect 19521 37207 19579 37213
rect 19702 37204 19708 37256
rect 19760 37204 19766 37256
rect 21821 37247 21879 37253
rect 21821 37213 21833 37247
rect 21867 37244 21879 37247
rect 23382 37244 23388 37256
rect 21867 37216 23388 37244
rect 21867 37213 21879 37216
rect 21821 37207 21879 37213
rect 23382 37204 23388 37216
rect 23440 37204 23446 37256
rect 26970 37244 26976 37256
rect 26931 37216 26976 37244
rect 26970 37204 26976 37216
rect 27028 37204 27034 37256
rect 27246 37244 27252 37256
rect 27207 37216 27252 37244
rect 27246 37204 27252 37216
rect 27304 37204 27310 37256
rect 28534 37244 28540 37256
rect 28495 37216 28540 37244
rect 28534 37204 28540 37216
rect 28592 37204 28598 37256
rect 28810 37244 28816 37256
rect 28771 37216 28816 37244
rect 28810 37204 28816 37216
rect 28868 37204 28874 37256
rect 31113 37247 31171 37253
rect 31113 37213 31125 37247
rect 31159 37244 31171 37247
rect 32125 37247 32183 37253
rect 32125 37244 32137 37247
rect 31159 37216 32137 37244
rect 31159 37213 31171 37216
rect 31113 37207 31171 37213
rect 32125 37213 32137 37216
rect 32171 37244 32183 37247
rect 32306 37244 32312 37256
rect 32171 37216 32312 37244
rect 32171 37213 32183 37216
rect 32125 37207 32183 37213
rect 32306 37204 32312 37216
rect 32364 37204 32370 37256
rect 33778 37204 33784 37256
rect 33836 37244 33842 37256
rect 33965 37247 34023 37253
rect 33965 37244 33977 37247
rect 33836 37216 33977 37244
rect 33836 37204 33842 37216
rect 33965 37213 33977 37216
rect 34011 37213 34023 37247
rect 34238 37244 34244 37256
rect 34199 37216 34244 37244
rect 33965 37207 34023 37213
rect 34238 37204 34244 37216
rect 34296 37204 34302 37256
rect 19935 37179 19993 37185
rect 19935 37145 19947 37179
rect 19981 37176 19993 37179
rect 23198 37176 23204 37188
rect 19981 37148 23204 37176
rect 19981 37145 19993 37148
rect 19935 37139 19993 37145
rect 23198 37136 23204 37148
rect 23256 37176 23262 37188
rect 23293 37179 23351 37185
rect 23293 37176 23305 37179
rect 23256 37148 23305 37176
rect 23256 37136 23262 37148
rect 23293 37145 23305 37148
rect 23339 37145 23351 37179
rect 23293 37139 23351 37145
rect 31570 37136 31576 37188
rect 31628 37176 31634 37188
rect 38396 37176 38424 37275
rect 38838 37272 38844 37284
rect 38896 37272 38902 37324
rect 39117 37247 39175 37253
rect 39117 37213 39129 37247
rect 39163 37244 39175 37247
rect 39945 37247 40003 37253
rect 39945 37244 39957 37247
rect 39163 37216 39957 37244
rect 39163 37213 39175 37216
rect 39117 37207 39175 37213
rect 39945 37213 39957 37216
rect 39991 37244 40003 37247
rect 40126 37244 40132 37256
rect 39991 37216 40132 37244
rect 39991 37213 40003 37216
rect 39945 37207 40003 37213
rect 40126 37204 40132 37216
rect 40184 37204 40190 37256
rect 41782 37244 41788 37256
rect 41743 37216 41788 37244
rect 41782 37204 41788 37216
rect 41840 37204 41846 37256
rect 42429 37247 42487 37253
rect 42429 37213 42441 37247
rect 42475 37244 42487 37247
rect 42610 37244 42616 37256
rect 42475 37216 42616 37244
rect 42475 37213 42487 37216
rect 42429 37207 42487 37213
rect 42610 37204 42616 37216
rect 42668 37204 42674 37256
rect 39022 37176 39028 37188
rect 31628 37148 39028 37176
rect 31628 37136 31634 37148
rect 39022 37136 39028 37148
rect 39080 37136 39086 37188
rect 19150 37108 19156 37120
rect 18472 37080 19156 37108
rect 18472 37068 18478 37080
rect 19150 37068 19156 37080
rect 19208 37068 19214 37120
rect 19242 37068 19248 37120
rect 19300 37108 19306 37120
rect 21726 37108 21732 37120
rect 19300 37080 21732 37108
rect 19300 37068 19306 37080
rect 21726 37068 21732 37080
rect 21784 37108 21790 37120
rect 24762 37108 24768 37120
rect 21784 37080 24768 37108
rect 21784 37068 21790 37080
rect 24762 37068 24768 37080
rect 24820 37068 24826 37120
rect 26694 37108 26700 37120
rect 26655 37080 26700 37108
rect 26694 37068 26700 37080
rect 26752 37068 26758 37120
rect 33686 37108 33692 37120
rect 33647 37080 33692 37108
rect 33686 37068 33692 37080
rect 33744 37068 33750 37120
rect 36814 37108 36820 37120
rect 36775 37080 36820 37108
rect 36814 37068 36820 37080
rect 36872 37068 36878 37120
rect 1104 37018 48852 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 48852 37018
rect 1104 36944 48852 36966
rect 12158 36904 12164 36916
rect 11348 36876 12164 36904
rect 11348 36777 11376 36876
rect 12158 36864 12164 36876
rect 12216 36864 12222 36916
rect 13446 36904 13452 36916
rect 13407 36876 13452 36904
rect 13446 36864 13452 36876
rect 13504 36864 13510 36916
rect 16022 36864 16028 36916
rect 16080 36904 16086 36916
rect 16117 36907 16175 36913
rect 16117 36904 16129 36907
rect 16080 36876 16129 36904
rect 16080 36864 16086 36876
rect 16117 36873 16129 36876
rect 16163 36873 16175 36907
rect 17034 36904 17040 36916
rect 16995 36876 17040 36904
rect 16117 36867 16175 36873
rect 17034 36864 17040 36876
rect 17092 36864 17098 36916
rect 18601 36907 18659 36913
rect 18601 36873 18613 36907
rect 18647 36904 18659 36907
rect 18782 36904 18788 36916
rect 18647 36876 18788 36904
rect 18647 36873 18659 36876
rect 18601 36867 18659 36873
rect 18782 36864 18788 36876
rect 18840 36864 18846 36916
rect 19702 36864 19708 36916
rect 19760 36904 19766 36916
rect 19889 36907 19947 36913
rect 19889 36904 19901 36907
rect 19760 36876 19901 36904
rect 19760 36864 19766 36876
rect 19889 36873 19901 36876
rect 19935 36873 19947 36907
rect 21818 36904 21824 36916
rect 21779 36876 21824 36904
rect 19889 36867 19947 36873
rect 13081 36839 13139 36845
rect 13081 36805 13093 36839
rect 13127 36836 13139 36839
rect 13262 36836 13268 36848
rect 13127 36808 13268 36836
rect 13127 36805 13139 36808
rect 13081 36799 13139 36805
rect 11333 36771 11391 36777
rect 11333 36737 11345 36771
rect 11379 36737 11391 36771
rect 11333 36731 11391 36737
rect 12596 36703 12654 36709
rect 12596 36669 12608 36703
rect 12642 36700 12654 36703
rect 13096 36700 13124 36799
rect 13262 36796 13268 36808
rect 13320 36836 13326 36848
rect 15749 36839 15807 36845
rect 13320 36808 13952 36836
rect 13320 36796 13326 36808
rect 13633 36771 13691 36777
rect 13633 36737 13645 36771
rect 13679 36768 13691 36771
rect 13814 36768 13820 36780
rect 13679 36740 13820 36768
rect 13679 36737 13691 36740
rect 13633 36731 13691 36737
rect 13814 36728 13820 36740
rect 13872 36728 13878 36780
rect 13924 36777 13952 36808
rect 15749 36805 15761 36839
rect 15795 36836 15807 36839
rect 15930 36836 15936 36848
rect 15795 36808 15936 36836
rect 15795 36805 15807 36808
rect 15749 36799 15807 36805
rect 15930 36796 15936 36808
rect 15988 36796 15994 36848
rect 19904 36836 19932 36867
rect 21818 36864 21824 36876
rect 21876 36864 21882 36916
rect 22925 36907 22983 36913
rect 22925 36873 22937 36907
rect 22971 36904 22983 36907
rect 23382 36904 23388 36916
rect 22971 36876 23388 36904
rect 22971 36873 22983 36876
rect 22925 36867 22983 36873
rect 23382 36864 23388 36876
rect 23440 36864 23446 36916
rect 24026 36864 24032 36916
rect 24084 36904 24090 36916
rect 24489 36907 24547 36913
rect 24489 36904 24501 36907
rect 24084 36876 24501 36904
rect 24084 36864 24090 36876
rect 24489 36873 24501 36876
rect 24535 36873 24547 36907
rect 24489 36867 24547 36873
rect 25915 36907 25973 36913
rect 25915 36873 25927 36907
rect 25961 36904 25973 36907
rect 26694 36904 26700 36916
rect 25961 36876 26700 36904
rect 25961 36873 25973 36876
rect 25915 36867 25973 36873
rect 26694 36864 26700 36876
rect 26752 36864 26758 36916
rect 30834 36864 30840 36916
rect 30892 36904 30898 36916
rect 31113 36907 31171 36913
rect 31113 36904 31125 36907
rect 30892 36876 31125 36904
rect 30892 36864 30898 36876
rect 31113 36873 31125 36876
rect 31159 36873 31171 36907
rect 32674 36904 32680 36916
rect 32635 36876 32680 36904
rect 31113 36867 31171 36873
rect 32674 36864 32680 36876
rect 32732 36864 32738 36916
rect 33778 36864 33784 36916
rect 33836 36904 33842 36916
rect 34241 36907 34299 36913
rect 34241 36904 34253 36907
rect 33836 36876 34253 36904
rect 33836 36864 33842 36876
rect 34241 36873 34253 36876
rect 34287 36873 34299 36907
rect 37458 36904 37464 36916
rect 34241 36867 34299 36873
rect 36372 36876 37464 36904
rect 26510 36836 26516 36848
rect 19904 36808 26516 36836
rect 26510 36796 26516 36808
rect 26568 36796 26574 36848
rect 26605 36839 26663 36845
rect 26605 36805 26617 36839
rect 26651 36836 26663 36839
rect 26786 36836 26792 36848
rect 26651 36808 26792 36836
rect 26651 36805 26663 36808
rect 26605 36799 26663 36805
rect 26786 36796 26792 36808
rect 26844 36836 26850 36848
rect 27062 36836 27068 36848
rect 26844 36808 27068 36836
rect 26844 36796 26850 36808
rect 27062 36796 27068 36808
rect 27120 36836 27126 36848
rect 28445 36839 28503 36845
rect 28445 36836 28457 36839
rect 27120 36808 28457 36836
rect 27120 36796 27126 36808
rect 28445 36805 28457 36808
rect 28491 36836 28503 36839
rect 28626 36836 28632 36848
rect 28491 36808 28632 36836
rect 28491 36805 28503 36808
rect 28445 36799 28503 36805
rect 28626 36796 28632 36808
rect 28684 36796 28690 36848
rect 32214 36836 32220 36848
rect 29794 36808 32220 36836
rect 13909 36771 13967 36777
rect 13909 36737 13921 36771
rect 13955 36768 13967 36771
rect 16758 36768 16764 36780
rect 13955 36740 16764 36768
rect 13955 36737 13967 36740
rect 13909 36731 13967 36737
rect 16758 36728 16764 36740
rect 16816 36728 16822 36780
rect 18690 36768 18696 36780
rect 18651 36740 18696 36768
rect 18690 36728 18696 36740
rect 18748 36728 18754 36780
rect 20530 36768 20536 36780
rect 20491 36740 20536 36768
rect 20530 36728 20536 36740
rect 20588 36728 20594 36780
rect 22554 36728 22560 36780
rect 22612 36768 22618 36780
rect 25133 36771 25191 36777
rect 25133 36768 25145 36771
rect 22612 36740 25145 36768
rect 22612 36728 22618 36740
rect 25133 36737 25145 36740
rect 25179 36737 25191 36771
rect 25133 36731 25191 36737
rect 25317 36771 25375 36777
rect 25317 36737 25329 36771
rect 25363 36768 25375 36771
rect 29794 36768 29822 36808
rect 32214 36796 32220 36808
rect 32272 36796 32278 36848
rect 33410 36796 33416 36848
rect 33468 36836 33474 36848
rect 33505 36839 33563 36845
rect 33505 36836 33517 36839
rect 33468 36808 33517 36836
rect 33468 36796 33474 36808
rect 33505 36805 33517 36808
rect 33551 36805 33563 36839
rect 33505 36799 33563 36805
rect 31386 36768 31392 36780
rect 25363 36740 29822 36768
rect 31347 36740 31392 36768
rect 25363 36737 25375 36740
rect 25317 36731 25375 36737
rect 12642 36672 13124 36700
rect 19613 36703 19671 36709
rect 12642 36669 12654 36672
rect 12596 36663 12654 36669
rect 19613 36669 19625 36703
rect 19659 36700 19671 36703
rect 20257 36703 20315 36709
rect 20257 36700 20269 36703
rect 19659 36672 20269 36700
rect 19659 36669 19671 36672
rect 19613 36663 19671 36669
rect 20257 36669 20269 36672
rect 20303 36669 20315 36703
rect 20257 36663 20315 36669
rect 13722 36632 13728 36644
rect 13683 36604 13728 36632
rect 13722 36592 13728 36604
rect 13780 36592 13786 36644
rect 14645 36635 14703 36641
rect 14645 36601 14657 36635
rect 14691 36632 14703 36635
rect 15194 36632 15200 36644
rect 14691 36604 15200 36632
rect 14691 36601 14703 36604
rect 14645 36595 14703 36601
rect 15194 36592 15200 36604
rect 15252 36592 15258 36644
rect 15289 36635 15347 36641
rect 15289 36601 15301 36635
rect 15335 36601 15347 36635
rect 15289 36595 15347 36601
rect 11149 36567 11207 36573
rect 11149 36533 11161 36567
rect 11195 36564 11207 36567
rect 11238 36564 11244 36576
rect 11195 36536 11244 36564
rect 11195 36533 11207 36536
rect 11149 36527 11207 36533
rect 11238 36524 11244 36536
rect 11296 36524 11302 36576
rect 11606 36524 11612 36576
rect 11664 36564 11670 36576
rect 12667 36567 12725 36573
rect 12667 36564 12679 36567
rect 11664 36536 12679 36564
rect 11664 36524 11670 36536
rect 12667 36533 12679 36536
rect 12713 36533 12725 36567
rect 12667 36527 12725 36533
rect 14458 36524 14464 36576
rect 14516 36564 14522 36576
rect 15013 36567 15071 36573
rect 15013 36564 15025 36567
rect 14516 36536 15025 36564
rect 14516 36524 14522 36536
rect 15013 36533 15025 36536
rect 15059 36564 15071 36567
rect 15304 36564 15332 36595
rect 18782 36592 18788 36644
rect 18840 36632 18846 36644
rect 19014 36635 19072 36641
rect 19014 36632 19026 36635
rect 18840 36604 19026 36632
rect 18840 36592 18846 36604
rect 19014 36601 19026 36604
rect 19060 36601 19072 36635
rect 19014 36595 19072 36601
rect 15059 36536 15332 36564
rect 15059 36533 15071 36536
rect 15013 36527 15071 36533
rect 16482 36524 16488 36576
rect 16540 36564 16546 36576
rect 16577 36567 16635 36573
rect 16577 36564 16589 36567
rect 16540 36536 16589 36564
rect 16540 36524 16546 36536
rect 16577 36533 16589 36536
rect 16623 36533 16635 36567
rect 16577 36527 16635 36533
rect 17402 36524 17408 36576
rect 17460 36564 17466 36576
rect 17773 36567 17831 36573
rect 17773 36564 17785 36567
rect 17460 36536 17785 36564
rect 17460 36524 17466 36536
rect 17773 36533 17785 36536
rect 17819 36564 17831 36567
rect 18138 36564 18144 36576
rect 17819 36536 18144 36564
rect 17819 36533 17831 36536
rect 17773 36527 17831 36533
rect 18138 36524 18144 36536
rect 18196 36524 18202 36576
rect 20272 36564 20300 36663
rect 21726 36660 21732 36712
rect 21784 36700 21790 36712
rect 22040 36703 22098 36709
rect 22040 36700 22052 36703
rect 21784 36672 22052 36700
rect 21784 36660 21790 36672
rect 22040 36669 22052 36672
rect 22086 36700 22098 36703
rect 22465 36703 22523 36709
rect 22465 36700 22477 36703
rect 22086 36672 22477 36700
rect 22086 36669 22098 36672
rect 22040 36663 22098 36669
rect 22465 36669 22477 36672
rect 22511 36669 22523 36703
rect 22465 36663 22523 36669
rect 23290 36660 23296 36712
rect 23348 36700 23354 36712
rect 23728 36703 23786 36709
rect 23728 36700 23740 36703
rect 23348 36672 23740 36700
rect 23348 36660 23354 36672
rect 23728 36669 23740 36672
rect 23774 36700 23786 36703
rect 24121 36703 24179 36709
rect 24121 36700 24133 36703
rect 23774 36672 24133 36700
rect 23774 36669 23786 36672
rect 23728 36663 23786 36669
rect 24121 36669 24133 36672
rect 24167 36669 24179 36703
rect 24121 36663 24179 36669
rect 24302 36660 24308 36712
rect 24360 36700 24366 36712
rect 24816 36703 24874 36709
rect 24816 36700 24828 36703
rect 24360 36672 24828 36700
rect 24360 36660 24366 36672
rect 24816 36669 24828 36672
rect 24862 36700 24874 36703
rect 25332 36700 25360 36731
rect 31386 36728 31392 36740
rect 31444 36728 31450 36780
rect 31662 36768 31668 36780
rect 31623 36740 31668 36768
rect 31662 36728 31668 36740
rect 31720 36728 31726 36780
rect 32950 36768 32956 36780
rect 32863 36740 32956 36768
rect 32950 36728 32956 36740
rect 33008 36768 33014 36780
rect 33686 36768 33692 36780
rect 33008 36740 33692 36768
rect 33008 36728 33014 36740
rect 33686 36728 33692 36740
rect 33744 36728 33750 36780
rect 35894 36768 35900 36780
rect 35452 36740 35900 36768
rect 35452 36712 35480 36740
rect 35894 36728 35900 36740
rect 35952 36768 35958 36780
rect 36372 36777 36400 36876
rect 37458 36864 37464 36876
rect 37516 36904 37522 36916
rect 38013 36907 38071 36913
rect 38013 36904 38025 36907
rect 37516 36876 38025 36904
rect 37516 36864 37522 36876
rect 38013 36873 38025 36876
rect 38059 36873 38071 36907
rect 38013 36867 38071 36873
rect 38335 36907 38393 36913
rect 38335 36873 38347 36907
rect 38381 36904 38393 36907
rect 38930 36904 38936 36916
rect 38381 36876 38936 36904
rect 38381 36873 38393 36876
rect 38335 36867 38393 36873
rect 36998 36836 37004 36848
rect 36648 36808 37004 36836
rect 36648 36777 36676 36808
rect 36998 36796 37004 36808
rect 37056 36796 37062 36848
rect 38028 36836 38056 36867
rect 38930 36864 38936 36876
rect 38988 36864 38994 36916
rect 39022 36864 39028 36916
rect 39080 36904 39086 36916
rect 41598 36904 41604 36916
rect 39080 36876 39125 36904
rect 41559 36876 41604 36904
rect 39080 36864 39086 36876
rect 41598 36864 41604 36876
rect 41656 36864 41662 36916
rect 41923 36907 41981 36913
rect 41923 36873 41935 36907
rect 41969 36904 41981 36907
rect 42518 36904 42524 36916
rect 41969 36876 42524 36904
rect 41969 36873 41981 36876
rect 41923 36867 41981 36873
rect 42518 36864 42524 36876
rect 42576 36864 42582 36916
rect 38838 36836 38844 36848
rect 38028 36808 38844 36836
rect 38838 36796 38844 36808
rect 38896 36796 38902 36848
rect 40911 36839 40969 36845
rect 40911 36805 40923 36839
rect 40957 36836 40969 36839
rect 41782 36836 41788 36848
rect 40957 36808 41788 36836
rect 40957 36805 40969 36808
rect 40911 36799 40969 36805
rect 41782 36796 41788 36808
rect 41840 36796 41846 36848
rect 36357 36771 36415 36777
rect 36357 36768 36369 36771
rect 35952 36740 36369 36768
rect 35952 36728 35958 36740
rect 36357 36737 36369 36740
rect 36403 36737 36415 36771
rect 36357 36731 36415 36737
rect 36633 36771 36691 36777
rect 36633 36737 36645 36771
rect 36679 36737 36691 36771
rect 36906 36768 36912 36780
rect 36867 36740 36912 36768
rect 36633 36731 36691 36737
rect 36906 36728 36912 36740
rect 36964 36728 36970 36780
rect 37274 36728 37280 36780
rect 37332 36768 37338 36780
rect 37332 36740 38367 36768
rect 37332 36728 37338 36740
rect 24862 36672 25360 36700
rect 25844 36703 25902 36709
rect 24862 36669 24874 36672
rect 24816 36663 24874 36669
rect 25844 36669 25856 36703
rect 25890 36700 25902 36703
rect 26053 36703 26111 36709
rect 26053 36700 26065 36703
rect 25890 36672 26065 36700
rect 25890 36669 25902 36672
rect 25844 36663 25902 36669
rect 26053 36669 26065 36672
rect 26099 36669 26111 36703
rect 26053 36663 26111 36669
rect 27522 36660 27528 36712
rect 27580 36700 27586 36712
rect 29549 36703 29607 36709
rect 27580 36672 27625 36700
rect 27580 36660 27586 36672
rect 29549 36669 29561 36703
rect 29595 36669 29607 36703
rect 34698 36700 34704 36712
rect 34611 36672 34704 36700
rect 29549 36663 29607 36669
rect 20625 36635 20683 36641
rect 20625 36601 20637 36635
rect 20671 36601 20683 36635
rect 21174 36632 21180 36644
rect 21135 36604 21180 36632
rect 20625 36595 20683 36601
rect 20640 36564 20668 36595
rect 21174 36592 21180 36604
rect 21232 36592 21238 36644
rect 23106 36592 23112 36644
rect 23164 36632 23170 36644
rect 23385 36635 23443 36641
rect 23385 36632 23397 36635
rect 23164 36604 23397 36632
rect 23164 36592 23170 36604
rect 23385 36601 23397 36604
rect 23431 36632 23443 36635
rect 24210 36632 24216 36644
rect 23431 36604 24216 36632
rect 23431 36601 23443 36604
rect 23385 36595 23443 36601
rect 24210 36592 24216 36604
rect 24268 36632 24274 36644
rect 24578 36632 24584 36644
rect 24268 36604 24584 36632
rect 24268 36592 24274 36604
rect 24578 36592 24584 36604
rect 24636 36592 24642 36644
rect 24903 36635 24961 36641
rect 24903 36601 24915 36635
rect 24949 36632 24961 36635
rect 26881 36635 26939 36641
rect 26881 36632 26893 36635
rect 24949 36604 26893 36632
rect 24949 36601 24961 36604
rect 24903 36595 24961 36601
rect 26881 36601 26893 36604
rect 26927 36601 26939 36635
rect 26881 36595 26939 36601
rect 26973 36635 27031 36641
rect 26973 36601 26985 36635
rect 27019 36632 27031 36635
rect 27062 36632 27068 36644
rect 27019 36604 27068 36632
rect 27019 36601 27031 36604
rect 26973 36595 27031 36601
rect 20272 36536 20668 36564
rect 21910 36524 21916 36576
rect 21968 36564 21974 36576
rect 22143 36567 22201 36573
rect 22143 36564 22155 36567
rect 21968 36536 22155 36564
rect 21968 36524 21974 36536
rect 22143 36533 22155 36536
rect 22189 36533 22201 36567
rect 22143 36527 22201 36533
rect 23566 36524 23572 36576
rect 23624 36564 23630 36576
rect 23799 36567 23857 36573
rect 23799 36564 23811 36567
rect 23624 36536 23811 36564
rect 23624 36524 23630 36536
rect 23799 36533 23811 36536
rect 23845 36533 23857 36567
rect 23799 36527 23857 36533
rect 25133 36567 25191 36573
rect 25133 36533 25145 36567
rect 25179 36564 25191 36567
rect 26053 36567 26111 36573
rect 26053 36564 26065 36567
rect 25179 36536 26065 36564
rect 25179 36533 25191 36536
rect 25133 36527 25191 36533
rect 26053 36533 26065 36536
rect 26099 36564 26111 36567
rect 26237 36567 26295 36573
rect 26237 36564 26249 36567
rect 26099 36536 26249 36564
rect 26099 36533 26111 36536
rect 26053 36527 26111 36533
rect 26237 36533 26249 36536
rect 26283 36564 26295 36567
rect 26786 36564 26792 36576
rect 26283 36536 26792 36564
rect 26283 36533 26295 36536
rect 26237 36527 26295 36533
rect 26786 36524 26792 36536
rect 26844 36524 26850 36576
rect 26896 36564 26924 36595
rect 27062 36592 27068 36604
rect 27120 36592 27126 36644
rect 27801 36567 27859 36573
rect 27801 36564 27813 36567
rect 26896 36536 27813 36564
rect 27801 36533 27813 36536
rect 27847 36533 27859 36567
rect 28994 36564 29000 36576
rect 28955 36536 29000 36564
rect 27801 36527 27859 36533
rect 28994 36524 29000 36536
rect 29052 36564 29058 36576
rect 29564 36564 29592 36663
rect 34698 36660 34704 36672
rect 34756 36700 34762 36712
rect 34885 36703 34943 36709
rect 34885 36700 34897 36703
rect 34756 36672 34897 36700
rect 34756 36660 34762 36672
rect 34885 36669 34897 36672
rect 34931 36669 34943 36703
rect 35434 36700 35440 36712
rect 35395 36672 35440 36700
rect 34885 36663 34943 36669
rect 35434 36660 35440 36672
rect 35492 36660 35498 36712
rect 35710 36660 35716 36712
rect 35768 36700 35774 36712
rect 35989 36703 36047 36709
rect 35989 36700 36001 36703
rect 35768 36672 36001 36700
rect 35768 36660 35774 36672
rect 35989 36669 36001 36672
rect 36035 36700 36047 36703
rect 36262 36700 36268 36712
rect 36035 36672 36268 36700
rect 36035 36669 36047 36672
rect 35989 36663 36047 36669
rect 36262 36660 36268 36672
rect 36320 36660 36326 36712
rect 38010 36660 38016 36712
rect 38068 36700 38074 36712
rect 38232 36703 38290 36709
rect 38232 36700 38244 36703
rect 38068 36672 38244 36700
rect 38068 36660 38074 36672
rect 38232 36669 38244 36672
rect 38278 36669 38290 36703
rect 38339 36700 38367 36740
rect 39260 36703 39318 36709
rect 39260 36700 39272 36703
rect 38339 36672 39272 36700
rect 38232 36663 38290 36669
rect 39260 36669 39272 36672
rect 39306 36700 39318 36703
rect 40840 36703 40898 36709
rect 39306 36672 39804 36700
rect 39306 36669 39318 36672
rect 39260 36663 39318 36669
rect 29638 36592 29644 36644
rect 29696 36632 29702 36644
rect 29870 36635 29928 36641
rect 29870 36632 29882 36635
rect 29696 36604 29882 36632
rect 29696 36592 29702 36604
rect 29870 36601 29882 36604
rect 29916 36601 29928 36635
rect 29870 36595 29928 36601
rect 30742 36592 30748 36644
rect 30800 36632 30806 36644
rect 30837 36635 30895 36641
rect 30837 36632 30849 36635
rect 30800 36604 30849 36632
rect 30800 36592 30806 36604
rect 30837 36601 30849 36604
rect 30883 36632 30895 36635
rect 30883 36604 31248 36632
rect 30883 36601 30895 36604
rect 30837 36595 30895 36601
rect 30466 36564 30472 36576
rect 29052 36536 29592 36564
rect 30427 36536 30472 36564
rect 29052 36524 29058 36536
rect 30466 36524 30472 36536
rect 30524 36524 30530 36576
rect 31220 36564 31248 36604
rect 31478 36592 31484 36644
rect 31536 36632 31542 36644
rect 31536 36604 31581 36632
rect 31536 36592 31542 36604
rect 32674 36592 32680 36644
rect 32732 36632 32738 36644
rect 33045 36635 33103 36641
rect 33045 36632 33057 36635
rect 32732 36604 33057 36632
rect 32732 36592 32738 36604
rect 33045 36601 33057 36604
rect 33091 36632 33103 36635
rect 33873 36635 33931 36641
rect 33873 36632 33885 36635
rect 33091 36604 33885 36632
rect 33091 36601 33103 36604
rect 33045 36595 33103 36601
rect 33873 36601 33885 36604
rect 33919 36601 33931 36635
rect 35618 36632 35624 36644
rect 35579 36604 35624 36632
rect 33873 36595 33931 36601
rect 35618 36592 35624 36604
rect 35676 36592 35682 36644
rect 36725 36635 36783 36641
rect 36725 36601 36737 36635
rect 36771 36632 36783 36635
rect 36814 36632 36820 36644
rect 36771 36604 36820 36632
rect 36771 36601 36783 36604
rect 36725 36595 36783 36601
rect 36814 36592 36820 36604
rect 36872 36592 36878 36644
rect 39776 36641 39804 36672
rect 40840 36669 40852 36703
rect 40886 36700 40898 36703
rect 41138 36700 41144 36712
rect 40886 36672 41144 36700
rect 40886 36669 40898 36672
rect 40840 36663 40898 36669
rect 41138 36660 41144 36672
rect 41196 36700 41202 36712
rect 41233 36703 41291 36709
rect 41233 36700 41245 36703
rect 41196 36672 41245 36700
rect 41196 36660 41202 36672
rect 41233 36669 41245 36672
rect 41279 36669 41291 36703
rect 41233 36663 41291 36669
rect 41690 36660 41696 36712
rect 41748 36700 41754 36712
rect 41820 36703 41878 36709
rect 41820 36700 41832 36703
rect 41748 36672 41832 36700
rect 41748 36660 41754 36672
rect 41820 36669 41832 36672
rect 41866 36700 41878 36703
rect 42245 36703 42303 36709
rect 42245 36700 42257 36703
rect 41866 36672 42257 36700
rect 41866 36669 41878 36672
rect 41820 36663 41878 36669
rect 42245 36669 42257 36672
rect 42291 36669 42303 36703
rect 42245 36663 42303 36669
rect 39347 36635 39405 36641
rect 39347 36632 39359 36635
rect 36924 36604 39359 36632
rect 31570 36564 31576 36576
rect 31220 36536 31576 36564
rect 31570 36524 31576 36536
rect 31628 36524 31634 36576
rect 31846 36524 31852 36576
rect 31904 36564 31910 36576
rect 32309 36567 32367 36573
rect 32309 36564 32321 36567
rect 31904 36536 32321 36564
rect 31904 36524 31910 36536
rect 32309 36533 32321 36536
rect 32355 36564 32367 36567
rect 32490 36564 32496 36576
rect 32355 36536 32496 36564
rect 32355 36533 32367 36536
rect 32309 36527 32367 36533
rect 32490 36524 32496 36536
rect 32548 36524 32554 36576
rect 33226 36524 33232 36576
rect 33284 36564 33290 36576
rect 36924 36564 36952 36604
rect 39347 36601 39359 36604
rect 39393 36601 39405 36635
rect 39347 36595 39405 36601
rect 39761 36635 39819 36641
rect 39761 36601 39773 36635
rect 39807 36632 39819 36635
rect 42334 36632 42340 36644
rect 39807 36604 42340 36632
rect 39807 36601 39819 36604
rect 39761 36595 39819 36601
rect 42334 36592 42340 36604
rect 42392 36592 42398 36644
rect 33284 36536 36952 36564
rect 33284 36524 33290 36536
rect 38010 36524 38016 36576
rect 38068 36564 38074 36576
rect 38657 36567 38715 36573
rect 38657 36564 38669 36567
rect 38068 36536 38669 36564
rect 38068 36524 38074 36536
rect 38657 36533 38669 36536
rect 38703 36533 38715 36567
rect 40034 36564 40040 36576
rect 39995 36536 40040 36564
rect 38657 36527 38715 36533
rect 40034 36524 40040 36536
rect 40092 36524 40098 36576
rect 1104 36474 48852 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 48852 36474
rect 1104 36400 48852 36422
rect 13633 36363 13691 36369
rect 13633 36329 13645 36363
rect 13679 36360 13691 36363
rect 13722 36360 13728 36372
rect 13679 36332 13728 36360
rect 13679 36329 13691 36332
rect 13633 36323 13691 36329
rect 13722 36320 13728 36332
rect 13780 36320 13786 36372
rect 13998 36360 14004 36372
rect 13959 36332 14004 36360
rect 13998 36320 14004 36332
rect 14056 36320 14062 36372
rect 15194 36320 15200 36372
rect 15252 36360 15258 36372
rect 15427 36363 15485 36369
rect 15427 36360 15439 36363
rect 15252 36332 15439 36360
rect 15252 36320 15258 36332
rect 15427 36329 15439 36332
rect 15473 36329 15485 36363
rect 15427 36323 15485 36329
rect 16298 36320 16304 36372
rect 16356 36360 16362 36372
rect 16761 36363 16819 36369
rect 16761 36360 16773 36363
rect 16356 36332 16773 36360
rect 16356 36320 16362 36332
rect 16761 36329 16773 36332
rect 16807 36360 16819 36363
rect 20530 36360 20536 36372
rect 16807 36332 18828 36360
rect 20491 36332 20536 36360
rect 16807 36329 16819 36332
rect 16761 36323 16819 36329
rect 18800 36304 18828 36332
rect 20530 36320 20536 36332
rect 20588 36360 20594 36372
rect 26329 36363 26387 36369
rect 20588 36332 22600 36360
rect 20588 36320 20594 36332
rect 12710 36292 12716 36304
rect 12671 36264 12716 36292
rect 12710 36252 12716 36264
rect 12768 36252 12774 36304
rect 13262 36292 13268 36304
rect 13223 36264 13268 36292
rect 13262 36252 13268 36264
rect 13320 36252 13326 36304
rect 18782 36252 18788 36304
rect 18840 36292 18846 36304
rect 18922 36295 18980 36301
rect 18922 36292 18934 36295
rect 18840 36264 18934 36292
rect 18840 36252 18846 36264
rect 18922 36261 18934 36264
rect 18968 36261 18980 36295
rect 19886 36292 19892 36304
rect 19847 36264 19892 36292
rect 18922 36255 18980 36261
rect 19886 36252 19892 36264
rect 19944 36252 19950 36304
rect 22005 36295 22063 36301
rect 22005 36261 22017 36295
rect 22051 36292 22063 36295
rect 22094 36292 22100 36304
rect 22051 36264 22100 36292
rect 22051 36261 22063 36264
rect 22005 36255 22063 36261
rect 22094 36252 22100 36264
rect 22152 36252 22158 36304
rect 22572 36301 22600 36332
rect 26329 36329 26341 36363
rect 26375 36360 26387 36363
rect 26835 36363 26893 36369
rect 26835 36360 26847 36363
rect 26375 36332 26847 36360
rect 26375 36329 26387 36332
rect 26329 36323 26387 36329
rect 26835 36329 26847 36332
rect 26881 36360 26893 36363
rect 26970 36360 26976 36372
rect 26881 36332 26976 36360
rect 26881 36329 26893 36332
rect 26835 36323 26893 36329
rect 26970 36320 26976 36332
rect 27028 36320 27034 36372
rect 27062 36320 27068 36372
rect 27120 36360 27126 36372
rect 27157 36363 27215 36369
rect 27157 36360 27169 36363
rect 27120 36332 27169 36360
rect 27120 36320 27126 36332
rect 27157 36329 27169 36332
rect 27203 36329 27215 36363
rect 27157 36323 27215 36329
rect 30466 36320 30472 36372
rect 30524 36360 30530 36372
rect 30742 36360 30748 36372
rect 30524 36332 30748 36360
rect 30524 36320 30530 36332
rect 30742 36320 30748 36332
rect 30800 36320 30806 36372
rect 32306 36360 32312 36372
rect 32267 36332 32312 36360
rect 32306 36320 32312 36332
rect 32364 36320 32370 36372
rect 35618 36360 35624 36372
rect 35579 36332 35624 36360
rect 35618 36320 35624 36332
rect 35676 36320 35682 36372
rect 36170 36360 36176 36372
rect 36131 36332 36176 36360
rect 36170 36320 36176 36332
rect 36228 36320 36234 36372
rect 36725 36363 36783 36369
rect 36725 36329 36737 36363
rect 36771 36360 36783 36363
rect 37734 36360 37740 36372
rect 36771 36332 37740 36360
rect 36771 36329 36783 36332
rect 36725 36323 36783 36329
rect 37734 36320 37740 36332
rect 37792 36360 37798 36372
rect 40126 36360 40132 36372
rect 37792 36332 37964 36360
rect 40087 36332 40132 36360
rect 37792 36320 37798 36332
rect 22557 36295 22615 36301
rect 22557 36261 22569 36295
rect 22603 36261 22615 36295
rect 22557 36255 22615 36261
rect 22738 36252 22744 36304
rect 22796 36292 22802 36304
rect 23014 36292 23020 36304
rect 22796 36264 23020 36292
rect 22796 36252 22802 36264
rect 23014 36252 23020 36264
rect 23072 36292 23078 36304
rect 28721 36295 28779 36301
rect 23072 36264 26775 36292
rect 23072 36252 23078 36264
rect 10410 36224 10416 36236
rect 10371 36196 10416 36224
rect 10410 36184 10416 36196
rect 10468 36184 10474 36236
rect 10870 36224 10876 36236
rect 10831 36196 10876 36224
rect 10870 36184 10876 36196
rect 10928 36184 10934 36236
rect 14090 36224 14096 36236
rect 14051 36196 14096 36224
rect 14090 36184 14096 36196
rect 14148 36184 14154 36236
rect 15197 36227 15255 36233
rect 15197 36193 15209 36227
rect 15243 36224 15255 36227
rect 15286 36224 15292 36236
rect 15243 36196 15292 36224
rect 15243 36193 15255 36196
rect 15197 36187 15255 36193
rect 15286 36184 15292 36196
rect 15344 36224 15350 36236
rect 15344 36196 17264 36224
rect 15344 36184 15350 36196
rect 10962 36156 10968 36168
rect 10923 36128 10968 36156
rect 10962 36116 10968 36128
rect 11020 36116 11026 36168
rect 12158 36116 12164 36168
rect 12216 36156 12222 36168
rect 12618 36156 12624 36168
rect 12216 36128 12624 36156
rect 12216 36116 12222 36128
rect 12618 36116 12624 36128
rect 12676 36116 12682 36168
rect 16390 36156 16396 36168
rect 16351 36128 16396 36156
rect 16390 36116 16396 36128
rect 16448 36116 16454 36168
rect 17236 36156 17264 36196
rect 17310 36184 17316 36236
rect 17368 36224 17374 36236
rect 18322 36224 18328 36236
rect 17368 36196 18328 36224
rect 17368 36184 17374 36196
rect 18322 36184 18328 36196
rect 18380 36224 18386 36236
rect 18601 36227 18659 36233
rect 18601 36224 18613 36227
rect 18380 36196 18613 36224
rect 18380 36184 18386 36196
rect 18601 36193 18613 36196
rect 18647 36193 18659 36227
rect 21726 36224 21732 36236
rect 18601 36187 18659 36193
rect 20916 36196 21732 36224
rect 20916 36156 20944 36196
rect 21726 36184 21732 36196
rect 21784 36184 21790 36236
rect 24029 36227 24087 36233
rect 24029 36193 24041 36227
rect 24075 36193 24087 36227
rect 24210 36224 24216 36236
rect 24171 36196 24216 36224
rect 24029 36187 24087 36193
rect 17236 36128 20944 36156
rect 20990 36116 20996 36168
rect 21048 36156 21054 36168
rect 21910 36156 21916 36168
rect 21048 36128 21916 36156
rect 21048 36116 21054 36128
rect 21910 36116 21916 36128
rect 21968 36116 21974 36168
rect 16482 36048 16488 36100
rect 16540 36088 16546 36100
rect 23382 36088 23388 36100
rect 16540 36060 23388 36088
rect 16540 36048 16546 36060
rect 23382 36048 23388 36060
rect 23440 36088 23446 36100
rect 24044 36088 24072 36187
rect 24210 36184 24216 36196
rect 24268 36184 24274 36236
rect 24762 36184 24768 36236
rect 24820 36224 24826 36236
rect 25406 36224 25412 36236
rect 25464 36233 25470 36236
rect 26747 36233 26775 36264
rect 28721 36261 28733 36295
rect 28767 36292 28779 36295
rect 28994 36292 29000 36304
rect 28767 36264 29000 36292
rect 28767 36261 28779 36264
rect 28721 36255 28779 36261
rect 28994 36252 29000 36264
rect 29052 36252 29058 36304
rect 29638 36252 29644 36304
rect 29696 36292 29702 36304
rect 29870 36295 29928 36301
rect 29870 36292 29882 36295
rect 29696 36264 29882 36292
rect 29696 36252 29702 36264
rect 29870 36261 29882 36264
rect 29916 36292 29928 36295
rect 31846 36292 31852 36304
rect 29916 36264 31852 36292
rect 29916 36261 29928 36264
rect 29870 36255 29928 36261
rect 31846 36252 31852 36264
rect 31904 36252 31910 36304
rect 32030 36252 32036 36304
rect 32088 36292 32094 36304
rect 32858 36292 32864 36304
rect 32088 36264 32864 36292
rect 32088 36252 32094 36264
rect 32858 36252 32864 36264
rect 32916 36252 32922 36304
rect 32953 36295 33011 36301
rect 32953 36261 32965 36295
rect 32999 36292 33011 36295
rect 33134 36292 33140 36304
rect 32999 36264 33140 36292
rect 32999 36261 33011 36264
rect 32953 36255 33011 36261
rect 33134 36252 33140 36264
rect 33192 36252 33198 36304
rect 37826 36292 37832 36304
rect 37787 36264 37832 36292
rect 37826 36252 37832 36264
rect 37884 36252 37890 36304
rect 37936 36301 37964 36332
rect 40126 36320 40132 36332
rect 40184 36320 40190 36372
rect 41230 36360 41236 36372
rect 40281 36332 41236 36360
rect 37921 36295 37979 36301
rect 37921 36261 37933 36295
rect 37967 36261 37979 36295
rect 37921 36255 37979 36261
rect 38010 36252 38016 36304
rect 38068 36292 38074 36304
rect 40281 36292 40309 36332
rect 41230 36320 41236 36332
rect 41288 36360 41294 36372
rect 41782 36360 41788 36372
rect 41288 36332 41460 36360
rect 41743 36332 41788 36360
rect 41288 36320 41294 36332
rect 40862 36292 40868 36304
rect 38068 36264 40309 36292
rect 40823 36264 40868 36292
rect 38068 36252 38074 36264
rect 40862 36252 40868 36264
rect 40920 36252 40926 36304
rect 41432 36301 41460 36332
rect 41782 36320 41788 36332
rect 41840 36320 41846 36372
rect 41417 36295 41475 36301
rect 41417 36261 41429 36295
rect 41463 36261 41475 36295
rect 41417 36255 41475 36261
rect 25464 36227 25502 36233
rect 24820 36196 25412 36224
rect 24820 36184 24826 36196
rect 25406 36184 25412 36196
rect 25490 36193 25502 36227
rect 25464 36187 25502 36193
rect 26732 36227 26790 36233
rect 26732 36193 26744 36227
rect 26778 36224 26790 36227
rect 27062 36224 27068 36236
rect 26778 36196 27068 36224
rect 26778 36193 26790 36196
rect 26732 36187 26790 36193
rect 25464 36184 25470 36187
rect 27062 36184 27068 36196
rect 27120 36184 27126 36236
rect 28261 36227 28319 36233
rect 28261 36193 28273 36227
rect 28307 36224 28319 36227
rect 28350 36224 28356 36236
rect 28307 36196 28356 36224
rect 28307 36193 28319 36196
rect 28261 36187 28319 36193
rect 28350 36184 28356 36196
rect 28408 36184 28414 36236
rect 28442 36184 28448 36236
rect 28500 36224 28506 36236
rect 29454 36224 29460 36236
rect 28500 36196 29460 36224
rect 28500 36184 28506 36196
rect 29454 36184 29460 36196
rect 29512 36224 29518 36236
rect 30006 36224 30012 36236
rect 29512 36196 30012 36224
rect 29512 36184 29518 36196
rect 30006 36184 30012 36196
rect 30064 36184 30070 36236
rect 30469 36227 30527 36233
rect 30469 36193 30481 36227
rect 30515 36224 30527 36227
rect 31297 36227 31355 36233
rect 31297 36224 31309 36227
rect 30515 36196 31309 36224
rect 30515 36193 30527 36196
rect 30469 36187 30527 36193
rect 31297 36193 31309 36196
rect 31343 36224 31355 36227
rect 31478 36224 31484 36236
rect 31343 36196 31484 36224
rect 31343 36193 31355 36196
rect 31297 36187 31355 36193
rect 31478 36184 31484 36196
rect 31536 36184 31542 36236
rect 34330 36224 34336 36236
rect 34291 36196 34336 36224
rect 34330 36184 34336 36196
rect 34388 36184 34394 36236
rect 39666 36224 39672 36236
rect 39627 36196 39672 36224
rect 39666 36184 39672 36196
rect 39724 36184 39730 36236
rect 24302 36156 24308 36168
rect 24263 36128 24308 36156
rect 24302 36116 24308 36128
rect 24360 36116 24366 36168
rect 25547 36159 25605 36165
rect 25547 36125 25559 36159
rect 25593 36156 25605 36159
rect 28534 36156 28540 36168
rect 25593 36128 28540 36156
rect 25593 36125 25605 36128
rect 25547 36119 25605 36125
rect 28534 36116 28540 36128
rect 28592 36156 28598 36168
rect 28997 36159 29055 36165
rect 28997 36156 29009 36159
rect 28592 36128 29009 36156
rect 28592 36116 28598 36128
rect 28997 36125 29009 36128
rect 29043 36125 29055 36159
rect 29546 36156 29552 36168
rect 29507 36128 29552 36156
rect 28997 36119 29055 36125
rect 29546 36116 29552 36128
rect 29604 36116 29610 36168
rect 33137 36159 33195 36165
rect 33137 36125 33149 36159
rect 33183 36125 33195 36159
rect 35802 36156 35808 36168
rect 35763 36128 35808 36156
rect 33137 36119 33195 36125
rect 28350 36088 28356 36100
rect 23440 36060 28356 36088
rect 23440 36048 23446 36060
rect 28350 36048 28356 36060
rect 28408 36048 28414 36100
rect 31386 36048 31392 36100
rect 31444 36088 31450 36100
rect 33152 36088 33180 36119
rect 35802 36116 35808 36128
rect 35860 36116 35866 36168
rect 38105 36159 38163 36165
rect 38105 36125 38117 36159
rect 38151 36125 38163 36159
rect 38105 36119 38163 36125
rect 40773 36159 40831 36165
rect 40773 36125 40785 36159
rect 40819 36156 40831 36159
rect 41690 36156 41696 36168
rect 40819 36128 41696 36156
rect 40819 36125 40831 36128
rect 40773 36119 40831 36125
rect 31444 36060 33180 36088
rect 31444 36048 31450 36060
rect 36906 36048 36912 36100
rect 36964 36088 36970 36100
rect 38120 36088 38148 36119
rect 41690 36116 41696 36128
rect 41748 36116 41754 36168
rect 38470 36088 38476 36100
rect 36964 36060 38476 36088
rect 36964 36048 36970 36060
rect 38470 36048 38476 36060
rect 38528 36048 38534 36100
rect 38764 36060 40908 36088
rect 12066 36020 12072 36032
rect 12027 35992 12072 36020
rect 12066 35980 12072 35992
rect 12124 35980 12130 36032
rect 14323 36023 14381 36029
rect 14323 35989 14335 36023
rect 14369 36020 14381 36023
rect 14642 36020 14648 36032
rect 14369 35992 14648 36020
rect 14369 35989 14381 35992
rect 14323 35983 14381 35989
rect 14642 35980 14648 35992
rect 14700 35980 14706 36032
rect 16574 35980 16580 36032
rect 16632 36020 16638 36032
rect 17313 36023 17371 36029
rect 17313 36020 17325 36023
rect 16632 35992 17325 36020
rect 16632 35980 16638 35992
rect 17313 35989 17325 35992
rect 17359 35989 17371 36023
rect 17313 35983 17371 35989
rect 18233 36023 18291 36029
rect 18233 35989 18245 36023
rect 18279 36020 18291 36023
rect 18414 36020 18420 36032
rect 18279 35992 18420 36020
rect 18279 35989 18291 35992
rect 18233 35983 18291 35989
rect 18414 35980 18420 35992
rect 18472 35980 18478 36032
rect 19518 36020 19524 36032
rect 19479 35992 19524 36020
rect 19518 35980 19524 35992
rect 19576 35980 19582 36032
rect 24762 36020 24768 36032
rect 24723 35992 24768 36020
rect 24762 35980 24768 35992
rect 24820 35980 24826 36032
rect 27706 36020 27712 36032
rect 27667 35992 27712 36020
rect 27706 35980 27712 35992
rect 27764 35980 27770 36032
rect 34471 36023 34529 36029
rect 34471 35989 34483 36023
rect 34517 36020 34529 36023
rect 34790 36020 34796 36032
rect 34517 35992 34796 36020
rect 34517 35989 34529 35992
rect 34471 35983 34529 35989
rect 34790 35980 34796 35992
rect 34848 35980 34854 36032
rect 34977 36023 35035 36029
rect 34977 35989 34989 36023
rect 35023 36020 35035 36023
rect 35434 36020 35440 36032
rect 35023 35992 35440 36020
rect 35023 35989 35035 35992
rect 34977 35983 35035 35989
rect 35434 35980 35440 35992
rect 35492 35980 35498 36032
rect 36998 35980 37004 36032
rect 37056 36020 37062 36032
rect 37093 36023 37151 36029
rect 37093 36020 37105 36023
rect 37056 35992 37105 36020
rect 37056 35980 37062 35992
rect 37093 35989 37105 35992
rect 37139 36020 37151 36023
rect 38764 36020 38792 36060
rect 37139 35992 38792 36020
rect 39807 36023 39865 36029
rect 37139 35989 37151 35992
rect 37093 35983 37151 35989
rect 39807 35989 39819 36023
rect 39853 36020 39865 36023
rect 40770 36020 40776 36032
rect 39853 35992 40776 36020
rect 39853 35989 39865 35992
rect 39807 35983 39865 35989
rect 40770 35980 40776 35992
rect 40828 35980 40834 36032
rect 40880 36020 40908 36060
rect 41414 36020 41420 36032
rect 40880 35992 41420 36020
rect 41414 35980 41420 35992
rect 41472 35980 41478 36032
rect 42337 36023 42395 36029
rect 42337 35989 42349 36023
rect 42383 36020 42395 36023
rect 42426 36020 42432 36032
rect 42383 35992 42432 36020
rect 42383 35989 42395 35992
rect 42337 35983 42395 35989
rect 42426 35980 42432 35992
rect 42484 35980 42490 36032
rect 1104 35930 48852 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 48852 35930
rect 1104 35856 48852 35878
rect 9674 35776 9680 35828
rect 9732 35816 9738 35828
rect 10410 35816 10416 35828
rect 9732 35788 10416 35816
rect 9732 35776 9738 35788
rect 10410 35776 10416 35788
rect 10468 35776 10474 35828
rect 10870 35776 10876 35828
rect 10928 35816 10934 35828
rect 11330 35816 11336 35828
rect 10928 35788 11336 35816
rect 10928 35776 10934 35788
rect 11330 35776 11336 35788
rect 11388 35816 11394 35828
rect 11793 35819 11851 35825
rect 11793 35816 11805 35819
rect 11388 35788 11805 35816
rect 11388 35776 11394 35788
rect 11793 35785 11805 35788
rect 11839 35785 11851 35819
rect 11793 35779 11851 35785
rect 13449 35819 13507 35825
rect 13449 35785 13461 35819
rect 13495 35816 13507 35819
rect 13722 35816 13728 35828
rect 13495 35788 13728 35816
rect 13495 35785 13507 35788
rect 13449 35779 13507 35785
rect 13722 35776 13728 35788
rect 13780 35776 13786 35828
rect 16298 35816 16304 35828
rect 16259 35788 16304 35816
rect 16298 35776 16304 35788
rect 16356 35776 16362 35828
rect 18322 35816 18328 35828
rect 18283 35788 18328 35816
rect 18322 35776 18328 35788
rect 18380 35776 18386 35828
rect 18782 35776 18788 35828
rect 18840 35816 18846 35828
rect 18969 35819 19027 35825
rect 18969 35816 18981 35819
rect 18840 35788 18981 35816
rect 18840 35776 18846 35788
rect 18969 35785 18981 35788
rect 19015 35785 19027 35819
rect 18969 35779 19027 35785
rect 19429 35819 19487 35825
rect 19429 35785 19441 35819
rect 19475 35816 19487 35819
rect 19518 35816 19524 35828
rect 19475 35788 19524 35816
rect 19475 35785 19487 35788
rect 19429 35779 19487 35785
rect 19518 35776 19524 35788
rect 19576 35776 19582 35828
rect 19886 35776 19892 35828
rect 19944 35816 19950 35828
rect 20990 35816 20996 35828
rect 19944 35788 20805 35816
rect 20951 35788 20996 35816
rect 19944 35776 19950 35788
rect 12526 35708 12532 35760
rect 12584 35708 12590 35760
rect 13998 35708 14004 35760
rect 14056 35748 14062 35760
rect 19904 35748 19932 35776
rect 14056 35720 14688 35748
rect 14056 35708 14062 35720
rect 12544 35680 12572 35708
rect 14090 35680 14096 35692
rect 11072 35652 12572 35680
rect 14051 35652 14096 35680
rect 11072 35621 11100 35652
rect 14090 35640 14096 35652
rect 14148 35640 14154 35692
rect 14366 35680 14372 35692
rect 14327 35652 14372 35680
rect 14366 35640 14372 35652
rect 14424 35640 14430 35692
rect 14660 35689 14688 35720
rect 19628 35720 19932 35748
rect 20777 35748 20805 35788
rect 20990 35776 20996 35788
rect 21048 35776 21054 35828
rect 23106 35816 23112 35828
rect 23067 35788 23112 35816
rect 23106 35776 23112 35788
rect 23164 35776 23170 35828
rect 23382 35816 23388 35828
rect 23343 35788 23388 35816
rect 23382 35776 23388 35788
rect 23440 35776 23446 35828
rect 24213 35819 24271 35825
rect 24213 35785 24225 35819
rect 24259 35816 24271 35819
rect 24670 35816 24676 35828
rect 24259 35788 24676 35816
rect 24259 35785 24271 35788
rect 24213 35779 24271 35785
rect 24670 35776 24676 35788
rect 24728 35776 24734 35828
rect 25406 35776 25412 35828
rect 25464 35816 25470 35828
rect 25501 35819 25559 35825
rect 25501 35816 25513 35819
rect 25464 35788 25513 35816
rect 25464 35776 25470 35788
rect 25501 35785 25513 35788
rect 25547 35785 25559 35819
rect 27062 35816 27068 35828
rect 27023 35788 27068 35816
rect 25501 35779 25559 35785
rect 27062 35776 27068 35788
rect 27120 35776 27126 35828
rect 27525 35819 27583 35825
rect 27525 35785 27537 35819
rect 27571 35816 27583 35819
rect 28442 35816 28448 35828
rect 27571 35788 28448 35816
rect 27571 35785 27583 35788
rect 27525 35779 27583 35785
rect 28442 35776 28448 35788
rect 28500 35776 28506 35828
rect 29089 35819 29147 35825
rect 29089 35785 29101 35819
rect 29135 35816 29147 35819
rect 29546 35816 29552 35828
rect 29135 35788 29552 35816
rect 29135 35785 29147 35788
rect 29089 35779 29147 35785
rect 29546 35776 29552 35788
rect 29604 35776 29610 35828
rect 29638 35776 29644 35828
rect 29696 35816 29702 35828
rect 30101 35819 30159 35825
rect 30101 35816 30113 35819
rect 29696 35788 30113 35816
rect 29696 35776 29702 35788
rect 30101 35785 30113 35788
rect 30147 35785 30159 35819
rect 30101 35779 30159 35785
rect 32490 35776 32496 35828
rect 32548 35816 32554 35828
rect 34330 35816 34336 35828
rect 32548 35788 34336 35816
rect 32548 35776 32554 35788
rect 34330 35776 34336 35788
rect 34388 35816 34394 35828
rect 36449 35819 36507 35825
rect 34388 35788 34468 35816
rect 34388 35776 34394 35788
rect 22465 35751 22523 35757
rect 22465 35748 22477 35751
rect 20777 35720 22477 35748
rect 14645 35683 14703 35689
rect 14645 35649 14657 35683
rect 14691 35649 14703 35683
rect 14645 35643 14703 35649
rect 15933 35683 15991 35689
rect 15933 35649 15945 35683
rect 15979 35680 15991 35683
rect 16574 35680 16580 35692
rect 15979 35652 16580 35680
rect 15979 35649 15991 35652
rect 15933 35643 15991 35649
rect 16574 35640 16580 35652
rect 16632 35640 16638 35692
rect 16758 35680 16764 35692
rect 16719 35652 16764 35680
rect 16758 35640 16764 35652
rect 16816 35640 16822 35692
rect 19628 35689 19656 35720
rect 22465 35717 22477 35720
rect 22511 35717 22523 35751
rect 28261 35751 28319 35757
rect 28261 35748 28273 35751
rect 22465 35711 22523 35717
rect 26160 35720 28273 35748
rect 26160 35692 26188 35720
rect 28261 35717 28273 35720
rect 28307 35748 28319 35751
rect 28810 35748 28816 35760
rect 28307 35720 28816 35748
rect 28307 35717 28319 35720
rect 28261 35711 28319 35717
rect 28810 35708 28816 35720
rect 28868 35708 28874 35760
rect 31573 35751 31631 35757
rect 31573 35748 31585 35751
rect 30668 35720 31585 35748
rect 19613 35683 19671 35689
rect 19613 35649 19625 35683
rect 19659 35649 19671 35683
rect 19886 35680 19892 35692
rect 19847 35652 19892 35680
rect 19613 35643 19671 35649
rect 19886 35640 19892 35652
rect 19944 35640 19950 35692
rect 21913 35683 21971 35689
rect 21913 35649 21925 35683
rect 21959 35680 21971 35683
rect 22002 35680 22008 35692
rect 21959 35652 22008 35680
rect 21959 35649 21971 35652
rect 21913 35643 21971 35649
rect 22002 35640 22008 35652
rect 22060 35680 22066 35692
rect 23566 35680 23572 35692
rect 22060 35652 23572 35680
rect 22060 35640 22066 35652
rect 23566 35640 23572 35652
rect 23624 35640 23630 35692
rect 24305 35683 24363 35689
rect 24305 35649 24317 35683
rect 24351 35680 24363 35683
rect 24762 35680 24768 35692
rect 24351 35652 24768 35680
rect 24351 35649 24363 35652
rect 24305 35643 24363 35649
rect 24762 35640 24768 35652
rect 24820 35640 24826 35692
rect 26142 35680 26148 35692
rect 26103 35652 26148 35680
rect 26142 35640 26148 35652
rect 26200 35640 26206 35692
rect 26418 35680 26424 35692
rect 26379 35652 26424 35680
rect 26418 35640 26424 35652
rect 26476 35640 26482 35692
rect 27709 35683 27767 35689
rect 27709 35649 27721 35683
rect 27755 35680 27767 35683
rect 28166 35680 28172 35692
rect 27755 35652 28172 35680
rect 27755 35649 27767 35652
rect 27709 35643 27767 35649
rect 28166 35640 28172 35652
rect 28224 35640 28230 35692
rect 28350 35640 28356 35692
rect 28408 35680 28414 35692
rect 28718 35680 28724 35692
rect 28408 35652 28724 35680
rect 28408 35640 28414 35652
rect 28718 35640 28724 35652
rect 28776 35640 28782 35692
rect 30668 35689 30696 35720
rect 31573 35717 31585 35720
rect 31619 35748 31631 35751
rect 32398 35748 32404 35760
rect 31619 35720 32404 35748
rect 31619 35717 31631 35720
rect 31573 35711 31631 35717
rect 32398 35708 32404 35720
rect 32456 35748 32462 35760
rect 34440 35757 34468 35788
rect 36449 35785 36461 35819
rect 36495 35816 36507 35819
rect 36814 35816 36820 35828
rect 36495 35788 36820 35816
rect 36495 35785 36507 35788
rect 36449 35779 36507 35785
rect 36814 35776 36820 35788
rect 36872 35776 36878 35828
rect 37734 35816 37740 35828
rect 37695 35788 37740 35816
rect 37734 35776 37740 35788
rect 37792 35776 37798 35828
rect 38378 35776 38384 35828
rect 38436 35816 38442 35828
rect 39666 35816 39672 35828
rect 38436 35788 39672 35816
rect 38436 35776 38442 35788
rect 39666 35776 39672 35788
rect 39724 35776 39730 35828
rect 41690 35816 41696 35828
rect 41651 35788 41696 35816
rect 41690 35776 41696 35788
rect 41748 35776 41754 35828
rect 34425 35751 34483 35757
rect 32456 35720 33272 35748
rect 32456 35708 32462 35720
rect 30653 35683 30711 35689
rect 30653 35649 30665 35683
rect 30699 35649 30711 35683
rect 31294 35680 31300 35692
rect 31207 35652 31300 35680
rect 30653 35643 30711 35649
rect 31294 35640 31300 35652
rect 31352 35680 31358 35692
rect 31662 35680 31668 35692
rect 31352 35652 31668 35680
rect 31352 35640 31358 35652
rect 31662 35640 31668 35652
rect 31720 35640 31726 35692
rect 32033 35683 32091 35689
rect 32033 35649 32045 35683
rect 32079 35680 32091 35683
rect 32953 35683 33011 35689
rect 32953 35680 32965 35683
rect 32079 35652 32965 35680
rect 32079 35649 32091 35652
rect 32033 35643 32091 35649
rect 32953 35649 32965 35652
rect 32999 35680 33011 35683
rect 33042 35680 33048 35692
rect 32999 35652 33048 35680
rect 32999 35649 33011 35652
rect 32953 35643 33011 35649
rect 33042 35640 33048 35652
rect 33100 35640 33106 35692
rect 33244 35689 33272 35720
rect 34425 35717 34437 35751
rect 34471 35748 34483 35751
rect 37274 35748 37280 35760
rect 34471 35720 37280 35748
rect 34471 35717 34483 35720
rect 34425 35711 34483 35717
rect 37274 35708 37280 35720
rect 37332 35708 37338 35760
rect 39209 35751 39267 35757
rect 39209 35748 39221 35751
rect 38212 35720 39221 35748
rect 33229 35683 33287 35689
rect 33229 35649 33241 35683
rect 33275 35649 33287 35683
rect 33229 35643 33287 35649
rect 35529 35683 35587 35689
rect 35529 35649 35541 35683
rect 35575 35680 35587 35683
rect 35618 35680 35624 35692
rect 35575 35652 35624 35680
rect 35575 35649 35587 35652
rect 35529 35643 35587 35649
rect 35618 35640 35624 35652
rect 35676 35640 35682 35692
rect 35802 35640 35808 35692
rect 35860 35680 35866 35692
rect 38212 35689 38240 35720
rect 39209 35717 39221 35720
rect 39255 35748 39267 35751
rect 39298 35748 39304 35760
rect 39255 35720 39304 35748
rect 39255 35717 39267 35720
rect 39209 35711 39267 35717
rect 39298 35708 39304 35720
rect 39356 35748 39362 35760
rect 39356 35720 42656 35748
rect 39356 35708 39362 35720
rect 42628 35692 42656 35720
rect 36725 35683 36783 35689
rect 36725 35680 36737 35683
rect 35860 35652 36737 35680
rect 35860 35640 35866 35652
rect 36725 35649 36737 35652
rect 36771 35649 36783 35683
rect 36725 35643 36783 35649
rect 38197 35683 38255 35689
rect 38197 35649 38209 35683
rect 38243 35649 38255 35683
rect 38470 35680 38476 35692
rect 38431 35652 38476 35680
rect 38197 35643 38255 35649
rect 38470 35640 38476 35652
rect 38528 35640 38534 35692
rect 40770 35680 40776 35692
rect 40731 35652 40776 35680
rect 40770 35640 40776 35652
rect 40828 35640 40834 35692
rect 41414 35680 41420 35692
rect 41375 35652 41420 35680
rect 41414 35640 41420 35652
rect 41472 35640 41478 35692
rect 42610 35680 42616 35692
rect 42571 35652 42616 35680
rect 42610 35640 42616 35652
rect 42668 35640 42674 35692
rect 10137 35615 10195 35621
rect 10137 35581 10149 35615
rect 10183 35612 10195 35615
rect 11057 35615 11115 35621
rect 11057 35612 11069 35615
rect 10183 35584 11069 35612
rect 10183 35581 10195 35584
rect 10137 35575 10195 35581
rect 11057 35581 11069 35584
rect 11103 35581 11115 35615
rect 11330 35612 11336 35624
rect 11291 35584 11336 35612
rect 11057 35575 11115 35581
rect 11330 35572 11336 35584
rect 11388 35572 11394 35624
rect 11517 35615 11575 35621
rect 11517 35581 11529 35615
rect 11563 35612 11575 35615
rect 12529 35615 12587 35621
rect 12529 35612 12541 35615
rect 11563 35584 12541 35612
rect 11563 35581 11575 35584
rect 11517 35575 11575 35581
rect 12529 35581 12541 35584
rect 12575 35612 12587 35615
rect 13725 35615 13783 35621
rect 13725 35612 13737 35615
rect 12575 35584 13737 35612
rect 12575 35581 12587 35584
rect 12529 35575 12587 35581
rect 13725 35581 13737 35584
rect 13771 35581 13783 35615
rect 29308 35615 29366 35621
rect 29308 35612 29320 35615
rect 13725 35575 13783 35581
rect 28644 35584 29320 35612
rect 11974 35504 11980 35556
rect 12032 35544 12038 35556
rect 12253 35547 12311 35553
rect 12253 35544 12265 35547
rect 12032 35516 12265 35544
rect 12032 35504 12038 35516
rect 12253 35513 12265 35516
rect 12299 35544 12311 35547
rect 12891 35547 12949 35553
rect 12891 35544 12903 35547
rect 12299 35516 12903 35544
rect 12299 35513 12311 35516
rect 12253 35507 12311 35513
rect 12891 35513 12903 35516
rect 12937 35544 12949 35547
rect 13354 35544 13360 35556
rect 12937 35516 13360 35544
rect 12937 35513 12949 35516
rect 12891 35507 12949 35513
rect 13354 35504 13360 35516
rect 13412 35504 13418 35556
rect 14458 35544 14464 35556
rect 14419 35516 14464 35544
rect 14458 35504 14464 35516
rect 14516 35504 14522 35556
rect 15930 35504 15936 35556
rect 15988 35544 15994 35556
rect 16485 35547 16543 35553
rect 16485 35544 16497 35547
rect 15988 35516 16497 35544
rect 15988 35504 15994 35516
rect 16485 35513 16497 35516
rect 16531 35513 16543 35547
rect 16485 35507 16543 35513
rect 15286 35476 15292 35488
rect 15247 35448 15292 35476
rect 15286 35436 15292 35448
rect 15344 35436 15350 35488
rect 16500 35476 16528 35507
rect 16574 35504 16580 35556
rect 16632 35544 16638 35556
rect 18509 35547 18567 35553
rect 16632 35516 16677 35544
rect 16632 35504 16638 35516
rect 18509 35513 18521 35547
rect 18555 35544 18567 35547
rect 18555 35516 19282 35544
rect 18555 35513 18567 35516
rect 18509 35507 18567 35513
rect 17405 35479 17463 35485
rect 17405 35476 17417 35479
rect 16500 35448 17417 35476
rect 17405 35445 17417 35448
rect 17451 35445 17463 35479
rect 19254 35476 19282 35516
rect 19702 35504 19708 35556
rect 19760 35544 19766 35556
rect 21361 35547 21419 35553
rect 19760 35516 19805 35544
rect 19760 35504 19766 35516
rect 21361 35513 21373 35547
rect 21407 35544 21419 35547
rect 21729 35547 21787 35553
rect 21729 35544 21741 35547
rect 21407 35516 21741 35544
rect 21407 35513 21419 35516
rect 21361 35507 21419 35513
rect 21729 35513 21741 35516
rect 21775 35544 21787 35547
rect 22005 35547 22063 35553
rect 22005 35544 22017 35547
rect 21775 35516 22017 35544
rect 21775 35513 21787 35516
rect 21729 35507 21787 35513
rect 22005 35513 22017 35516
rect 22051 35544 22063 35547
rect 22094 35544 22100 35556
rect 22051 35516 22100 35544
rect 22051 35513 22063 35516
rect 22005 35507 22063 35513
rect 22094 35504 22100 35516
rect 22152 35504 22158 35556
rect 26237 35547 26295 35553
rect 26237 35513 26249 35547
rect 26283 35513 26295 35547
rect 26237 35507 26295 35513
rect 22370 35476 22376 35488
rect 19254 35448 22376 35476
rect 17405 35439 17463 35445
rect 22370 35436 22376 35448
rect 22428 35436 22434 35488
rect 24670 35476 24676 35488
rect 24631 35448 24676 35476
rect 24670 35436 24676 35448
rect 24728 35436 24734 35488
rect 25222 35476 25228 35488
rect 25183 35448 25228 35476
rect 25222 35436 25228 35448
rect 25280 35436 25286 35488
rect 25866 35476 25872 35488
rect 25827 35448 25872 35476
rect 25866 35436 25872 35448
rect 25924 35476 25930 35488
rect 26252 35476 26280 35507
rect 27706 35504 27712 35556
rect 27764 35544 27770 35556
rect 27801 35547 27859 35553
rect 27801 35544 27813 35547
rect 27764 35516 27813 35544
rect 27764 35504 27770 35516
rect 27801 35513 27813 35516
rect 27847 35513 27859 35547
rect 27801 35507 27859 35513
rect 25924 35448 26280 35476
rect 25924 35436 25930 35448
rect 26510 35436 26516 35488
rect 26568 35476 26574 35488
rect 28644 35476 28672 35584
rect 29308 35581 29320 35584
rect 29354 35612 29366 35615
rect 29730 35612 29736 35624
rect 29354 35584 29736 35612
rect 29354 35581 29366 35584
rect 29308 35575 29366 35581
rect 29730 35572 29736 35584
rect 29788 35572 29794 35624
rect 30742 35504 30748 35556
rect 30800 35544 30806 35556
rect 32401 35547 32459 35553
rect 30800 35516 30845 35544
rect 30800 35504 30806 35516
rect 32401 35513 32413 35547
rect 32447 35544 32459 35547
rect 32769 35547 32827 35553
rect 32769 35544 32781 35547
rect 32447 35516 32781 35544
rect 32447 35513 32459 35516
rect 32401 35507 32459 35513
rect 32769 35513 32781 35516
rect 32815 35544 32827 35547
rect 33045 35547 33103 35553
rect 33045 35544 33057 35547
rect 32815 35516 33057 35544
rect 32815 35513 32827 35516
rect 32769 35507 32827 35513
rect 33045 35513 33057 35516
rect 33091 35544 33103 35547
rect 33134 35544 33140 35556
rect 33091 35516 33140 35544
rect 33091 35513 33103 35516
rect 33045 35507 33103 35513
rect 33134 35504 33140 35516
rect 33192 35504 33198 35556
rect 35437 35547 35495 35553
rect 35437 35513 35449 35547
rect 35483 35544 35495 35547
rect 35891 35547 35949 35553
rect 35891 35544 35903 35547
rect 35483 35516 35903 35544
rect 35483 35513 35495 35516
rect 35437 35507 35495 35513
rect 35891 35513 35903 35516
rect 35937 35544 35949 35547
rect 36170 35544 36176 35556
rect 35937 35516 36176 35544
rect 35937 35513 35949 35516
rect 35891 35507 35949 35513
rect 36170 35504 36176 35516
rect 36228 35504 36234 35556
rect 38289 35547 38347 35553
rect 38289 35513 38301 35547
rect 38335 35513 38347 35547
rect 38289 35507 38347 35513
rect 40313 35547 40371 35553
rect 40313 35513 40325 35547
rect 40359 35544 40371 35547
rect 40862 35544 40868 35556
rect 40359 35516 40868 35544
rect 40359 35513 40371 35516
rect 40313 35507 40371 35513
rect 26568 35448 28672 35476
rect 26568 35436 26574 35448
rect 28718 35436 28724 35488
rect 28776 35476 28782 35488
rect 29411 35479 29469 35485
rect 29411 35476 29423 35479
rect 28776 35448 29423 35476
rect 28776 35436 28782 35448
rect 29411 35445 29423 35448
rect 29457 35445 29469 35479
rect 29411 35439 29469 35445
rect 37461 35479 37519 35485
rect 37461 35445 37473 35479
rect 37507 35476 37519 35479
rect 38304 35476 38332 35507
rect 40862 35504 40868 35516
rect 40920 35504 40926 35556
rect 42337 35547 42395 35553
rect 42337 35513 42349 35547
rect 42383 35513 42395 35547
rect 42337 35507 42395 35513
rect 38654 35476 38660 35488
rect 37507 35448 38660 35476
rect 37507 35445 37519 35448
rect 37461 35439 37519 35445
rect 38654 35436 38660 35448
rect 38712 35436 38718 35488
rect 42058 35476 42064 35488
rect 42019 35448 42064 35476
rect 42058 35436 42064 35448
rect 42116 35476 42122 35488
rect 42352 35476 42380 35507
rect 42426 35504 42432 35556
rect 42484 35544 42490 35556
rect 42484 35516 42529 35544
rect 42484 35504 42490 35516
rect 42116 35448 42380 35476
rect 42116 35436 42122 35448
rect 1104 35386 48852 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 48852 35386
rect 1104 35312 48852 35334
rect 10505 35275 10563 35281
rect 10505 35241 10517 35275
rect 10551 35272 10563 35275
rect 10870 35272 10876 35284
rect 10551 35244 10876 35272
rect 10551 35241 10563 35244
rect 10505 35235 10563 35241
rect 10870 35232 10876 35244
rect 10928 35232 10934 35284
rect 12158 35272 12164 35284
rect 12119 35244 12164 35272
rect 12158 35232 12164 35244
rect 12216 35232 12222 35284
rect 12529 35275 12587 35281
rect 12529 35241 12541 35275
rect 12575 35272 12587 35275
rect 12710 35272 12716 35284
rect 12575 35244 12716 35272
rect 12575 35241 12587 35244
rect 12529 35235 12587 35241
rect 12710 35232 12716 35244
rect 12768 35272 12774 35284
rect 13541 35275 13599 35281
rect 13541 35272 13553 35275
rect 12768 35244 13553 35272
rect 12768 35232 12774 35244
rect 13541 35241 13553 35244
rect 13587 35241 13599 35275
rect 13541 35235 13599 35241
rect 14366 35232 14372 35284
rect 14424 35272 14430 35284
rect 14645 35275 14703 35281
rect 14645 35272 14657 35275
rect 14424 35244 14657 35272
rect 14424 35232 14430 35244
rect 14645 35241 14657 35244
rect 14691 35241 14703 35275
rect 14645 35235 14703 35241
rect 16390 35232 16396 35284
rect 16448 35272 16454 35284
rect 16761 35275 16819 35281
rect 16761 35272 16773 35275
rect 16448 35244 16773 35272
rect 16448 35232 16454 35244
rect 16761 35241 16773 35244
rect 16807 35272 16819 35275
rect 17405 35275 17463 35281
rect 17405 35272 17417 35275
rect 16807 35244 17417 35272
rect 16807 35241 16819 35244
rect 16761 35235 16819 35241
rect 17405 35241 17417 35244
rect 17451 35241 17463 35275
rect 22002 35272 22008 35284
rect 21963 35244 22008 35272
rect 17405 35235 17463 35241
rect 22002 35232 22008 35244
rect 22060 35232 22066 35284
rect 23106 35232 23112 35284
rect 23164 35272 23170 35284
rect 23842 35272 23848 35284
rect 23164 35244 23848 35272
rect 23164 35232 23170 35244
rect 23842 35232 23848 35244
rect 23900 35232 23906 35284
rect 24670 35272 24676 35284
rect 24631 35244 24676 35272
rect 24670 35232 24676 35244
rect 24728 35232 24734 35284
rect 25225 35275 25283 35281
rect 25225 35241 25237 35275
rect 25271 35272 25283 35275
rect 25866 35272 25872 35284
rect 25271 35244 25872 35272
rect 25271 35241 25283 35244
rect 25225 35235 25283 35241
rect 25866 35232 25872 35244
rect 25924 35232 25930 35284
rect 26142 35272 26148 35284
rect 26103 35244 26148 35272
rect 26142 35232 26148 35244
rect 26200 35232 26206 35284
rect 27338 35272 27344 35284
rect 27251 35244 27344 35272
rect 11235 35207 11293 35213
rect 11235 35173 11247 35207
rect 11281 35204 11293 35207
rect 11974 35204 11980 35216
rect 11281 35176 11980 35204
rect 11281 35173 11293 35176
rect 11235 35167 11293 35173
rect 11974 35164 11980 35176
rect 12032 35164 12038 35216
rect 12983 35207 13041 35213
rect 12983 35173 12995 35207
rect 13029 35204 13041 35207
rect 13354 35204 13360 35216
rect 13029 35176 13360 35204
rect 13029 35173 13041 35176
rect 12983 35167 13041 35173
rect 13354 35164 13360 35176
rect 13412 35164 13418 35216
rect 15654 35164 15660 35216
rect 15712 35204 15718 35216
rect 15927 35207 15985 35213
rect 15927 35204 15939 35207
rect 15712 35176 15939 35204
rect 15712 35164 15718 35176
rect 15927 35173 15939 35176
rect 15973 35204 15985 35207
rect 16298 35204 16304 35216
rect 15973 35176 16304 35204
rect 15973 35173 15985 35176
rect 15927 35167 15985 35173
rect 16298 35164 16304 35176
rect 16356 35164 16362 35216
rect 19334 35164 19340 35216
rect 19392 35204 19398 35216
rect 19429 35207 19487 35213
rect 19429 35204 19441 35207
rect 19392 35176 19441 35204
rect 19392 35164 19398 35176
rect 19429 35173 19441 35176
rect 19475 35173 19487 35207
rect 21082 35204 21088 35216
rect 21043 35176 21088 35204
rect 19429 35167 19487 35173
rect 21082 35164 21088 35176
rect 21140 35164 21146 35216
rect 22094 35164 22100 35216
rect 22152 35204 22158 35216
rect 22649 35207 22707 35213
rect 22649 35204 22661 35207
rect 22152 35176 22661 35204
rect 22152 35164 22158 35176
rect 22649 35173 22661 35176
rect 22695 35173 22707 35207
rect 22649 35167 22707 35173
rect 25406 35164 25412 35216
rect 25464 35204 25470 35216
rect 25593 35207 25651 35213
rect 25593 35204 25605 35207
rect 25464 35176 25605 35204
rect 25464 35164 25470 35176
rect 25593 35173 25605 35176
rect 25639 35204 25651 35207
rect 27154 35204 27160 35216
rect 25639 35176 27160 35204
rect 25639 35173 25651 35176
rect 25593 35167 25651 35173
rect 27154 35164 27160 35176
rect 27212 35164 27218 35216
rect 27264 35213 27292 35244
rect 27338 35232 27344 35244
rect 27396 35272 27402 35284
rect 27706 35272 27712 35284
rect 27396 35244 27712 35272
rect 27396 35232 27402 35244
rect 27706 35232 27712 35244
rect 27764 35232 27770 35284
rect 32858 35272 32864 35284
rect 32819 35244 32864 35272
rect 32858 35232 32864 35244
rect 32916 35232 32922 35284
rect 37553 35275 37611 35281
rect 37553 35241 37565 35275
rect 37599 35272 37611 35275
rect 37826 35272 37832 35284
rect 37599 35244 37832 35272
rect 37599 35241 37611 35244
rect 37553 35235 37611 35241
rect 37826 35232 37832 35244
rect 37884 35232 37890 35284
rect 38654 35272 38660 35284
rect 38615 35244 38660 35272
rect 38654 35232 38660 35244
rect 38712 35232 38718 35284
rect 40497 35275 40555 35281
rect 40497 35241 40509 35275
rect 40543 35241 40555 35275
rect 40497 35235 40555 35241
rect 27249 35207 27307 35213
rect 27249 35173 27261 35207
rect 27295 35173 27307 35207
rect 27249 35167 27307 35173
rect 29546 35164 29552 35216
rect 29604 35204 29610 35216
rect 29641 35207 29699 35213
rect 29641 35204 29653 35207
rect 29604 35176 29653 35204
rect 29604 35164 29610 35176
rect 29641 35173 29653 35176
rect 29687 35173 29699 35207
rect 33134 35204 33140 35216
rect 33095 35176 33140 35204
rect 29641 35167 29699 35173
rect 33134 35164 33140 35176
rect 33192 35164 33198 35216
rect 35253 35207 35311 35213
rect 35253 35173 35265 35207
rect 35299 35204 35311 35207
rect 35802 35204 35808 35216
rect 35299 35176 35808 35204
rect 35299 35173 35311 35176
rect 35253 35167 35311 35173
rect 35802 35164 35808 35176
rect 35860 35164 35866 35216
rect 35897 35207 35955 35213
rect 35897 35173 35909 35207
rect 35943 35204 35955 35207
rect 36170 35204 36176 35216
rect 35943 35176 36176 35204
rect 35943 35173 35955 35176
rect 35897 35167 35955 35173
rect 36170 35164 36176 35176
rect 36228 35204 36234 35216
rect 37918 35204 37924 35216
rect 36228 35176 37924 35204
rect 36228 35164 36234 35176
rect 37918 35164 37924 35176
rect 37976 35204 37982 35216
rect 38099 35207 38157 35213
rect 38099 35204 38111 35207
rect 37976 35176 38111 35204
rect 37976 35164 37982 35176
rect 38099 35173 38111 35176
rect 38145 35204 38157 35207
rect 39939 35207 39997 35213
rect 39939 35204 39951 35207
rect 38145 35176 39951 35204
rect 38145 35173 38157 35176
rect 38099 35167 38157 35173
rect 39939 35173 39951 35176
rect 39985 35173 39997 35207
rect 40512 35204 40540 35235
rect 40770 35232 40776 35284
rect 40828 35272 40834 35284
rect 41141 35275 41199 35281
rect 41141 35272 41153 35275
rect 40828 35244 41153 35272
rect 40828 35232 40834 35244
rect 41141 35241 41153 35244
rect 41187 35241 41199 35275
rect 41141 35235 41199 35241
rect 40862 35204 40868 35216
rect 40512 35176 40868 35204
rect 39939 35167 39997 35173
rect 40862 35164 40868 35176
rect 40920 35204 40926 35216
rect 41506 35204 41512 35216
rect 40920 35176 41512 35204
rect 40920 35164 40926 35176
rect 41506 35164 41512 35176
rect 41564 35204 41570 35216
rect 42426 35204 42432 35216
rect 41564 35176 42432 35204
rect 41564 35164 41570 35176
rect 42426 35164 42432 35176
rect 42484 35164 42490 35216
rect 10873 35139 10931 35145
rect 10873 35105 10885 35139
rect 10919 35136 10931 35139
rect 10962 35136 10968 35148
rect 10919 35108 10968 35136
rect 10919 35105 10931 35108
rect 10873 35099 10931 35105
rect 10962 35096 10968 35108
rect 11020 35096 11026 35148
rect 11793 35139 11851 35145
rect 11793 35105 11805 35139
rect 11839 35136 11851 35139
rect 12066 35136 12072 35148
rect 11839 35108 12072 35136
rect 11839 35105 11851 35108
rect 11793 35099 11851 35105
rect 12066 35096 12072 35108
rect 12124 35136 12130 35148
rect 14369 35139 14427 35145
rect 14369 35136 14381 35139
rect 12124 35108 14381 35136
rect 12124 35096 12130 35108
rect 14369 35105 14381 35108
rect 14415 35136 14427 35139
rect 14458 35136 14464 35148
rect 14415 35108 14464 35136
rect 14415 35105 14427 35108
rect 14369 35099 14427 35105
rect 14458 35096 14464 35108
rect 14516 35096 14522 35148
rect 17310 35136 17316 35148
rect 17271 35108 17316 35136
rect 17310 35096 17316 35108
rect 17368 35096 17374 35148
rect 17770 35136 17776 35148
rect 17731 35108 17776 35136
rect 17770 35096 17776 35108
rect 17828 35096 17834 35148
rect 24302 35136 24308 35148
rect 24263 35108 24308 35136
rect 24302 35096 24308 35108
rect 24360 35096 24366 35148
rect 28994 35136 29000 35148
rect 28955 35108 29000 35136
rect 28994 35096 29000 35108
rect 29052 35096 29058 35148
rect 29454 35136 29460 35148
rect 29415 35108 29460 35136
rect 29454 35096 29460 35108
rect 29512 35096 29518 35148
rect 30466 35136 30472 35148
rect 30427 35108 30472 35136
rect 30466 35096 30472 35108
rect 30524 35096 30530 35148
rect 30929 35139 30987 35145
rect 30929 35105 30941 35139
rect 30975 35105 30987 35139
rect 34514 35136 34520 35148
rect 34475 35108 34520 35136
rect 30929 35099 30987 35105
rect 12434 35028 12440 35080
rect 12492 35068 12498 35080
rect 12621 35071 12679 35077
rect 12621 35068 12633 35071
rect 12492 35040 12633 35068
rect 12492 35028 12498 35040
rect 12621 35037 12633 35040
rect 12667 35037 12679 35071
rect 15562 35068 15568 35080
rect 15523 35040 15568 35068
rect 12621 35031 12679 35037
rect 15562 35028 15568 35040
rect 15620 35028 15626 35080
rect 19153 35071 19211 35077
rect 19153 35037 19165 35071
rect 19199 35068 19211 35071
rect 19337 35071 19395 35077
rect 19337 35068 19349 35071
rect 19199 35040 19349 35068
rect 19199 35037 19211 35040
rect 19153 35031 19211 35037
rect 19337 35037 19349 35040
rect 19383 35068 19395 35071
rect 19426 35068 19432 35080
rect 19383 35040 19432 35068
rect 19383 35037 19395 35040
rect 19337 35031 19395 35037
rect 19426 35028 19432 35040
rect 19484 35028 19490 35080
rect 19613 35071 19671 35077
rect 19613 35037 19625 35071
rect 19659 35037 19671 35071
rect 20990 35068 20996 35080
rect 20951 35040 20996 35068
rect 19613 35031 19671 35037
rect 18046 34960 18052 35012
rect 18104 35000 18110 35012
rect 19628 35000 19656 35031
rect 20990 35028 20996 35040
rect 21048 35068 21054 35080
rect 21048 35040 22186 35068
rect 21048 35028 21054 35040
rect 19886 35000 19892 35012
rect 18104 34972 19892 35000
rect 18104 34960 18110 34972
rect 19886 34960 19892 34972
rect 19944 35000 19950 35012
rect 21174 35000 21180 35012
rect 19944 34972 21180 35000
rect 19944 34960 19950 34972
rect 21174 34960 21180 34972
rect 21232 35000 21238 35012
rect 21545 35003 21603 35009
rect 21545 35000 21557 35003
rect 21232 34972 21557 35000
rect 21232 34960 21238 34972
rect 21545 34969 21557 34972
rect 21591 34969 21603 35003
rect 22158 35000 22186 35040
rect 22370 35028 22376 35080
rect 22428 35068 22434 35080
rect 22557 35071 22615 35077
rect 22557 35068 22569 35071
rect 22428 35040 22569 35068
rect 22428 35028 22434 35040
rect 22557 35037 22569 35040
rect 22603 35037 22615 35071
rect 22557 35031 22615 35037
rect 22833 35071 22891 35077
rect 22833 35037 22845 35071
rect 22879 35068 22891 35071
rect 23658 35068 23664 35080
rect 22879 35040 23664 35068
rect 22879 35037 22891 35040
rect 22833 35031 22891 35037
rect 22848 35000 22876 35031
rect 23658 35028 23664 35040
rect 23716 35028 23722 35080
rect 27154 35068 27160 35080
rect 27067 35040 27160 35068
rect 27154 35028 27160 35040
rect 27212 35068 27218 35080
rect 28718 35068 28724 35080
rect 27212 35040 28724 35068
rect 27212 35028 27218 35040
rect 28718 35028 28724 35040
rect 28776 35028 28782 35080
rect 29472 35068 29500 35096
rect 30558 35068 30564 35080
rect 29472 35040 30564 35068
rect 30558 35028 30564 35040
rect 30616 35068 30622 35080
rect 30944 35068 30972 35099
rect 34514 35096 34520 35108
rect 34572 35096 34578 35148
rect 35069 35139 35127 35145
rect 35069 35105 35081 35139
rect 35115 35136 35127 35139
rect 35434 35136 35440 35148
rect 35115 35108 35440 35136
rect 35115 35105 35127 35108
rect 35069 35099 35127 35105
rect 35434 35096 35440 35108
rect 35492 35096 35498 35148
rect 35986 35096 35992 35148
rect 36044 35136 36050 35148
rect 36081 35139 36139 35145
rect 36081 35136 36093 35139
rect 36044 35108 36093 35136
rect 36044 35096 36050 35108
rect 36081 35105 36093 35108
rect 36127 35105 36139 35139
rect 36081 35099 36139 35105
rect 36541 35139 36599 35145
rect 36541 35105 36553 35139
rect 36587 35105 36599 35139
rect 36541 35099 36599 35105
rect 42061 35139 42119 35145
rect 42061 35105 42073 35139
rect 42107 35136 42119 35139
rect 42150 35136 42156 35148
rect 42107 35108 42156 35136
rect 42107 35105 42119 35108
rect 42061 35099 42119 35105
rect 31202 35068 31208 35080
rect 30616 35040 30972 35068
rect 31163 35040 31208 35068
rect 30616 35028 30622 35040
rect 31202 35028 31208 35040
rect 31260 35028 31266 35080
rect 33042 35068 33048 35080
rect 33003 35040 33048 35068
rect 33042 35028 33048 35040
rect 33100 35028 33106 35080
rect 33410 35068 33416 35080
rect 33371 35040 33416 35068
rect 33410 35028 33416 35040
rect 33468 35028 33474 35080
rect 35452 35068 35480 35096
rect 36556 35068 36584 35099
rect 35452 35040 36584 35068
rect 36817 35071 36875 35077
rect 36817 35037 36829 35071
rect 36863 35068 36875 35071
rect 37737 35071 37795 35077
rect 37737 35068 37749 35071
rect 36863 35040 37749 35068
rect 36863 35037 36875 35040
rect 36817 35031 36875 35037
rect 37737 35037 37749 35040
rect 37783 35068 37795 35071
rect 38102 35068 38108 35080
rect 37783 35040 38108 35068
rect 37783 35037 37795 35040
rect 37737 35031 37795 35037
rect 38102 35028 38108 35040
rect 38160 35028 38166 35080
rect 39574 35068 39580 35080
rect 39535 35040 39580 35068
rect 39574 35028 39580 35040
rect 39632 35028 39638 35080
rect 41414 35068 41420 35080
rect 41375 35040 41420 35068
rect 41414 35028 41420 35040
rect 41472 35028 41478 35080
rect 22158 34972 22876 35000
rect 21545 34963 21603 34969
rect 27246 34960 27252 35012
rect 27304 35000 27310 35012
rect 27709 35003 27767 35009
rect 27709 35000 27721 35003
rect 27304 34972 27721 35000
rect 27304 34960 27310 34972
rect 27709 34969 27721 34972
rect 27755 34969 27767 35003
rect 32398 35000 32404 35012
rect 32311 34972 32404 35000
rect 27709 34963 27767 34969
rect 32398 34960 32404 34972
rect 32456 35000 32462 35012
rect 33428 35000 33456 35028
rect 37182 35000 37188 35012
rect 32456 34972 33456 35000
rect 37095 34972 37188 35000
rect 32456 34960 32462 34972
rect 37182 34960 37188 34972
rect 37240 35000 37246 35012
rect 42076 35000 42104 35099
rect 42150 35096 42156 35108
rect 42208 35096 42214 35148
rect 37240 34972 42104 35000
rect 37240 34960 37246 34972
rect 16482 34932 16488 34944
rect 16443 34904 16488 34932
rect 16482 34892 16488 34904
rect 16540 34892 16546 34944
rect 23842 34932 23848 34944
rect 23803 34904 23848 34932
rect 23842 34892 23848 34904
rect 23900 34892 23906 34944
rect 28166 34932 28172 34944
rect 28127 34904 28172 34932
rect 28166 34892 28172 34904
rect 28224 34892 28230 34944
rect 1104 34842 48852 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 48852 34842
rect 1104 34768 48852 34790
rect 11701 34731 11759 34737
rect 11701 34697 11713 34731
rect 11747 34728 11759 34731
rect 11974 34728 11980 34740
rect 11747 34700 11980 34728
rect 11747 34697 11759 34700
rect 11701 34691 11759 34697
rect 11974 34688 11980 34700
rect 12032 34688 12038 34740
rect 13081 34731 13139 34737
rect 13081 34697 13093 34731
rect 13127 34728 13139 34731
rect 13446 34728 13452 34740
rect 13127 34700 13452 34728
rect 13127 34697 13139 34700
rect 13081 34691 13139 34697
rect 11333 34595 11391 34601
rect 11333 34561 11345 34595
rect 11379 34592 11391 34595
rect 12161 34595 12219 34601
rect 12161 34592 12173 34595
rect 11379 34564 12173 34592
rect 11379 34561 11391 34564
rect 11333 34555 11391 34561
rect 12161 34561 12173 34564
rect 12207 34592 12219 34595
rect 12434 34592 12440 34604
rect 12207 34564 12440 34592
rect 12207 34561 12219 34564
rect 12161 34555 12219 34561
rect 12434 34552 12440 34564
rect 12492 34552 12498 34604
rect 13096 34536 13124 34691
rect 13446 34688 13452 34700
rect 13504 34688 13510 34740
rect 14090 34728 14096 34740
rect 14051 34700 14096 34728
rect 14090 34688 14096 34700
rect 14148 34688 14154 34740
rect 14458 34728 14464 34740
rect 14419 34700 14464 34728
rect 14458 34688 14464 34700
rect 14516 34688 14522 34740
rect 14550 34688 14556 34740
rect 14608 34728 14614 34740
rect 17770 34728 17776 34740
rect 14608 34700 17776 34728
rect 14608 34688 14614 34700
rect 17770 34688 17776 34700
rect 17828 34688 17834 34740
rect 18598 34728 18604 34740
rect 18559 34700 18604 34728
rect 18598 34688 18604 34700
rect 18656 34688 18662 34740
rect 18782 34688 18788 34740
rect 18840 34728 18846 34740
rect 19245 34731 19303 34737
rect 19245 34728 19257 34731
rect 18840 34700 19257 34728
rect 18840 34688 18846 34700
rect 19245 34697 19257 34700
rect 19291 34728 19303 34731
rect 19429 34731 19487 34737
rect 19429 34728 19441 34731
rect 19291 34700 19441 34728
rect 19291 34697 19303 34700
rect 19245 34691 19303 34697
rect 19429 34697 19441 34700
rect 19475 34697 19487 34731
rect 19429 34691 19487 34697
rect 20533 34731 20591 34737
rect 20533 34697 20545 34731
rect 20579 34728 20591 34731
rect 20993 34731 21051 34737
rect 20993 34728 21005 34731
rect 20579 34700 21005 34728
rect 20579 34697 20591 34700
rect 20533 34691 20591 34697
rect 20993 34697 21005 34700
rect 21039 34728 21051 34731
rect 21082 34728 21088 34740
rect 21039 34700 21088 34728
rect 21039 34697 21051 34700
rect 20993 34691 21051 34697
rect 21082 34688 21088 34700
rect 21140 34688 21146 34740
rect 22370 34688 22376 34740
rect 22428 34728 22434 34740
rect 22925 34731 22983 34737
rect 22925 34728 22937 34731
rect 22428 34700 22937 34728
rect 22428 34688 22434 34700
rect 22925 34697 22937 34700
rect 22971 34697 22983 34731
rect 22925 34691 22983 34697
rect 24670 34688 24676 34740
rect 24728 34728 24734 34740
rect 24765 34731 24823 34737
rect 24765 34728 24777 34731
rect 24728 34700 24777 34728
rect 24728 34688 24734 34700
rect 24765 34697 24777 34700
rect 24811 34697 24823 34731
rect 25222 34728 25228 34740
rect 25183 34700 25228 34728
rect 24765 34691 24823 34697
rect 25222 34688 25228 34700
rect 25280 34688 25286 34740
rect 25332 34700 27752 34728
rect 13354 34660 13360 34672
rect 13267 34632 13360 34660
rect 13354 34620 13360 34632
rect 13412 34660 13418 34672
rect 15654 34660 15660 34672
rect 13412 34632 15660 34660
rect 13412 34620 13418 34632
rect 15654 34620 15660 34632
rect 15712 34620 15718 34672
rect 16758 34660 16764 34672
rect 16719 34632 16764 34660
rect 16758 34620 16764 34632
rect 16816 34620 16822 34672
rect 17310 34620 17316 34672
rect 17368 34660 17374 34672
rect 23385 34663 23443 34669
rect 23385 34660 23397 34663
rect 17368 34632 23397 34660
rect 17368 34620 17374 34632
rect 23385 34629 23397 34632
rect 23431 34629 23443 34663
rect 25332 34660 25360 34700
rect 23385 34623 23443 34629
rect 23768 34632 25360 34660
rect 27724 34660 27752 34700
rect 28166 34688 28172 34740
rect 28224 34728 28230 34740
rect 29411 34731 29469 34737
rect 29411 34728 29423 34731
rect 28224 34700 29423 34728
rect 28224 34688 28230 34700
rect 29411 34697 29423 34700
rect 29457 34697 29469 34731
rect 32582 34728 32588 34740
rect 29411 34691 29469 34697
rect 29794 34700 32588 34728
rect 28350 34660 28356 34672
rect 27724 34632 28356 34660
rect 14642 34592 14648 34604
rect 14603 34564 14648 34592
rect 14642 34552 14648 34564
rect 14700 34552 14706 34604
rect 15289 34595 15347 34601
rect 15289 34561 15301 34595
rect 15335 34592 15347 34595
rect 15378 34592 15384 34604
rect 15335 34564 15384 34592
rect 15335 34561 15347 34564
rect 15289 34555 15347 34561
rect 15378 34552 15384 34564
rect 15436 34592 15442 34604
rect 16209 34595 16267 34601
rect 16209 34592 16221 34595
rect 15436 34564 16221 34592
rect 15436 34552 15442 34564
rect 16209 34561 16221 34564
rect 16255 34592 16267 34595
rect 16666 34592 16672 34604
rect 16255 34564 16672 34592
rect 16255 34561 16267 34564
rect 16209 34555 16267 34561
rect 16666 34552 16672 34564
rect 16724 34552 16730 34604
rect 17770 34592 17776 34604
rect 17683 34564 17776 34592
rect 17770 34552 17776 34564
rect 17828 34592 17834 34604
rect 19150 34592 19156 34604
rect 17828 34564 19156 34592
rect 17828 34552 17834 34564
rect 19150 34552 19156 34564
rect 19208 34552 19214 34604
rect 19426 34552 19432 34604
rect 19484 34592 19490 34604
rect 22281 34595 22339 34601
rect 22281 34592 22293 34595
rect 19484 34564 22293 34592
rect 19484 34552 19490 34564
rect 22281 34561 22293 34564
rect 22327 34561 22339 34595
rect 22281 34555 22339 34561
rect 10597 34527 10655 34533
rect 10597 34493 10609 34527
rect 10643 34493 10655 34527
rect 10597 34487 10655 34493
rect 10612 34400 10640 34487
rect 10870 34484 10876 34536
rect 10928 34524 10934 34536
rect 11057 34527 11115 34533
rect 11057 34524 11069 34527
rect 10928 34496 11069 34524
rect 10928 34484 10934 34496
rect 11057 34493 11069 34496
rect 11103 34493 11115 34527
rect 11057 34487 11115 34493
rect 12596 34527 12654 34533
rect 12596 34493 12608 34527
rect 12642 34524 12654 34527
rect 13078 34524 13084 34536
rect 12642 34496 13084 34524
rect 12642 34493 12654 34496
rect 12596 34487 12654 34493
rect 13078 34484 13084 34496
rect 13136 34484 13142 34536
rect 13608 34527 13666 34533
rect 13608 34493 13620 34527
rect 13654 34524 13666 34527
rect 14090 34524 14096 34536
rect 13654 34496 14096 34524
rect 13654 34493 13666 34496
rect 13608 34487 13666 34493
rect 14090 34484 14096 34496
rect 14148 34484 14154 34536
rect 18116 34527 18174 34533
rect 18116 34493 18128 34527
rect 18162 34524 18174 34527
rect 18598 34524 18604 34536
rect 18162 34496 18604 34524
rect 18162 34493 18174 34496
rect 18116 34487 18174 34493
rect 18598 34484 18604 34496
rect 18656 34484 18662 34536
rect 19613 34527 19671 34533
rect 19613 34493 19625 34527
rect 19659 34524 19671 34527
rect 20070 34524 20076 34536
rect 19659 34496 20076 34524
rect 19659 34493 19671 34496
rect 19613 34487 19671 34493
rect 20070 34484 20076 34496
rect 20128 34484 20134 34536
rect 23400 34524 23428 34623
rect 23768 34533 23796 34632
rect 28350 34620 28356 34632
rect 28408 34660 28414 34672
rect 28994 34660 29000 34672
rect 28408 34632 29000 34660
rect 28408 34620 28414 34632
rect 28994 34620 29000 34632
rect 29052 34660 29058 34672
rect 29794 34660 29822 34700
rect 32582 34688 32588 34700
rect 32640 34688 32646 34740
rect 33042 34688 33048 34740
rect 33100 34728 33106 34740
rect 33321 34731 33379 34737
rect 33321 34728 33333 34731
rect 33100 34700 33333 34728
rect 33100 34688 33106 34700
rect 33321 34697 33333 34700
rect 33367 34697 33379 34731
rect 38102 34728 38108 34740
rect 33321 34691 33379 34697
rect 35176 34700 37964 34728
rect 38063 34700 38108 34728
rect 35176 34660 35204 34700
rect 36630 34660 36636 34672
rect 29052 34632 29822 34660
rect 31312 34632 32720 34660
rect 29052 34620 29058 34632
rect 31312 34604 31340 34632
rect 24489 34595 24547 34601
rect 24489 34561 24501 34595
rect 24535 34592 24547 34595
rect 24762 34592 24768 34604
rect 24535 34564 24768 34592
rect 24535 34561 24547 34564
rect 24489 34555 24547 34561
rect 24762 34552 24768 34564
rect 24820 34552 24826 34604
rect 25406 34592 25412 34604
rect 25367 34564 25412 34592
rect 25406 34552 25412 34564
rect 25464 34552 25470 34604
rect 26053 34595 26111 34601
rect 26053 34561 26065 34595
rect 26099 34592 26111 34595
rect 26418 34592 26424 34604
rect 26099 34564 26424 34592
rect 26099 34561 26111 34564
rect 26053 34555 26111 34561
rect 26418 34552 26424 34564
rect 26476 34552 26482 34604
rect 26697 34595 26755 34601
rect 26697 34561 26709 34595
rect 26743 34592 26755 34595
rect 27338 34592 27344 34604
rect 26743 34564 27344 34592
rect 26743 34561 26755 34564
rect 26697 34555 26755 34561
rect 27338 34552 27344 34564
rect 27396 34552 27402 34604
rect 27522 34552 27528 34604
rect 27580 34592 27586 34604
rect 27617 34595 27675 34601
rect 27617 34592 27629 34595
rect 27580 34564 27629 34592
rect 27580 34552 27586 34564
rect 27617 34561 27629 34564
rect 27663 34561 27675 34595
rect 27617 34555 27675 34561
rect 28534 34552 28540 34604
rect 28592 34592 28598 34604
rect 28629 34595 28687 34601
rect 28629 34592 28641 34595
rect 28592 34564 28641 34592
rect 28592 34552 28598 34564
rect 28629 34561 28641 34564
rect 28675 34592 28687 34595
rect 29454 34592 29460 34604
rect 28675 34564 29460 34592
rect 28675 34561 28687 34564
rect 28629 34555 28687 34561
rect 29454 34552 29460 34564
rect 29512 34552 29518 34604
rect 31294 34592 31300 34604
rect 31255 34564 31300 34592
rect 31294 34552 31300 34564
rect 31352 34552 31358 34604
rect 31665 34595 31723 34601
rect 31665 34561 31677 34595
rect 31711 34592 31723 34595
rect 31754 34592 31760 34604
rect 31711 34564 31760 34592
rect 31711 34561 31723 34564
rect 31665 34555 31723 34561
rect 23753 34527 23811 34533
rect 23753 34524 23765 34527
rect 23400 34496 23765 34524
rect 23753 34493 23765 34496
rect 23799 34493 23811 34527
rect 23753 34487 23811 34493
rect 23842 34484 23848 34536
rect 23900 34524 23906 34536
rect 24305 34527 24363 34533
rect 24305 34524 24317 34527
rect 23900 34496 24317 34524
rect 23900 34484 23906 34496
rect 24305 34493 24317 34496
rect 24351 34524 24363 34527
rect 24946 34524 24952 34536
rect 24351 34496 24952 34524
rect 24351 34493 24363 34496
rect 24305 34487 24363 34493
rect 24946 34484 24952 34496
rect 25004 34484 25010 34536
rect 29340 34527 29398 34533
rect 29340 34524 29352 34527
rect 28966 34496 29352 34524
rect 14458 34416 14464 34468
rect 14516 34456 14522 34468
rect 14737 34459 14795 34465
rect 14737 34456 14749 34459
rect 14516 34428 14749 34456
rect 14516 34416 14522 34428
rect 14737 34425 14749 34428
rect 14783 34425 14795 34459
rect 14737 34419 14795 34425
rect 16301 34459 16359 34465
rect 16301 34425 16313 34459
rect 16347 34456 16359 34459
rect 16482 34456 16488 34468
rect 16347 34428 16488 34456
rect 16347 34425 16359 34428
rect 16301 34419 16359 34425
rect 10505 34391 10563 34397
rect 10505 34357 10517 34391
rect 10551 34388 10563 34391
rect 10594 34388 10600 34400
rect 10551 34360 10600 34388
rect 10551 34357 10563 34360
rect 10505 34351 10563 34357
rect 10594 34348 10600 34360
rect 10652 34348 10658 34400
rect 12667 34391 12725 34397
rect 12667 34357 12679 34391
rect 12713 34388 12725 34391
rect 12894 34388 12900 34400
rect 12713 34360 12900 34388
rect 12713 34357 12725 34360
rect 12667 34351 12725 34357
rect 12894 34348 12900 34360
rect 12952 34348 12958 34400
rect 13679 34391 13737 34397
rect 13679 34357 13691 34391
rect 13725 34388 13737 34391
rect 13906 34388 13912 34400
rect 13725 34360 13912 34388
rect 13725 34357 13737 34360
rect 13679 34351 13737 34357
rect 13906 34348 13912 34360
rect 13964 34348 13970 34400
rect 16025 34391 16083 34397
rect 16025 34357 16037 34391
rect 16071 34388 16083 34391
rect 16316 34388 16344 34419
rect 16482 34416 16488 34428
rect 16540 34416 16546 34468
rect 19242 34456 19248 34468
rect 19155 34428 19248 34456
rect 19242 34416 19248 34428
rect 19300 34456 19306 34468
rect 19426 34456 19432 34468
rect 19300 34428 19432 34456
rect 19300 34416 19306 34428
rect 19426 34416 19432 34428
rect 19484 34456 19490 34468
rect 19934 34459 19992 34465
rect 19934 34456 19946 34459
rect 19484 34428 19946 34456
rect 19484 34416 19490 34428
rect 19934 34425 19946 34428
rect 19980 34425 19992 34459
rect 19934 34419 19992 34425
rect 21453 34459 21511 34465
rect 21453 34425 21465 34459
rect 21499 34456 21511 34459
rect 22002 34456 22008 34468
rect 21499 34428 22008 34456
rect 21499 34425 21511 34428
rect 21453 34419 21511 34425
rect 22002 34416 22008 34428
rect 22060 34416 22066 34468
rect 22094 34416 22100 34468
rect 22152 34456 22158 34468
rect 25501 34459 25559 34465
rect 22152 34428 22197 34456
rect 22152 34416 22158 34428
rect 25501 34425 25513 34459
rect 25547 34425 25559 34459
rect 25501 34419 25559 34425
rect 27249 34459 27307 34465
rect 27249 34425 27261 34459
rect 27295 34425 27307 34459
rect 27249 34419 27307 34425
rect 16071 34360 16344 34388
rect 16071 34357 16083 34360
rect 16025 34351 16083 34357
rect 16574 34348 16580 34400
rect 16632 34388 16638 34400
rect 17310 34388 17316 34400
rect 16632 34360 17316 34388
rect 16632 34348 16638 34360
rect 17310 34348 17316 34360
rect 17368 34348 17374 34400
rect 17770 34348 17776 34400
rect 17828 34388 17834 34400
rect 18187 34391 18245 34397
rect 18187 34388 18199 34391
rect 17828 34360 18199 34388
rect 17828 34348 17834 34360
rect 18187 34357 18199 34360
rect 18233 34357 18245 34391
rect 18187 34351 18245 34357
rect 19153 34391 19211 34397
rect 19153 34357 19165 34391
rect 19199 34388 19211 34391
rect 19334 34388 19340 34400
rect 19199 34360 19340 34388
rect 19199 34357 19211 34360
rect 19153 34351 19211 34357
rect 19334 34348 19340 34360
rect 19392 34348 19398 34400
rect 21821 34391 21879 34397
rect 21821 34357 21833 34391
rect 21867 34388 21879 34391
rect 22112 34388 22140 34416
rect 21867 34360 22140 34388
rect 21867 34357 21879 34360
rect 21821 34351 21879 34357
rect 25222 34348 25228 34400
rect 25280 34388 25286 34400
rect 25516 34388 25544 34419
rect 26970 34388 26976 34400
rect 25280 34360 25544 34388
rect 26931 34360 26976 34388
rect 25280 34348 25286 34360
rect 26970 34348 26976 34360
rect 27028 34388 27034 34400
rect 27264 34388 27292 34419
rect 27338 34416 27344 34468
rect 27396 34456 27402 34468
rect 27396 34428 27441 34456
rect 27396 34416 27402 34428
rect 27706 34416 27712 34468
rect 27764 34456 27770 34468
rect 28966 34456 28994 34496
rect 29340 34493 29352 34496
rect 29386 34524 29398 34527
rect 29386 34496 29868 34524
rect 29386 34493 29398 34496
rect 29340 34487 29398 34493
rect 27764 34428 28994 34456
rect 27764 34416 27770 34428
rect 27028 34360 27292 34388
rect 27356 34388 27384 34416
rect 29840 34400 29868 34496
rect 30466 34456 30472 34468
rect 30427 34428 30472 34456
rect 30466 34416 30472 34428
rect 30524 34416 30530 34468
rect 30653 34459 30711 34465
rect 30653 34425 30665 34459
rect 30699 34425 30711 34459
rect 30653 34419 30711 34425
rect 28169 34391 28227 34397
rect 28169 34388 28181 34391
rect 27356 34360 28181 34388
rect 27028 34348 27034 34360
rect 28169 34357 28181 34360
rect 28215 34357 28227 34391
rect 29822 34388 29828 34400
rect 29783 34360 29828 34388
rect 28169 34351 28227 34357
rect 29822 34348 29828 34360
rect 29880 34348 29886 34400
rect 30668 34388 30696 34419
rect 30742 34416 30748 34468
rect 30800 34456 30806 34468
rect 30800 34428 30845 34456
rect 30800 34416 30806 34428
rect 31680 34388 31708 34555
rect 31754 34552 31760 34564
rect 31812 34552 31818 34604
rect 32398 34592 32404 34604
rect 32359 34564 32404 34592
rect 32398 34552 32404 34564
rect 32456 34552 32462 34604
rect 32692 34601 32720 34632
rect 33106 34632 35204 34660
rect 35268 34632 36636 34660
rect 32677 34595 32735 34601
rect 32677 34561 32689 34595
rect 32723 34592 32735 34595
rect 33106 34592 33134 34632
rect 32723 34564 33134 34592
rect 32723 34561 32735 34564
rect 32677 34555 32735 34561
rect 35268 34533 35296 34632
rect 36630 34620 36636 34632
rect 36688 34620 36694 34672
rect 37936 34660 37964 34700
rect 38102 34688 38108 34700
rect 38160 34688 38166 34740
rect 41417 34731 41475 34737
rect 41417 34697 41429 34731
rect 41463 34728 41475 34731
rect 41506 34728 41512 34740
rect 41463 34700 41512 34728
rect 41463 34697 41475 34700
rect 41417 34691 41475 34697
rect 41506 34688 41512 34700
rect 41564 34688 41570 34740
rect 41690 34688 41696 34740
rect 41748 34728 41754 34740
rect 41831 34731 41889 34737
rect 41831 34728 41843 34731
rect 41748 34700 41843 34728
rect 41748 34688 41754 34700
rect 41831 34697 41843 34700
rect 41877 34697 41889 34731
rect 41831 34691 41889 34697
rect 41966 34660 41972 34672
rect 37936 34632 41972 34660
rect 41966 34620 41972 34632
rect 42024 34620 42030 34672
rect 35526 34592 35532 34604
rect 35487 34564 35532 34592
rect 35526 34552 35532 34564
rect 35584 34552 35590 34604
rect 36446 34552 36452 34604
rect 36504 34592 36510 34604
rect 36906 34592 36912 34604
rect 36504 34564 36912 34592
rect 36504 34552 36510 34564
rect 36906 34552 36912 34564
rect 36964 34552 36970 34604
rect 37829 34595 37887 34601
rect 37829 34561 37841 34595
rect 37875 34592 37887 34595
rect 37918 34592 37924 34604
rect 37875 34564 37924 34592
rect 37875 34561 37887 34564
rect 37829 34555 37887 34561
rect 37918 34552 37924 34564
rect 37976 34552 37982 34604
rect 39574 34592 39580 34604
rect 39487 34564 39580 34592
rect 39574 34552 39580 34564
rect 39632 34592 39638 34604
rect 40221 34595 40279 34601
rect 40221 34592 40233 34595
rect 39632 34564 40233 34592
rect 39632 34552 39638 34564
rect 40221 34561 40233 34564
rect 40267 34561 40279 34595
rect 40221 34555 40279 34561
rect 40681 34595 40739 34601
rect 40681 34561 40693 34595
rect 40727 34592 40739 34595
rect 42058 34592 42064 34604
rect 40727 34564 42064 34592
rect 40727 34561 40739 34564
rect 40681 34555 40739 34561
rect 42058 34552 42064 34564
rect 42116 34552 42122 34604
rect 34701 34527 34759 34533
rect 34701 34493 34713 34527
rect 34747 34524 34759 34527
rect 35253 34527 35311 34533
rect 35253 34524 35265 34527
rect 34747 34496 35265 34524
rect 34747 34493 34759 34496
rect 34701 34487 34759 34493
rect 35253 34493 35265 34496
rect 35299 34493 35311 34527
rect 35434 34524 35440 34536
rect 35395 34496 35440 34524
rect 35253 34487 35311 34493
rect 35434 34484 35440 34496
rect 35492 34484 35498 34536
rect 38841 34527 38899 34533
rect 38841 34493 38853 34527
rect 38887 34493 38899 34527
rect 39298 34524 39304 34536
rect 39259 34496 39304 34524
rect 38841 34487 38899 34493
rect 32493 34459 32551 34465
rect 32493 34425 32505 34459
rect 32539 34425 32551 34459
rect 32493 34419 32551 34425
rect 32122 34388 32128 34400
rect 30668 34360 31708 34388
rect 32083 34360 32128 34388
rect 32122 34348 32128 34360
rect 32180 34388 32186 34400
rect 32508 34388 32536 34419
rect 32582 34416 32588 34468
rect 32640 34456 32646 34468
rect 34333 34459 34391 34465
rect 34333 34456 34345 34459
rect 32640 34428 34345 34456
rect 32640 34416 32646 34428
rect 34333 34425 34345 34428
rect 34379 34456 34391 34459
rect 34514 34456 34520 34468
rect 34379 34428 34520 34456
rect 34379 34425 34391 34428
rect 34333 34419 34391 34425
rect 34514 34416 34520 34428
rect 34572 34456 34578 34468
rect 35894 34456 35900 34468
rect 34572 34428 35900 34456
rect 34572 34416 34578 34428
rect 35894 34416 35900 34428
rect 35952 34416 35958 34468
rect 36633 34459 36691 34465
rect 36633 34425 36645 34459
rect 36679 34425 36691 34459
rect 36633 34419 36691 34425
rect 32180 34360 32536 34388
rect 32180 34348 32186 34360
rect 33134 34348 33140 34400
rect 33192 34388 33198 34400
rect 33689 34391 33747 34397
rect 33689 34388 33701 34391
rect 33192 34360 33701 34388
rect 33192 34348 33198 34360
rect 33689 34357 33701 34360
rect 33735 34357 33747 34391
rect 33689 34351 33747 34357
rect 35986 34348 35992 34400
rect 36044 34388 36050 34400
rect 36081 34391 36139 34397
rect 36081 34388 36093 34391
rect 36044 34360 36093 34388
rect 36044 34348 36050 34360
rect 36081 34357 36093 34360
rect 36127 34357 36139 34391
rect 36648 34388 36676 34419
rect 36722 34416 36728 34468
rect 36780 34456 36786 34468
rect 38654 34456 38660 34468
rect 36780 34428 36825 34456
rect 38615 34428 38660 34456
rect 36780 34416 36786 34428
rect 38654 34416 38660 34428
rect 38712 34456 38718 34468
rect 38856 34456 38884 34487
rect 39298 34484 39304 34496
rect 39356 34484 39362 34536
rect 41760 34527 41818 34533
rect 41760 34493 41772 34527
rect 41806 34524 41818 34527
rect 41806 34496 42288 34524
rect 41806 34493 41818 34496
rect 41760 34487 41818 34493
rect 38712 34428 38884 34456
rect 38712 34416 38718 34428
rect 42260 34400 42288 34496
rect 42426 34484 42432 34536
rect 42484 34524 42490 34536
rect 42740 34527 42798 34533
rect 42740 34524 42752 34527
rect 42484 34496 42752 34524
rect 42484 34484 42490 34496
rect 42740 34493 42752 34496
rect 42786 34524 42798 34527
rect 43165 34527 43223 34533
rect 43165 34524 43177 34527
rect 42786 34496 43177 34524
rect 42786 34493 42798 34496
rect 42740 34487 42798 34493
rect 43165 34493 43177 34496
rect 43211 34493 43223 34527
rect 43165 34487 43223 34493
rect 37182 34388 37188 34400
rect 36648 34360 37188 34388
rect 36081 34351 36139 34357
rect 37182 34348 37188 34360
rect 37240 34348 37246 34400
rect 39945 34391 40003 34397
rect 39945 34357 39957 34391
rect 39991 34388 40003 34391
rect 40126 34388 40132 34400
rect 39991 34360 40132 34388
rect 39991 34357 40003 34360
rect 39945 34351 40003 34357
rect 40126 34348 40132 34360
rect 40184 34348 40190 34400
rect 42242 34388 42248 34400
rect 42203 34360 42248 34388
rect 42242 34348 42248 34360
rect 42300 34348 42306 34400
rect 42334 34348 42340 34400
rect 42392 34388 42398 34400
rect 42843 34391 42901 34397
rect 42843 34388 42855 34391
rect 42392 34360 42855 34388
rect 42392 34348 42398 34360
rect 42843 34357 42855 34360
rect 42889 34357 42901 34391
rect 42843 34351 42901 34357
rect 1104 34298 48852 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 48852 34298
rect 1104 34224 48852 34246
rect 10962 34184 10968 34196
rect 10923 34156 10968 34184
rect 10962 34144 10968 34156
rect 11020 34144 11026 34196
rect 14642 34184 14648 34196
rect 14603 34156 14648 34184
rect 14642 34144 14648 34156
rect 14700 34144 14706 34196
rect 15562 34184 15568 34196
rect 15371 34156 15568 34184
rect 10689 34119 10747 34125
rect 10689 34085 10701 34119
rect 10735 34116 10747 34119
rect 10870 34116 10876 34128
rect 10735 34088 10876 34116
rect 10735 34085 10747 34088
rect 10689 34079 10747 34085
rect 10870 34076 10876 34088
rect 10928 34076 10934 34128
rect 14369 34119 14427 34125
rect 14369 34085 14381 34119
rect 14415 34116 14427 34119
rect 15371 34116 15399 34156
rect 15562 34144 15568 34156
rect 15620 34184 15626 34196
rect 16301 34187 16359 34193
rect 16301 34184 16313 34187
rect 15620 34156 16313 34184
rect 15620 34144 15626 34156
rect 16301 34153 16313 34156
rect 16347 34153 16359 34187
rect 16666 34184 16672 34196
rect 16627 34156 16672 34184
rect 16301 34147 16359 34153
rect 16666 34144 16672 34156
rect 16724 34144 16730 34196
rect 19242 34184 19248 34196
rect 19203 34156 19248 34184
rect 19242 34144 19248 34156
rect 19300 34144 19306 34196
rect 19334 34144 19340 34196
rect 19392 34184 19398 34196
rect 19797 34187 19855 34193
rect 19797 34184 19809 34187
rect 19392 34156 19809 34184
rect 19392 34144 19398 34156
rect 19797 34153 19809 34156
rect 19843 34153 19855 34187
rect 20070 34184 20076 34196
rect 20031 34156 20076 34184
rect 19797 34147 19855 34153
rect 20070 34144 20076 34156
rect 20128 34144 20134 34196
rect 20990 34144 20996 34196
rect 21048 34184 21054 34196
rect 21085 34187 21143 34193
rect 21085 34184 21097 34187
rect 21048 34156 21097 34184
rect 21048 34144 21054 34156
rect 21085 34153 21097 34156
rect 21131 34153 21143 34187
rect 21818 34184 21824 34196
rect 21779 34156 21824 34184
rect 21085 34147 21143 34153
rect 21818 34144 21824 34156
rect 21876 34144 21882 34196
rect 22094 34144 22100 34196
rect 22152 34184 22158 34196
rect 22373 34187 22431 34193
rect 22373 34184 22385 34187
rect 22152 34156 22385 34184
rect 22152 34144 22158 34156
rect 22373 34153 22385 34156
rect 22419 34184 22431 34187
rect 22649 34187 22707 34193
rect 22649 34184 22661 34187
rect 22419 34156 22661 34184
rect 22419 34153 22431 34156
rect 22373 34147 22431 34153
rect 22649 34153 22661 34156
rect 22695 34153 22707 34187
rect 24302 34184 24308 34196
rect 24263 34156 24308 34184
rect 22649 34147 22707 34153
rect 24302 34144 24308 34156
rect 24360 34144 24366 34196
rect 27065 34187 27123 34193
rect 27065 34153 27077 34187
rect 27111 34184 27123 34187
rect 27154 34184 27160 34196
rect 27111 34156 27160 34184
rect 27111 34153 27123 34156
rect 27065 34147 27123 34153
rect 27154 34144 27160 34156
rect 27212 34144 27218 34196
rect 30377 34187 30435 34193
rect 30377 34153 30389 34187
rect 30423 34184 30435 34187
rect 30742 34184 30748 34196
rect 30423 34156 30748 34184
rect 30423 34153 30435 34156
rect 30377 34147 30435 34153
rect 30742 34144 30748 34156
rect 30800 34184 30806 34196
rect 31021 34187 31079 34193
rect 31021 34184 31033 34187
rect 30800 34156 31033 34184
rect 30800 34144 30806 34156
rect 31021 34153 31033 34156
rect 31067 34153 31079 34187
rect 31021 34147 31079 34153
rect 33042 34144 33048 34196
rect 33100 34184 33106 34196
rect 33873 34187 33931 34193
rect 33873 34184 33885 34187
rect 33100 34156 33885 34184
rect 33100 34144 33106 34156
rect 33873 34153 33885 34156
rect 33919 34153 33931 34187
rect 33873 34147 33931 34153
rect 36449 34187 36507 34193
rect 36449 34153 36461 34187
rect 36495 34184 36507 34187
rect 36722 34184 36728 34196
rect 36495 34156 36728 34184
rect 36495 34153 36507 34156
rect 36449 34147 36507 34153
rect 36722 34144 36728 34156
rect 36780 34184 36786 34196
rect 37093 34187 37151 34193
rect 37093 34184 37105 34187
rect 36780 34156 37105 34184
rect 36780 34144 36786 34156
rect 37093 34153 37105 34156
rect 37139 34153 37151 34187
rect 41414 34184 41420 34196
rect 41375 34156 41420 34184
rect 37093 34147 37151 34153
rect 41414 34144 41420 34156
rect 41472 34184 41478 34196
rect 42334 34184 42340 34196
rect 41472 34156 42340 34184
rect 41472 34144 41478 34156
rect 42334 34144 42340 34156
rect 42392 34144 42398 34196
rect 15470 34116 15476 34128
rect 14415 34088 15399 34116
rect 15431 34088 15476 34116
rect 14415 34085 14427 34088
rect 14369 34079 14427 34085
rect 15470 34076 15476 34088
rect 15528 34076 15534 34128
rect 23845 34119 23903 34125
rect 23845 34085 23857 34119
rect 23891 34116 23903 34119
rect 26970 34116 26976 34128
rect 23891 34088 26976 34116
rect 23891 34085 23903 34088
rect 23845 34079 23903 34085
rect 26970 34076 26976 34088
rect 27028 34076 27034 34128
rect 27338 34116 27344 34128
rect 27299 34088 27344 34116
rect 27338 34076 27344 34088
rect 27396 34076 27402 34128
rect 29638 34076 29644 34128
rect 29696 34116 29702 34128
rect 29778 34119 29836 34125
rect 29778 34116 29790 34119
rect 29696 34088 29790 34116
rect 29696 34076 29702 34088
rect 29778 34085 29790 34088
rect 29824 34085 29836 34119
rect 29778 34079 29836 34085
rect 30558 34076 30564 34128
rect 30616 34116 30622 34128
rect 30653 34119 30711 34125
rect 30653 34116 30665 34119
rect 30616 34088 30665 34116
rect 30616 34076 30622 34088
rect 30653 34085 30665 34088
rect 30699 34085 30711 34119
rect 30653 34079 30711 34085
rect 32306 34076 32312 34128
rect 32364 34116 32370 34128
rect 32446 34119 32504 34125
rect 32446 34116 32458 34119
rect 32364 34088 32458 34116
rect 32364 34076 32370 34088
rect 32446 34085 32458 34088
rect 32492 34085 32504 34119
rect 32446 34079 32504 34085
rect 35891 34119 35949 34125
rect 35891 34085 35903 34119
rect 35937 34116 35949 34119
rect 36538 34116 36544 34128
rect 35937 34088 36544 34116
rect 35937 34085 35949 34088
rect 35891 34079 35949 34085
rect 36538 34076 36544 34088
rect 36596 34116 36602 34128
rect 37918 34116 37924 34128
rect 36596 34088 37924 34116
rect 36596 34076 36602 34088
rect 37918 34076 37924 34088
rect 37976 34076 37982 34128
rect 38194 34116 38200 34128
rect 38073 34088 38200 34116
rect 11882 34048 11888 34060
rect 11843 34020 11888 34048
rect 11882 34008 11888 34020
rect 11940 34008 11946 34060
rect 13722 34048 13728 34060
rect 13683 34020 13728 34048
rect 13722 34008 13728 34020
rect 13780 34008 13786 34060
rect 14090 34008 14096 34060
rect 14148 34048 14154 34060
rect 14185 34051 14243 34057
rect 14185 34048 14197 34051
rect 14148 34020 14197 34048
rect 14148 34008 14154 34020
rect 14185 34017 14197 34020
rect 14231 34048 14243 34051
rect 14550 34048 14556 34060
rect 14231 34020 14556 34048
rect 14231 34017 14243 34020
rect 14185 34011 14243 34017
rect 14550 34008 14556 34020
rect 14608 34008 14614 34060
rect 16920 34051 16978 34057
rect 16920 34017 16932 34051
rect 16966 34048 16978 34051
rect 17494 34048 17500 34060
rect 16966 34020 17500 34048
rect 16966 34017 16978 34020
rect 16920 34011 16978 34017
rect 17494 34008 17500 34020
rect 17552 34008 17558 34060
rect 17932 34051 17990 34057
rect 17932 34017 17944 34051
rect 17978 34048 17990 34051
rect 18046 34048 18052 34060
rect 17978 34020 18052 34048
rect 17978 34017 17990 34020
rect 17932 34011 17990 34017
rect 18046 34008 18052 34020
rect 18104 34008 18110 34060
rect 24857 34051 24915 34057
rect 24857 34017 24869 34051
rect 24903 34017 24915 34051
rect 24857 34011 24915 34017
rect 15378 33980 15384 33992
rect 15339 33952 15384 33980
rect 15378 33940 15384 33952
rect 15436 33940 15442 33992
rect 18874 33980 18880 33992
rect 18835 33952 18880 33980
rect 18874 33940 18880 33952
rect 18932 33940 18938 33992
rect 21450 33980 21456 33992
rect 21411 33952 21456 33980
rect 21450 33940 21456 33952
rect 21508 33940 21514 33992
rect 24872 33980 24900 34011
rect 24946 34008 24952 34060
rect 25004 34048 25010 34060
rect 25317 34051 25375 34057
rect 25317 34048 25329 34051
rect 25004 34020 25329 34048
rect 25004 34008 25010 34020
rect 25317 34017 25329 34020
rect 25363 34017 25375 34051
rect 25682 34048 25688 34060
rect 25317 34011 25375 34017
rect 25424 34020 25688 34048
rect 25424 33980 25452 34020
rect 25682 34008 25688 34020
rect 25740 34008 25746 34060
rect 31202 34008 31208 34060
rect 31260 34048 31266 34060
rect 32125 34051 32183 34057
rect 32125 34048 32137 34051
rect 31260 34020 32137 34048
rect 31260 34008 31266 34020
rect 32125 34017 32137 34020
rect 32171 34048 32183 34051
rect 33870 34048 33876 34060
rect 32171 34020 33876 34048
rect 32171 34017 32183 34020
rect 32125 34011 32183 34017
rect 33870 34008 33876 34020
rect 33928 34008 33934 34060
rect 35618 34008 35624 34060
rect 35676 34048 35682 34060
rect 38073 34057 38101 34088
rect 38194 34076 38200 34088
rect 38252 34076 38258 34128
rect 38654 34076 38660 34128
rect 38712 34116 38718 34128
rect 38712 34088 41736 34116
rect 38712 34076 38718 34088
rect 41708 34060 41736 34088
rect 38059 34051 38117 34057
rect 38059 34048 38071 34051
rect 35676 34020 38071 34048
rect 35676 34008 35682 34020
rect 38059 34017 38071 34020
rect 38105 34017 38117 34051
rect 39022 34048 39028 34060
rect 38983 34020 39028 34048
rect 38059 34011 38117 34017
rect 39022 34008 39028 34020
rect 39080 34008 39086 34060
rect 39390 34008 39396 34060
rect 39448 34048 39454 34060
rect 39485 34051 39543 34057
rect 39485 34048 39497 34051
rect 39448 34020 39497 34048
rect 39448 34008 39454 34020
rect 39485 34017 39497 34020
rect 39531 34017 39543 34051
rect 39485 34011 39543 34017
rect 40310 34008 40316 34060
rect 40368 34048 40374 34060
rect 40624 34051 40682 34057
rect 40624 34048 40636 34051
rect 40368 34020 40636 34048
rect 40368 34008 40374 34020
rect 40624 34017 40636 34020
rect 40670 34017 40682 34051
rect 41690 34048 41696 34060
rect 41603 34020 41696 34048
rect 40624 34011 40682 34017
rect 41690 34008 41696 34020
rect 41748 34008 41754 34060
rect 42150 34048 42156 34060
rect 42111 34020 42156 34048
rect 42150 34008 42156 34020
rect 42208 34008 42214 34060
rect 25590 33980 25596 33992
rect 24872 33952 25452 33980
rect 25551 33952 25596 33980
rect 25590 33940 25596 33952
rect 25648 33940 25654 33992
rect 27249 33983 27307 33989
rect 27249 33949 27261 33983
rect 27295 33980 27307 33983
rect 27614 33980 27620 33992
rect 27295 33952 27620 33980
rect 27295 33949 27307 33952
rect 27249 33943 27307 33949
rect 27614 33940 27620 33952
rect 27672 33940 27678 33992
rect 29454 33980 29460 33992
rect 29415 33952 29460 33980
rect 29454 33940 29460 33952
rect 29512 33940 29518 33992
rect 35526 33980 35532 33992
rect 35487 33952 35532 33980
rect 35526 33940 35532 33952
rect 35584 33940 35590 33992
rect 38151 33983 38209 33989
rect 38151 33949 38163 33983
rect 38197 33980 38209 33983
rect 38470 33980 38476 33992
rect 38197 33952 38476 33980
rect 38197 33949 38209 33952
rect 38151 33943 38209 33949
rect 38470 33940 38476 33952
rect 38528 33940 38534 33992
rect 39758 33980 39764 33992
rect 39719 33952 39764 33980
rect 39758 33940 39764 33952
rect 39816 33940 39822 33992
rect 42429 33983 42487 33989
rect 42429 33949 42441 33983
rect 42475 33980 42487 33983
rect 42610 33980 42616 33992
rect 42475 33952 42616 33980
rect 42475 33949 42487 33952
rect 42429 33943 42487 33949
rect 42610 33940 42616 33952
rect 42668 33940 42674 33992
rect 15930 33912 15936 33924
rect 15891 33884 15936 33912
rect 15930 33872 15936 33884
rect 15988 33872 15994 33924
rect 16758 33872 16764 33924
rect 16816 33912 16822 33924
rect 18003 33915 18061 33921
rect 18003 33912 18015 33915
rect 16816 33884 18015 33912
rect 16816 33872 16822 33884
rect 18003 33881 18015 33884
rect 18049 33881 18061 33915
rect 18003 33875 18061 33881
rect 22186 33872 22192 33924
rect 22244 33912 22250 33924
rect 23290 33912 23296 33924
rect 22244 33884 23296 33912
rect 22244 33872 22250 33884
rect 23290 33872 23296 33884
rect 23348 33912 23354 33924
rect 27706 33912 27712 33924
rect 23348 33884 27712 33912
rect 23348 33872 23354 33884
rect 27706 33872 27712 33884
rect 27764 33872 27770 33924
rect 27798 33872 27804 33924
rect 27856 33912 27862 33924
rect 27856 33884 27901 33912
rect 27856 33872 27862 33884
rect 31754 33872 31760 33924
rect 31812 33912 31818 33924
rect 33318 33912 33324 33924
rect 31812 33884 33324 33912
rect 31812 33872 31818 33884
rect 33318 33872 33324 33884
rect 33376 33872 33382 33924
rect 34514 33912 34520 33924
rect 34475 33884 34520 33912
rect 34514 33872 34520 33884
rect 34572 33912 34578 33924
rect 34977 33915 35035 33921
rect 34977 33912 34989 33915
rect 34572 33884 34989 33912
rect 34572 33872 34578 33884
rect 34977 33881 34989 33884
rect 35023 33912 35035 33915
rect 35434 33912 35440 33924
rect 35023 33884 35440 33912
rect 35023 33881 35035 33884
rect 34977 33875 35035 33881
rect 35434 33872 35440 33884
rect 35492 33912 35498 33924
rect 36725 33915 36783 33921
rect 36725 33912 36737 33915
rect 35492 33884 36737 33912
rect 35492 33872 35498 33884
rect 36725 33881 36737 33884
rect 36771 33912 36783 33915
rect 38841 33915 38899 33921
rect 38841 33912 38853 33915
rect 36771 33884 38853 33912
rect 36771 33881 36783 33884
rect 36725 33875 36783 33881
rect 38841 33881 38853 33884
rect 38887 33912 38899 33915
rect 39298 33912 39304 33924
rect 38887 33884 39304 33912
rect 38887 33881 38899 33884
rect 38841 33875 38899 33881
rect 39298 33872 39304 33884
rect 39356 33872 39362 33924
rect 12023 33847 12081 33853
rect 12023 33813 12035 33847
rect 12069 33844 12081 33847
rect 12437 33847 12495 33853
rect 12437 33844 12449 33847
rect 12069 33816 12449 33844
rect 12069 33813 12081 33816
rect 12023 33807 12081 33813
rect 12437 33813 12449 33816
rect 12483 33844 12495 33847
rect 12526 33844 12532 33856
rect 12483 33816 12532 33844
rect 12483 33813 12495 33816
rect 12437 33807 12495 33813
rect 12526 33804 12532 33816
rect 12584 33804 12590 33856
rect 16991 33847 17049 33853
rect 16991 33813 17003 33847
rect 17037 33844 17049 33847
rect 17862 33844 17868 33856
rect 17037 33816 17868 33844
rect 17037 33813 17049 33816
rect 16991 33807 17049 33813
rect 17862 33804 17868 33816
rect 17920 33804 17926 33856
rect 18414 33844 18420 33856
rect 18375 33816 18420 33844
rect 18414 33804 18420 33816
rect 18472 33804 18478 33856
rect 22922 33804 22928 33856
rect 22980 33844 22986 33856
rect 27522 33844 27528 33856
rect 22980 33816 27528 33844
rect 22980 33804 22986 33816
rect 27522 33804 27528 33816
rect 27580 33804 27586 33856
rect 33042 33844 33048 33856
rect 33003 33816 33048 33844
rect 33042 33804 33048 33816
rect 33100 33804 33106 33856
rect 37918 33804 37924 33856
rect 37976 33844 37982 33856
rect 40770 33853 40776 33856
rect 38473 33847 38531 33853
rect 38473 33844 38485 33847
rect 37976 33816 38485 33844
rect 37976 33804 37982 33816
rect 38473 33813 38485 33816
rect 38519 33813 38531 33847
rect 38473 33807 38531 33813
rect 40497 33847 40555 33853
rect 40497 33813 40509 33847
rect 40543 33844 40555 33847
rect 40727 33847 40776 33853
rect 40727 33844 40739 33847
rect 40543 33816 40739 33844
rect 40543 33813 40555 33816
rect 40497 33807 40555 33813
rect 40727 33813 40739 33816
rect 40773 33813 40776 33847
rect 40727 33807 40776 33813
rect 40770 33804 40776 33807
rect 40828 33804 40834 33856
rect 43622 33844 43628 33856
rect 43583 33816 43628 33844
rect 43622 33804 43628 33816
rect 43680 33804 43686 33856
rect 1104 33754 48852 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 48852 33754
rect 1104 33680 48852 33702
rect 10502 33640 10508 33652
rect 10463 33612 10508 33640
rect 10502 33600 10508 33612
rect 10560 33600 10566 33652
rect 11882 33640 11888 33652
rect 11843 33612 11888 33640
rect 11882 33600 11888 33612
rect 11940 33600 11946 33652
rect 13722 33640 13728 33652
rect 13683 33612 13728 33640
rect 13722 33600 13728 33612
rect 13780 33640 13786 33652
rect 14090 33640 14096 33652
rect 13780 33600 13814 33640
rect 14051 33612 14096 33640
rect 14090 33600 14096 33612
rect 14148 33600 14154 33652
rect 15378 33600 15384 33652
rect 15436 33640 15442 33652
rect 16022 33640 16028 33652
rect 15436 33612 16028 33640
rect 15436 33600 15442 33612
rect 16022 33600 16028 33612
rect 16080 33600 16086 33652
rect 17494 33640 17500 33652
rect 17455 33612 17500 33640
rect 17494 33600 17500 33612
rect 17552 33600 17558 33652
rect 17865 33643 17923 33649
rect 17865 33609 17877 33643
rect 17911 33640 17923 33643
rect 17954 33640 17960 33652
rect 17911 33612 17960 33640
rect 17911 33609 17923 33612
rect 17865 33603 17923 33609
rect 17954 33600 17960 33612
rect 18012 33600 18018 33652
rect 19426 33640 19432 33652
rect 19387 33612 19432 33640
rect 19426 33600 19432 33612
rect 19484 33640 19490 33652
rect 20346 33640 20352 33652
rect 19484 33612 20352 33640
rect 19484 33600 19490 33612
rect 20346 33600 20352 33612
rect 20404 33640 20410 33652
rect 21818 33640 21824 33652
rect 20404 33612 21824 33640
rect 20404 33600 20410 33612
rect 21818 33600 21824 33612
rect 21876 33640 21882 33652
rect 21913 33643 21971 33649
rect 21913 33640 21925 33643
rect 21876 33612 21925 33640
rect 21876 33600 21882 33612
rect 21913 33609 21925 33612
rect 21959 33609 21971 33643
rect 21913 33603 21971 33609
rect 22002 33600 22008 33652
rect 22060 33640 22066 33652
rect 22603 33643 22661 33649
rect 22603 33640 22615 33643
rect 22060 33612 22615 33640
rect 22060 33600 22066 33612
rect 22603 33609 22615 33612
rect 22649 33609 22661 33643
rect 25593 33643 25651 33649
rect 25593 33640 25605 33643
rect 22603 33603 22661 33609
rect 23446 33612 25605 33640
rect 13786 33572 13814 33600
rect 23446 33572 23474 33612
rect 25593 33609 25605 33612
rect 25639 33640 25651 33643
rect 25682 33640 25688 33652
rect 25639 33612 25688 33640
rect 25639 33609 25651 33612
rect 25593 33603 25651 33609
rect 25682 33600 25688 33612
rect 25740 33600 25746 33652
rect 26973 33643 27031 33649
rect 26973 33609 26985 33643
rect 27019 33640 27031 33643
rect 27338 33640 27344 33652
rect 27019 33612 27344 33640
rect 27019 33609 27031 33612
rect 26973 33603 27031 33609
rect 27338 33600 27344 33612
rect 27396 33600 27402 33652
rect 27614 33640 27620 33652
rect 27575 33612 27620 33640
rect 27614 33600 27620 33612
rect 27672 33640 27678 33652
rect 27939 33643 27997 33649
rect 27939 33640 27951 33643
rect 27672 33612 27951 33640
rect 27672 33600 27678 33612
rect 27939 33609 27951 33612
rect 27985 33609 27997 33643
rect 27939 33603 27997 33609
rect 29638 33600 29644 33652
rect 29696 33640 29702 33652
rect 30285 33643 30343 33649
rect 30285 33640 30297 33643
rect 29696 33612 30297 33640
rect 29696 33600 29702 33612
rect 30285 33609 30297 33612
rect 30331 33640 30343 33643
rect 30374 33640 30380 33652
rect 30331 33612 30380 33640
rect 30331 33609 30343 33612
rect 30285 33603 30343 33609
rect 30374 33600 30380 33612
rect 30432 33640 30438 33652
rect 30837 33643 30895 33649
rect 30837 33640 30849 33643
rect 30432 33612 30849 33640
rect 30432 33600 30438 33612
rect 30837 33609 30849 33612
rect 30883 33640 30895 33643
rect 30929 33643 30987 33649
rect 30929 33640 30941 33643
rect 30883 33612 30941 33640
rect 30883 33609 30895 33612
rect 30837 33603 30895 33609
rect 30929 33609 30941 33612
rect 30975 33609 30987 33643
rect 30929 33603 30987 33609
rect 32033 33643 32091 33649
rect 32033 33609 32045 33643
rect 32079 33640 32091 33643
rect 32122 33640 32128 33652
rect 32079 33612 32128 33640
rect 32079 33609 32091 33612
rect 32033 33603 32091 33609
rect 32122 33600 32128 33612
rect 32180 33600 32186 33652
rect 32769 33643 32827 33649
rect 32769 33609 32781 33643
rect 32815 33640 32827 33643
rect 33042 33640 33048 33652
rect 32815 33612 33048 33640
rect 32815 33609 32827 33612
rect 32769 33603 32827 33609
rect 27798 33572 27804 33584
rect 13786 33544 18368 33572
rect 12526 33504 12532 33516
rect 12487 33476 12532 33504
rect 12526 33464 12532 33476
rect 12584 33464 12590 33516
rect 13906 33464 13912 33516
rect 13964 33504 13970 33516
rect 14734 33504 14740 33516
rect 13964 33476 14740 33504
rect 13964 33464 13970 33476
rect 14734 33464 14740 33476
rect 14792 33464 14798 33516
rect 18340 33448 18368 33544
rect 21192 33544 23474 33572
rect 24596 33544 27804 33572
rect 18874 33464 18880 33516
rect 18932 33504 18938 33516
rect 19061 33507 19119 33513
rect 19061 33504 19073 33507
rect 18932 33476 19073 33504
rect 18932 33464 18938 33476
rect 19061 33473 19073 33476
rect 19107 33504 19119 33507
rect 19705 33507 19763 33513
rect 19705 33504 19717 33507
rect 19107 33476 19717 33504
rect 19107 33473 19119 33476
rect 19061 33467 19119 33473
rect 19705 33473 19717 33476
rect 19751 33473 19763 33507
rect 19705 33467 19763 33473
rect 21192 33448 21220 33544
rect 21450 33464 21456 33516
rect 21508 33504 21514 33516
rect 24596 33513 24624 33544
rect 27798 33532 27804 33544
rect 27856 33532 27862 33584
rect 21637 33507 21695 33513
rect 21637 33504 21649 33507
rect 21508 33476 21649 33504
rect 21508 33464 21514 33476
rect 21637 33473 21649 33476
rect 21683 33504 21695 33507
rect 22281 33507 22339 33513
rect 22281 33504 22293 33507
rect 21683 33476 22293 33504
rect 21683 33473 21695 33476
rect 21637 33467 21695 33473
rect 22281 33473 22293 33476
rect 22327 33473 22339 33507
rect 22281 33467 22339 33473
rect 24029 33507 24087 33513
rect 24029 33473 24041 33507
rect 24075 33504 24087 33507
rect 24581 33507 24639 33513
rect 24581 33504 24593 33507
rect 24075 33476 24593 33504
rect 24075 33473 24087 33476
rect 24029 33467 24087 33473
rect 24581 33473 24593 33476
rect 24627 33473 24639 33507
rect 24581 33467 24639 33473
rect 24670 33464 24676 33516
rect 24728 33504 24734 33516
rect 24728 33476 25544 33504
rect 24728 33464 24734 33476
rect 10502 33396 10508 33448
rect 10560 33436 10566 33448
rect 10597 33439 10655 33445
rect 10597 33436 10609 33439
rect 10560 33408 10609 33436
rect 10560 33396 10566 33408
rect 10597 33405 10609 33408
rect 10643 33405 10655 33439
rect 10597 33399 10655 33405
rect 10962 33396 10968 33448
rect 11020 33436 11026 33448
rect 11057 33439 11115 33445
rect 11057 33436 11069 33439
rect 11020 33408 11069 33436
rect 11020 33396 11026 33408
rect 11057 33405 11069 33408
rect 11103 33405 11115 33439
rect 11057 33399 11115 33405
rect 17012 33439 17070 33445
rect 17012 33405 17024 33439
rect 17058 33436 17070 33439
rect 17954 33436 17960 33448
rect 17058 33408 17960 33436
rect 17058 33405 17070 33408
rect 17012 33399 17070 33405
rect 17954 33396 17960 33408
rect 18012 33396 18018 33448
rect 18322 33436 18328 33448
rect 18235 33408 18328 33436
rect 18322 33396 18328 33408
rect 18380 33396 18386 33448
rect 18414 33396 18420 33448
rect 18472 33436 18478 33448
rect 18785 33439 18843 33445
rect 18785 33436 18797 33439
rect 18472 33408 18797 33436
rect 18472 33396 18478 33408
rect 18785 33405 18797 33408
rect 18831 33436 18843 33439
rect 20809 33439 20867 33445
rect 18831 33408 19288 33436
rect 18831 33405 18843 33408
rect 18785 33399 18843 33405
rect 19260 33380 19288 33408
rect 20809 33405 20821 33439
rect 20855 33436 20867 33439
rect 21174 33436 21180 33448
rect 20855 33408 21180 33436
rect 20855 33405 20867 33408
rect 20809 33399 20867 33405
rect 21174 33396 21180 33408
rect 21232 33396 21238 33448
rect 21361 33439 21419 33445
rect 21361 33405 21373 33439
rect 21407 33436 21419 33439
rect 21726 33436 21732 33448
rect 21407 33408 21732 33436
rect 21407 33405 21419 33408
rect 21361 33399 21419 33405
rect 11333 33371 11391 33377
rect 11333 33337 11345 33371
rect 11379 33368 11391 33371
rect 11422 33368 11428 33380
rect 11379 33340 11428 33368
rect 11379 33337 11391 33340
rect 11333 33331 11391 33337
rect 11422 33328 11428 33340
rect 11480 33328 11486 33380
rect 12621 33371 12679 33377
rect 12621 33337 12633 33371
rect 12667 33368 12679 33371
rect 12710 33368 12716 33380
rect 12667 33340 12716 33368
rect 12667 33337 12679 33340
rect 12621 33331 12679 33337
rect 12710 33328 12716 33340
rect 12768 33328 12774 33380
rect 13170 33368 13176 33380
rect 13131 33340 13176 33368
rect 13170 33328 13176 33340
rect 13228 33328 13234 33380
rect 14829 33371 14887 33377
rect 14829 33337 14841 33371
rect 14875 33337 14887 33371
rect 15378 33368 15384 33380
rect 15339 33340 15384 33368
rect 14829 33331 14887 33337
rect 14550 33300 14556 33312
rect 14463 33272 14556 33300
rect 14550 33260 14556 33272
rect 14608 33300 14614 33312
rect 14844 33300 14872 33331
rect 15378 33328 15384 33340
rect 15436 33328 15442 33380
rect 19242 33328 19248 33380
rect 19300 33368 19306 33380
rect 20441 33371 20499 33377
rect 20441 33368 20453 33371
rect 19300 33340 20453 33368
rect 19300 33328 19306 33340
rect 20441 33337 20453 33340
rect 20487 33368 20499 33371
rect 21376 33368 21404 33399
rect 21726 33396 21732 33408
rect 21784 33396 21790 33448
rect 22532 33439 22590 33445
rect 22532 33405 22544 33439
rect 22578 33436 22590 33439
rect 22922 33436 22928 33448
rect 22578 33408 22928 33436
rect 22578 33405 22590 33408
rect 22532 33399 22590 33405
rect 22922 33396 22928 33408
rect 22980 33396 22986 33448
rect 25516 33436 25544 33476
rect 25590 33464 25596 33516
rect 25648 33504 25654 33516
rect 26050 33504 26056 33516
rect 25648 33476 26056 33504
rect 25648 33464 25654 33476
rect 26050 33464 26056 33476
rect 26108 33464 26114 33516
rect 25869 33439 25927 33445
rect 25869 33436 25881 33439
rect 25516 33408 25881 33436
rect 25869 33405 25881 33408
rect 25915 33436 25927 33439
rect 25915 33408 26417 33436
rect 25915 33405 25927 33408
rect 25869 33399 25927 33405
rect 20487 33340 21404 33368
rect 24673 33371 24731 33377
rect 20487 33337 20499 33340
rect 20441 33331 20499 33337
rect 24673 33337 24685 33371
rect 24719 33337 24731 33371
rect 25222 33368 25228 33380
rect 25183 33340 25228 33368
rect 24673 33331 24731 33337
rect 14608 33272 14872 33300
rect 14608 33260 14614 33272
rect 14918 33260 14924 33312
rect 14976 33300 14982 33312
rect 15470 33300 15476 33312
rect 14976 33272 15476 33300
rect 14976 33260 14982 33272
rect 15470 33260 15476 33272
rect 15528 33300 15534 33312
rect 15657 33303 15715 33309
rect 15657 33300 15669 33303
rect 15528 33272 15669 33300
rect 15528 33260 15534 33272
rect 15657 33269 15669 33272
rect 15703 33269 15715 33303
rect 15657 33263 15715 33269
rect 16942 33260 16948 33312
rect 17000 33300 17006 33312
rect 17083 33303 17141 33309
rect 17083 33300 17095 33303
rect 17000 33272 17095 33300
rect 17000 33260 17006 33272
rect 17083 33269 17095 33272
rect 17129 33269 17141 33303
rect 24394 33300 24400 33312
rect 24307 33272 24400 33300
rect 17083 33263 17141 33269
rect 24394 33260 24400 33272
rect 24452 33300 24458 33312
rect 24688 33300 24716 33331
rect 25222 33328 25228 33340
rect 25280 33328 25286 33380
rect 26389 33377 26417 33408
rect 27522 33396 27528 33448
rect 27580 33436 27586 33448
rect 27836 33439 27894 33445
rect 27836 33436 27848 33439
rect 27580 33408 27848 33436
rect 27580 33396 27586 33408
rect 27836 33405 27848 33408
rect 27882 33436 27894 33439
rect 28258 33436 28264 33448
rect 27882 33408 28264 33436
rect 27882 33405 27894 33408
rect 27836 33399 27894 33405
rect 28258 33396 28264 33408
rect 28316 33396 28322 33448
rect 28626 33396 28632 33448
rect 28684 33436 28690 33448
rect 29089 33439 29147 33445
rect 29089 33436 29101 33439
rect 28684 33408 29101 33436
rect 28684 33396 28690 33408
rect 29089 33405 29101 33408
rect 29135 33436 29147 33439
rect 29549 33439 29607 33445
rect 29549 33436 29561 33439
rect 29135 33408 29561 33436
rect 29135 33405 29147 33408
rect 29089 33399 29147 33405
rect 29549 33405 29561 33408
rect 29595 33405 29607 33439
rect 29549 33399 29607 33405
rect 29825 33439 29883 33445
rect 29825 33405 29837 33439
rect 29871 33436 29883 33439
rect 30558 33436 30564 33448
rect 29871 33408 30564 33436
rect 29871 33405 29883 33408
rect 29825 33399 29883 33405
rect 30558 33396 30564 33408
rect 30616 33396 30622 33448
rect 31110 33436 31116 33448
rect 31071 33408 31116 33436
rect 31110 33396 31116 33408
rect 31168 33396 31174 33448
rect 32784 33436 32812 33603
rect 33042 33600 33048 33612
rect 33100 33600 33106 33652
rect 33870 33640 33876 33652
rect 33831 33612 33876 33640
rect 33870 33600 33876 33612
rect 33928 33600 33934 33652
rect 35526 33600 35532 33652
rect 35584 33640 35590 33652
rect 36265 33643 36323 33649
rect 36265 33640 36277 33643
rect 35584 33612 36277 33640
rect 35584 33600 35590 33612
rect 36265 33609 36277 33612
rect 36311 33609 36323 33643
rect 36265 33603 36323 33609
rect 38194 33600 38200 33652
rect 38252 33640 38258 33652
rect 38841 33643 38899 33649
rect 38841 33640 38853 33643
rect 38252 33612 38853 33640
rect 38252 33600 38258 33612
rect 38841 33609 38853 33612
rect 38887 33609 38899 33643
rect 38841 33603 38899 33609
rect 39022 33600 39028 33652
rect 39080 33640 39086 33652
rect 39209 33643 39267 33649
rect 39209 33640 39221 33643
rect 39080 33612 39221 33640
rect 39080 33600 39086 33612
rect 39209 33609 39221 33612
rect 39255 33609 39267 33643
rect 39209 33603 39267 33609
rect 40034 33600 40040 33652
rect 40092 33640 40098 33652
rect 40310 33640 40316 33652
rect 40092 33612 40316 33640
rect 40092 33600 40098 33612
rect 40310 33600 40316 33612
rect 40368 33600 40374 33652
rect 40589 33643 40647 33649
rect 40589 33609 40601 33643
rect 40635 33640 40647 33643
rect 41506 33640 41512 33652
rect 40635 33612 41512 33640
rect 40635 33609 40647 33612
rect 40589 33603 40647 33609
rect 41506 33600 41512 33612
rect 41564 33600 41570 33652
rect 41690 33640 41696 33652
rect 41651 33612 41696 33640
rect 41690 33600 41696 33612
rect 41748 33600 41754 33652
rect 42150 33640 42156 33652
rect 42111 33612 42156 33640
rect 42150 33600 42156 33612
rect 42208 33600 42214 33652
rect 37458 33532 37464 33584
rect 37516 33572 37522 33584
rect 39531 33575 39589 33581
rect 39531 33572 39543 33575
rect 37516 33544 39543 33572
rect 37516 33532 37522 33544
rect 39531 33541 39543 33544
rect 39577 33541 39589 33575
rect 41325 33575 41383 33581
rect 41325 33572 41337 33575
rect 39531 33535 39589 33541
rect 39960 33544 41337 33572
rect 33318 33504 33324 33516
rect 33279 33476 33324 33504
rect 33318 33464 33324 33476
rect 33376 33464 33382 33516
rect 36078 33464 36084 33516
rect 36136 33504 36142 33516
rect 36955 33507 37013 33513
rect 36136 33476 36895 33504
rect 36136 33464 36142 33476
rect 32692 33408 32812 33436
rect 35856 33439 35914 33445
rect 26374 33371 26432 33377
rect 26374 33337 26386 33371
rect 26420 33337 26432 33371
rect 26374 33331 26432 33337
rect 28721 33371 28779 33377
rect 28721 33337 28733 33371
rect 28767 33368 28779 33371
rect 30837 33371 30895 33377
rect 28767 33340 29500 33368
rect 28767 33337 28779 33340
rect 28721 33331 28779 33337
rect 29472 33312 29500 33340
rect 30837 33337 30849 33371
rect 30883 33368 30895 33371
rect 31434 33371 31492 33377
rect 31434 33368 31446 33371
rect 30883 33340 31446 33368
rect 30883 33337 30895 33340
rect 30837 33331 30895 33337
rect 31434 33337 31446 33340
rect 31480 33368 31492 33371
rect 32306 33368 32312 33380
rect 31480 33340 32312 33368
rect 31480 33337 31492 33340
rect 31434 33331 31492 33337
rect 32306 33328 32312 33340
rect 32364 33328 32370 33380
rect 24452 33272 24716 33300
rect 24452 33260 24458 33272
rect 29454 33260 29460 33312
rect 29512 33300 29518 33312
rect 29549 33303 29607 33309
rect 29549 33300 29561 33303
rect 29512 33272 29561 33300
rect 29512 33260 29518 33272
rect 29549 33269 29561 33272
rect 29595 33269 29607 33303
rect 32692 33300 32720 33408
rect 35856 33405 35868 33439
rect 35902 33436 35914 33439
rect 36446 33436 36452 33448
rect 35902 33408 36452 33436
rect 35902 33405 35914 33408
rect 35856 33399 35914 33405
rect 36446 33396 36452 33408
rect 36504 33436 36510 33448
rect 36867 33445 36895 33476
rect 36955 33473 36967 33507
rect 37001 33504 37013 33507
rect 37918 33504 37924 33516
rect 37001 33476 37924 33504
rect 37001 33473 37013 33476
rect 36955 33467 37013 33473
rect 37918 33464 37924 33476
rect 37976 33464 37982 33516
rect 38286 33464 38292 33516
rect 38344 33504 38350 33516
rect 38565 33507 38623 33513
rect 38565 33504 38577 33507
rect 38344 33476 38577 33504
rect 38344 33464 38350 33476
rect 38565 33473 38577 33476
rect 38611 33504 38623 33507
rect 39960 33504 39988 33544
rect 41325 33541 41337 33544
rect 41371 33572 41383 33575
rect 44174 33572 44180 33584
rect 41371 33544 44180 33572
rect 41371 33541 41383 33544
rect 41325 33535 41383 33541
rect 44174 33532 44180 33544
rect 44232 33532 44238 33584
rect 40770 33504 40776 33516
rect 38611 33476 39988 33504
rect 40731 33476 40776 33504
rect 38611 33473 38623 33476
rect 38565 33467 38623 33473
rect 40770 33464 40776 33476
rect 40828 33464 40834 33516
rect 43622 33504 43628 33516
rect 43583 33476 43628 33504
rect 43622 33464 43628 33476
rect 43680 33464 43686 33516
rect 36633 33439 36691 33445
rect 36633 33436 36645 33439
rect 36504 33408 36645 33436
rect 36504 33396 36510 33408
rect 36633 33405 36645 33408
rect 36679 33405 36691 33439
rect 36633 33399 36691 33405
rect 36852 33439 36910 33445
rect 36852 33405 36864 33439
rect 36898 33436 36910 33439
rect 37277 33439 37335 33445
rect 37277 33436 37289 33439
rect 36898 33408 37289 33436
rect 36898 33405 36910 33408
rect 36852 33399 36910 33405
rect 37277 33405 37289 33408
rect 37323 33436 37335 33439
rect 37642 33436 37648 33448
rect 37323 33408 37648 33436
rect 37323 33405 37335 33408
rect 37277 33399 37335 33405
rect 37642 33396 37648 33408
rect 37700 33396 37706 33448
rect 39206 33396 39212 33448
rect 39264 33436 39270 33448
rect 39428 33439 39486 33445
rect 39428 33436 39440 33439
rect 39264 33408 39440 33436
rect 39264 33396 39270 33408
rect 39428 33405 39440 33408
rect 39474 33436 39486 33439
rect 39853 33439 39911 33445
rect 39853 33436 39865 33439
rect 39474 33408 39865 33436
rect 39474 33405 39486 33408
rect 39428 33399 39486 33405
rect 39853 33405 39865 33408
rect 39899 33436 39911 33439
rect 40589 33439 40647 33445
rect 40589 33436 40601 33439
rect 39899 33408 40601 33436
rect 39899 33405 39911 33408
rect 39853 33399 39911 33405
rect 40589 33405 40601 33408
rect 40635 33405 40647 33439
rect 40589 33399 40647 33405
rect 41966 33396 41972 33448
rect 42024 33436 42030 33448
rect 42280 33439 42338 33445
rect 42280 33436 42292 33439
rect 42024 33408 42292 33436
rect 42024 33396 42030 33408
rect 42280 33405 42292 33408
rect 42326 33436 42338 33439
rect 42705 33439 42763 33445
rect 42705 33436 42717 33439
rect 42326 33408 42717 33436
rect 42326 33405 42338 33408
rect 42280 33399 42338 33405
rect 42705 33405 42717 33408
rect 42751 33405 42763 33439
rect 42705 33399 42763 33405
rect 32766 33328 32772 33380
rect 32824 33368 32830 33380
rect 32942 33371 33000 33377
rect 32942 33368 32954 33371
rect 32824 33340 32954 33368
rect 32824 33328 32830 33340
rect 32942 33337 32954 33340
rect 32988 33337 33000 33371
rect 32942 33331 33000 33337
rect 33054 33371 33112 33377
rect 33054 33337 33066 33371
rect 33100 33368 33112 33371
rect 33100 33337 33134 33368
rect 33054 33331 33134 33337
rect 33106 33300 33134 33331
rect 34606 33328 34612 33380
rect 34664 33368 34670 33380
rect 35943 33371 36001 33377
rect 35943 33368 35955 33371
rect 34664 33340 35955 33368
rect 34664 33328 34670 33340
rect 35943 33337 35955 33340
rect 35989 33337 36001 33371
rect 35943 33331 36001 33337
rect 38013 33371 38071 33377
rect 38013 33337 38025 33371
rect 38059 33337 38071 33371
rect 38013 33331 38071 33337
rect 32692 33272 33134 33300
rect 35621 33303 35679 33309
rect 29549 33263 29607 33269
rect 35621 33269 35633 33303
rect 35667 33300 35679 33303
rect 36538 33300 36544 33312
rect 35667 33272 36544 33300
rect 35667 33269 35679 33272
rect 35621 33263 35679 33269
rect 36538 33260 36544 33272
rect 36596 33260 36602 33312
rect 37737 33303 37795 33309
rect 37737 33269 37749 33303
rect 37783 33300 37795 33303
rect 38028 33300 38056 33331
rect 40862 33328 40868 33380
rect 40920 33368 40926 33380
rect 42383 33371 42441 33377
rect 42383 33368 42395 33371
rect 40920 33340 40965 33368
rect 41575 33340 42395 33368
rect 40920 33328 40926 33340
rect 38102 33300 38108 33312
rect 37783 33272 38108 33300
rect 37783 33269 37795 33272
rect 37737 33263 37795 33269
rect 38102 33260 38108 33272
rect 38160 33260 38166 33312
rect 40494 33260 40500 33312
rect 40552 33300 40558 33312
rect 41575 33300 41603 33340
rect 42383 33337 42395 33340
rect 42429 33337 42441 33371
rect 42383 33331 42441 33337
rect 43441 33371 43499 33377
rect 43441 33337 43453 33371
rect 43487 33368 43499 33371
rect 43717 33371 43775 33377
rect 43717 33368 43729 33371
rect 43487 33340 43729 33368
rect 43487 33337 43499 33340
rect 43441 33331 43499 33337
rect 43717 33337 43729 33340
rect 43763 33368 43775 33371
rect 44082 33368 44088 33380
rect 43763 33340 44088 33368
rect 43763 33337 43775 33340
rect 43717 33331 43775 33337
rect 44082 33328 44088 33340
rect 44140 33328 44146 33380
rect 44266 33368 44272 33380
rect 44227 33340 44272 33368
rect 44266 33328 44272 33340
rect 44324 33328 44330 33380
rect 40552 33272 41603 33300
rect 40552 33260 40558 33272
rect 1104 33210 48852 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 48852 33210
rect 1104 33136 48852 33158
rect 14734 33096 14740 33108
rect 14695 33068 14740 33096
rect 14734 33056 14740 33068
rect 14792 33056 14798 33108
rect 15427 33099 15485 33105
rect 15427 33065 15439 33099
rect 15473 33096 15485 33099
rect 16022 33096 16028 33108
rect 15473 33068 16028 33096
rect 15473 33065 15485 33068
rect 15427 33059 15485 33065
rect 16022 33056 16028 33068
rect 16080 33056 16086 33108
rect 18046 33096 18052 33108
rect 18007 33068 18052 33096
rect 18046 33056 18052 33068
rect 18104 33056 18110 33108
rect 24394 33096 24400 33108
rect 24355 33068 24400 33096
rect 24394 33056 24400 33068
rect 24452 33056 24458 33108
rect 24946 33096 24952 33108
rect 24907 33068 24952 33096
rect 24946 33056 24952 33068
rect 25004 33056 25010 33108
rect 26050 33096 26056 33108
rect 26011 33068 26056 33096
rect 26050 33056 26056 33068
rect 26108 33056 26114 33108
rect 32214 33096 32220 33108
rect 32175 33068 32220 33096
rect 32214 33056 32220 33068
rect 32272 33056 32278 33108
rect 33226 33096 33232 33108
rect 33187 33068 33232 33096
rect 33226 33056 33232 33068
rect 33284 33056 33290 33108
rect 34790 33056 34796 33108
rect 34848 33096 34854 33108
rect 34885 33099 34943 33105
rect 34885 33096 34897 33099
rect 34848 33068 34897 33096
rect 34848 33056 34854 33068
rect 34885 33065 34897 33068
rect 34931 33065 34943 33099
rect 34885 33059 34943 33065
rect 36538 33056 36544 33108
rect 36596 33096 36602 33108
rect 37826 33096 37832 33108
rect 36596 33068 37832 33096
rect 36596 33056 36602 33068
rect 37826 33056 37832 33068
rect 37884 33096 37890 33108
rect 37884 33068 38101 33096
rect 37884 33056 37890 33068
rect 11511 33031 11569 33037
rect 11511 32997 11523 33031
rect 11557 33028 11569 33031
rect 11974 33028 11980 33040
rect 11557 33000 11980 33028
rect 11557 32997 11569 33000
rect 11511 32991 11569 32997
rect 11974 32988 11980 33000
rect 12032 32988 12038 33040
rect 12894 32988 12900 33040
rect 12952 33028 12958 33040
rect 13446 33028 13452 33040
rect 12952 33000 13452 33028
rect 12952 32988 12958 33000
rect 13446 32988 13452 33000
rect 13504 32988 13510 33040
rect 13538 32988 13544 33040
rect 13596 33028 13602 33040
rect 14550 33028 14556 33040
rect 13596 33000 14556 33028
rect 13596 32988 13602 33000
rect 14550 32988 14556 33000
rect 14608 32988 14614 33040
rect 17123 33031 17181 33037
rect 17123 32997 17135 33031
rect 17169 33028 17181 33031
rect 17494 33028 17500 33040
rect 17169 33000 17500 33028
rect 17169 32997 17181 33000
rect 17123 32991 17181 32997
rect 17494 32988 17500 33000
rect 17552 32988 17558 33040
rect 18877 33031 18935 33037
rect 18877 32997 18889 33031
rect 18923 33028 18935 33031
rect 19242 33028 19248 33040
rect 18923 33000 19248 33028
rect 18923 32997 18935 33000
rect 18877 32991 18935 32997
rect 19242 32988 19248 33000
rect 19300 33028 19306 33040
rect 19705 33031 19763 33037
rect 19300 33000 19472 33028
rect 19300 32988 19306 33000
rect 15356 32963 15414 32969
rect 15356 32929 15368 32963
rect 15402 32960 15414 32963
rect 15746 32960 15752 32972
rect 15402 32932 15752 32960
rect 15402 32929 15414 32932
rect 15356 32923 15414 32929
rect 15746 32920 15752 32932
rect 15804 32920 15810 32972
rect 19058 32960 19064 32972
rect 19019 32932 19064 32960
rect 19058 32920 19064 32932
rect 19116 32920 19122 32972
rect 19444 32969 19472 33000
rect 19705 32997 19717 33031
rect 19751 33028 19763 33031
rect 20070 33028 20076 33040
rect 19751 33000 20076 33028
rect 19751 32997 19763 33000
rect 19705 32991 19763 32997
rect 20070 32988 20076 33000
rect 20128 32988 20134 33040
rect 20346 32988 20352 33040
rect 20404 33028 20410 33040
rect 23106 33028 23112 33040
rect 20404 33000 23112 33028
rect 20404 32988 20410 33000
rect 23106 32988 23112 33000
rect 23164 33028 23170 33040
rect 23839 33031 23897 33037
rect 23839 33028 23851 33031
rect 23164 33000 23851 33028
rect 23164 32988 23170 33000
rect 23839 32997 23851 33000
rect 23885 33028 23897 33031
rect 24762 33028 24768 33040
rect 23885 33000 24768 33028
rect 23885 32997 23897 33000
rect 23839 32991 23897 32997
rect 24762 32988 24768 33000
rect 24820 32988 24826 33040
rect 26418 32988 26424 33040
rect 26476 33028 26482 33040
rect 26697 33031 26755 33037
rect 26697 33028 26709 33031
rect 26476 33000 26709 33028
rect 26476 32988 26482 33000
rect 26697 32997 26709 33000
rect 26743 32997 26755 33031
rect 28810 33028 28816 33040
rect 28771 33000 28816 33028
rect 26697 32991 26755 32997
rect 28810 32988 28816 33000
rect 28868 32988 28874 33040
rect 29822 32988 29828 33040
rect 29880 33028 29886 33040
rect 34057 33031 34115 33037
rect 34057 33028 34069 33031
rect 29880 33000 34069 33028
rect 29880 32988 29886 33000
rect 34057 32997 34069 33000
rect 34103 33028 34115 33031
rect 34330 33028 34336 33040
rect 34103 33000 34336 33028
rect 34103 32997 34115 33000
rect 34057 32991 34115 32997
rect 34330 32988 34336 33000
rect 34388 32988 34394 33040
rect 38073 33037 38101 33068
rect 39390 33056 39396 33108
rect 39448 33096 39454 33108
rect 42058 33096 42064 33108
rect 39448 33068 42064 33096
rect 39448 33056 39454 33068
rect 42058 33056 42064 33068
rect 42116 33056 42122 33108
rect 43622 33056 43628 33108
rect 43680 33096 43686 33108
rect 43717 33099 43775 33105
rect 43717 33096 43729 33099
rect 43680 33068 43729 33096
rect 43680 33056 43686 33068
rect 43717 33065 43729 33068
rect 43763 33065 43775 33099
rect 43717 33059 43775 33065
rect 44082 33056 44088 33108
rect 44140 33096 44146 33108
rect 44269 33099 44327 33105
rect 44269 33096 44281 33099
rect 44140 33068 44281 33096
rect 44140 33056 44146 33068
rect 44269 33065 44281 33068
rect 44315 33065 44327 33099
rect 44269 33059 44327 33065
rect 38058 33031 38116 33037
rect 38058 32997 38070 33031
rect 38104 32997 38116 33031
rect 38058 32991 38116 32997
rect 38562 32988 38568 33040
rect 38620 33028 38626 33040
rect 38930 33028 38936 33040
rect 38620 33000 38936 33028
rect 38620 32988 38626 33000
rect 38930 32988 38936 33000
rect 38988 32988 38994 33040
rect 39850 32988 39856 33040
rect 39908 33028 39914 33040
rect 40126 33037 40132 33040
rect 40082 33031 40132 33037
rect 40082 33028 40094 33031
rect 39908 33000 40094 33028
rect 39908 32988 39914 33000
rect 40082 32997 40094 33000
rect 40128 32997 40132 33031
rect 40082 32991 40132 32997
rect 40126 32988 40132 32991
rect 40184 32988 40190 33040
rect 40862 32988 40868 33040
rect 40920 33028 40926 33040
rect 41693 33031 41751 33037
rect 41693 33028 41705 33031
rect 40920 33000 41705 33028
rect 40920 32988 40926 33000
rect 41693 32997 41705 33000
rect 41739 32997 41751 33031
rect 41693 32991 41751 32997
rect 19429 32963 19487 32969
rect 19429 32929 19441 32963
rect 19475 32929 19487 32963
rect 19429 32923 19487 32929
rect 22189 32963 22247 32969
rect 22189 32929 22201 32963
rect 22235 32960 22247 32963
rect 22278 32960 22284 32972
rect 22235 32932 22284 32960
rect 22235 32929 22247 32932
rect 22189 32923 22247 32929
rect 22278 32920 22284 32932
rect 22336 32920 22342 32972
rect 22462 32960 22468 32972
rect 22423 32932 22468 32960
rect 22462 32920 22468 32932
rect 22520 32920 22526 32972
rect 25133 32963 25191 32969
rect 25133 32929 25145 32963
rect 25179 32960 25191 32963
rect 25222 32960 25228 32972
rect 25179 32932 25228 32960
rect 25179 32929 25191 32932
rect 25133 32923 25191 32929
rect 25222 32920 25228 32932
rect 25280 32920 25286 32972
rect 28074 32960 28080 32972
rect 28035 32932 28080 32960
rect 28074 32920 28080 32932
rect 28132 32920 28138 32972
rect 28258 32920 28264 32972
rect 28316 32960 28322 32972
rect 30466 32960 30472 32972
rect 28316 32932 28994 32960
rect 30427 32932 30472 32960
rect 28316 32920 28322 32932
rect 10134 32892 10140 32904
rect 10095 32864 10140 32892
rect 10134 32852 10140 32864
rect 10192 32852 10198 32904
rect 11149 32895 11207 32901
rect 11149 32861 11161 32895
rect 11195 32892 11207 32895
rect 11422 32892 11428 32904
rect 11195 32864 11428 32892
rect 11195 32861 11207 32864
rect 11149 32855 11207 32861
rect 11422 32852 11428 32864
rect 11480 32852 11486 32904
rect 13722 32892 13728 32904
rect 13683 32864 13728 32892
rect 13722 32852 13728 32864
rect 13780 32852 13786 32904
rect 16761 32895 16819 32901
rect 16761 32861 16773 32895
rect 16807 32892 16819 32895
rect 17034 32892 17040 32904
rect 16807 32864 17040 32892
rect 16807 32861 16819 32864
rect 16761 32855 16819 32861
rect 17034 32852 17040 32864
rect 17092 32852 17098 32904
rect 22649 32895 22707 32901
rect 22649 32861 22661 32895
rect 22695 32892 22707 32895
rect 23290 32892 23296 32904
rect 22695 32864 23296 32892
rect 22695 32861 22707 32864
rect 22649 32855 22707 32861
rect 23290 32852 23296 32864
rect 23348 32892 23354 32904
rect 23477 32895 23535 32901
rect 23477 32892 23489 32895
rect 23348 32864 23489 32892
rect 23348 32852 23354 32864
rect 23477 32861 23489 32864
rect 23523 32861 23535 32895
rect 23477 32855 23535 32861
rect 26605 32895 26663 32901
rect 26605 32861 26617 32895
rect 26651 32861 26663 32895
rect 26878 32892 26884 32904
rect 26839 32864 26884 32892
rect 26605 32855 26663 32861
rect 26326 32784 26332 32836
rect 26384 32824 26390 32836
rect 26620 32824 26648 32855
rect 26878 32852 26884 32864
rect 26936 32852 26942 32904
rect 28445 32895 28503 32901
rect 28445 32861 28457 32895
rect 28491 32892 28503 32895
rect 28626 32892 28632 32904
rect 28491 32864 28632 32892
rect 28491 32861 28503 32864
rect 28445 32855 28503 32861
rect 28626 32852 28632 32864
rect 28684 32852 28690 32904
rect 27430 32824 27436 32836
rect 26384 32796 27436 32824
rect 26384 32784 26390 32796
rect 27430 32784 27436 32796
rect 27488 32784 27494 32836
rect 28353 32827 28411 32833
rect 28353 32824 28365 32827
rect 28000 32796 28365 32824
rect 28000 32768 28028 32796
rect 28353 32793 28365 32796
rect 28399 32793 28411 32827
rect 28966 32824 28994 32932
rect 30466 32920 30472 32932
rect 30524 32920 30530 32972
rect 30742 32960 30748 32972
rect 30703 32932 30748 32960
rect 30742 32920 30748 32932
rect 30800 32920 30806 32972
rect 30929 32963 30987 32969
rect 30929 32929 30941 32963
rect 30975 32960 30987 32963
rect 31110 32960 31116 32972
rect 30975 32932 31116 32960
rect 30975 32929 30987 32932
rect 30929 32923 30987 32929
rect 31110 32920 31116 32932
rect 31168 32960 31174 32972
rect 31205 32963 31263 32969
rect 31205 32960 31217 32963
rect 31168 32932 31217 32960
rect 31168 32920 31174 32932
rect 31205 32929 31217 32932
rect 31251 32929 31263 32963
rect 31205 32923 31263 32929
rect 32122 32920 32128 32972
rect 32180 32960 32186 32972
rect 32401 32963 32459 32969
rect 32401 32960 32413 32963
rect 32180 32932 32413 32960
rect 32180 32920 32186 32932
rect 32401 32929 32413 32932
rect 32447 32960 32459 32963
rect 32490 32960 32496 32972
rect 32447 32932 32496 32960
rect 32447 32929 32459 32932
rect 32401 32923 32459 32929
rect 32490 32920 32496 32932
rect 32548 32920 32554 32972
rect 32674 32960 32680 32972
rect 32635 32932 32680 32960
rect 32674 32920 32680 32932
rect 32732 32920 32738 32972
rect 36262 32960 36268 32972
rect 36223 32932 36268 32960
rect 36262 32920 36268 32932
rect 36320 32920 36326 32972
rect 36538 32960 36544 32972
rect 36499 32932 36544 32960
rect 36538 32920 36544 32932
rect 36596 32960 36602 32972
rect 39025 32963 39083 32969
rect 39025 32960 39037 32963
rect 36596 32932 39037 32960
rect 36596 32920 36602 32932
rect 39025 32929 39037 32932
rect 39071 32960 39083 32963
rect 39390 32960 39396 32972
rect 39071 32932 39396 32960
rect 39071 32929 39083 32932
rect 39025 32923 39083 32929
rect 39390 32920 39396 32932
rect 39448 32920 39454 32972
rect 42610 32920 42616 32972
rect 42668 32960 42674 32972
rect 43349 32963 43407 32969
rect 43349 32960 43361 32963
rect 42668 32932 43361 32960
rect 42668 32920 42674 32932
rect 43349 32929 43361 32932
rect 43395 32929 43407 32963
rect 43349 32923 43407 32929
rect 32306 32852 32312 32904
rect 32364 32892 32370 32904
rect 35986 32892 35992 32904
rect 32364 32864 35992 32892
rect 32364 32852 32370 32864
rect 35986 32852 35992 32864
rect 36044 32892 36050 32904
rect 36722 32892 36728 32904
rect 36044 32864 36728 32892
rect 36044 32852 36050 32864
rect 36722 32852 36728 32864
rect 36780 32852 36786 32904
rect 36817 32895 36875 32901
rect 36817 32861 36829 32895
rect 36863 32892 36875 32895
rect 37182 32892 37188 32904
rect 36863 32864 37188 32892
rect 36863 32861 36875 32864
rect 36817 32855 36875 32861
rect 37182 32852 37188 32864
rect 37240 32892 37246 32904
rect 37737 32895 37795 32901
rect 37737 32892 37749 32895
rect 37240 32864 37749 32892
rect 37240 32852 37246 32864
rect 37737 32861 37749 32864
rect 37783 32861 37795 32895
rect 39758 32892 39764 32904
rect 39719 32864 39764 32892
rect 37737 32855 37795 32861
rect 39758 32852 39764 32864
rect 39816 32852 39822 32904
rect 41598 32892 41604 32904
rect 41559 32864 41604 32892
rect 41598 32852 41604 32864
rect 41656 32852 41662 32904
rect 42245 32895 42303 32901
rect 42245 32861 42257 32895
rect 42291 32892 42303 32895
rect 42978 32892 42984 32904
rect 42291 32864 42984 32892
rect 42291 32861 42303 32864
rect 42245 32855 42303 32861
rect 42978 32852 42984 32864
rect 43036 32852 43042 32904
rect 45094 32892 45100 32904
rect 45055 32864 45100 32892
rect 45094 32852 45100 32864
rect 45152 32852 45158 32904
rect 32398 32824 32404 32836
rect 28966 32796 32404 32824
rect 28353 32787 28411 32793
rect 32398 32784 32404 32796
rect 32456 32784 32462 32836
rect 38102 32784 38108 32836
rect 38160 32824 38166 32836
rect 38562 32824 38568 32836
rect 38160 32796 38568 32824
rect 38160 32784 38166 32796
rect 38562 32784 38568 32796
rect 38620 32824 38626 32836
rect 38657 32827 38715 32833
rect 38657 32824 38669 32827
rect 38620 32796 38669 32824
rect 38620 32784 38626 32796
rect 38657 32793 38669 32796
rect 38703 32793 38715 32827
rect 42150 32824 42156 32836
rect 38657 32787 38715 32793
rect 39821 32796 42156 32824
rect 10686 32756 10692 32768
rect 10647 32728 10692 32756
rect 10686 32716 10692 32728
rect 10744 32756 10750 32768
rect 10962 32756 10968 32768
rect 10744 32728 10968 32756
rect 10744 32716 10750 32728
rect 10962 32716 10968 32728
rect 11020 32716 11026 32768
rect 12069 32759 12127 32765
rect 12069 32725 12081 32759
rect 12115 32756 12127 32759
rect 12526 32756 12532 32768
rect 12115 32728 12532 32756
rect 12115 32725 12127 32728
rect 12069 32719 12127 32725
rect 12526 32716 12532 32728
rect 12584 32716 12590 32768
rect 17678 32756 17684 32768
rect 17639 32728 17684 32756
rect 17678 32716 17684 32728
rect 17736 32716 17742 32768
rect 18322 32756 18328 32768
rect 18283 32728 18328 32756
rect 18322 32716 18328 32728
rect 18380 32716 18386 32768
rect 21361 32759 21419 32765
rect 21361 32725 21373 32759
rect 21407 32756 21419 32759
rect 21542 32756 21548 32768
rect 21407 32728 21548 32756
rect 21407 32725 21419 32728
rect 21361 32719 21419 32725
rect 21542 32716 21548 32728
rect 21600 32716 21606 32768
rect 23566 32716 23572 32768
rect 23624 32756 23630 32768
rect 25363 32759 25421 32765
rect 25363 32756 25375 32759
rect 23624 32728 25375 32756
rect 23624 32716 23630 32728
rect 25363 32725 25375 32728
rect 25409 32725 25421 32759
rect 25682 32756 25688 32768
rect 25643 32728 25688 32756
rect 25363 32719 25421 32725
rect 25682 32716 25688 32728
rect 25740 32716 25746 32768
rect 27709 32759 27767 32765
rect 27709 32725 27721 32759
rect 27755 32756 27767 32759
rect 27982 32756 27988 32768
rect 27755 32728 27988 32756
rect 27755 32725 27767 32728
rect 27709 32719 27767 32725
rect 27982 32716 27988 32728
rect 28040 32716 28046 32768
rect 28258 32765 28264 32768
rect 28242 32759 28264 32765
rect 28242 32725 28254 32759
rect 28242 32719 28264 32725
rect 28258 32716 28264 32719
rect 28316 32716 28322 32768
rect 28442 32716 28448 32768
rect 28500 32756 28506 32768
rect 29273 32759 29331 32765
rect 29273 32756 29285 32759
rect 28500 32728 29285 32756
rect 28500 32716 28506 32728
rect 29273 32725 29285 32728
rect 29319 32725 29331 32759
rect 29273 32719 29331 32725
rect 29917 32759 29975 32765
rect 29917 32725 29929 32759
rect 29963 32756 29975 32759
rect 30006 32756 30012 32768
rect 29963 32728 30012 32756
rect 29963 32725 29975 32728
rect 29917 32719 29975 32725
rect 30006 32716 30012 32728
rect 30064 32716 30070 32768
rect 31570 32756 31576 32768
rect 31531 32728 31576 32756
rect 31570 32716 31576 32728
rect 31628 32716 31634 32768
rect 34287 32759 34345 32765
rect 34287 32725 34299 32759
rect 34333 32756 34345 32759
rect 36078 32756 36084 32768
rect 34333 32728 36084 32756
rect 34333 32725 34345 32728
rect 34287 32719 34345 32725
rect 36078 32716 36084 32728
rect 36136 32716 36142 32768
rect 37550 32716 37556 32768
rect 37608 32756 37614 32768
rect 39821 32756 39849 32796
rect 42150 32784 42156 32796
rect 42208 32784 42214 32836
rect 37608 32728 39849 32756
rect 40681 32759 40739 32765
rect 37608 32716 37614 32728
rect 40681 32725 40693 32759
rect 40727 32756 40739 32759
rect 40862 32756 40868 32768
rect 40727 32728 40868 32756
rect 40727 32725 40739 32728
rect 40681 32719 40739 32725
rect 40862 32716 40868 32728
rect 40920 32756 40926 32768
rect 40957 32759 41015 32765
rect 40957 32756 40969 32759
rect 40920 32728 40969 32756
rect 40920 32716 40926 32728
rect 40957 32725 40969 32728
rect 41003 32725 41015 32759
rect 40957 32719 41015 32725
rect 41046 32716 41052 32768
rect 41104 32756 41110 32768
rect 41325 32759 41383 32765
rect 41325 32756 41337 32759
rect 41104 32728 41337 32756
rect 41104 32716 41110 32728
rect 41325 32725 41337 32728
rect 41371 32725 41383 32759
rect 41325 32719 41383 32725
rect 1104 32666 48852 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 48852 32666
rect 1104 32592 48852 32614
rect 10134 32512 10140 32564
rect 10192 32552 10198 32564
rect 12161 32555 12219 32561
rect 12161 32552 12173 32555
rect 10192 32524 12173 32552
rect 10192 32512 10198 32524
rect 12161 32521 12173 32524
rect 12207 32552 12219 32555
rect 12207 32524 12572 32552
rect 12207 32521 12219 32524
rect 12161 32515 12219 32521
rect 10505 32487 10563 32493
rect 10505 32453 10517 32487
rect 10551 32484 10563 32487
rect 11885 32487 11943 32493
rect 11885 32484 11897 32487
rect 10551 32456 11897 32484
rect 10551 32453 10563 32456
rect 10505 32447 10563 32453
rect 10137 32351 10195 32357
rect 10137 32317 10149 32351
rect 10183 32348 10195 32351
rect 10502 32348 10508 32360
rect 10183 32320 10508 32348
rect 10183 32317 10195 32320
rect 10137 32311 10195 32317
rect 10502 32308 10508 32320
rect 10560 32348 10566 32360
rect 10597 32351 10655 32357
rect 10597 32348 10609 32351
rect 10560 32320 10609 32348
rect 10560 32308 10566 32320
rect 10597 32317 10609 32320
rect 10643 32317 10655 32351
rect 10597 32311 10655 32317
rect 10974 32289 11002 32456
rect 11885 32453 11897 32456
rect 11931 32484 11943 32487
rect 11974 32484 11980 32496
rect 11931 32456 11980 32484
rect 11931 32453 11943 32456
rect 11885 32447 11943 32453
rect 11974 32444 11980 32456
rect 12032 32444 12038 32496
rect 12544 32425 12572 32524
rect 13446 32512 13452 32564
rect 13504 32552 13510 32564
rect 13817 32555 13875 32561
rect 13817 32552 13829 32555
rect 13504 32524 13829 32552
rect 13504 32512 13510 32524
rect 13817 32521 13829 32524
rect 13863 32521 13875 32555
rect 17494 32552 17500 32564
rect 17407 32524 17500 32552
rect 13817 32515 13875 32521
rect 17494 32512 17500 32524
rect 17552 32552 17558 32564
rect 20346 32552 20352 32564
rect 17552 32524 20352 32552
rect 17552 32512 17558 32524
rect 20346 32512 20352 32524
rect 20404 32512 20410 32564
rect 21726 32552 21732 32564
rect 21687 32524 21732 32552
rect 21726 32512 21732 32524
rect 21784 32512 21790 32564
rect 22462 32512 22468 32564
rect 22520 32552 22526 32564
rect 22649 32555 22707 32561
rect 22649 32552 22661 32555
rect 22520 32524 22661 32552
rect 22520 32512 22526 32524
rect 22649 32521 22661 32524
rect 22695 32521 22707 32555
rect 22649 32515 22707 32521
rect 22833 32555 22891 32561
rect 22833 32521 22845 32555
rect 22879 32552 22891 32555
rect 23826 32555 23884 32561
rect 23826 32552 23838 32555
rect 22879 32524 23838 32552
rect 22879 32521 22891 32524
rect 22833 32515 22891 32521
rect 23826 32521 23838 32524
rect 23872 32552 23884 32555
rect 24026 32552 24032 32564
rect 23872 32524 24032 32552
rect 23872 32521 23884 32524
rect 23826 32515 23884 32521
rect 13538 32484 13544 32496
rect 13499 32456 13544 32484
rect 13538 32444 13544 32456
rect 13596 32444 13602 32496
rect 21542 32484 21548 32496
rect 15856 32456 18460 32484
rect 15856 32428 15884 32456
rect 12529 32419 12587 32425
rect 12529 32385 12541 32419
rect 12575 32385 12587 32419
rect 13170 32416 13176 32428
rect 13131 32388 13176 32416
rect 12529 32379 12587 32385
rect 13170 32376 13176 32388
rect 13228 32376 13234 32428
rect 15378 32416 15384 32428
rect 15339 32388 15384 32416
rect 15378 32376 15384 32388
rect 15436 32416 15442 32428
rect 15838 32416 15844 32428
rect 15436 32388 15844 32416
rect 15436 32376 15442 32388
rect 15838 32376 15844 32388
rect 15896 32376 15902 32428
rect 16482 32416 16488 32428
rect 16395 32388 16488 32416
rect 16482 32376 16488 32388
rect 16540 32416 16546 32428
rect 17770 32416 17776 32428
rect 16540 32388 17776 32416
rect 16540 32376 16546 32388
rect 17770 32376 17776 32388
rect 17828 32376 17834 32428
rect 18432 32425 18460 32456
rect 20364 32456 21548 32484
rect 18417 32419 18475 32425
rect 18417 32385 18429 32419
rect 18463 32416 18475 32419
rect 18782 32416 18788 32428
rect 18463 32388 18788 32416
rect 18463 32385 18475 32388
rect 18417 32379 18475 32385
rect 18782 32376 18788 32388
rect 18840 32376 18846 32428
rect 19886 32376 19892 32428
rect 19944 32416 19950 32428
rect 20364 32425 20392 32456
rect 21542 32444 21548 32456
rect 21600 32444 21606 32496
rect 20349 32419 20407 32425
rect 20349 32416 20361 32419
rect 19944 32388 20361 32416
rect 19944 32376 19950 32388
rect 20349 32385 20361 32388
rect 20395 32385 20407 32419
rect 20349 32379 20407 32385
rect 20990 32376 20996 32428
rect 21048 32416 21054 32428
rect 21637 32419 21695 32425
rect 21637 32416 21649 32419
rect 21048 32388 21649 32416
rect 21048 32376 21054 32388
rect 21637 32385 21649 32388
rect 21683 32385 21695 32419
rect 21637 32379 21695 32385
rect 11517 32351 11575 32357
rect 11517 32317 11529 32351
rect 11563 32317 11575 32351
rect 11517 32311 11575 32317
rect 10959 32283 11017 32289
rect 10959 32249 10971 32283
rect 11005 32249 11017 32283
rect 11532 32280 11560 32311
rect 18874 32308 18880 32360
rect 18932 32348 18938 32360
rect 19521 32351 19579 32357
rect 19521 32348 19533 32351
rect 18932 32320 19533 32348
rect 18932 32308 18938 32320
rect 19521 32317 19533 32320
rect 19567 32348 19579 32351
rect 20254 32348 20260 32360
rect 19567 32320 20260 32348
rect 19567 32317 19579 32320
rect 19521 32311 19579 32317
rect 20254 32308 20260 32320
rect 20312 32308 20318 32360
rect 20809 32351 20867 32357
rect 20809 32317 20821 32351
rect 20855 32348 20867 32351
rect 21416 32351 21474 32357
rect 21416 32348 21428 32351
rect 20855 32320 21428 32348
rect 20855 32317 20867 32320
rect 20809 32311 20867 32317
rect 21416 32317 21428 32320
rect 21462 32348 21474 32351
rect 21726 32348 21732 32360
rect 21462 32320 21732 32348
rect 21462 32317 21474 32320
rect 21416 32311 21474 32317
rect 21726 32308 21732 32320
rect 21784 32348 21790 32360
rect 22664 32348 22692 32515
rect 24026 32512 24032 32524
rect 24084 32512 24090 32564
rect 24305 32555 24363 32561
rect 24305 32521 24317 32555
rect 24351 32552 24363 32555
rect 24946 32552 24952 32564
rect 24351 32524 24952 32552
rect 24351 32521 24363 32524
rect 24305 32515 24363 32521
rect 23106 32484 23112 32496
rect 23067 32456 23112 32484
rect 23106 32444 23112 32456
rect 23164 32444 23170 32496
rect 23934 32484 23940 32496
rect 23895 32456 23940 32484
rect 23934 32444 23940 32456
rect 23992 32444 23998 32496
rect 22738 32376 22744 32428
rect 22796 32416 22802 32428
rect 23477 32419 23535 32425
rect 23477 32416 23489 32419
rect 22796 32388 23489 32416
rect 22796 32376 22802 32388
rect 23477 32385 23489 32388
rect 23523 32416 23535 32419
rect 24029 32419 24087 32425
rect 24029 32416 24041 32419
rect 23523 32388 24041 32416
rect 23523 32385 23535 32388
rect 23477 32379 23535 32385
rect 24029 32385 24041 32388
rect 24075 32385 24087 32419
rect 24029 32379 24087 32385
rect 24320 32348 24348 32515
rect 24946 32512 24952 32524
rect 25004 32512 25010 32564
rect 27893 32555 27951 32561
rect 27893 32521 27905 32555
rect 27939 32552 27951 32555
rect 27982 32552 27988 32564
rect 27939 32524 27988 32552
rect 27939 32521 27951 32524
rect 27893 32515 27951 32521
rect 27982 32512 27988 32524
rect 28040 32552 28046 32564
rect 28997 32555 29055 32561
rect 28997 32552 29009 32555
rect 28040 32524 29009 32552
rect 28040 32512 28046 32524
rect 28997 32521 29009 32524
rect 29043 32521 29055 32555
rect 28997 32515 29055 32521
rect 32674 32512 32680 32564
rect 32732 32552 32738 32564
rect 32769 32555 32827 32561
rect 32769 32552 32781 32555
rect 32732 32524 32781 32552
rect 32732 32512 32738 32524
rect 32769 32521 32781 32524
rect 32815 32521 32827 32555
rect 32769 32515 32827 32521
rect 34054 32512 34060 32564
rect 34112 32552 34118 32564
rect 34241 32555 34299 32561
rect 34241 32552 34253 32555
rect 34112 32524 34253 32552
rect 34112 32512 34118 32524
rect 34241 32521 34253 32524
rect 34287 32552 34299 32555
rect 34330 32552 34336 32564
rect 34287 32524 34336 32552
rect 34287 32521 34299 32524
rect 34241 32515 34299 32521
rect 34330 32512 34336 32524
rect 34388 32512 34394 32564
rect 37182 32552 37188 32564
rect 37143 32524 37188 32552
rect 37182 32512 37188 32524
rect 37240 32512 37246 32564
rect 37826 32552 37832 32564
rect 37787 32524 37832 32552
rect 37826 32512 37832 32524
rect 37884 32512 37890 32564
rect 39758 32512 39764 32564
rect 39816 32552 39822 32564
rect 40129 32555 40187 32561
rect 40129 32552 40141 32555
rect 39816 32524 40141 32552
rect 39816 32512 39822 32524
rect 40129 32521 40141 32524
rect 40175 32521 40187 32555
rect 42610 32552 42616 32564
rect 42571 32524 42616 32552
rect 40129 32515 40187 32521
rect 42610 32512 42616 32524
rect 42668 32512 42674 32564
rect 43622 32552 43628 32564
rect 42766 32524 43628 32552
rect 29457 32487 29515 32493
rect 29457 32484 29469 32487
rect 28966 32456 29469 32484
rect 25130 32376 25136 32428
rect 25188 32416 25194 32428
rect 25225 32419 25283 32425
rect 25225 32416 25237 32419
rect 25188 32388 25237 32416
rect 25188 32376 25194 32388
rect 25225 32385 25237 32388
rect 25271 32416 25283 32419
rect 25682 32416 25688 32428
rect 25271 32388 25688 32416
rect 25271 32385 25283 32388
rect 25225 32379 25283 32385
rect 25682 32376 25688 32388
rect 25740 32376 25746 32428
rect 27430 32376 27436 32428
rect 27488 32416 27494 32428
rect 27985 32419 28043 32425
rect 27985 32416 27997 32419
rect 27488 32388 27997 32416
rect 27488 32376 27494 32388
rect 27985 32385 27997 32388
rect 28031 32385 28043 32419
rect 27985 32379 28043 32385
rect 27764 32351 27822 32357
rect 27764 32348 27776 32351
rect 21784 32320 22462 32348
rect 22664 32320 24348 32348
rect 26712 32320 27776 32348
rect 21784 32308 21790 32320
rect 12618 32280 12624 32292
rect 11532 32252 12624 32280
rect 10959 32243 11017 32249
rect 12618 32240 12624 32252
rect 12676 32280 12682 32292
rect 13538 32280 13544 32292
rect 12676 32252 13544 32280
rect 12676 32240 12682 32252
rect 13538 32240 13544 32252
rect 13596 32240 13602 32292
rect 14734 32280 14740 32292
rect 14695 32252 14740 32280
rect 14734 32240 14740 32252
rect 14792 32240 14798 32292
rect 14826 32240 14832 32292
rect 14884 32280 14890 32292
rect 16301 32283 16359 32289
rect 14884 32252 14929 32280
rect 14884 32240 14890 32252
rect 16301 32249 16313 32283
rect 16347 32280 16359 32283
rect 16577 32283 16635 32289
rect 16577 32280 16589 32283
rect 16347 32252 16589 32280
rect 16347 32249 16359 32252
rect 16301 32243 16359 32249
rect 16577 32249 16589 32252
rect 16623 32249 16635 32283
rect 17126 32280 17132 32292
rect 17087 32252 17132 32280
rect 16577 32243 16635 32249
rect 14553 32215 14611 32221
rect 14553 32181 14565 32215
rect 14599 32212 14611 32215
rect 14844 32212 14872 32240
rect 15746 32212 15752 32224
rect 14599 32184 14872 32212
rect 15707 32184 15752 32212
rect 14599 32181 14611 32184
rect 14553 32175 14611 32181
rect 15746 32172 15752 32184
rect 15804 32172 15810 32224
rect 16592 32212 16620 32243
rect 17126 32240 17132 32252
rect 17184 32240 17190 32292
rect 17678 32280 17684 32292
rect 17236 32252 17684 32280
rect 17236 32224 17264 32252
rect 17678 32240 17684 32252
rect 17736 32280 17742 32292
rect 17773 32283 17831 32289
rect 17773 32280 17785 32283
rect 17736 32252 17785 32280
rect 17736 32240 17742 32252
rect 17773 32249 17785 32252
rect 17819 32249 17831 32283
rect 17773 32243 17831 32249
rect 17218 32212 17224 32224
rect 16592 32184 17224 32212
rect 17218 32172 17224 32184
rect 17276 32172 17282 32224
rect 17788 32212 17816 32243
rect 17862 32240 17868 32292
rect 17920 32280 17926 32292
rect 18138 32280 18144 32292
rect 17920 32252 18144 32280
rect 17920 32240 17926 32252
rect 18138 32240 18144 32252
rect 18196 32240 18202 32292
rect 18233 32283 18291 32289
rect 18233 32249 18245 32283
rect 18279 32249 18291 32283
rect 18233 32243 18291 32249
rect 21269 32283 21327 32289
rect 21269 32249 21281 32283
rect 21315 32249 21327 32283
rect 22434 32280 22462 32320
rect 22833 32283 22891 32289
rect 22833 32280 22845 32283
rect 22434 32252 22845 32280
rect 21269 32243 21327 32249
rect 22833 32249 22845 32252
rect 22879 32249 22891 32283
rect 22833 32243 22891 32249
rect 18248 32212 18276 32243
rect 17788 32184 18276 32212
rect 19058 32172 19064 32224
rect 19116 32212 19122 32224
rect 19153 32215 19211 32221
rect 19153 32212 19165 32215
rect 19116 32184 19165 32212
rect 19116 32172 19122 32184
rect 19153 32181 19165 32184
rect 19199 32212 19211 32215
rect 19978 32212 19984 32224
rect 19199 32184 19984 32212
rect 19199 32181 19211 32184
rect 19153 32175 19211 32181
rect 19978 32172 19984 32184
rect 20036 32172 20042 32224
rect 20990 32172 20996 32224
rect 21048 32212 21054 32224
rect 21085 32215 21143 32221
rect 21085 32212 21097 32215
rect 21048 32184 21097 32212
rect 21048 32172 21054 32184
rect 21085 32181 21097 32184
rect 21131 32181 21143 32215
rect 21284 32212 21312 32243
rect 23106 32240 23112 32292
rect 23164 32280 23170 32292
rect 23661 32283 23719 32289
rect 23661 32280 23673 32283
rect 23164 32252 23673 32280
rect 23164 32240 23170 32252
rect 23661 32249 23673 32252
rect 23707 32280 23719 32283
rect 24673 32283 24731 32289
rect 24673 32280 24685 32283
rect 23707 32252 24685 32280
rect 23707 32249 23719 32252
rect 23661 32243 23719 32249
rect 24673 32249 24685 32252
rect 24719 32280 24731 32283
rect 26602 32280 26608 32292
rect 24719 32252 26608 32280
rect 24719 32249 24731 32252
rect 24673 32243 24731 32249
rect 26602 32240 26608 32252
rect 26660 32240 26666 32292
rect 26712 32224 26740 32320
rect 27764 32317 27776 32320
rect 27810 32348 27822 32351
rect 28258 32348 28264 32360
rect 27810 32320 28264 32348
rect 27810 32317 27822 32320
rect 27764 32311 27822 32317
rect 28258 32308 28264 32320
rect 28316 32348 28322 32360
rect 28966 32348 28994 32456
rect 29457 32453 29469 32456
rect 29503 32453 29515 32487
rect 37844 32484 37872 32512
rect 39850 32484 39856 32496
rect 37844 32456 39856 32484
rect 29457 32447 29515 32453
rect 39850 32444 39856 32456
rect 39908 32484 39914 32496
rect 42766 32484 42794 32524
rect 43622 32512 43628 32524
rect 43680 32512 43686 32564
rect 44821 32555 44879 32561
rect 44821 32521 44833 32555
rect 44867 32552 44879 32555
rect 45094 32552 45100 32564
rect 44867 32524 45100 32552
rect 44867 32521 44879 32524
rect 44821 32515 44879 32521
rect 44358 32484 44364 32496
rect 39908 32456 42794 32484
rect 44319 32456 44364 32484
rect 39908 32444 39914 32456
rect 44358 32444 44364 32456
rect 44416 32444 44422 32496
rect 29917 32419 29975 32425
rect 29917 32385 29929 32419
rect 29963 32416 29975 32419
rect 31570 32416 31576 32428
rect 29963 32388 31576 32416
rect 29963 32385 29975 32388
rect 29917 32379 29975 32385
rect 31570 32376 31576 32388
rect 31628 32376 31634 32428
rect 32766 32416 32772 32428
rect 31680 32388 32772 32416
rect 31294 32348 31300 32360
rect 28316 32320 28994 32348
rect 31207 32320 31300 32348
rect 28316 32308 28322 32320
rect 31294 32308 31300 32320
rect 31352 32348 31358 32360
rect 31680 32357 31708 32388
rect 32766 32376 32772 32388
rect 32824 32376 32830 32428
rect 34790 32376 34796 32428
rect 34848 32416 34854 32428
rect 34977 32419 35035 32425
rect 34977 32416 34989 32419
rect 34848 32388 34989 32416
rect 34848 32376 34854 32388
rect 34977 32385 34989 32388
rect 35023 32385 35035 32419
rect 35434 32416 35440 32428
rect 35395 32388 35440 32416
rect 34977 32379 35035 32385
rect 35434 32376 35440 32388
rect 35492 32376 35498 32428
rect 38470 32416 38476 32428
rect 38431 32388 38476 32416
rect 38470 32376 38476 32388
rect 38528 32376 38534 32428
rect 39117 32419 39175 32425
rect 39117 32385 39129 32419
rect 39163 32416 39175 32419
rect 41138 32416 41144 32428
rect 39163 32388 41144 32416
rect 39163 32385 39175 32388
rect 39117 32379 39175 32385
rect 41138 32376 41144 32388
rect 41196 32376 41202 32428
rect 43809 32419 43867 32425
rect 43809 32385 43821 32419
rect 43855 32416 43867 32419
rect 44836 32416 44864 32515
rect 45094 32512 45100 32524
rect 45152 32512 45158 32564
rect 43855 32388 44864 32416
rect 43855 32385 43867 32388
rect 43809 32379 43867 32385
rect 31665 32351 31723 32357
rect 31665 32348 31677 32351
rect 31352 32320 31677 32348
rect 31352 32308 31358 32320
rect 31665 32317 31677 32320
rect 31711 32317 31723 32351
rect 31938 32348 31944 32360
rect 31851 32320 31944 32348
rect 31665 32311 31723 32317
rect 31938 32308 31944 32320
rect 31996 32348 32002 32360
rect 32674 32348 32680 32360
rect 31996 32320 32680 32348
rect 31996 32308 32002 32320
rect 32674 32308 32680 32320
rect 32732 32308 32738 32360
rect 37436 32351 37494 32357
rect 37436 32317 37448 32351
rect 37482 32348 37494 32351
rect 37482 32320 38056 32348
rect 37482 32317 37494 32320
rect 37436 32311 37494 32317
rect 27157 32283 27215 32289
rect 27157 32249 27169 32283
rect 27203 32280 27215 32283
rect 27522 32280 27528 32292
rect 27203 32252 27528 32280
rect 27203 32249 27215 32252
rect 27157 32243 27215 32249
rect 27522 32240 27528 32252
rect 27580 32280 27586 32292
rect 27617 32283 27675 32289
rect 27617 32280 27629 32283
rect 27580 32252 27629 32280
rect 27580 32240 27586 32252
rect 27617 32249 27629 32252
rect 27663 32249 27675 32283
rect 27617 32243 27675 32249
rect 28353 32283 28411 32289
rect 28353 32249 28365 32283
rect 28399 32280 28411 32283
rect 29914 32280 29920 32292
rect 28399 32252 29920 32280
rect 28399 32249 28411 32252
rect 28353 32243 28411 32249
rect 29914 32240 29920 32252
rect 29972 32240 29978 32292
rect 30006 32240 30012 32292
rect 30064 32280 30070 32292
rect 30558 32280 30564 32292
rect 30064 32252 30109 32280
rect 30519 32252 30564 32280
rect 30064 32240 30070 32252
rect 30558 32240 30564 32252
rect 30616 32240 30622 32292
rect 32122 32280 32128 32292
rect 32083 32252 32128 32280
rect 32122 32240 32128 32252
rect 32180 32240 32186 32292
rect 35069 32283 35127 32289
rect 35069 32280 35081 32283
rect 34624 32252 35081 32280
rect 21358 32212 21364 32224
rect 21284 32184 21364 32212
rect 21085 32175 21143 32181
rect 21358 32172 21364 32184
rect 21416 32172 21422 32224
rect 22278 32212 22284 32224
rect 22239 32184 22284 32212
rect 22278 32172 22284 32184
rect 22336 32172 22342 32224
rect 24762 32172 24768 32224
rect 24820 32212 24826 32224
rect 25133 32215 25191 32221
rect 25133 32212 25145 32215
rect 24820 32184 25145 32212
rect 24820 32172 24826 32184
rect 25133 32181 25145 32184
rect 25179 32212 25191 32215
rect 25593 32215 25651 32221
rect 25593 32212 25605 32215
rect 25179 32184 25605 32212
rect 25179 32181 25191 32184
rect 25133 32175 25191 32181
rect 25593 32181 25605 32184
rect 25639 32181 25651 32215
rect 25593 32175 25651 32181
rect 26145 32215 26203 32221
rect 26145 32181 26157 32215
rect 26191 32212 26203 32215
rect 26418 32212 26424 32224
rect 26191 32184 26424 32212
rect 26191 32181 26203 32184
rect 26145 32175 26203 32181
rect 26418 32172 26424 32184
rect 26476 32172 26482 32224
rect 26694 32212 26700 32224
rect 26655 32184 26700 32212
rect 26694 32172 26700 32184
rect 26752 32172 26758 32224
rect 27430 32212 27436 32224
rect 27391 32184 27436 32212
rect 27430 32172 27436 32184
rect 27488 32172 27494 32224
rect 27798 32172 27804 32224
rect 27856 32212 27862 32224
rect 28626 32212 28632 32224
rect 27856 32184 28632 32212
rect 27856 32172 27862 32184
rect 28626 32172 28632 32184
rect 28684 32172 28690 32224
rect 30466 32172 30472 32224
rect 30524 32212 30530 32224
rect 30929 32215 30987 32221
rect 30929 32212 30941 32215
rect 30524 32184 30941 32212
rect 30524 32172 30530 32184
rect 30929 32181 30941 32184
rect 30975 32212 30987 32215
rect 32306 32212 32312 32224
rect 30975 32184 32312 32212
rect 30975 32181 30987 32184
rect 30929 32175 30987 32181
rect 32306 32172 32312 32184
rect 32364 32172 32370 32224
rect 32493 32215 32551 32221
rect 32493 32181 32505 32215
rect 32539 32212 32551 32215
rect 32582 32212 32588 32224
rect 32539 32184 32588 32212
rect 32539 32181 32551 32184
rect 32493 32175 32551 32181
rect 32582 32172 32588 32184
rect 32640 32172 32646 32224
rect 32953 32215 33011 32221
rect 32953 32181 32965 32215
rect 32999 32212 33011 32215
rect 33042 32212 33048 32224
rect 32999 32184 33048 32212
rect 32999 32181 33011 32184
rect 32953 32175 33011 32181
rect 33042 32172 33048 32184
rect 33100 32172 33106 32224
rect 34514 32172 34520 32224
rect 34572 32212 34578 32224
rect 34624 32221 34652 32252
rect 35069 32249 35081 32252
rect 35115 32249 35127 32283
rect 35069 32243 35127 32249
rect 38028 32224 38056 32320
rect 42150 32308 42156 32360
rect 42208 32348 42214 32360
rect 42740 32351 42798 32357
rect 42740 32348 42752 32351
rect 42208 32320 42752 32348
rect 42208 32308 42214 32320
rect 42740 32317 42752 32320
rect 42786 32348 42798 32351
rect 43165 32351 43223 32357
rect 43165 32348 43177 32351
rect 42786 32320 43177 32348
rect 42786 32317 42798 32320
rect 42740 32311 42798 32317
rect 43165 32317 43177 32320
rect 43211 32317 43223 32351
rect 43165 32311 43223 32317
rect 38562 32280 38568 32292
rect 38523 32252 38568 32280
rect 38562 32240 38568 32252
rect 38620 32240 38626 32292
rect 41046 32280 41052 32292
rect 41007 32252 41052 32280
rect 41046 32240 41052 32252
rect 41104 32240 41110 32292
rect 41141 32283 41199 32289
rect 41141 32249 41153 32283
rect 41187 32249 41199 32283
rect 41690 32280 41696 32292
rect 41651 32252 41696 32280
rect 41141 32243 41199 32249
rect 34609 32215 34667 32221
rect 34609 32212 34621 32215
rect 34572 32184 34621 32212
rect 34572 32172 34578 32184
rect 34609 32181 34621 32184
rect 34655 32181 34667 32215
rect 34609 32175 34667 32181
rect 36173 32215 36231 32221
rect 36173 32181 36185 32215
rect 36219 32212 36231 32215
rect 36262 32212 36268 32224
rect 36219 32184 36268 32212
rect 36219 32181 36231 32184
rect 36173 32175 36231 32181
rect 36262 32172 36268 32184
rect 36320 32172 36326 32224
rect 36538 32212 36544 32224
rect 36451 32184 36544 32212
rect 36538 32172 36544 32184
rect 36596 32212 36602 32224
rect 36814 32212 36820 32224
rect 36596 32184 36820 32212
rect 36596 32172 36602 32184
rect 36814 32172 36820 32184
rect 36872 32172 36878 32224
rect 37507 32215 37565 32221
rect 37507 32181 37519 32215
rect 37553 32212 37565 32215
rect 37734 32212 37740 32224
rect 37553 32184 37740 32212
rect 37553 32181 37565 32184
rect 37507 32175 37565 32181
rect 37734 32172 37740 32184
rect 37792 32172 37798 32224
rect 38010 32172 38016 32224
rect 38068 32212 38074 32224
rect 38197 32215 38255 32221
rect 38197 32212 38209 32215
rect 38068 32184 38209 32212
rect 38068 32172 38074 32184
rect 38197 32181 38209 32184
rect 38243 32181 38255 32215
rect 38580 32212 38608 32240
rect 39393 32215 39451 32221
rect 39393 32212 39405 32215
rect 38580 32184 39405 32212
rect 38197 32175 38255 32181
rect 39393 32181 39405 32184
rect 39439 32181 39451 32215
rect 40862 32212 40868 32224
rect 40823 32184 40868 32212
rect 39393 32175 39451 32181
rect 40862 32172 40868 32184
rect 40920 32212 40926 32224
rect 41156 32212 41184 32243
rect 41690 32240 41696 32252
rect 41748 32240 41754 32292
rect 43901 32283 43959 32289
rect 43901 32249 43913 32283
rect 43947 32280 43959 32283
rect 44082 32280 44088 32292
rect 43947 32252 44088 32280
rect 43947 32249 43959 32252
rect 43901 32243 43959 32249
rect 44082 32240 44088 32252
rect 44140 32240 44146 32292
rect 41969 32215 42027 32221
rect 41969 32212 41981 32215
rect 40920 32184 41981 32212
rect 40920 32172 40926 32184
rect 41969 32181 41981 32184
rect 42015 32181 42027 32215
rect 41969 32175 42027 32181
rect 42843 32215 42901 32221
rect 42843 32181 42855 32215
rect 42889 32212 42901 32215
rect 43622 32212 43628 32224
rect 42889 32184 43628 32212
rect 42889 32181 42901 32184
rect 42843 32175 42901 32181
rect 43622 32172 43628 32184
rect 43680 32172 43686 32224
rect 1104 32122 48852 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 48852 32122
rect 1104 32048 48852 32070
rect 10502 32008 10508 32020
rect 10463 31980 10508 32008
rect 10502 31968 10508 31980
rect 10560 31968 10566 32020
rect 11422 32008 11428 32020
rect 11383 31980 11428 32008
rect 11422 31968 11428 31980
rect 11480 31968 11486 32020
rect 12618 32008 12624 32020
rect 12579 31980 12624 32008
rect 12618 31968 12624 31980
rect 12676 31968 12682 32020
rect 12989 32011 13047 32017
rect 12989 31977 13001 32011
rect 13035 32008 13047 32011
rect 13170 32008 13176 32020
rect 13035 31980 13176 32008
rect 13035 31977 13047 31980
rect 12989 31971 13047 31977
rect 13170 31968 13176 31980
rect 13228 31968 13234 32020
rect 16482 32008 16488 32020
rect 16443 31980 16488 32008
rect 16482 31968 16488 31980
rect 16540 31968 16546 32020
rect 18230 32008 18236 32020
rect 18143 31980 18236 32008
rect 18230 31968 18236 31980
rect 18288 32008 18294 32020
rect 18874 32008 18880 32020
rect 18288 31980 18880 32008
rect 18288 31968 18294 31980
rect 18874 31968 18880 31980
rect 18932 31968 18938 32020
rect 20070 32008 20076 32020
rect 19260 31980 20076 32008
rect 12526 31900 12532 31952
rect 12584 31940 12590 31952
rect 13265 31943 13323 31949
rect 13265 31940 13277 31943
rect 12584 31912 13277 31940
rect 12584 31900 12590 31912
rect 13265 31909 13277 31912
rect 13311 31940 13323 31943
rect 13446 31940 13452 31952
rect 13311 31912 13452 31940
rect 13311 31909 13323 31912
rect 13265 31903 13323 31909
rect 13446 31900 13452 31912
rect 13504 31940 13510 31952
rect 14826 31940 14832 31952
rect 13504 31912 14832 31940
rect 13504 31900 13510 31912
rect 14826 31900 14832 31912
rect 14884 31900 14890 31952
rect 15470 31940 15476 31952
rect 15431 31912 15476 31940
rect 15470 31900 15476 31912
rect 15528 31900 15534 31952
rect 16942 31900 16948 31952
rect 17000 31940 17006 31952
rect 17129 31943 17187 31949
rect 17129 31940 17141 31943
rect 17000 31912 17141 31940
rect 17000 31900 17006 31912
rect 17129 31909 17141 31912
rect 17175 31909 17187 31943
rect 17129 31903 17187 31909
rect 17218 31900 17224 31952
rect 17276 31940 17282 31952
rect 19260 31949 19288 31980
rect 20070 31968 20076 31980
rect 20128 32008 20134 32020
rect 23106 32008 23112 32020
rect 20128 31980 23112 32008
rect 20128 31968 20134 31980
rect 23106 31968 23112 31980
rect 23164 31968 23170 32020
rect 23290 32008 23296 32020
rect 23251 31980 23296 32008
rect 23290 31968 23296 31980
rect 23348 31968 23354 32020
rect 23753 32011 23811 32017
rect 23753 32008 23765 32011
rect 23446 31980 23765 32008
rect 23446 31952 23474 31980
rect 23753 31977 23765 31980
rect 23799 32008 23811 32011
rect 23934 32008 23940 32020
rect 23799 31980 23940 32008
rect 23799 31977 23811 31980
rect 23753 31971 23811 31977
rect 23934 31968 23940 31980
rect 23992 31968 23998 32020
rect 24026 31968 24032 32020
rect 24084 32008 24090 32020
rect 24084 31980 24129 32008
rect 24084 31968 24090 31980
rect 25222 31968 25228 32020
rect 25280 32008 25286 32020
rect 25777 32011 25835 32017
rect 25777 32008 25789 32011
rect 25280 31980 25789 32008
rect 25280 31968 25286 31980
rect 25777 31977 25789 31980
rect 25823 31977 25835 32011
rect 26326 32008 26332 32020
rect 26287 31980 26332 32008
rect 25777 31971 25835 31977
rect 26326 31968 26332 31980
rect 26384 31968 26390 32020
rect 26418 31968 26424 32020
rect 26476 32008 26482 32020
rect 26973 32011 27031 32017
rect 26973 32008 26985 32011
rect 26476 31980 26985 32008
rect 26476 31968 26482 31980
rect 26973 31977 26985 31980
rect 27019 31977 27031 32011
rect 30742 32008 30748 32020
rect 30703 31980 30748 32008
rect 26973 31971 27031 31977
rect 30742 31968 30748 31980
rect 30800 31968 30806 32020
rect 31481 32011 31539 32017
rect 31481 31977 31493 32011
rect 31527 32008 31539 32011
rect 31938 32008 31944 32020
rect 31527 31980 31944 32008
rect 31527 31977 31539 31980
rect 31481 31971 31539 31977
rect 31938 31968 31944 31980
rect 31996 31968 32002 32020
rect 32490 32008 32496 32020
rect 32451 31980 32496 32008
rect 32490 31968 32496 31980
rect 32548 31968 32554 32020
rect 38470 31968 38476 32020
rect 38528 32008 38534 32020
rect 38933 32011 38991 32017
rect 38933 32008 38945 32011
rect 38528 31980 38945 32008
rect 38528 31968 38534 31980
rect 38933 31977 38945 31980
rect 38979 31977 38991 32011
rect 38933 31971 38991 31977
rect 39807 32011 39865 32017
rect 39807 31977 39819 32011
rect 39853 32008 39865 32011
rect 41598 32008 41604 32020
rect 39853 31980 41604 32008
rect 39853 31977 39865 31980
rect 39807 31971 39865 31977
rect 41598 31968 41604 31980
rect 41656 32008 41662 32020
rect 41693 32011 41751 32017
rect 41693 32008 41705 32011
rect 41656 31980 41705 32008
rect 41656 31968 41662 31980
rect 41693 31977 41705 31980
rect 41739 31977 41751 32011
rect 41693 31971 41751 31977
rect 43714 31968 43720 32020
rect 43772 32008 43778 32020
rect 45143 32011 45201 32017
rect 45143 32008 45155 32011
rect 43772 31980 45155 32008
rect 43772 31968 43778 31980
rect 45143 31977 45155 31980
rect 45189 31977 45201 32011
rect 45143 31971 45201 31977
rect 18785 31943 18843 31949
rect 17276 31912 17321 31940
rect 17276 31900 17282 31912
rect 18785 31909 18797 31943
rect 18831 31940 18843 31943
rect 19245 31943 19303 31949
rect 19245 31940 19257 31943
rect 18831 31912 19257 31940
rect 18831 31909 18843 31912
rect 18785 31903 18843 31909
rect 19245 31909 19257 31912
rect 19291 31909 19303 31943
rect 19245 31903 19303 31909
rect 21542 31900 21548 31952
rect 21600 31940 21606 31952
rect 23446 31940 23480 31952
rect 21600 31912 23480 31940
rect 21600 31900 21606 31912
rect 9674 31832 9680 31884
rect 9732 31872 9738 31884
rect 10410 31872 10416 31884
rect 9732 31844 10416 31872
rect 9732 31832 9738 31844
rect 10410 31832 10416 31844
rect 10468 31832 10474 31884
rect 10686 31832 10692 31884
rect 10744 31872 10750 31884
rect 10873 31875 10931 31881
rect 10873 31872 10885 31875
rect 10744 31844 10885 31872
rect 10744 31832 10750 31844
rect 10873 31841 10885 31844
rect 10919 31841 10931 31875
rect 10873 31835 10931 31841
rect 12120 31875 12178 31881
rect 12120 31841 12132 31875
rect 12166 31872 12178 31875
rect 12342 31872 12348 31884
rect 12166 31844 12348 31872
rect 12166 31841 12178 31844
rect 12120 31835 12178 31841
rect 12342 31832 12348 31844
rect 12400 31872 12406 31884
rect 12986 31872 12992 31884
rect 12400 31844 12992 31872
rect 12400 31832 12406 31844
rect 12986 31832 12992 31844
rect 13044 31832 13050 31884
rect 19334 31832 19340 31884
rect 19392 31872 19398 31884
rect 19981 31875 20039 31881
rect 19981 31872 19993 31875
rect 19392 31844 19993 31872
rect 19392 31832 19398 31844
rect 19981 31841 19993 31844
rect 20027 31841 20039 31875
rect 19981 31835 20039 31841
rect 20806 31832 20812 31884
rect 20864 31872 20870 31884
rect 21120 31875 21178 31881
rect 21120 31872 21132 31875
rect 20864 31844 21132 31872
rect 20864 31832 20870 31844
rect 21120 31841 21132 31844
rect 21166 31872 21178 31875
rect 22186 31872 22192 31884
rect 21166 31844 22192 31872
rect 21166 31841 21178 31844
rect 21120 31835 21178 31841
rect 22186 31832 22192 31844
rect 22244 31832 22250 31884
rect 22388 31881 22416 31912
rect 23474 31900 23480 31912
rect 23532 31900 23538 31952
rect 24854 31940 24860 31952
rect 24412 31912 24860 31940
rect 22373 31875 22431 31881
rect 22373 31841 22385 31875
rect 22419 31841 22431 31875
rect 22646 31872 22652 31884
rect 22607 31844 22652 31872
rect 22373 31835 22431 31841
rect 22646 31832 22652 31844
rect 22704 31832 22710 31884
rect 24412 31881 24440 31912
rect 24854 31900 24860 31912
rect 24912 31900 24918 31952
rect 25130 31940 25136 31952
rect 25091 31912 25136 31940
rect 25130 31900 25136 31912
rect 25188 31900 25194 31952
rect 26602 31900 26608 31952
rect 26660 31940 26666 31952
rect 28074 31940 28080 31952
rect 26660 31912 28080 31940
rect 26660 31900 26666 31912
rect 28074 31900 28080 31912
rect 28132 31940 28138 31952
rect 28442 31940 28448 31952
rect 28132 31912 28279 31940
rect 28403 31912 28448 31940
rect 28132 31900 28138 31912
rect 24397 31875 24455 31881
rect 24397 31841 24409 31875
rect 24443 31841 24455 31875
rect 24397 31835 24455 31841
rect 24486 31832 24492 31884
rect 24544 31872 24550 31884
rect 24946 31872 24952 31884
rect 24544 31844 24952 31872
rect 24544 31832 24550 31844
rect 24946 31832 24952 31844
rect 25004 31832 25010 31884
rect 26418 31872 26424 31884
rect 26379 31844 26424 31872
rect 26418 31832 26424 31844
rect 26476 31832 26482 31884
rect 27522 31832 27528 31884
rect 27580 31872 27586 31884
rect 27709 31875 27767 31881
rect 27709 31872 27721 31875
rect 27580 31844 27721 31872
rect 27580 31832 27586 31844
rect 27709 31841 27721 31844
rect 27755 31841 27767 31875
rect 28251 31872 28279 31912
rect 28442 31900 28448 31912
rect 28500 31900 28506 31952
rect 29917 31943 29975 31949
rect 29917 31909 29929 31943
rect 29963 31940 29975 31943
rect 30006 31940 30012 31952
rect 29963 31912 30012 31940
rect 29963 31909 29975 31912
rect 29917 31903 29975 31909
rect 30006 31900 30012 31912
rect 30064 31900 30070 31952
rect 34514 31900 34520 31952
rect 34572 31940 34578 31952
rect 34609 31943 34667 31949
rect 34609 31940 34621 31943
rect 34572 31912 34621 31940
rect 34572 31900 34578 31912
rect 34609 31909 34621 31912
rect 34655 31909 34667 31943
rect 36078 31940 36084 31952
rect 36039 31912 36084 31940
rect 34609 31903 34667 31909
rect 36078 31900 36084 31912
rect 36136 31900 36142 31952
rect 36170 31900 36176 31952
rect 36228 31940 36234 31952
rect 36228 31912 36273 31940
rect 36228 31900 36234 31912
rect 37734 31900 37740 31952
rect 37792 31940 37798 31952
rect 38013 31943 38071 31949
rect 38013 31940 38025 31943
rect 37792 31912 38025 31940
rect 37792 31900 37798 31912
rect 38013 31909 38025 31912
rect 38059 31909 38071 31943
rect 38013 31903 38071 31909
rect 38102 31900 38108 31952
rect 38160 31940 38166 31952
rect 38160 31912 38205 31940
rect 38160 31900 38166 31912
rect 40310 31900 40316 31952
rect 40368 31940 40374 31952
rect 40862 31940 40868 31952
rect 40368 31912 40868 31940
rect 40368 31900 40374 31912
rect 40862 31900 40868 31912
rect 40920 31900 40926 31952
rect 43625 31943 43683 31949
rect 43625 31909 43637 31943
rect 43671 31940 43683 31943
rect 43990 31940 43996 31952
rect 43671 31912 43996 31940
rect 43671 31909 43683 31912
rect 43625 31903 43683 31909
rect 43990 31900 43996 31912
rect 44048 31900 44054 31952
rect 28721 31875 28779 31881
rect 28721 31872 28733 31875
rect 28251 31844 28733 31872
rect 27709 31835 27767 31841
rect 28721 31841 28733 31844
rect 28767 31841 28779 31875
rect 28721 31835 28779 31841
rect 38930 31832 38936 31884
rect 38988 31872 38994 31884
rect 39736 31875 39794 31881
rect 39736 31872 39748 31875
rect 38988 31844 39748 31872
rect 38988 31832 38994 31844
rect 39736 31841 39748 31844
rect 39782 31872 39794 31875
rect 39850 31872 39856 31884
rect 39782 31844 39856 31872
rect 39782 31841 39794 31844
rect 39736 31835 39794 31841
rect 39850 31832 39856 31844
rect 39908 31832 39914 31884
rect 42242 31872 42248 31884
rect 42203 31844 42248 31872
rect 42242 31832 42248 31844
rect 42300 31832 42306 31884
rect 45005 31875 45063 31881
rect 45005 31841 45017 31875
rect 45051 31872 45063 31875
rect 45094 31872 45100 31884
rect 45051 31844 45100 31872
rect 45051 31841 45063 31844
rect 45005 31835 45063 31841
rect 45094 31832 45100 31844
rect 45152 31832 45158 31884
rect 12207 31807 12265 31813
rect 12207 31773 12219 31807
rect 12253 31804 12265 31807
rect 13173 31807 13231 31813
rect 13173 31804 13185 31807
rect 12253 31776 13185 31804
rect 12253 31773 12265 31776
rect 12207 31767 12265 31773
rect 13173 31773 13185 31776
rect 13219 31804 13231 31807
rect 13814 31804 13820 31816
rect 13219 31776 13820 31804
rect 13219 31773 13231 31776
rect 13173 31767 13231 31773
rect 13814 31764 13820 31776
rect 13872 31764 13878 31816
rect 15378 31804 15384 31816
rect 15339 31776 15384 31804
rect 15378 31764 15384 31776
rect 15436 31764 15442 31816
rect 17405 31807 17463 31813
rect 17405 31773 17417 31807
rect 17451 31773 17463 31807
rect 19610 31804 19616 31816
rect 19571 31776 19616 31804
rect 17405 31767 17463 31773
rect 13722 31736 13728 31748
rect 13683 31708 13728 31736
rect 13722 31696 13728 31708
rect 13780 31696 13786 31748
rect 15930 31736 15936 31748
rect 15891 31708 15936 31736
rect 15930 31696 15936 31708
rect 15988 31736 15994 31748
rect 17420 31736 17448 31767
rect 19610 31764 19616 31776
rect 19668 31804 19674 31816
rect 20990 31804 20996 31816
rect 19668 31776 20996 31804
rect 19668 31764 19674 31776
rect 20990 31764 20996 31776
rect 21048 31764 21054 31816
rect 22465 31807 22523 31813
rect 22465 31773 22477 31807
rect 22511 31804 22523 31807
rect 26694 31804 26700 31816
rect 22511 31776 26700 31804
rect 22511 31773 22523 31776
rect 22465 31767 22523 31773
rect 26694 31764 26700 31776
rect 26752 31804 26758 31816
rect 27154 31804 27160 31816
rect 26752 31776 27160 31804
rect 26752 31764 26758 31776
rect 27154 31764 27160 31776
rect 27212 31804 27218 31816
rect 27212 31776 27568 31804
rect 27212 31764 27218 31776
rect 17494 31736 17500 31748
rect 15988 31708 17500 31736
rect 15988 31696 15994 31708
rect 17494 31696 17500 31708
rect 17552 31696 17558 31748
rect 19153 31739 19211 31745
rect 19153 31705 19165 31739
rect 19199 31736 19211 31739
rect 19521 31739 19579 31745
rect 19521 31736 19533 31739
rect 19199 31708 19533 31736
rect 19199 31705 19211 31708
rect 19153 31699 19211 31705
rect 19521 31705 19533 31708
rect 19567 31736 19579 31739
rect 19886 31736 19892 31748
rect 19567 31708 19892 31736
rect 19567 31705 19579 31708
rect 19521 31699 19579 31705
rect 19886 31696 19892 31708
rect 19944 31696 19950 31748
rect 21223 31739 21281 31745
rect 21223 31705 21235 31739
rect 21269 31736 21281 31739
rect 26326 31736 26332 31748
rect 21269 31708 26332 31736
rect 21269 31705 21281 31708
rect 21223 31699 21281 31705
rect 26326 31696 26332 31708
rect 26384 31696 26390 31748
rect 12986 31628 12992 31680
rect 13044 31668 13050 31680
rect 14645 31671 14703 31677
rect 14645 31668 14657 31671
rect 13044 31640 14657 31668
rect 13044 31628 13050 31640
rect 14645 31637 14657 31640
rect 14691 31668 14703 31671
rect 14734 31668 14740 31680
rect 14691 31640 14740 31668
rect 14691 31637 14703 31640
rect 14645 31631 14703 31637
rect 14734 31628 14740 31640
rect 14792 31628 14798 31680
rect 16853 31671 16911 31677
rect 16853 31637 16865 31671
rect 16899 31668 16911 31671
rect 17034 31668 17040 31680
rect 16899 31640 17040 31668
rect 16899 31637 16911 31640
rect 16853 31631 16911 31637
rect 17034 31628 17040 31640
rect 17092 31628 17098 31680
rect 19426 31677 19432 31680
rect 19410 31671 19432 31677
rect 19410 31637 19422 31671
rect 19410 31631 19432 31637
rect 19426 31628 19432 31631
rect 19484 31628 19490 31680
rect 20346 31668 20352 31680
rect 20307 31640 20352 31668
rect 20346 31628 20352 31640
rect 20404 31668 20410 31680
rect 21358 31668 21364 31680
rect 20404 31640 21364 31668
rect 20404 31628 20410 31640
rect 21358 31628 21364 31640
rect 21416 31668 21422 31680
rect 21545 31671 21603 31677
rect 21545 31668 21557 31671
rect 21416 31640 21557 31668
rect 21416 31628 21422 31640
rect 21545 31637 21557 31640
rect 21591 31637 21603 31671
rect 25406 31668 25412 31680
rect 25367 31640 25412 31668
rect 21545 31631 21603 31637
rect 25406 31628 25412 31640
rect 25464 31628 25470 31680
rect 25866 31628 25872 31680
rect 25924 31668 25930 31680
rect 26651 31671 26709 31677
rect 26651 31668 26663 31671
rect 25924 31640 26663 31668
rect 25924 31628 25930 31640
rect 26651 31637 26663 31640
rect 26697 31637 26709 31671
rect 27540 31668 27568 31776
rect 27798 31764 27804 31816
rect 27856 31804 27862 31816
rect 28077 31807 28135 31813
rect 28077 31804 28089 31807
rect 27856 31776 28089 31804
rect 27856 31764 27862 31776
rect 28077 31773 28089 31776
rect 28123 31773 28135 31807
rect 28077 31767 28135 31773
rect 29546 31764 29552 31816
rect 29604 31804 29610 31816
rect 29825 31807 29883 31813
rect 29825 31804 29837 31807
rect 29604 31776 29837 31804
rect 29604 31764 29610 31776
rect 29825 31773 29837 31776
rect 29871 31773 29883 31807
rect 32122 31804 32128 31816
rect 32035 31776 32128 31804
rect 29825 31767 29883 31773
rect 32122 31764 32128 31776
rect 32180 31804 32186 31816
rect 32674 31804 32680 31816
rect 32180 31776 32680 31804
rect 32180 31764 32186 31776
rect 32674 31764 32680 31776
rect 32732 31764 32738 31816
rect 33962 31764 33968 31816
rect 34020 31804 34026 31816
rect 34517 31807 34575 31813
rect 34517 31804 34529 31807
rect 34020 31776 34529 31804
rect 34020 31764 34026 31776
rect 34517 31773 34529 31776
rect 34563 31773 34575 31807
rect 34517 31767 34575 31773
rect 34793 31807 34851 31813
rect 34793 31773 34805 31807
rect 34839 31773 34851 31807
rect 34793 31767 34851 31773
rect 27617 31739 27675 31745
rect 27617 31705 27629 31739
rect 27663 31736 27675 31739
rect 28166 31736 28172 31748
rect 27663 31708 28172 31736
rect 27663 31705 27675 31708
rect 27617 31699 27675 31705
rect 28166 31696 28172 31708
rect 28224 31696 28230 31748
rect 30282 31696 30288 31748
rect 30340 31736 30346 31748
rect 30377 31739 30435 31745
rect 30377 31736 30389 31739
rect 30340 31708 30389 31736
rect 30340 31696 30346 31708
rect 30377 31705 30389 31708
rect 30423 31736 30435 31739
rect 34808 31736 34836 31767
rect 35250 31764 35256 31816
rect 35308 31804 35314 31816
rect 36357 31807 36415 31813
rect 36357 31804 36369 31807
rect 35308 31776 36369 31804
rect 35308 31764 35314 31776
rect 36357 31773 36369 31776
rect 36403 31773 36415 31807
rect 38378 31804 38384 31816
rect 38339 31776 38384 31804
rect 36357 31767 36415 31773
rect 38378 31764 38384 31776
rect 38436 31764 38442 31816
rect 40770 31804 40776 31816
rect 40731 31776 40776 31804
rect 40770 31764 40776 31776
rect 40828 31764 40834 31816
rect 41138 31804 41144 31816
rect 41099 31776 41144 31804
rect 41138 31764 41144 31776
rect 41196 31764 41202 31816
rect 42383 31807 42441 31813
rect 42383 31773 42395 31807
rect 42429 31804 42441 31807
rect 42610 31804 42616 31816
rect 42429 31776 42616 31804
rect 42429 31773 42441 31776
rect 42383 31767 42441 31773
rect 42610 31764 42616 31776
rect 42668 31804 42674 31816
rect 43533 31807 43591 31813
rect 43533 31804 43545 31807
rect 42668 31776 43545 31804
rect 42668 31764 42674 31776
rect 43533 31773 43545 31776
rect 43579 31773 43591 31807
rect 44174 31804 44180 31816
rect 44087 31776 44180 31804
rect 43533 31767 43591 31773
rect 44174 31764 44180 31776
rect 44232 31804 44238 31816
rect 45278 31804 45284 31816
rect 44232 31776 45284 31804
rect 44232 31764 44238 31776
rect 45278 31764 45284 31776
rect 45336 31764 45342 31816
rect 35342 31736 35348 31748
rect 30423 31708 35348 31736
rect 30423 31705 30435 31708
rect 30377 31699 30435 31705
rect 35342 31696 35348 31708
rect 35400 31696 35406 31748
rect 44082 31696 44088 31748
rect 44140 31736 44146 31748
rect 44453 31739 44511 31745
rect 44453 31736 44465 31739
rect 44140 31708 44465 31736
rect 44140 31696 44146 31708
rect 44453 31705 44465 31708
rect 44499 31705 44511 31739
rect 44453 31699 44511 31705
rect 27847 31671 27905 31677
rect 27847 31668 27859 31671
rect 27540 31640 27859 31668
rect 26651 31631 26709 31637
rect 27847 31637 27859 31640
rect 27893 31637 27905 31671
rect 27982 31668 27988 31680
rect 27943 31640 27988 31668
rect 27847 31631 27905 31637
rect 27982 31628 27988 31640
rect 28040 31628 28046 31680
rect 29270 31668 29276 31680
rect 29231 31640 29276 31668
rect 29270 31628 29276 31640
rect 29328 31628 29334 31680
rect 32858 31628 32864 31680
rect 32916 31668 32922 31680
rect 33045 31671 33103 31677
rect 33045 31668 33057 31671
rect 32916 31640 33057 31668
rect 32916 31628 32922 31640
rect 33045 31637 33057 31640
rect 33091 31637 33103 31671
rect 33045 31631 33103 31637
rect 34790 31628 34796 31680
rect 34848 31668 34854 31680
rect 35437 31671 35495 31677
rect 35437 31668 35449 31671
rect 34848 31640 35449 31668
rect 34848 31628 34854 31640
rect 35437 31637 35449 31640
rect 35483 31637 35495 31671
rect 35437 31631 35495 31637
rect 41138 31628 41144 31680
rect 41196 31668 41202 31680
rect 44266 31668 44272 31680
rect 41196 31640 44272 31668
rect 41196 31628 41202 31640
rect 44266 31628 44272 31640
rect 44324 31628 44330 31680
rect 1104 31578 48852 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 48852 31578
rect 1104 31504 48852 31526
rect 11471 31467 11529 31473
rect 11471 31433 11483 31467
rect 11517 31464 11529 31467
rect 12986 31464 12992 31476
rect 11517 31436 12992 31464
rect 11517 31433 11529 31436
rect 11471 31427 11529 31433
rect 12986 31424 12992 31436
rect 13044 31424 13050 31476
rect 13446 31464 13452 31476
rect 13407 31436 13452 31464
rect 13446 31424 13452 31436
rect 13504 31424 13510 31476
rect 13814 31424 13820 31476
rect 13872 31464 13878 31476
rect 15381 31467 15439 31473
rect 13872 31436 13917 31464
rect 13872 31424 13878 31436
rect 15381 31433 15393 31467
rect 15427 31464 15439 31467
rect 15470 31464 15476 31476
rect 15427 31436 15476 31464
rect 15427 31433 15439 31436
rect 15381 31427 15439 31433
rect 15470 31424 15476 31436
rect 15528 31424 15534 31476
rect 17218 31424 17224 31476
rect 17276 31464 17282 31476
rect 17405 31467 17463 31473
rect 17405 31464 17417 31467
rect 17276 31436 17417 31464
rect 17276 31424 17282 31436
rect 17405 31433 17417 31436
rect 17451 31433 17463 31467
rect 17405 31427 17463 31433
rect 19150 31424 19156 31476
rect 19208 31464 19214 31476
rect 19981 31467 20039 31473
rect 19981 31464 19993 31467
rect 19208 31436 19993 31464
rect 19208 31424 19214 31436
rect 19981 31433 19993 31436
rect 20027 31433 20039 31467
rect 19981 31427 20039 31433
rect 21637 31467 21695 31473
rect 21637 31433 21649 31467
rect 21683 31464 21695 31467
rect 21726 31464 21732 31476
rect 21683 31436 21732 31464
rect 21683 31433 21695 31436
rect 21637 31427 21695 31433
rect 21726 31424 21732 31436
rect 21784 31424 21790 31476
rect 23017 31467 23075 31473
rect 23017 31433 23029 31467
rect 23063 31464 23075 31467
rect 23474 31464 23480 31476
rect 23063 31436 23480 31464
rect 23063 31433 23075 31436
rect 23017 31427 23075 31433
rect 23474 31424 23480 31436
rect 23532 31424 23538 31476
rect 26418 31424 26424 31476
rect 26476 31464 26482 31476
rect 26605 31467 26663 31473
rect 26605 31464 26617 31467
rect 26476 31436 26617 31464
rect 26476 31424 26482 31436
rect 26605 31433 26617 31436
rect 26651 31433 26663 31467
rect 26605 31427 26663 31433
rect 30006 31424 30012 31476
rect 30064 31464 30070 31476
rect 30193 31467 30251 31473
rect 30193 31464 30205 31467
rect 30064 31436 30205 31464
rect 30064 31424 30070 31436
rect 30193 31433 30205 31436
rect 30239 31464 30251 31467
rect 30469 31467 30527 31473
rect 30469 31464 30481 31467
rect 30239 31436 30481 31464
rect 30239 31433 30251 31436
rect 30193 31427 30251 31433
rect 30469 31433 30481 31436
rect 30515 31433 30527 31467
rect 30469 31427 30527 31433
rect 31159 31467 31217 31473
rect 31159 31433 31171 31467
rect 31205 31464 31217 31467
rect 31570 31464 31576 31476
rect 31205 31436 31576 31464
rect 31205 31433 31217 31436
rect 31159 31427 31217 31433
rect 31570 31424 31576 31436
rect 31628 31424 31634 31476
rect 32858 31424 32864 31476
rect 32916 31464 32922 31476
rect 34241 31467 34299 31473
rect 34241 31464 34253 31467
rect 32916 31436 34253 31464
rect 32916 31424 32922 31436
rect 34241 31433 34253 31436
rect 34287 31464 34299 31467
rect 34514 31464 34520 31476
rect 34287 31436 34520 31464
rect 34287 31433 34299 31436
rect 34241 31427 34299 31433
rect 34514 31424 34520 31436
rect 34572 31424 34578 31476
rect 35894 31424 35900 31476
rect 35952 31464 35958 31476
rect 36633 31467 36691 31473
rect 36633 31464 36645 31467
rect 35952 31436 36645 31464
rect 35952 31424 35958 31436
rect 36633 31433 36645 31436
rect 36679 31433 36691 31467
rect 36633 31427 36691 31433
rect 38013 31467 38071 31473
rect 38013 31433 38025 31467
rect 38059 31464 38071 31467
rect 38102 31464 38108 31476
rect 38059 31436 38108 31464
rect 38059 31433 38071 31436
rect 38013 31427 38071 31433
rect 13630 31396 13636 31408
rect 11716 31368 13636 31396
rect 11400 31263 11458 31269
rect 11400 31229 11412 31263
rect 11446 31260 11458 31263
rect 11716 31260 11744 31368
rect 13630 31356 13636 31368
rect 13688 31356 13694 31408
rect 16114 31356 16120 31408
rect 16172 31396 16178 31408
rect 17773 31399 17831 31405
rect 17773 31396 17785 31399
rect 16172 31368 17785 31396
rect 16172 31356 16178 31368
rect 17773 31365 17785 31368
rect 17819 31365 17831 31399
rect 17773 31359 17831 31365
rect 12526 31328 12532 31340
rect 12439 31300 12532 31328
rect 12526 31288 12532 31300
rect 12584 31328 12590 31340
rect 13170 31328 13176 31340
rect 12584 31300 13176 31328
rect 12584 31288 12590 31300
rect 13170 31288 13176 31300
rect 13228 31288 13234 31340
rect 14599 31331 14657 31337
rect 14599 31297 14611 31331
rect 14645 31328 14657 31331
rect 15378 31328 15384 31340
rect 14645 31300 15384 31328
rect 14645 31297 14657 31300
rect 14599 31291 14657 31297
rect 15378 31288 15384 31300
rect 15436 31328 15442 31340
rect 15657 31331 15715 31337
rect 15657 31328 15669 31331
rect 15436 31300 15669 31328
rect 15436 31288 15442 31300
rect 15657 31297 15669 31300
rect 15703 31297 15715 31331
rect 17034 31328 17040 31340
rect 16995 31300 17040 31328
rect 15657 31291 15715 31297
rect 17034 31288 17040 31300
rect 17092 31288 17098 31340
rect 17788 31328 17816 31359
rect 19610 31356 19616 31408
rect 19668 31356 19674 31408
rect 19794 31396 19800 31408
rect 19755 31368 19800 31396
rect 19794 31356 19800 31368
rect 19852 31356 19858 31408
rect 20806 31396 20812 31408
rect 20767 31368 20812 31396
rect 20806 31356 20812 31368
rect 20864 31356 20870 31408
rect 20990 31356 20996 31408
rect 21048 31396 21054 31408
rect 22557 31399 22615 31405
rect 22557 31396 22569 31399
rect 21048 31368 22569 31396
rect 21048 31356 21054 31368
rect 22557 31365 22569 31368
rect 22603 31396 22615 31399
rect 22646 31396 22652 31408
rect 22603 31368 22652 31396
rect 22603 31365 22615 31368
rect 22557 31359 22615 31365
rect 22646 31356 22652 31368
rect 22704 31356 22710 31408
rect 27430 31396 27436 31408
rect 23860 31368 27436 31396
rect 18969 31331 19027 31337
rect 18969 31328 18981 31331
rect 17788 31300 18981 31328
rect 11446 31232 11744 31260
rect 11446 31229 11458 31232
rect 11400 31223 11458 31229
rect 11716 31136 11744 31232
rect 14512 31263 14570 31269
rect 14512 31229 14524 31263
rect 14558 31260 14570 31263
rect 15286 31260 15292 31272
rect 14558 31232 15292 31260
rect 14558 31229 14570 31232
rect 14512 31223 14570 31229
rect 12621 31195 12679 31201
rect 12621 31161 12633 31195
rect 12667 31192 12679 31195
rect 12802 31192 12808 31204
rect 12667 31164 12808 31192
rect 12667 31161 12679 31164
rect 12621 31155 12679 31161
rect 12802 31152 12808 31164
rect 12860 31152 12866 31204
rect 12894 31152 12900 31204
rect 12952 31192 12958 31204
rect 13173 31195 13231 31201
rect 13173 31192 13185 31195
rect 12952 31164 13185 31192
rect 12952 31152 12958 31164
rect 13173 31161 13185 31164
rect 13219 31161 13231 31195
rect 13173 31155 13231 31161
rect 14936 31136 14964 31232
rect 15286 31220 15292 31232
rect 15344 31220 15350 31272
rect 16393 31263 16451 31269
rect 16393 31229 16405 31263
rect 16439 31229 16451 31263
rect 16393 31223 16451 31229
rect 16301 31195 16359 31201
rect 16301 31161 16313 31195
rect 16347 31192 16359 31195
rect 16408 31192 16436 31223
rect 16482 31220 16488 31272
rect 16540 31260 16546 31272
rect 16853 31263 16911 31269
rect 16853 31260 16865 31263
rect 16540 31232 16865 31260
rect 16540 31220 16546 31232
rect 16853 31229 16865 31232
rect 16899 31229 16911 31263
rect 16853 31223 16911 31229
rect 18141 31263 18199 31269
rect 18141 31229 18153 31263
rect 18187 31260 18199 31263
rect 18230 31260 18236 31272
rect 18187 31232 18236 31260
rect 18187 31229 18199 31232
rect 18141 31223 18199 31229
rect 18230 31220 18236 31232
rect 18288 31220 18294 31272
rect 18340 31269 18368 31300
rect 18969 31297 18981 31300
rect 19015 31328 19027 31331
rect 19337 31331 19395 31337
rect 19337 31328 19349 31331
rect 19015 31300 19349 31328
rect 19015 31297 19027 31300
rect 18969 31291 19027 31297
rect 19337 31297 19349 31300
rect 19383 31328 19395 31331
rect 19628 31328 19656 31356
rect 19889 31331 19947 31337
rect 19889 31328 19901 31331
rect 19383 31300 19901 31328
rect 19383 31297 19395 31300
rect 19337 31291 19395 31297
rect 19889 31297 19901 31300
rect 19935 31297 19947 31331
rect 19889 31291 19947 31297
rect 18325 31263 18383 31269
rect 18325 31229 18337 31263
rect 18371 31229 18383 31263
rect 18325 31223 18383 31229
rect 19426 31220 19432 31272
rect 19484 31260 19490 31272
rect 19668 31263 19726 31269
rect 19668 31260 19680 31263
rect 19484 31232 19680 31260
rect 19484 31220 19490 31232
rect 19668 31229 19680 31232
rect 19714 31260 19726 31263
rect 20438 31260 20444 31272
rect 19714 31232 20444 31260
rect 19714 31229 19726 31232
rect 19668 31223 19726 31229
rect 20438 31220 20444 31232
rect 20496 31220 20502 31272
rect 20898 31220 20904 31272
rect 20956 31260 20962 31272
rect 23860 31269 23888 31368
rect 27430 31356 27436 31368
rect 27488 31356 27494 31408
rect 34532 31396 34560 31424
rect 35989 31399 36047 31405
rect 35989 31396 36001 31399
rect 34532 31368 36001 31396
rect 35989 31365 36001 31368
rect 36035 31396 36047 31399
rect 36170 31396 36176 31408
rect 36035 31368 36176 31396
rect 36035 31365 36047 31368
rect 35989 31359 36047 31365
rect 36170 31356 36176 31368
rect 36228 31356 36234 31408
rect 25317 31331 25375 31337
rect 25317 31297 25329 31331
rect 25363 31328 25375 31331
rect 25774 31328 25780 31340
rect 25363 31300 25780 31328
rect 25363 31297 25375 31300
rect 25317 31291 25375 31297
rect 25774 31288 25780 31300
rect 25832 31288 25838 31340
rect 27982 31328 27988 31340
rect 27632 31300 27988 31328
rect 21545 31263 21603 31269
rect 21545 31260 21557 31263
rect 20956 31232 21557 31260
rect 20956 31220 20962 31232
rect 21545 31229 21557 31232
rect 21591 31260 21603 31263
rect 22189 31263 22247 31269
rect 22189 31260 22201 31263
rect 21591 31232 22201 31260
rect 21591 31229 21603 31232
rect 21545 31223 21603 31229
rect 22189 31229 22201 31232
rect 22235 31229 22247 31263
rect 22189 31223 22247 31229
rect 23477 31263 23535 31269
rect 23477 31229 23489 31263
rect 23523 31260 23535 31263
rect 23845 31263 23903 31269
rect 23845 31260 23857 31263
rect 23523 31232 23857 31260
rect 23523 31229 23535 31232
rect 23477 31223 23535 31229
rect 23845 31229 23857 31232
rect 23891 31229 23903 31263
rect 24946 31260 24952 31272
rect 24907 31232 24952 31260
rect 23845 31223 23903 31229
rect 24946 31220 24952 31232
rect 25004 31220 25010 31272
rect 27632 31204 27660 31300
rect 27982 31288 27988 31300
rect 28040 31288 28046 31340
rect 28353 31331 28411 31337
rect 28353 31297 28365 31331
rect 28399 31328 28411 31331
rect 29270 31328 29276 31340
rect 28399 31300 29276 31328
rect 28399 31297 28411 31300
rect 28353 31291 28411 31297
rect 29270 31288 29276 31300
rect 29328 31288 29334 31340
rect 32125 31331 32183 31337
rect 32125 31297 32137 31331
rect 32171 31328 32183 31331
rect 32214 31328 32220 31340
rect 32171 31300 32220 31328
rect 32171 31297 32183 31300
rect 32125 31291 32183 31297
rect 32214 31288 32220 31300
rect 32272 31288 32278 31340
rect 34238 31288 34244 31340
rect 34296 31328 34302 31340
rect 35158 31328 35164 31340
rect 34296 31300 35164 31328
rect 34296 31288 34302 31300
rect 35158 31288 35164 31300
rect 35216 31288 35222 31340
rect 35434 31328 35440 31340
rect 35395 31300 35440 31328
rect 35434 31288 35440 31300
rect 35492 31288 35498 31340
rect 27893 31263 27951 31269
rect 27893 31229 27905 31263
rect 27939 31229 27951 31263
rect 28166 31260 28172 31272
rect 28079 31232 28172 31260
rect 27893 31223 27951 31229
rect 17402 31192 17408 31204
rect 16347 31164 17408 31192
rect 16347 31161 16359 31164
rect 16301 31155 16359 31161
rect 17402 31152 17408 31164
rect 17460 31192 17466 31204
rect 17862 31192 17868 31204
rect 17460 31164 17868 31192
rect 17460 31152 17466 31164
rect 17862 31152 17868 31164
rect 17920 31152 17926 31204
rect 18693 31195 18751 31201
rect 18693 31161 18705 31195
rect 18739 31192 18751 31195
rect 19150 31192 19156 31204
rect 18739 31164 19156 31192
rect 18739 31161 18751 31164
rect 18693 31155 18751 31161
rect 19150 31152 19156 31164
rect 19208 31152 19214 31204
rect 19521 31195 19579 31201
rect 19521 31161 19533 31195
rect 19567 31192 19579 31195
rect 20346 31192 20352 31204
rect 19567 31164 20352 31192
rect 19567 31161 19579 31164
rect 19521 31155 19579 31161
rect 20346 31152 20352 31164
rect 20404 31152 20410 31204
rect 21269 31195 21327 31201
rect 21269 31161 21281 31195
rect 21315 31192 21327 31195
rect 21361 31195 21419 31201
rect 21361 31192 21373 31195
rect 21315 31164 21373 31192
rect 21315 31161 21327 31164
rect 21269 31155 21327 31161
rect 21361 31161 21373 31164
rect 21407 31192 21419 31195
rect 23661 31195 23719 31201
rect 23661 31192 23673 31195
rect 21407 31164 23673 31192
rect 21407 31161 21419 31164
rect 21361 31155 21419 31161
rect 23661 31161 23673 31164
rect 23707 31192 23719 31195
rect 24581 31195 24639 31201
rect 24581 31192 24593 31195
rect 23707 31164 24593 31192
rect 23707 31161 23719 31164
rect 23661 31155 23719 31161
rect 24581 31161 24593 31164
rect 24627 31192 24639 31195
rect 25406 31192 25412 31204
rect 24627 31164 25268 31192
rect 25367 31164 25412 31192
rect 24627 31161 24639 31164
rect 24581 31155 24639 31161
rect 10410 31124 10416 31136
rect 10371 31096 10416 31124
rect 10410 31084 10416 31096
rect 10468 31084 10474 31136
rect 10686 31084 10692 31136
rect 10744 31124 10750 31136
rect 10781 31127 10839 31133
rect 10781 31124 10793 31127
rect 10744 31096 10793 31124
rect 10744 31084 10750 31096
rect 10781 31093 10793 31096
rect 10827 31093 10839 31127
rect 10781 31087 10839 31093
rect 11698 31084 11704 31136
rect 11756 31124 11762 31136
rect 11793 31127 11851 31133
rect 11793 31124 11805 31127
rect 11756 31096 11805 31124
rect 11756 31084 11762 31096
rect 11793 31093 11805 31096
rect 11839 31093 11851 31127
rect 11793 31087 11851 31093
rect 12253 31127 12311 31133
rect 12253 31093 12265 31127
rect 12299 31124 12311 31127
rect 12342 31124 12348 31136
rect 12299 31096 12348 31124
rect 12299 31093 12311 31096
rect 12253 31087 12311 31093
rect 12342 31084 12348 31096
rect 12400 31124 12406 31136
rect 13078 31124 13084 31136
rect 12400 31096 13084 31124
rect 12400 31084 12406 31096
rect 13078 31084 13084 31096
rect 13136 31084 13142 31136
rect 14918 31124 14924 31136
rect 14879 31096 14924 31124
rect 14918 31084 14924 31096
rect 14976 31084 14982 31136
rect 18966 31084 18972 31136
rect 19024 31124 19030 31136
rect 22278 31124 22284 31136
rect 19024 31096 22284 31124
rect 19024 31084 19030 31096
rect 22278 31084 22284 31096
rect 22336 31084 22342 31136
rect 23934 31124 23940 31136
rect 23895 31096 23940 31124
rect 23934 31084 23940 31096
rect 23992 31084 23998 31136
rect 25240 31124 25268 31164
rect 25406 31152 25412 31164
rect 25464 31152 25470 31204
rect 25958 31192 25964 31204
rect 25919 31164 25964 31192
rect 25958 31152 25964 31164
rect 26016 31152 26022 31204
rect 27157 31195 27215 31201
rect 27157 31161 27169 31195
rect 27203 31192 27215 31195
rect 27614 31192 27620 31204
rect 27203 31164 27620 31192
rect 27203 31161 27215 31164
rect 27157 31155 27215 31161
rect 27614 31152 27620 31164
rect 27672 31152 27678 31204
rect 27908 31192 27936 31223
rect 28166 31220 28172 31232
rect 28224 31260 28230 31272
rect 28626 31260 28632 31272
rect 28224 31232 28632 31260
rect 28224 31220 28230 31232
rect 28626 31220 28632 31232
rect 28684 31220 28690 31272
rect 30926 31260 30932 31272
rect 30887 31232 30932 31260
rect 30926 31220 30932 31232
rect 30984 31260 30990 31272
rect 31056 31263 31114 31269
rect 31056 31260 31068 31263
rect 30984 31232 31068 31260
rect 30984 31220 30990 31232
rect 31056 31229 31068 31232
rect 31102 31229 31114 31263
rect 36648 31260 36676 31427
rect 38102 31424 38108 31436
rect 38160 31424 38166 31476
rect 40310 31464 40316 31476
rect 40271 31436 40316 31464
rect 40310 31424 40316 31436
rect 40368 31424 40374 31476
rect 41046 31424 41052 31476
rect 41104 31464 41110 31476
rect 41647 31467 41705 31473
rect 41647 31464 41659 31467
rect 41104 31436 41659 31464
rect 41104 31424 41110 31436
rect 41647 31433 41659 31436
rect 41693 31433 41705 31467
rect 42610 31464 42616 31476
rect 42571 31436 42616 31464
rect 41647 31427 41705 31433
rect 42610 31424 42616 31436
rect 42668 31424 42674 31476
rect 43073 31467 43131 31473
rect 43073 31433 43085 31467
rect 43119 31464 43131 31467
rect 43441 31467 43499 31473
rect 43441 31464 43453 31467
rect 43119 31436 43453 31464
rect 43119 31433 43131 31436
rect 43073 31427 43131 31433
rect 43441 31433 43453 31436
rect 43487 31464 43499 31467
rect 43714 31464 43720 31476
rect 43487 31436 43720 31464
rect 43487 31433 43499 31436
rect 43441 31427 43499 31433
rect 43714 31424 43720 31436
rect 43772 31464 43778 31476
rect 44082 31464 44088 31476
rect 43772 31436 44088 31464
rect 43772 31424 43778 31436
rect 44082 31424 44088 31436
rect 44140 31424 44146 31476
rect 40586 31356 40592 31408
rect 40644 31396 40650 31408
rect 40862 31396 40868 31408
rect 40644 31368 40868 31396
rect 40644 31356 40650 31368
rect 40862 31356 40868 31368
rect 40920 31356 40926 31408
rect 42978 31356 42984 31408
rect 43036 31396 43042 31408
rect 44177 31399 44235 31405
rect 44177 31396 44189 31399
rect 43036 31368 44189 31396
rect 43036 31356 43042 31368
rect 44177 31365 44189 31368
rect 44223 31365 44235 31399
rect 44177 31359 44235 31365
rect 37366 31328 37372 31340
rect 37327 31300 37372 31328
rect 37366 31288 37372 31300
rect 37424 31288 37430 31340
rect 43622 31328 43628 31340
rect 38304 31300 39344 31328
rect 43583 31300 43628 31328
rect 36817 31263 36875 31269
rect 36817 31260 36829 31263
rect 36648 31232 36829 31260
rect 31056 31223 31114 31229
rect 36817 31229 36829 31232
rect 36863 31229 36875 31263
rect 36817 31223 36875 31229
rect 36906 31220 36912 31272
rect 36964 31260 36970 31272
rect 38304 31269 38332 31300
rect 39316 31269 39344 31300
rect 43622 31288 43628 31300
rect 43680 31328 43686 31340
rect 44545 31331 44603 31337
rect 44545 31328 44557 31331
rect 43680 31300 44557 31328
rect 43680 31288 43686 31300
rect 44545 31297 44557 31300
rect 44591 31297 44603 31331
rect 44545 31291 44603 31297
rect 37277 31263 37335 31269
rect 37277 31260 37289 31263
rect 36964 31232 37289 31260
rect 36964 31220 36970 31232
rect 37277 31229 37289 31232
rect 37323 31260 37335 31263
rect 38289 31263 38347 31269
rect 38289 31260 38301 31263
rect 37323 31232 38301 31260
rect 37323 31229 37335 31232
rect 37277 31223 37335 31229
rect 38289 31229 38301 31232
rect 38335 31229 38347 31263
rect 38289 31223 38347 31229
rect 38841 31263 38899 31269
rect 38841 31229 38853 31263
rect 38887 31229 38899 31263
rect 38841 31223 38899 31229
rect 39301 31263 39359 31269
rect 39301 31229 39313 31263
rect 39347 31229 39359 31263
rect 39942 31260 39948 31272
rect 39301 31223 39359 31229
rect 39408 31232 39948 31260
rect 32490 31201 32496 31204
rect 29635 31195 29693 31201
rect 27908 31164 28764 31192
rect 28736 31136 28764 31164
rect 29635 31161 29647 31195
rect 29681 31161 29693 31195
rect 32446 31195 32496 31201
rect 32446 31192 32458 31195
rect 29635 31155 29693 31161
rect 31956 31164 32458 31192
rect 26234 31124 26240 31136
rect 25240 31096 26240 31124
rect 26234 31084 26240 31096
rect 26292 31084 26298 31136
rect 27525 31127 27583 31133
rect 27525 31093 27537 31127
rect 27571 31124 27583 31127
rect 27706 31124 27712 31136
rect 27571 31096 27712 31124
rect 27571 31093 27583 31096
rect 27525 31087 27583 31093
rect 27706 31084 27712 31096
rect 27764 31084 27770 31136
rect 28718 31124 28724 31136
rect 28679 31096 28724 31124
rect 28718 31084 28724 31096
rect 28776 31084 28782 31136
rect 28994 31124 29000 31136
rect 28955 31096 29000 31124
rect 28994 31084 29000 31096
rect 29052 31124 29058 31136
rect 29650 31124 29678 31155
rect 30374 31124 30380 31136
rect 29052 31096 30380 31124
rect 29052 31084 29058 31096
rect 30374 31084 30380 31096
rect 30432 31124 30438 31136
rect 31956 31133 31984 31164
rect 32446 31161 32458 31164
rect 32492 31161 32496 31195
rect 32446 31155 32496 31161
rect 32490 31152 32496 31155
rect 32548 31152 32554 31204
rect 34609 31195 34667 31201
rect 34609 31192 34621 31195
rect 33428 31164 34621 31192
rect 33428 31136 33456 31164
rect 34609 31161 34621 31164
rect 34655 31192 34667 31195
rect 34698 31192 34704 31204
rect 34655 31164 34704 31192
rect 34655 31161 34667 31164
rect 34609 31155 34667 31161
rect 34698 31152 34704 31164
rect 34756 31152 34762 31204
rect 34790 31152 34796 31204
rect 34848 31192 34854 31204
rect 34977 31195 35035 31201
rect 34977 31192 34989 31195
rect 34848 31164 34989 31192
rect 34848 31152 34854 31164
rect 34977 31161 34989 31164
rect 35023 31161 35035 31195
rect 34977 31155 35035 31161
rect 35069 31195 35127 31201
rect 35069 31161 35081 31195
rect 35115 31161 35127 31195
rect 35069 31155 35127 31161
rect 31573 31127 31631 31133
rect 31573 31124 31585 31127
rect 30432 31096 31585 31124
rect 30432 31084 30438 31096
rect 31573 31093 31585 31096
rect 31619 31124 31631 31127
rect 31941 31127 31999 31133
rect 31941 31124 31953 31127
rect 31619 31096 31953 31124
rect 31619 31093 31631 31096
rect 31573 31087 31631 31093
rect 31941 31093 31953 31096
rect 31987 31093 31999 31127
rect 31941 31087 31999 31093
rect 33045 31127 33103 31133
rect 33045 31093 33057 31127
rect 33091 31124 33103 31127
rect 33410 31124 33416 31136
rect 33091 31096 33416 31124
rect 33091 31093 33103 31096
rect 33045 31087 33103 31093
rect 33410 31084 33416 31096
rect 33468 31084 33474 31136
rect 33962 31124 33968 31136
rect 33923 31096 33968 31124
rect 33962 31084 33968 31096
rect 34020 31084 34026 31136
rect 34716 31124 34744 31152
rect 35084 31124 35112 31155
rect 35158 31152 35164 31204
rect 35216 31192 35222 31204
rect 38657 31195 38715 31201
rect 38657 31192 38669 31195
rect 35216 31164 38669 31192
rect 35216 31152 35222 31164
rect 38657 31161 38669 31164
rect 38703 31192 38715 31195
rect 38856 31192 38884 31223
rect 38703 31164 38884 31192
rect 38703 31161 38715 31164
rect 38657 31155 38715 31161
rect 34716 31096 35112 31124
rect 35526 31084 35532 31136
rect 35584 31124 35590 31136
rect 39408 31124 39436 31232
rect 39942 31220 39948 31232
rect 40000 31260 40006 31272
rect 40310 31260 40316 31272
rect 40000 31232 40316 31260
rect 40000 31220 40006 31232
rect 40310 31220 40316 31232
rect 40368 31260 40374 31272
rect 40532 31263 40590 31269
rect 40532 31260 40544 31263
rect 40368 31232 40544 31260
rect 40368 31220 40374 31232
rect 40532 31229 40544 31232
rect 40578 31260 40590 31263
rect 40957 31263 41015 31269
rect 40957 31260 40969 31263
rect 40578 31232 40969 31260
rect 40578 31229 40590 31232
rect 40532 31223 40590 31229
rect 40957 31229 40969 31232
rect 41003 31229 41015 31263
rect 41544 31263 41602 31269
rect 41544 31260 41556 31263
rect 40957 31223 41015 31229
rect 41340 31232 41556 31260
rect 39574 31192 39580 31204
rect 39535 31164 39580 31192
rect 39574 31152 39580 31164
rect 39632 31152 39638 31204
rect 40635 31195 40693 31201
rect 40635 31161 40647 31195
rect 40681 31192 40693 31195
rect 40770 31192 40776 31204
rect 40681 31164 40776 31192
rect 40681 31161 40693 31164
rect 40635 31155 40693 31161
rect 40770 31152 40776 31164
rect 40828 31192 40834 31204
rect 41230 31192 41236 31204
rect 40828 31164 41236 31192
rect 40828 31152 40834 31164
rect 41230 31152 41236 31164
rect 41288 31152 41294 31204
rect 39850 31124 39856 31136
rect 35584 31096 39436 31124
rect 39811 31096 39856 31124
rect 35584 31084 35590 31096
rect 39850 31084 39856 31096
rect 39908 31084 39914 31136
rect 40862 31084 40868 31136
rect 40920 31124 40926 31136
rect 41340 31133 41368 31232
rect 41544 31229 41556 31232
rect 41590 31229 41602 31263
rect 41544 31223 41602 31229
rect 44726 31220 44732 31272
rect 44784 31260 44790 31272
rect 45094 31260 45100 31272
rect 44784 31232 45100 31260
rect 44784 31220 44790 31232
rect 45094 31220 45100 31232
rect 45152 31220 45158 31272
rect 43714 31192 43720 31204
rect 43675 31164 43720 31192
rect 43714 31152 43720 31164
rect 43772 31152 43778 31204
rect 41325 31127 41383 31133
rect 41325 31124 41337 31127
rect 40920 31096 41337 31124
rect 40920 31084 40926 31096
rect 41325 31093 41337 31096
rect 41371 31093 41383 31127
rect 42334 31124 42340 31136
rect 42295 31096 42340 31124
rect 41325 31087 41383 31093
rect 42334 31084 42340 31096
rect 42392 31084 42398 31136
rect 1104 31034 48852 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 48852 31034
rect 1104 30960 48852 30982
rect 13722 30920 13728 30932
rect 13683 30892 13728 30920
rect 13722 30880 13728 30892
rect 13780 30920 13786 30932
rect 13780 30892 16068 30920
rect 13780 30880 13786 30892
rect 11974 30852 11980 30864
rect 11935 30824 11980 30852
rect 11974 30812 11980 30824
rect 12032 30812 12038 30864
rect 12526 30852 12532 30864
rect 12487 30824 12532 30852
rect 12526 30812 12532 30824
rect 12584 30812 12590 30864
rect 15470 30852 15476 30864
rect 15431 30824 15476 30852
rect 15470 30812 15476 30824
rect 15528 30812 15534 30864
rect 16040 30861 16068 30892
rect 16942 30880 16948 30932
rect 17000 30920 17006 30932
rect 17037 30923 17095 30929
rect 17037 30920 17049 30923
rect 17000 30892 17049 30920
rect 17000 30880 17006 30892
rect 17037 30889 17049 30892
rect 17083 30889 17095 30923
rect 17037 30883 17095 30889
rect 18138 30880 18144 30932
rect 18196 30920 18202 30932
rect 18417 30923 18475 30929
rect 18417 30920 18429 30923
rect 18196 30892 18429 30920
rect 18196 30880 18202 30892
rect 18417 30889 18429 30892
rect 18463 30889 18475 30923
rect 19058 30920 19064 30932
rect 19019 30892 19064 30920
rect 18417 30883 18475 30889
rect 19058 30880 19064 30892
rect 19116 30880 19122 30932
rect 20438 30920 20444 30932
rect 20351 30892 20444 30920
rect 20438 30880 20444 30892
rect 20496 30920 20502 30932
rect 23934 30920 23940 30932
rect 20496 30892 23940 30920
rect 20496 30880 20502 30892
rect 23934 30880 23940 30892
rect 23992 30880 23998 30932
rect 24486 30920 24492 30932
rect 24447 30892 24492 30920
rect 24486 30880 24492 30892
rect 24544 30880 24550 30932
rect 28258 30880 28264 30932
rect 28316 30920 28322 30932
rect 28445 30923 28503 30929
rect 28445 30920 28457 30923
rect 28316 30892 28457 30920
rect 28316 30880 28322 30892
rect 28445 30889 28457 30892
rect 28491 30889 28503 30923
rect 28445 30883 28503 30889
rect 30006 30880 30012 30932
rect 30064 30920 30070 30932
rect 30064 30892 30236 30920
rect 30064 30880 30070 30892
rect 16025 30855 16083 30861
rect 16025 30821 16037 30855
rect 16071 30852 16083 30855
rect 17126 30852 17132 30864
rect 16071 30824 17132 30852
rect 16071 30821 16083 30824
rect 16025 30815 16083 30821
rect 17126 30812 17132 30824
rect 17184 30812 17190 30864
rect 17586 30852 17592 30864
rect 17547 30824 17592 30852
rect 17586 30812 17592 30824
rect 17644 30812 17650 30864
rect 18877 30855 18935 30861
rect 18877 30821 18889 30855
rect 18923 30852 18935 30855
rect 20456 30852 20484 30880
rect 22922 30852 22928 30864
rect 18923 30824 20484 30852
rect 22883 30824 22928 30852
rect 18923 30821 18935 30824
rect 18877 30815 18935 30821
rect 22922 30812 22928 30824
rect 22980 30812 22986 30864
rect 24857 30855 24915 30861
rect 24857 30821 24869 30855
rect 24903 30852 24915 30855
rect 24946 30852 24952 30864
rect 24903 30824 24952 30852
rect 24903 30821 24915 30824
rect 24857 30815 24915 30821
rect 24946 30812 24952 30824
rect 25004 30812 25010 30864
rect 25409 30855 25467 30861
rect 25409 30821 25421 30855
rect 25455 30852 25467 30855
rect 25958 30852 25964 30864
rect 25455 30824 25964 30852
rect 25455 30821 25467 30824
rect 25409 30815 25467 30821
rect 25958 30812 25964 30824
rect 26016 30812 26022 30864
rect 30208 30861 30236 30892
rect 32214 30880 32220 30932
rect 32272 30920 32278 30932
rect 32309 30923 32367 30929
rect 32309 30920 32321 30923
rect 32272 30892 32321 30920
rect 32272 30880 32278 30892
rect 32309 30889 32321 30892
rect 32355 30889 32367 30923
rect 32674 30920 32680 30932
rect 32635 30892 32680 30920
rect 32309 30883 32367 30889
rect 32674 30880 32680 30892
rect 32732 30880 32738 30932
rect 32858 30880 32864 30932
rect 32916 30920 32922 30932
rect 32916 30892 33180 30920
rect 32916 30880 32922 30892
rect 30193 30855 30251 30861
rect 30193 30821 30205 30855
rect 30239 30852 30251 30855
rect 30466 30852 30472 30864
rect 30239 30824 30472 30852
rect 30239 30821 30251 30824
rect 30193 30815 30251 30821
rect 30466 30812 30472 30824
rect 30524 30812 30530 30864
rect 33042 30852 33048 30864
rect 33003 30824 33048 30852
rect 33042 30812 33048 30824
rect 33100 30812 33106 30864
rect 33152 30861 33180 30892
rect 33318 30880 33324 30932
rect 33376 30920 33382 30932
rect 36219 30923 36277 30929
rect 36219 30920 36231 30923
rect 33376 30892 36231 30920
rect 33376 30880 33382 30892
rect 36219 30889 36231 30892
rect 36265 30889 36277 30923
rect 36219 30883 36277 30889
rect 37734 30880 37740 30932
rect 37792 30920 37798 30932
rect 37921 30923 37979 30929
rect 37921 30920 37933 30923
rect 37792 30892 37933 30920
rect 37792 30880 37798 30892
rect 37921 30889 37933 30892
rect 37967 30889 37979 30923
rect 41230 30920 41236 30932
rect 41191 30892 41236 30920
rect 37921 30883 37979 30889
rect 41230 30880 41236 30892
rect 41288 30880 41294 30932
rect 41690 30920 41696 30932
rect 41651 30892 41696 30920
rect 41690 30880 41696 30892
rect 41748 30880 41754 30932
rect 42383 30923 42441 30929
rect 42383 30889 42395 30923
rect 42429 30920 42441 30923
rect 42429 30892 45048 30920
rect 42429 30889 42441 30892
rect 42383 30883 42441 30889
rect 45020 30864 45048 30892
rect 33137 30855 33195 30861
rect 33137 30821 33149 30855
rect 33183 30821 33195 30855
rect 34698 30852 34704 30864
rect 34659 30824 34704 30852
rect 33137 30815 33195 30821
rect 34698 30812 34704 30824
rect 34756 30812 34762 30864
rect 35250 30852 35256 30864
rect 35211 30824 35256 30852
rect 35250 30812 35256 30824
rect 35308 30812 35314 30864
rect 35986 30852 35992 30864
rect 35947 30824 35992 30852
rect 35986 30812 35992 30824
rect 36044 30812 36050 30864
rect 36814 30852 36820 30864
rect 36775 30824 36820 30852
rect 36814 30812 36820 30824
rect 36872 30812 36878 30864
rect 38470 30852 38476 30864
rect 38431 30824 38476 30852
rect 38470 30812 38476 30824
rect 38528 30812 38534 30864
rect 40402 30852 40408 30864
rect 40363 30824 40408 30852
rect 40402 30812 40408 30824
rect 40460 30812 40466 30864
rect 40678 30812 40684 30864
rect 40736 30852 40742 30864
rect 43533 30855 43591 30861
rect 40736 30824 42323 30852
rect 40736 30812 40742 30824
rect 42295 30796 42323 30824
rect 43533 30821 43545 30855
rect 43579 30852 43591 30855
rect 43898 30852 43904 30864
rect 43579 30824 43904 30852
rect 43579 30821 43591 30824
rect 43533 30815 43591 30821
rect 43898 30812 43904 30824
rect 43956 30812 43962 30864
rect 44085 30855 44143 30861
rect 44085 30821 44097 30855
rect 44131 30852 44143 30855
rect 44266 30852 44272 30864
rect 44131 30824 44272 30852
rect 44131 30821 44143 30824
rect 44085 30815 44143 30821
rect 44266 30812 44272 30824
rect 44324 30812 44330 30864
rect 45002 30852 45008 30864
rect 44915 30824 45008 30852
rect 45002 30812 45008 30824
rect 45060 30812 45066 30864
rect 45094 30812 45100 30864
rect 45152 30852 45158 30864
rect 45152 30824 45197 30852
rect 45152 30812 45158 30824
rect 10502 30784 10508 30796
rect 10463 30756 10508 30784
rect 10502 30744 10508 30756
rect 10560 30744 10566 30796
rect 10686 30784 10692 30796
rect 10647 30756 10692 30784
rect 10686 30744 10692 30756
rect 10744 30744 10750 30796
rect 13630 30744 13636 30796
rect 13688 30784 13694 30796
rect 14236 30787 14294 30793
rect 14236 30784 14248 30787
rect 13688 30756 14248 30784
rect 13688 30744 13694 30756
rect 14236 30753 14248 30756
rect 14282 30784 14294 30787
rect 14642 30784 14648 30796
rect 14282 30756 14648 30784
rect 14282 30753 14294 30756
rect 14236 30747 14294 30753
rect 14642 30744 14648 30756
rect 14700 30744 14706 30796
rect 18322 30744 18328 30796
rect 18380 30784 18386 30796
rect 18966 30784 18972 30796
rect 18380 30756 18972 30784
rect 18380 30744 18386 30756
rect 18966 30744 18972 30756
rect 19024 30744 19030 30796
rect 19426 30784 19432 30796
rect 19076 30756 19432 30784
rect 10778 30716 10784 30728
rect 10739 30688 10784 30716
rect 10778 30676 10784 30688
rect 10836 30676 10842 30728
rect 11882 30716 11888 30728
rect 11843 30688 11888 30716
rect 11882 30676 11888 30688
rect 11940 30676 11946 30728
rect 14323 30719 14381 30725
rect 14323 30685 14335 30719
rect 14369 30716 14381 30719
rect 15010 30716 15016 30728
rect 14369 30688 15016 30716
rect 14369 30685 14381 30688
rect 14323 30679 14381 30685
rect 15010 30676 15016 30688
rect 15068 30716 15074 30728
rect 15381 30719 15439 30725
rect 15381 30716 15393 30719
rect 15068 30688 15393 30716
rect 15068 30676 15074 30688
rect 15381 30685 15393 30688
rect 15427 30685 15439 30719
rect 17494 30716 17500 30728
rect 17455 30688 17500 30716
rect 15381 30679 15439 30685
rect 17494 30676 17500 30688
rect 17552 30676 17558 30728
rect 18049 30651 18107 30657
rect 18049 30648 18061 30651
rect 16040 30620 18061 30648
rect 12802 30580 12808 30592
rect 12763 30552 12808 30580
rect 12802 30540 12808 30552
rect 12860 30540 12866 30592
rect 14366 30540 14372 30592
rect 14424 30580 14430 30592
rect 16040 30580 16068 30620
rect 18049 30617 18061 30620
rect 18095 30648 18107 30651
rect 18966 30648 18972 30660
rect 18095 30620 18972 30648
rect 18095 30617 18107 30620
rect 18049 30611 18107 30617
rect 18966 30608 18972 30620
rect 19024 30608 19030 30660
rect 16390 30580 16396 30592
rect 14424 30552 16068 30580
rect 16351 30552 16396 30580
rect 14424 30540 14430 30552
rect 16390 30540 16396 30552
rect 16448 30580 16454 30592
rect 19076 30580 19104 30756
rect 19426 30744 19432 30756
rect 19484 30744 19490 30796
rect 19886 30744 19892 30796
rect 19944 30784 19950 30796
rect 19981 30787 20039 30793
rect 19981 30784 19993 30787
rect 19944 30756 19993 30784
rect 19944 30744 19950 30756
rect 19981 30753 19993 30756
rect 20027 30753 20039 30787
rect 19981 30747 20039 30753
rect 20622 30744 20628 30796
rect 20680 30784 20686 30796
rect 21174 30784 21180 30796
rect 20680 30756 21180 30784
rect 20680 30744 20686 30756
rect 21174 30744 21180 30756
rect 21232 30744 21238 30796
rect 21634 30784 21640 30796
rect 21595 30756 21640 30784
rect 21634 30744 21640 30756
rect 21692 30744 21698 30796
rect 27065 30787 27123 30793
rect 27065 30753 27077 30787
rect 27111 30784 27123 30787
rect 27522 30784 27528 30796
rect 27111 30756 27528 30784
rect 27111 30753 27123 30756
rect 27065 30747 27123 30753
rect 21913 30719 21971 30725
rect 21913 30685 21925 30719
rect 21959 30716 21971 30719
rect 22186 30716 22192 30728
rect 21959 30688 22192 30716
rect 21959 30685 21971 30688
rect 21913 30679 21971 30685
rect 22186 30676 22192 30688
rect 22244 30676 22250 30728
rect 22646 30676 22652 30728
rect 22704 30716 22710 30728
rect 22833 30719 22891 30725
rect 22833 30716 22845 30719
rect 22704 30688 22845 30716
rect 22704 30676 22710 30688
rect 22833 30685 22845 30688
rect 22879 30685 22891 30719
rect 22833 30679 22891 30685
rect 23474 30676 23480 30728
rect 23532 30716 23538 30728
rect 24118 30716 24124 30728
rect 23532 30688 23577 30716
rect 24031 30688 24124 30716
rect 23532 30676 23538 30688
rect 24118 30676 24124 30688
rect 24176 30716 24182 30728
rect 24765 30719 24823 30725
rect 24765 30716 24777 30719
rect 24176 30688 24777 30716
rect 24176 30676 24182 30688
rect 24765 30685 24777 30688
rect 24811 30685 24823 30719
rect 24765 30679 24823 30685
rect 20346 30608 20352 30660
rect 20404 30648 20410 30660
rect 27080 30648 27108 30747
rect 27522 30744 27528 30756
rect 27580 30784 27586 30796
rect 28077 30787 28135 30793
rect 28077 30784 28089 30787
rect 27580 30756 28089 30784
rect 27580 30744 27586 30756
rect 28077 30753 28089 30756
rect 28123 30753 28135 30787
rect 28077 30747 28135 30753
rect 28997 30787 29055 30793
rect 28997 30753 29009 30787
rect 29043 30784 29055 30787
rect 29086 30784 29092 30796
rect 29043 30756 29092 30784
rect 29043 30753 29055 30756
rect 28997 30747 29055 30753
rect 29086 30744 29092 30756
rect 29144 30744 29150 30796
rect 36148 30787 36206 30793
rect 36148 30753 36160 30787
rect 36194 30784 36206 30787
rect 36354 30784 36360 30796
rect 36194 30756 36360 30784
rect 36194 30753 36206 30756
rect 36148 30747 36206 30753
rect 36354 30744 36360 30756
rect 36412 30744 36418 30796
rect 42242 30784 42248 30796
rect 42300 30793 42323 30796
rect 42300 30787 42338 30793
rect 42190 30756 42248 30784
rect 42242 30744 42248 30756
rect 42326 30753 42338 30787
rect 42300 30747 42338 30753
rect 42300 30744 42306 30747
rect 27430 30716 27436 30728
rect 27391 30688 27436 30716
rect 27430 30676 27436 30688
rect 27488 30676 27494 30728
rect 27801 30719 27859 30725
rect 27801 30685 27813 30719
rect 27847 30716 27859 30719
rect 28626 30716 28632 30728
rect 27847 30688 28632 30716
rect 27847 30685 27859 30688
rect 27801 30679 27859 30685
rect 28626 30676 28632 30688
rect 28684 30676 28690 30728
rect 30098 30716 30104 30728
rect 30059 30688 30104 30716
rect 30098 30676 30104 30688
rect 30156 30676 30162 30728
rect 30745 30719 30803 30725
rect 30745 30685 30757 30719
rect 30791 30716 30803 30719
rect 30834 30716 30840 30728
rect 30791 30688 30840 30716
rect 30791 30685 30803 30688
rect 30745 30679 30803 30685
rect 30834 30676 30840 30688
rect 30892 30676 30898 30728
rect 33226 30716 33232 30728
rect 32461 30688 33232 30716
rect 20404 30620 27108 30648
rect 20404 30608 20410 30620
rect 29546 30608 29552 30660
rect 29604 30648 29610 30660
rect 29733 30651 29791 30657
rect 29733 30648 29745 30651
rect 29604 30620 29745 30648
rect 29604 30608 29610 30620
rect 29733 30617 29745 30620
rect 29779 30617 29791 30651
rect 29733 30611 29791 30617
rect 30558 30608 30564 30660
rect 30616 30648 30622 30660
rect 32461 30648 32489 30688
rect 33226 30676 33232 30688
rect 33284 30716 33290 30728
rect 33502 30716 33508 30728
rect 33284 30688 33508 30716
rect 33284 30676 33290 30688
rect 33502 30676 33508 30688
rect 33560 30676 33566 30728
rect 33686 30716 33692 30728
rect 33647 30688 33692 30716
rect 33686 30676 33692 30688
rect 33744 30676 33750 30728
rect 34425 30719 34483 30725
rect 34425 30685 34437 30719
rect 34471 30716 34483 30719
rect 34609 30719 34667 30725
rect 34609 30716 34621 30719
rect 34471 30688 34621 30716
rect 34471 30685 34483 30688
rect 34425 30679 34483 30685
rect 34609 30685 34621 30688
rect 34655 30716 34667 30719
rect 37458 30716 37464 30728
rect 34655 30688 37464 30716
rect 34655 30685 34667 30688
rect 34609 30679 34667 30685
rect 37458 30676 37464 30688
rect 37516 30676 37522 30728
rect 38378 30716 38384 30728
rect 38339 30688 38384 30716
rect 38378 30676 38384 30688
rect 38436 30676 38442 30728
rect 38562 30676 38568 30728
rect 38620 30716 38626 30728
rect 38657 30719 38715 30725
rect 38657 30716 38669 30719
rect 38620 30688 38669 30716
rect 38620 30676 38626 30688
rect 38657 30685 38669 30688
rect 38703 30685 38715 30719
rect 38657 30679 38715 30685
rect 40313 30719 40371 30725
rect 40313 30685 40325 30719
rect 40359 30716 40371 30719
rect 40770 30716 40776 30728
rect 40359 30688 40776 30716
rect 40359 30685 40371 30688
rect 40313 30679 40371 30685
rect 30616 30620 32489 30648
rect 30616 30608 30622 30620
rect 32950 30608 32956 30660
rect 33008 30648 33014 30660
rect 33704 30648 33732 30676
rect 33008 30620 33732 30648
rect 38672 30648 38700 30679
rect 40770 30676 40776 30688
rect 40828 30716 40834 30728
rect 41138 30716 41144 30728
rect 40828 30688 41144 30716
rect 40828 30676 40834 30688
rect 41138 30676 41144 30688
rect 41196 30676 41202 30728
rect 43438 30716 43444 30728
rect 43399 30688 43444 30716
rect 43438 30676 43444 30688
rect 43496 30676 43502 30728
rect 45278 30716 45284 30728
rect 45239 30688 45284 30716
rect 45278 30676 45284 30688
rect 45336 30676 45342 30728
rect 40865 30651 40923 30657
rect 40865 30648 40877 30651
rect 38672 30620 40877 30648
rect 33008 30608 33014 30620
rect 40865 30617 40877 30620
rect 40911 30648 40923 30651
rect 41874 30648 41880 30660
rect 40911 30620 41880 30648
rect 40911 30617 40923 30620
rect 40865 30611 40923 30617
rect 41874 30608 41880 30620
rect 41932 30608 41938 30660
rect 16448 30552 19104 30580
rect 16448 30540 16454 30552
rect 21818 30540 21824 30592
rect 21876 30580 21882 30592
rect 22189 30583 22247 30589
rect 22189 30580 22201 30583
rect 21876 30552 22201 30580
rect 21876 30540 21882 30552
rect 22189 30549 22201 30552
rect 22235 30549 22247 30583
rect 25774 30580 25780 30592
rect 25735 30552 25780 30580
rect 22189 30543 22247 30549
rect 25774 30540 25780 30552
rect 25832 30540 25838 30592
rect 27062 30540 27068 30592
rect 27120 30580 27126 30592
rect 27203 30583 27261 30589
rect 27203 30580 27215 30583
rect 27120 30552 27215 30580
rect 27120 30540 27126 30552
rect 27203 30549 27215 30552
rect 27249 30549 27261 30583
rect 27203 30543 27261 30549
rect 27341 30583 27399 30589
rect 27341 30549 27353 30583
rect 27387 30580 27399 30583
rect 27614 30580 27620 30592
rect 27387 30552 27620 30580
rect 27387 30549 27399 30552
rect 27341 30543 27399 30549
rect 27614 30540 27620 30552
rect 27672 30540 27678 30592
rect 29135 30583 29193 30589
rect 29135 30549 29147 30583
rect 29181 30580 29193 30583
rect 29638 30580 29644 30592
rect 29181 30552 29644 30580
rect 29181 30549 29193 30552
rect 29135 30543 29193 30549
rect 29638 30540 29644 30552
rect 29696 30540 29702 30592
rect 30926 30540 30932 30592
rect 30984 30580 30990 30592
rect 31021 30583 31079 30589
rect 31021 30580 31033 30583
rect 30984 30552 31033 30580
rect 30984 30540 30990 30552
rect 31021 30549 31033 30552
rect 31067 30549 31079 30583
rect 31021 30543 31079 30549
rect 35250 30540 35256 30592
rect 35308 30580 35314 30592
rect 35529 30583 35587 30589
rect 35529 30580 35541 30583
rect 35308 30552 35541 30580
rect 35308 30540 35314 30552
rect 35529 30549 35541 30552
rect 35575 30549 35587 30583
rect 35529 30543 35587 30549
rect 41690 30540 41696 30592
rect 41748 30580 41754 30592
rect 44266 30580 44272 30592
rect 41748 30552 44272 30580
rect 41748 30540 41754 30552
rect 44266 30540 44272 30552
rect 44324 30540 44330 30592
rect 44450 30580 44456 30592
rect 44411 30552 44456 30580
rect 44450 30540 44456 30552
rect 44508 30540 44514 30592
rect 1104 30490 48852 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 48852 30490
rect 1104 30416 48852 30438
rect 11517 30379 11575 30385
rect 11517 30345 11529 30379
rect 11563 30376 11575 30379
rect 12802 30376 12808 30388
rect 11563 30348 12808 30376
rect 11563 30345 11575 30348
rect 11517 30339 11575 30345
rect 12802 30336 12808 30348
rect 12860 30336 12866 30388
rect 13173 30379 13231 30385
rect 13173 30345 13185 30379
rect 13219 30376 13231 30379
rect 13354 30376 13360 30388
rect 13219 30348 13360 30376
rect 13219 30345 13231 30348
rect 13173 30339 13231 30345
rect 13354 30336 13360 30348
rect 13412 30376 13418 30388
rect 14274 30376 14280 30388
rect 13412 30348 14280 30376
rect 13412 30336 13418 30348
rect 14274 30336 14280 30348
rect 14332 30336 14338 30388
rect 14642 30376 14648 30388
rect 14603 30348 14648 30376
rect 14642 30336 14648 30348
rect 14700 30336 14706 30388
rect 17310 30376 17316 30388
rect 17271 30348 17316 30376
rect 17310 30336 17316 30348
rect 17368 30336 17374 30388
rect 17586 30376 17592 30388
rect 17547 30348 17592 30376
rect 17586 30336 17592 30348
rect 17644 30336 17650 30388
rect 19426 30336 19432 30388
rect 19484 30376 19490 30388
rect 19981 30379 20039 30385
rect 19981 30376 19993 30379
rect 19484 30348 19993 30376
rect 19484 30336 19490 30348
rect 19981 30345 19993 30348
rect 20027 30345 20039 30379
rect 20622 30376 20628 30388
rect 20583 30348 20628 30376
rect 19981 30339 20039 30345
rect 20622 30336 20628 30348
rect 20680 30336 20686 30388
rect 20947 30379 21005 30385
rect 20947 30345 20959 30379
rect 20993 30376 21005 30379
rect 22646 30376 22652 30388
rect 20993 30348 22652 30376
rect 20993 30345 21005 30348
rect 20947 30339 21005 30345
rect 22646 30336 22652 30348
rect 22704 30336 22710 30388
rect 22741 30379 22799 30385
rect 22741 30345 22753 30379
rect 22787 30376 22799 30379
rect 22922 30376 22928 30388
rect 22787 30348 22928 30376
rect 22787 30345 22799 30348
rect 22741 30339 22799 30345
rect 22922 30336 22928 30348
rect 22980 30376 22986 30388
rect 23017 30379 23075 30385
rect 23017 30376 23029 30379
rect 22980 30348 23029 30376
rect 22980 30336 22986 30348
rect 23017 30345 23029 30348
rect 23063 30345 23075 30379
rect 23017 30339 23075 30345
rect 23799 30379 23857 30385
rect 23799 30345 23811 30379
rect 23845 30376 23857 30379
rect 24118 30376 24124 30388
rect 23845 30348 24124 30376
rect 23845 30345 23857 30348
rect 23799 30339 23857 30345
rect 24118 30336 24124 30348
rect 24176 30336 24182 30388
rect 25777 30379 25835 30385
rect 25777 30345 25789 30379
rect 25823 30376 25835 30379
rect 25866 30376 25872 30388
rect 25823 30348 25872 30376
rect 25823 30345 25835 30348
rect 25777 30339 25835 30345
rect 9723 30311 9781 30317
rect 9723 30277 9735 30311
rect 9769 30308 9781 30311
rect 11882 30308 11888 30320
rect 9769 30280 11888 30308
rect 9769 30277 9781 30280
rect 9723 30271 9781 30277
rect 11882 30268 11888 30280
rect 11940 30308 11946 30320
rect 12161 30311 12219 30317
rect 12161 30308 12173 30311
rect 11940 30280 12173 30308
rect 11940 30268 11946 30280
rect 12161 30277 12173 30280
rect 12207 30277 12219 30311
rect 14921 30311 14979 30317
rect 14921 30308 14933 30311
rect 12161 30271 12219 30277
rect 12360 30280 14933 30308
rect 10597 30243 10655 30249
rect 10597 30209 10609 30243
rect 10643 30240 10655 30243
rect 10778 30240 10784 30252
rect 10643 30212 10784 30240
rect 10643 30209 10655 30212
rect 10597 30203 10655 30209
rect 10778 30200 10784 30212
rect 10836 30200 10842 30252
rect 11790 30240 11796 30252
rect 11703 30212 11796 30240
rect 11790 30200 11796 30212
rect 11848 30240 11854 30252
rect 11974 30240 11980 30252
rect 11848 30212 11980 30240
rect 11848 30200 11854 30212
rect 11974 30200 11980 30212
rect 12032 30240 12038 30252
rect 12360 30240 12388 30280
rect 14921 30277 14933 30280
rect 14967 30308 14979 30311
rect 15013 30311 15071 30317
rect 15013 30308 15025 30311
rect 14967 30280 15025 30308
rect 14967 30277 14979 30280
rect 14921 30271 14979 30277
rect 15013 30277 15025 30280
rect 15059 30277 15071 30311
rect 15838 30308 15844 30320
rect 15799 30280 15844 30308
rect 15013 30271 15071 30277
rect 15838 30268 15844 30280
rect 15896 30268 15902 30320
rect 21637 30311 21695 30317
rect 21637 30277 21649 30311
rect 21683 30277 21695 30311
rect 22664 30308 22692 30336
rect 23385 30311 23443 30317
rect 23385 30308 23397 30311
rect 22664 30280 23397 30308
rect 21637 30271 21695 30277
rect 23385 30277 23397 30280
rect 23431 30277 23443 30311
rect 23385 30271 23443 30277
rect 12032 30212 12388 30240
rect 12759 30243 12817 30249
rect 12032 30200 12038 30212
rect 12759 30209 12771 30243
rect 12805 30240 12817 30243
rect 15289 30243 15347 30249
rect 15289 30240 15301 30243
rect 12805 30212 15301 30240
rect 12805 30209 12817 30212
rect 12759 30203 12817 30209
rect 15289 30209 15301 30212
rect 15335 30240 15347 30243
rect 16577 30243 16635 30249
rect 16577 30240 16589 30243
rect 15335 30212 16589 30240
rect 15335 30209 15347 30212
rect 15289 30203 15347 30209
rect 16577 30209 16589 30212
rect 16623 30209 16635 30243
rect 16577 30203 16635 30209
rect 18785 30243 18843 30249
rect 18785 30209 18797 30243
rect 18831 30240 18843 30243
rect 19058 30240 19064 30252
rect 18831 30212 19064 30240
rect 18831 30209 18843 30212
rect 18785 30203 18843 30209
rect 19058 30200 19064 30212
rect 19116 30200 19122 30252
rect 9652 30175 9710 30181
rect 9652 30141 9664 30175
rect 9698 30172 9710 30175
rect 11238 30172 11244 30184
rect 9698 30144 11244 30172
rect 9698 30141 9710 30144
rect 9652 30135 9710 30141
rect 10060 30048 10088 30144
rect 11238 30132 11244 30144
rect 11296 30132 11302 30184
rect 12672 30175 12730 30181
rect 12672 30141 12684 30175
rect 12718 30172 12730 30175
rect 13354 30172 13360 30184
rect 12718 30144 13360 30172
rect 12718 30141 12730 30144
rect 12672 30135 12730 30141
rect 13354 30132 13360 30144
rect 13412 30132 13418 30184
rect 14366 30132 14372 30184
rect 14424 30172 14430 30184
rect 16828 30175 16886 30181
rect 14424 30144 14469 30172
rect 14424 30132 14430 30144
rect 16828 30141 16840 30175
rect 16874 30172 16886 30175
rect 17310 30172 17316 30184
rect 16874 30144 17316 30172
rect 16874 30141 16886 30144
rect 16828 30135 16886 30141
rect 17310 30132 17316 30144
rect 17368 30132 17374 30184
rect 17678 30132 17684 30184
rect 17736 30172 17742 30184
rect 19886 30172 19892 30184
rect 17736 30144 19892 30172
rect 17736 30132 17742 30144
rect 19886 30132 19892 30144
rect 19944 30172 19950 30184
rect 20876 30175 20934 30181
rect 20876 30172 20888 30175
rect 19944 30144 20888 30172
rect 19944 30132 19950 30144
rect 20876 30141 20888 30144
rect 20922 30172 20934 30175
rect 21358 30172 21364 30184
rect 20922 30144 21364 30172
rect 20922 30141 20934 30144
rect 20876 30135 20934 30141
rect 21358 30132 21364 30144
rect 21416 30132 21422 30184
rect 10505 30107 10563 30113
rect 10505 30073 10517 30107
rect 10551 30104 10563 30107
rect 10959 30107 11017 30113
rect 10959 30104 10971 30107
rect 10551 30076 10971 30104
rect 10551 30073 10563 30076
rect 10505 30067 10563 30073
rect 10959 30073 10971 30076
rect 11005 30104 11017 30107
rect 11330 30104 11336 30116
rect 11005 30076 11336 30104
rect 11005 30073 11017 30076
rect 10959 30067 11017 30073
rect 11330 30064 11336 30076
rect 11388 30064 11394 30116
rect 13722 30104 13728 30116
rect 13683 30076 13728 30104
rect 13722 30064 13728 30076
rect 13780 30064 13786 30116
rect 13814 30064 13820 30116
rect 13872 30104 13878 30116
rect 14921 30107 14979 30113
rect 13872 30076 13917 30104
rect 13872 30064 13878 30076
rect 14921 30073 14933 30107
rect 14967 30104 14979 30107
rect 15381 30107 15439 30113
rect 15381 30104 15393 30107
rect 14967 30076 15393 30104
rect 14967 30073 14979 30076
rect 14921 30067 14979 30073
rect 15381 30073 15393 30076
rect 15427 30104 15439 30107
rect 15470 30104 15476 30116
rect 15427 30076 15476 30104
rect 15427 30073 15439 30076
rect 15381 30067 15439 30073
rect 15470 30064 15476 30076
rect 15528 30064 15534 30116
rect 18506 30064 18512 30116
rect 18564 30104 18570 30116
rect 18693 30107 18751 30113
rect 18693 30104 18705 30107
rect 18564 30076 18705 30104
rect 18564 30064 18570 30076
rect 18693 30073 18705 30076
rect 18739 30104 18751 30107
rect 19147 30107 19205 30113
rect 19147 30104 19159 30107
rect 18739 30076 19159 30104
rect 18739 30073 18751 30076
rect 18693 30067 18751 30073
rect 19147 30073 19159 30076
rect 19193 30104 19205 30107
rect 21652 30104 21680 30271
rect 24765 30243 24823 30249
rect 24765 30209 24777 30243
rect 24811 30240 24823 30243
rect 25792 30240 25820 30339
rect 25866 30336 25872 30348
rect 25924 30336 25930 30388
rect 25961 30379 26019 30385
rect 25961 30345 25973 30379
rect 26007 30376 26019 30379
rect 28307 30379 28365 30385
rect 26007 30348 28279 30376
rect 26007 30345 26019 30348
rect 25961 30339 26019 30345
rect 24811 30212 25820 30240
rect 25884 30280 26464 30308
rect 24811 30209 24823 30212
rect 24765 30203 24823 30209
rect 21818 30172 21824 30184
rect 21779 30144 21824 30172
rect 21818 30132 21824 30144
rect 21876 30132 21882 30184
rect 23569 30175 23627 30181
rect 23569 30141 23581 30175
rect 23615 30172 23627 30175
rect 23750 30172 23756 30184
rect 23615 30144 23756 30172
rect 23615 30141 23627 30144
rect 23569 30135 23627 30141
rect 23750 30132 23756 30144
rect 23808 30132 23814 30184
rect 25409 30175 25467 30181
rect 25409 30141 25421 30175
rect 25455 30172 25467 30175
rect 25590 30172 25596 30184
rect 25455 30144 25596 30172
rect 25455 30141 25467 30144
rect 25409 30135 25467 30141
rect 25590 30132 25596 30144
rect 25648 30172 25654 30184
rect 25884 30172 25912 30280
rect 26326 30240 26332 30252
rect 26287 30212 26332 30240
rect 26326 30200 26332 30212
rect 26384 30200 26390 30252
rect 26436 30240 26464 30280
rect 26605 30243 26663 30249
rect 26605 30240 26617 30243
rect 26436 30212 26617 30240
rect 26605 30209 26617 30212
rect 26651 30209 26663 30243
rect 26605 30203 26663 30209
rect 28251 30181 28279 30348
rect 28307 30345 28319 30379
rect 28353 30376 28365 30379
rect 29546 30376 29552 30388
rect 28353 30348 29552 30376
rect 28353 30345 28365 30348
rect 28307 30339 28365 30345
rect 29546 30336 29552 30348
rect 29604 30336 29610 30388
rect 29779 30379 29837 30385
rect 29779 30345 29791 30379
rect 29825 30376 29837 30379
rect 30098 30376 30104 30388
rect 29825 30348 30104 30376
rect 29825 30345 29837 30348
rect 29779 30339 29837 30345
rect 30098 30336 30104 30348
rect 30156 30336 30162 30388
rect 30466 30376 30472 30388
rect 30427 30348 30472 30376
rect 30466 30336 30472 30348
rect 30524 30336 30530 30388
rect 32677 30379 32735 30385
rect 32677 30345 32689 30379
rect 32723 30376 32735 30379
rect 32858 30376 32864 30388
rect 32723 30348 32864 30376
rect 32723 30345 32735 30348
rect 32677 30339 32735 30345
rect 32858 30336 32864 30348
rect 32916 30336 32922 30388
rect 33042 30376 33048 30388
rect 33003 30348 33048 30376
rect 33042 30336 33048 30348
rect 33100 30336 33106 30388
rect 36173 30379 36231 30385
rect 36173 30345 36185 30379
rect 36219 30376 36231 30379
rect 36354 30376 36360 30388
rect 36219 30348 36360 30376
rect 36219 30345 36231 30348
rect 36173 30339 36231 30345
rect 36354 30336 36360 30348
rect 36412 30336 36418 30388
rect 37277 30379 37335 30385
rect 37277 30345 37289 30379
rect 37323 30376 37335 30379
rect 37826 30376 37832 30388
rect 37323 30348 37832 30376
rect 37323 30345 37335 30348
rect 37277 30339 37335 30345
rect 37826 30336 37832 30348
rect 37884 30336 37890 30388
rect 38289 30379 38347 30385
rect 38289 30345 38301 30379
rect 38335 30376 38347 30379
rect 38470 30376 38476 30388
rect 38335 30348 38476 30376
rect 38335 30345 38347 30348
rect 38289 30339 38347 30345
rect 38470 30336 38476 30348
rect 38528 30376 38534 30388
rect 38565 30379 38623 30385
rect 38565 30376 38577 30379
rect 38528 30348 38577 30376
rect 38528 30336 38534 30348
rect 38565 30345 38577 30348
rect 38611 30345 38623 30379
rect 38565 30339 38623 30345
rect 40313 30379 40371 30385
rect 40313 30345 40325 30379
rect 40359 30376 40371 30379
rect 40402 30376 40408 30388
rect 40359 30348 40408 30376
rect 40359 30345 40371 30348
rect 40313 30339 40371 30345
rect 40402 30336 40408 30348
rect 40460 30336 40466 30388
rect 42843 30379 42901 30385
rect 40512 30348 42794 30376
rect 29638 30268 29644 30320
rect 29696 30308 29702 30320
rect 29696 30280 33134 30308
rect 29696 30268 29702 30280
rect 29086 30240 29092 30252
rect 28999 30212 29092 30240
rect 29086 30200 29092 30212
rect 29144 30240 29150 30252
rect 30190 30240 30196 30252
rect 29144 30212 30196 30240
rect 29144 30200 29150 30212
rect 30190 30200 30196 30212
rect 30248 30200 30254 30252
rect 30834 30240 30840 30252
rect 30747 30212 30840 30240
rect 30834 30200 30840 30212
rect 30892 30240 30898 30252
rect 31294 30240 31300 30252
rect 30892 30212 31300 30240
rect 30892 30200 30898 30212
rect 31294 30200 31300 30212
rect 31352 30200 31358 30252
rect 33106 30240 33134 30280
rect 33962 30268 33968 30320
rect 34020 30308 34026 30320
rect 34020 30280 38102 30308
rect 34020 30268 34026 30280
rect 34977 30243 35035 30249
rect 34977 30240 34989 30243
rect 33106 30212 34989 30240
rect 34977 30209 34989 30212
rect 35023 30240 35035 30243
rect 35250 30240 35256 30252
rect 35023 30212 35256 30240
rect 35023 30209 35035 30212
rect 34977 30203 35035 30209
rect 35250 30200 35256 30212
rect 35308 30200 35314 30252
rect 35342 30200 35348 30252
rect 35400 30240 35406 30252
rect 37366 30240 37372 30252
rect 35400 30212 35445 30240
rect 37327 30212 37372 30240
rect 35400 30200 35406 30212
rect 37366 30200 37372 30212
rect 37424 30200 37430 30252
rect 38074 30240 38102 30280
rect 38378 30268 38384 30320
rect 38436 30308 38442 30320
rect 39025 30311 39083 30317
rect 39025 30308 39037 30311
rect 38436 30280 39037 30308
rect 38436 30268 38442 30280
rect 39025 30277 39037 30280
rect 39071 30308 39083 30311
rect 40512 30308 40540 30348
rect 39071 30280 40540 30308
rect 39071 30277 39083 30280
rect 39025 30271 39083 30277
rect 41506 30268 41512 30320
rect 41564 30308 41570 30320
rect 42242 30308 42248 30320
rect 41564 30280 41920 30308
rect 42203 30280 42248 30308
rect 41564 30268 41570 30280
rect 39255 30243 39313 30249
rect 39255 30240 39267 30243
rect 38074 30212 39267 30240
rect 39255 30209 39267 30212
rect 39301 30209 39313 30243
rect 39255 30203 39313 30209
rect 41233 30243 41291 30249
rect 41233 30209 41245 30243
rect 41279 30240 41291 30243
rect 41690 30240 41696 30252
rect 41279 30212 41696 30240
rect 41279 30209 41291 30212
rect 41233 30203 41291 30209
rect 41690 30200 41696 30212
rect 41748 30200 41754 30252
rect 25648 30144 25912 30172
rect 28236 30175 28294 30181
rect 25648 30132 25654 30144
rect 28236 30141 28248 30175
rect 28282 30172 28294 30175
rect 28282 30144 28764 30172
rect 28282 30141 28294 30144
rect 28236 30135 28294 30141
rect 22142 30107 22200 30113
rect 22142 30104 22154 30107
rect 19193 30076 22154 30104
rect 19193 30073 19205 30076
rect 19147 30067 19205 30073
rect 22142 30073 22154 30076
rect 22188 30104 22200 30107
rect 22462 30104 22468 30116
rect 22188 30076 22468 30104
rect 22188 30073 22200 30076
rect 22142 30067 22200 30073
rect 22462 30064 22468 30076
rect 22520 30064 22526 30116
rect 22922 30064 22928 30116
rect 22980 30104 22986 30116
rect 24489 30107 24547 30113
rect 24489 30104 24501 30107
rect 22980 30076 24501 30104
rect 22980 30064 22986 30076
rect 24489 30073 24501 30076
rect 24535 30104 24547 30107
rect 24857 30107 24915 30113
rect 24857 30104 24869 30107
rect 24535 30076 24869 30104
rect 24535 30073 24547 30076
rect 24489 30067 24547 30073
rect 24857 30073 24869 30076
rect 24903 30104 24915 30107
rect 24946 30104 24952 30116
rect 24903 30076 24952 30104
rect 24903 30073 24915 30076
rect 24857 30067 24915 30073
rect 24946 30064 24952 30076
rect 25004 30064 25010 30116
rect 25961 30107 26019 30113
rect 25961 30104 25973 30107
rect 25193 30076 25973 30104
rect 9490 30036 9496 30048
rect 9451 30008 9496 30036
rect 9490 29996 9496 30008
rect 9548 29996 9554 30048
rect 10042 30036 10048 30048
rect 10003 30008 10048 30036
rect 10042 29996 10048 30008
rect 10100 29996 10106 30048
rect 13541 30039 13599 30045
rect 13541 30005 13553 30039
rect 13587 30036 13599 30039
rect 13832 30036 13860 30064
rect 13587 30008 13860 30036
rect 15488 30036 15516 30064
rect 16209 30039 16267 30045
rect 16209 30036 16221 30039
rect 15488 30008 16221 30036
rect 13587 30005 13599 30008
rect 13541 29999 13599 30005
rect 16209 30005 16221 30008
rect 16255 30005 16267 30039
rect 16209 29999 16267 30005
rect 16298 29996 16304 30048
rect 16356 30036 16362 30048
rect 16899 30039 16957 30045
rect 16899 30036 16911 30039
rect 16356 30008 16911 30036
rect 16356 29996 16362 30008
rect 16899 30005 16911 30008
rect 16945 30005 16957 30039
rect 18322 30036 18328 30048
rect 18283 30008 18328 30036
rect 16899 29999 16957 30005
rect 18322 29996 18328 30008
rect 18380 29996 18386 30048
rect 18874 29996 18880 30048
rect 18932 30036 18938 30048
rect 19705 30039 19763 30045
rect 19705 30036 19717 30039
rect 18932 30008 19717 30036
rect 18932 29996 18938 30008
rect 19705 30005 19717 30008
rect 19751 30005 19763 30039
rect 19705 29999 19763 30005
rect 23750 29996 23756 30048
rect 23808 30036 23814 30048
rect 24213 30039 24271 30045
rect 24213 30036 24225 30039
rect 23808 30008 24225 30036
rect 23808 29996 23814 30008
rect 24213 30005 24225 30008
rect 24259 30036 24271 30039
rect 25193 30036 25221 30076
rect 25961 30073 25973 30076
rect 26007 30073 26019 30107
rect 25961 30067 26019 30073
rect 26421 30107 26479 30113
rect 26421 30073 26433 30107
rect 26467 30073 26479 30107
rect 26421 30067 26479 30073
rect 24259 30008 25221 30036
rect 24259 30005 24271 30008
rect 24213 29999 24271 30005
rect 25406 29996 25412 30048
rect 25464 30036 25470 30048
rect 26053 30039 26111 30045
rect 26053 30036 26065 30039
rect 25464 30008 26065 30036
rect 25464 29996 25470 30008
rect 26053 30005 26065 30008
rect 26099 30036 26111 30039
rect 26436 30036 26464 30067
rect 26099 30008 26464 30036
rect 27341 30039 27399 30045
rect 26099 30005 26111 30008
rect 26053 29999 26111 30005
rect 27341 30005 27353 30039
rect 27387 30036 27399 30039
rect 27430 30036 27436 30048
rect 27387 30008 27436 30036
rect 27387 30005 27399 30008
rect 27341 29999 27399 30005
rect 27430 29996 27436 30008
rect 27488 29996 27494 30048
rect 27614 30036 27620 30048
rect 27575 30008 27620 30036
rect 27614 29996 27620 30008
rect 27672 29996 27678 30048
rect 28736 30045 28764 30144
rect 29546 30132 29552 30184
rect 29604 30172 29610 30184
rect 29676 30175 29734 30181
rect 29676 30172 29688 30175
rect 29604 30144 29688 30172
rect 29604 30132 29610 30144
rect 29676 30141 29688 30144
rect 29722 30172 29734 30175
rect 30006 30172 30012 30184
rect 29722 30144 30012 30172
rect 29722 30141 29734 30144
rect 29676 30135 29734 30141
rect 30006 30132 30012 30144
rect 30064 30172 30070 30184
rect 30101 30175 30159 30181
rect 30101 30172 30113 30175
rect 30064 30144 30113 30172
rect 30064 30132 30070 30144
rect 30101 30141 30113 30144
rect 30147 30141 30159 30175
rect 30101 30135 30159 30141
rect 39022 30132 39028 30184
rect 39080 30172 39086 30184
rect 39152 30175 39210 30181
rect 39152 30172 39164 30175
rect 39080 30144 39164 30172
rect 39080 30132 39086 30144
rect 39152 30141 39164 30144
rect 39198 30172 39210 30175
rect 39577 30175 39635 30181
rect 39577 30172 39589 30175
rect 39198 30144 39589 30172
rect 39198 30141 39210 30144
rect 39152 30135 39210 30141
rect 39577 30141 39589 30144
rect 39623 30141 39635 30175
rect 41892 30172 41920 30280
rect 42242 30268 42248 30280
rect 42300 30268 42306 30320
rect 42766 30308 42794 30348
rect 42843 30345 42855 30379
rect 42889 30376 42901 30379
rect 43438 30376 43444 30388
rect 42889 30348 43444 30376
rect 42889 30345 42901 30348
rect 42843 30339 42901 30345
rect 43438 30336 43444 30348
rect 43496 30336 43502 30388
rect 44450 30336 44456 30388
rect 44508 30376 44514 30388
rect 46247 30379 46305 30385
rect 46247 30376 46259 30379
rect 44508 30348 46259 30376
rect 44508 30336 44514 30348
rect 46247 30345 46259 30348
rect 46293 30345 46305 30379
rect 46566 30376 46572 30388
rect 46527 30348 46572 30376
rect 46247 30339 46305 30345
rect 46566 30336 46572 30348
rect 46624 30336 46630 30388
rect 42978 30308 42984 30320
rect 42766 30280 42984 30308
rect 42978 30268 42984 30280
rect 43036 30268 43042 30320
rect 44358 30308 44364 30320
rect 44319 30280 44364 30308
rect 44358 30268 44364 30280
rect 44416 30268 44422 30320
rect 42260 30240 42288 30268
rect 43622 30240 43628 30252
rect 42260 30212 43628 30240
rect 43622 30200 43628 30212
rect 43680 30200 43686 30252
rect 43809 30243 43867 30249
rect 43809 30209 43821 30243
rect 43855 30240 43867 30243
rect 44468 30240 44496 30336
rect 45002 30268 45008 30320
rect 45060 30308 45066 30320
rect 45465 30311 45523 30317
rect 45465 30308 45477 30311
rect 45060 30280 45477 30308
rect 45060 30268 45066 30280
rect 45465 30277 45477 30280
rect 45511 30277 45523 30311
rect 45465 30271 45523 30277
rect 43855 30212 44496 30240
rect 44821 30243 44879 30249
rect 43855 30209 43867 30212
rect 43809 30203 43867 30209
rect 44821 30209 44833 30243
rect 44867 30240 44879 30243
rect 45094 30240 45100 30252
rect 44867 30212 45100 30240
rect 44867 30209 44879 30212
rect 44821 30203 44879 30209
rect 45094 30200 45100 30212
rect 45152 30200 45158 30252
rect 42794 30181 42800 30184
rect 42772 30175 42800 30181
rect 42772 30172 42784 30175
rect 41892 30144 42784 30172
rect 39577 30135 39635 30141
rect 42772 30141 42784 30144
rect 42852 30172 42858 30184
rect 43165 30175 43223 30181
rect 43165 30172 43177 30175
rect 42852 30144 43177 30172
rect 42772 30135 42800 30141
rect 42794 30132 42800 30135
rect 42852 30132 42858 30144
rect 43165 30141 43177 30144
rect 43211 30141 43223 30175
rect 43165 30135 43223 30141
rect 44450 30132 44456 30184
rect 44508 30172 44514 30184
rect 46176 30175 46234 30181
rect 46176 30172 46188 30175
rect 44508 30144 46188 30172
rect 44508 30132 44514 30144
rect 46176 30141 46188 30144
rect 46222 30172 46234 30175
rect 46566 30172 46572 30184
rect 46222 30144 46572 30172
rect 46222 30141 46234 30144
rect 46176 30135 46234 30141
rect 46566 30132 46572 30144
rect 46624 30132 46630 30184
rect 30926 30064 30932 30116
rect 30984 30104 30990 30116
rect 31481 30107 31539 30113
rect 30984 30076 31029 30104
rect 30984 30064 30990 30076
rect 31481 30073 31493 30107
rect 31527 30073 31539 30107
rect 33318 30104 33324 30116
rect 33279 30076 33324 30104
rect 31481 30067 31539 30073
rect 28721 30039 28779 30045
rect 28721 30005 28733 30039
rect 28767 30036 28779 30039
rect 28810 30036 28816 30048
rect 28767 30008 28816 30036
rect 28767 30005 28779 30008
rect 28721 29999 28779 30005
rect 28810 29996 28816 30008
rect 28868 29996 28874 30048
rect 31386 29996 31392 30048
rect 31444 30036 31450 30048
rect 31496 30036 31524 30067
rect 33318 30064 33324 30076
rect 33376 30064 33382 30116
rect 33410 30064 33416 30116
rect 33468 30104 33474 30116
rect 33468 30076 33513 30104
rect 33468 30064 33474 30076
rect 33686 30064 33692 30116
rect 33744 30104 33750 30116
rect 33965 30107 34023 30113
rect 33965 30104 33977 30107
rect 33744 30076 33977 30104
rect 33744 30064 33750 30076
rect 33965 30073 33977 30076
rect 34011 30104 34023 30107
rect 34330 30104 34336 30116
rect 34011 30076 34336 30104
rect 34011 30073 34023 30076
rect 33965 30067 34023 30073
rect 34330 30064 34336 30076
rect 34388 30064 34394 30116
rect 35069 30107 35127 30113
rect 35069 30073 35081 30107
rect 35115 30073 35127 30107
rect 35069 30067 35127 30073
rect 37731 30107 37789 30113
rect 37731 30073 37743 30107
rect 37777 30104 37789 30107
rect 37826 30104 37832 30116
rect 37777 30076 37832 30104
rect 37777 30073 37789 30076
rect 37731 30067 37789 30073
rect 31444 30008 31524 30036
rect 33428 30036 33456 30064
rect 34517 30039 34575 30045
rect 34517 30036 34529 30039
rect 33428 30008 34529 30036
rect 31444 29996 31450 30008
rect 34517 30005 34529 30008
rect 34563 30036 34575 30039
rect 34974 30036 34980 30048
rect 34563 30008 34980 30036
rect 34563 30005 34575 30008
rect 34517 29999 34575 30005
rect 34974 29996 34980 30008
rect 35032 30036 35038 30048
rect 35084 30036 35112 30067
rect 37826 30064 37832 30076
rect 37884 30064 37890 30116
rect 41322 30064 41328 30116
rect 41380 30104 41386 30116
rect 41874 30104 41880 30116
rect 41380 30076 41425 30104
rect 41835 30076 41880 30104
rect 41380 30064 41386 30076
rect 41874 30064 41880 30076
rect 41932 30064 41938 30116
rect 43625 30107 43683 30113
rect 43625 30073 43637 30107
rect 43671 30104 43683 30107
rect 43898 30104 43904 30116
rect 43671 30076 43904 30104
rect 43671 30073 43683 30076
rect 43625 30067 43683 30073
rect 43898 30064 43904 30076
rect 43956 30064 43962 30116
rect 35032 30008 35112 30036
rect 41049 30039 41107 30045
rect 35032 29996 35038 30008
rect 41049 30005 41061 30039
rect 41095 30036 41107 30039
rect 41340 30036 41368 30064
rect 41095 30008 41368 30036
rect 41095 30005 41107 30008
rect 41049 29999 41107 30005
rect 1104 29946 48852 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 48852 29946
rect 1104 29872 48852 29894
rect 10413 29835 10471 29841
rect 10413 29801 10425 29835
rect 10459 29832 10471 29835
rect 10502 29832 10508 29844
rect 10459 29804 10508 29832
rect 10459 29801 10471 29804
rect 10413 29795 10471 29801
rect 10502 29792 10508 29804
rect 10560 29792 10566 29844
rect 10778 29832 10784 29844
rect 10739 29804 10784 29832
rect 10778 29792 10784 29804
rect 10836 29792 10842 29844
rect 11790 29832 11796 29844
rect 11751 29804 11796 29832
rect 11790 29792 11796 29804
rect 11848 29792 11854 29844
rect 13814 29792 13820 29844
rect 13872 29832 13878 29844
rect 13909 29835 13967 29841
rect 13909 29832 13921 29835
rect 13872 29804 13921 29832
rect 13872 29792 13878 29804
rect 13909 29801 13921 29804
rect 13955 29801 13967 29835
rect 15010 29832 15016 29844
rect 14971 29804 15016 29832
rect 13909 29795 13967 29801
rect 15010 29792 15016 29804
rect 15068 29792 15074 29844
rect 17310 29832 17316 29844
rect 15304 29804 17316 29832
rect 11235 29767 11293 29773
rect 11235 29733 11247 29767
rect 11281 29764 11293 29767
rect 11330 29764 11336 29776
rect 11281 29736 11336 29764
rect 11281 29733 11293 29736
rect 11235 29727 11293 29733
rect 11330 29724 11336 29736
rect 11388 29724 11394 29776
rect 13351 29767 13409 29773
rect 13351 29733 13363 29767
rect 13397 29764 13409 29767
rect 13446 29764 13452 29776
rect 13397 29736 13452 29764
rect 13397 29733 13409 29736
rect 13351 29727 13409 29733
rect 13446 29724 13452 29736
rect 13504 29764 13510 29776
rect 15304 29764 15332 29804
rect 17310 29792 17316 29804
rect 17368 29792 17374 29844
rect 17586 29792 17592 29844
rect 17644 29832 17650 29844
rect 17865 29835 17923 29841
rect 17865 29832 17877 29835
rect 17644 29804 17877 29832
rect 17644 29792 17650 29804
rect 17865 29801 17877 29804
rect 17911 29801 17923 29835
rect 17865 29795 17923 29801
rect 18601 29835 18659 29841
rect 18601 29801 18613 29835
rect 18647 29832 18659 29835
rect 19058 29832 19064 29844
rect 18647 29804 19064 29832
rect 18647 29801 18659 29804
rect 18601 29795 18659 29801
rect 19058 29792 19064 29804
rect 19116 29792 19122 29844
rect 22462 29792 22468 29844
rect 22520 29832 22526 29844
rect 22557 29835 22615 29841
rect 22557 29832 22569 29835
rect 22520 29804 22569 29832
rect 22520 29792 22526 29804
rect 22557 29801 22569 29804
rect 22603 29801 22615 29835
rect 22557 29795 22615 29801
rect 23109 29835 23167 29841
rect 23109 29801 23121 29835
rect 23155 29832 23167 29835
rect 24946 29832 24952 29844
rect 23155 29804 24164 29832
rect 24907 29804 24952 29832
rect 23155 29801 23167 29804
rect 23109 29795 23167 29801
rect 24136 29776 24164 29804
rect 24946 29792 24952 29804
rect 25004 29792 25010 29844
rect 25406 29792 25412 29844
rect 25464 29832 25470 29844
rect 25501 29835 25559 29841
rect 25501 29832 25513 29835
rect 25464 29804 25513 29832
rect 25464 29792 25470 29804
rect 25501 29801 25513 29804
rect 25547 29801 25559 29835
rect 25501 29795 25559 29801
rect 25774 29792 25780 29844
rect 25832 29832 25838 29844
rect 26651 29835 26709 29841
rect 26651 29832 26663 29835
rect 25832 29804 26663 29832
rect 25832 29792 25838 29804
rect 26651 29801 26663 29804
rect 26697 29801 26709 29835
rect 27522 29832 27528 29844
rect 27483 29804 27528 29832
rect 26651 29795 26709 29801
rect 27522 29792 27528 29804
rect 27580 29792 27586 29844
rect 30098 29832 30104 29844
rect 30059 29804 30104 29832
rect 30098 29792 30104 29804
rect 30156 29792 30162 29844
rect 33318 29792 33324 29844
rect 33376 29832 33382 29844
rect 33597 29835 33655 29841
rect 33597 29832 33609 29835
rect 33376 29804 33609 29832
rect 33376 29792 33382 29804
rect 33597 29801 33609 29804
rect 33643 29801 33655 29835
rect 34974 29832 34980 29844
rect 34935 29804 34980 29832
rect 33597 29795 33655 29801
rect 34974 29792 34980 29804
rect 35032 29792 35038 29844
rect 36630 29792 36636 29844
rect 36688 29832 36694 29844
rect 37001 29835 37059 29841
rect 37001 29832 37013 29835
rect 36688 29804 37013 29832
rect 36688 29792 36694 29804
rect 37001 29801 37013 29804
rect 37047 29801 37059 29835
rect 37366 29832 37372 29844
rect 37327 29804 37372 29832
rect 37001 29795 37059 29801
rect 37366 29792 37372 29804
rect 37424 29792 37430 29844
rect 40402 29832 40408 29844
rect 40363 29804 40408 29832
rect 40402 29792 40408 29804
rect 40460 29792 40466 29844
rect 40770 29832 40776 29844
rect 40731 29804 40776 29832
rect 40770 29792 40776 29804
rect 40828 29792 40834 29844
rect 41322 29792 41328 29844
rect 41380 29832 41386 29844
rect 42153 29835 42211 29841
rect 42153 29832 42165 29835
rect 41380 29804 42165 29832
rect 41380 29792 41386 29804
rect 42153 29801 42165 29804
rect 42199 29801 42211 29835
rect 43717 29835 43775 29841
rect 43717 29832 43729 29835
rect 42153 29795 42211 29801
rect 42766 29804 43729 29832
rect 15470 29764 15476 29776
rect 13504 29736 15332 29764
rect 15431 29736 15476 29764
rect 13504 29724 13510 29736
rect 15470 29724 15476 29736
rect 15528 29724 15534 29776
rect 17494 29724 17500 29776
rect 17552 29764 17558 29776
rect 18141 29767 18199 29773
rect 18141 29764 18153 29767
rect 17552 29736 18153 29764
rect 17552 29724 17558 29736
rect 18141 29733 18153 29736
rect 18187 29733 18199 29767
rect 18874 29764 18880 29776
rect 18835 29736 18880 29764
rect 18141 29727 18199 29733
rect 18874 29724 18880 29736
rect 18932 29724 18938 29776
rect 24118 29764 24124 29776
rect 24031 29736 24124 29764
rect 24118 29724 24124 29736
rect 24176 29764 24182 29776
rect 25424 29764 25452 29792
rect 26326 29764 26332 29776
rect 24176 29736 25452 29764
rect 26287 29736 26332 29764
rect 24176 29724 24182 29736
rect 26326 29724 26332 29736
rect 26384 29724 26390 29776
rect 30374 29764 30380 29776
rect 30335 29736 30380 29764
rect 30374 29724 30380 29736
rect 30432 29724 30438 29776
rect 31938 29724 31944 29776
rect 31996 29764 32002 29776
rect 31996 29736 32327 29764
rect 31996 29724 32002 29736
rect 12894 29696 12900 29708
rect 9876 29668 12900 29696
rect 9876 29640 9904 29668
rect 12894 29656 12900 29668
rect 12952 29696 12958 29708
rect 14366 29696 14372 29708
rect 12952 29668 14372 29696
rect 12952 29656 12958 29668
rect 14366 29656 14372 29668
rect 14424 29656 14430 29708
rect 21082 29656 21088 29708
rect 21140 29696 21146 29708
rect 21212 29699 21270 29705
rect 21212 29696 21224 29699
rect 21140 29668 21224 29696
rect 21140 29656 21146 29668
rect 21212 29665 21224 29668
rect 21258 29665 21270 29699
rect 21212 29659 21270 29665
rect 21315 29699 21373 29705
rect 21315 29665 21327 29699
rect 21361 29696 21373 29699
rect 26421 29699 26479 29705
rect 21361 29668 23474 29696
rect 21361 29665 21373 29668
rect 21315 29659 21373 29665
rect 9769 29631 9827 29637
rect 9769 29597 9781 29631
rect 9815 29628 9827 29631
rect 9858 29628 9864 29640
rect 9815 29600 9864 29628
rect 9815 29597 9827 29600
rect 9769 29591 9827 29597
rect 9858 29588 9864 29600
rect 9916 29588 9922 29640
rect 10870 29628 10876 29640
rect 10831 29600 10876 29628
rect 10870 29588 10876 29600
rect 10928 29588 10934 29640
rect 12986 29628 12992 29640
rect 12947 29600 12992 29628
rect 12986 29588 12992 29600
rect 13044 29588 13050 29640
rect 14642 29588 14648 29640
rect 14700 29628 14706 29640
rect 15381 29631 15439 29637
rect 15381 29628 15393 29631
rect 14700 29600 15393 29628
rect 14700 29588 14706 29600
rect 15381 29597 15393 29600
rect 15427 29628 15439 29631
rect 16298 29628 16304 29640
rect 15427 29600 16304 29628
rect 15427 29597 15439 29600
rect 15381 29591 15439 29597
rect 16298 29588 16304 29600
rect 16356 29588 16362 29640
rect 16942 29628 16948 29640
rect 16903 29600 16948 29628
rect 16942 29588 16948 29600
rect 17000 29588 17006 29640
rect 18782 29628 18788 29640
rect 18743 29600 18788 29628
rect 18782 29588 18788 29600
rect 18840 29588 18846 29640
rect 18966 29588 18972 29640
rect 19024 29628 19030 29640
rect 19061 29631 19119 29637
rect 19061 29628 19073 29631
rect 19024 29600 19073 29628
rect 19024 29588 19030 29600
rect 19061 29597 19073 29600
rect 19107 29597 19119 29631
rect 22186 29628 22192 29640
rect 22147 29600 22192 29628
rect 19061 29591 19119 29597
rect 22186 29588 22192 29600
rect 22244 29588 22250 29640
rect 23446 29628 23474 29668
rect 26421 29665 26433 29699
rect 26467 29696 26479 29699
rect 26602 29696 26608 29708
rect 26467 29668 26608 29696
rect 26467 29665 26479 29668
rect 26421 29659 26479 29665
rect 26602 29656 26608 29668
rect 26660 29656 26666 29708
rect 28350 29696 28356 29708
rect 28311 29668 28356 29696
rect 28350 29656 28356 29668
rect 28408 29656 28414 29708
rect 28718 29696 28724 29708
rect 28679 29668 28724 29696
rect 28718 29656 28724 29668
rect 28776 29656 28782 29708
rect 31478 29656 31484 29708
rect 31536 29696 31542 29708
rect 32122 29696 32128 29708
rect 31536 29668 32128 29696
rect 31536 29656 31542 29668
rect 32122 29656 32128 29668
rect 32180 29656 32186 29708
rect 32299 29696 32327 29736
rect 32490 29724 32496 29776
rect 32548 29764 32554 29776
rect 34057 29767 34115 29773
rect 34057 29764 34069 29767
rect 32548 29736 34069 29764
rect 32548 29724 32554 29736
rect 34057 29733 34069 29736
rect 34103 29733 34115 29767
rect 34057 29727 34115 29733
rect 34146 29724 34152 29776
rect 34204 29764 34210 29776
rect 34204 29736 34249 29764
rect 34204 29724 34210 29736
rect 37826 29724 37832 29776
rect 37884 29764 37890 29776
rect 38058 29767 38116 29773
rect 38058 29764 38070 29767
rect 37884 29736 38070 29764
rect 37884 29724 37890 29736
rect 38058 29733 38070 29736
rect 38104 29764 38116 29767
rect 39390 29764 39396 29776
rect 38104 29736 39396 29764
rect 38104 29733 38116 29736
rect 38058 29727 38116 29733
rect 39390 29724 39396 29736
rect 39448 29764 39454 29776
rect 39806 29767 39864 29773
rect 39806 29764 39818 29767
rect 39448 29736 39818 29764
rect 39448 29724 39454 29736
rect 39806 29733 39818 29736
rect 39852 29733 39864 29767
rect 39806 29727 39864 29733
rect 41138 29724 41144 29776
rect 41196 29764 41202 29776
rect 41554 29767 41612 29773
rect 41554 29764 41566 29767
rect 41196 29736 41566 29764
rect 41196 29724 41202 29736
rect 41554 29733 41566 29736
rect 41600 29764 41612 29767
rect 42766 29764 42794 29804
rect 43717 29801 43729 29804
rect 43763 29801 43775 29835
rect 43717 29795 43775 29801
rect 43898 29792 43904 29844
rect 43956 29832 43962 29844
rect 44269 29835 44327 29841
rect 44269 29832 44281 29835
rect 43956 29804 44281 29832
rect 43956 29792 43962 29804
rect 44269 29801 44281 29804
rect 44315 29832 44327 29835
rect 45094 29832 45100 29844
rect 44315 29804 45100 29832
rect 44315 29801 44327 29804
rect 44269 29795 44327 29801
rect 45094 29792 45100 29804
rect 45152 29792 45158 29844
rect 41600 29736 42794 29764
rect 43165 29767 43223 29773
rect 41600 29733 41612 29736
rect 41554 29727 41612 29733
rect 43165 29733 43177 29767
rect 43211 29764 43223 29767
rect 43438 29764 43444 29776
rect 43211 29736 43444 29764
rect 43211 29733 43223 29736
rect 43165 29727 43223 29733
rect 43438 29724 43444 29736
rect 43496 29724 43502 29776
rect 32582 29696 32588 29708
rect 32299 29668 32588 29696
rect 32582 29656 32588 29668
rect 32640 29656 32646 29708
rect 33321 29699 33379 29705
rect 33321 29665 33333 29699
rect 33367 29696 33379 29699
rect 33410 29696 33416 29708
rect 33367 29668 33416 29696
rect 33367 29665 33379 29668
rect 33321 29659 33379 29665
rect 33410 29656 33416 29668
rect 33468 29656 33474 29708
rect 35526 29696 35532 29708
rect 35487 29668 35532 29696
rect 35526 29656 35532 29668
rect 35584 29656 35590 29708
rect 36446 29656 36452 29708
rect 36504 29696 36510 29708
rect 36576 29699 36634 29705
rect 36576 29696 36588 29699
rect 36504 29668 36588 29696
rect 36504 29656 36510 29668
rect 36576 29665 36588 29668
rect 36622 29696 36634 29699
rect 39485 29699 39543 29705
rect 36622 29668 39436 29696
rect 36622 29665 36634 29668
rect 36576 29659 36634 29665
rect 24026 29628 24032 29640
rect 23446 29600 24032 29628
rect 24026 29588 24032 29600
rect 24084 29588 24090 29640
rect 24305 29631 24363 29637
rect 24305 29597 24317 29631
rect 24351 29597 24363 29631
rect 24305 29591 24363 29597
rect 28905 29631 28963 29637
rect 28905 29597 28917 29631
rect 28951 29628 28963 29631
rect 29178 29628 29184 29640
rect 28951 29600 29184 29628
rect 28951 29597 28963 29600
rect 28905 29591 28963 29597
rect 15930 29560 15936 29572
rect 15891 29532 15936 29560
rect 15930 29520 15936 29532
rect 15988 29520 15994 29572
rect 23290 29520 23296 29572
rect 23348 29560 23354 29572
rect 23474 29560 23480 29572
rect 23348 29532 23480 29560
rect 23348 29520 23354 29532
rect 23474 29520 23480 29532
rect 23532 29560 23538 29572
rect 24320 29560 24348 29591
rect 29178 29588 29184 29600
rect 29236 29588 29242 29640
rect 30282 29628 30288 29640
rect 30243 29600 30288 29628
rect 30282 29588 30288 29600
rect 30340 29588 30346 29640
rect 30561 29631 30619 29637
rect 30561 29597 30573 29631
rect 30607 29628 30619 29631
rect 31386 29628 31392 29640
rect 30607 29600 31392 29628
rect 30607 29597 30619 29600
rect 30561 29591 30619 29597
rect 23532 29532 24348 29560
rect 23532 29520 23538 29532
rect 25222 29520 25228 29572
rect 25280 29560 25286 29572
rect 27062 29560 27068 29572
rect 25280 29532 27068 29560
rect 25280 29520 25286 29532
rect 27062 29520 27068 29532
rect 27120 29520 27126 29572
rect 28442 29520 28448 29572
rect 28500 29560 28506 29572
rect 30576 29560 30604 29591
rect 31386 29588 31392 29600
rect 31444 29588 31450 29640
rect 32861 29631 32919 29637
rect 32861 29597 32873 29631
rect 32907 29628 32919 29631
rect 33042 29628 33048 29640
rect 32907 29600 33048 29628
rect 32907 29597 32919 29600
rect 32861 29591 32919 29597
rect 33042 29588 33048 29600
rect 33100 29588 33106 29640
rect 34330 29628 34336 29640
rect 34291 29600 34336 29628
rect 34330 29588 34336 29600
rect 34388 29588 34394 29640
rect 37734 29628 37740 29640
rect 37695 29600 37740 29628
rect 37734 29588 37740 29600
rect 37792 29588 37798 29640
rect 39408 29628 39436 29668
rect 39485 29665 39497 29699
rect 39531 29696 39543 29699
rect 39574 29696 39580 29708
rect 39531 29668 39580 29696
rect 39531 29665 39543 29668
rect 39485 29659 39543 29665
rect 39574 29656 39580 29668
rect 39632 29656 39638 29708
rect 45094 29696 45100 29708
rect 45055 29668 45100 29696
rect 45094 29656 45100 29668
rect 45152 29656 45158 29708
rect 39850 29628 39856 29640
rect 39408 29600 39856 29628
rect 39850 29588 39856 29600
rect 39908 29588 39914 29640
rect 41230 29628 41236 29640
rect 41191 29600 41236 29628
rect 41230 29588 41236 29600
rect 41288 29588 41294 29640
rect 43346 29628 43352 29640
rect 43307 29600 43352 29628
rect 43346 29588 43352 29600
rect 43404 29588 43410 29640
rect 31294 29560 31300 29572
rect 28500 29532 30604 29560
rect 31207 29532 31300 29560
rect 28500 29520 28506 29532
rect 31294 29520 31300 29532
rect 31352 29560 31358 29572
rect 35434 29560 35440 29572
rect 31352 29532 35440 29560
rect 31352 29520 31358 29532
rect 35434 29520 35440 29532
rect 35492 29520 35498 29572
rect 9999 29495 10057 29501
rect 9999 29461 10011 29495
rect 10045 29492 10057 29495
rect 10134 29492 10140 29504
rect 10045 29464 10140 29492
rect 10045 29461 10057 29464
rect 9999 29455 10057 29461
rect 10134 29452 10140 29464
rect 10192 29452 10198 29504
rect 12526 29492 12532 29504
rect 12487 29464 12532 29492
rect 12526 29452 12532 29464
rect 12584 29452 12590 29504
rect 20257 29495 20315 29501
rect 20257 29461 20269 29495
rect 20303 29492 20315 29495
rect 20438 29492 20444 29504
rect 20303 29464 20444 29492
rect 20303 29461 20315 29464
rect 20257 29455 20315 29461
rect 20438 29452 20444 29464
rect 20496 29452 20502 29504
rect 21634 29492 21640 29504
rect 21595 29464 21640 29492
rect 21634 29452 21640 29464
rect 21692 29492 21698 29504
rect 22005 29495 22063 29501
rect 22005 29492 22017 29495
rect 21692 29464 22017 29492
rect 21692 29452 21698 29464
rect 22005 29461 22017 29464
rect 22051 29461 22063 29495
rect 29270 29492 29276 29504
rect 29231 29464 29276 29492
rect 22005 29455 22063 29461
rect 29270 29452 29276 29464
rect 29328 29452 29334 29504
rect 35342 29492 35348 29504
rect 35303 29464 35348 29492
rect 35342 29452 35348 29464
rect 35400 29452 35406 29504
rect 35667 29495 35725 29501
rect 35667 29461 35679 29495
rect 35713 29492 35725 29495
rect 35894 29492 35900 29504
rect 35713 29464 35900 29492
rect 35713 29461 35725 29464
rect 35667 29455 35725 29461
rect 35894 29452 35900 29464
rect 35952 29452 35958 29504
rect 35986 29452 35992 29504
rect 36044 29492 36050 29504
rect 36679 29495 36737 29501
rect 36679 29492 36691 29495
rect 36044 29464 36691 29492
rect 36044 29452 36050 29464
rect 36679 29461 36691 29464
rect 36725 29461 36737 29495
rect 38654 29492 38660 29504
rect 38615 29464 38660 29492
rect 36679 29455 36737 29461
rect 38654 29452 38660 29464
rect 38712 29452 38718 29504
rect 44818 29452 44824 29504
rect 44876 29492 44882 29504
rect 45235 29495 45293 29501
rect 45235 29492 45247 29495
rect 44876 29464 45247 29492
rect 44876 29452 44882 29464
rect 45235 29461 45247 29464
rect 45281 29461 45293 29495
rect 45235 29455 45293 29461
rect 1104 29402 48852 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 48852 29402
rect 1104 29328 48852 29350
rect 10137 29291 10195 29297
rect 10137 29257 10149 29291
rect 10183 29288 10195 29291
rect 10226 29288 10232 29300
rect 10183 29260 10232 29288
rect 10183 29257 10195 29260
rect 10137 29251 10195 29257
rect 10226 29248 10232 29260
rect 10284 29248 10290 29300
rect 12253 29291 12311 29297
rect 12253 29257 12265 29291
rect 12299 29288 12311 29291
rect 12434 29288 12440 29300
rect 12299 29260 12440 29288
rect 12299 29257 12311 29260
rect 12253 29251 12311 29257
rect 12434 29248 12440 29260
rect 12492 29248 12498 29300
rect 13446 29288 13452 29300
rect 13407 29260 13452 29288
rect 13446 29248 13452 29260
rect 13504 29248 13510 29300
rect 14642 29288 14648 29300
rect 14603 29260 14648 29288
rect 14642 29248 14648 29260
rect 14700 29248 14706 29300
rect 15470 29248 15476 29300
rect 15528 29288 15534 29300
rect 15565 29291 15623 29297
rect 15565 29288 15577 29291
rect 15528 29260 15577 29288
rect 15528 29248 15534 29260
rect 15565 29257 15577 29260
rect 15611 29257 15623 29291
rect 15565 29251 15623 29257
rect 18414 29248 18420 29300
rect 18472 29288 18478 29300
rect 18509 29291 18567 29297
rect 18509 29288 18521 29291
rect 18472 29260 18521 29288
rect 18472 29248 18478 29260
rect 18509 29257 18521 29260
rect 18555 29257 18567 29291
rect 18874 29288 18880 29300
rect 18835 29260 18880 29288
rect 18509 29251 18567 29257
rect 18874 29248 18880 29260
rect 18932 29248 18938 29300
rect 19150 29248 19156 29300
rect 19208 29288 19214 29300
rect 19613 29291 19671 29297
rect 19613 29288 19625 29291
rect 19208 29260 19625 29288
rect 19208 29248 19214 29260
rect 19613 29257 19625 29260
rect 19659 29288 19671 29291
rect 20303 29291 20361 29297
rect 20303 29288 20315 29291
rect 19659 29260 20315 29288
rect 19659 29257 19671 29260
rect 19613 29251 19671 29257
rect 20303 29257 20315 29260
rect 20349 29288 20361 29291
rect 22557 29291 22615 29297
rect 22557 29288 22569 29291
rect 20349 29260 22569 29288
rect 20349 29257 20361 29260
rect 20303 29251 20361 29257
rect 22557 29257 22569 29260
rect 22603 29257 22615 29291
rect 22557 29251 22615 29257
rect 24026 29248 24032 29300
rect 24084 29288 24090 29300
rect 24305 29291 24363 29297
rect 24305 29288 24317 29291
rect 24084 29260 24317 29288
rect 24084 29248 24090 29260
rect 24305 29257 24317 29260
rect 24351 29257 24363 29291
rect 24305 29251 24363 29257
rect 28261 29291 28319 29297
rect 28261 29257 28273 29291
rect 28307 29288 28319 29291
rect 28350 29288 28356 29300
rect 28307 29260 28356 29288
rect 28307 29257 28319 29260
rect 28261 29251 28319 29257
rect 28350 29248 28356 29260
rect 28408 29248 28414 29300
rect 28629 29291 28687 29297
rect 28629 29257 28641 29291
rect 28675 29288 28687 29291
rect 28718 29288 28724 29300
rect 28675 29260 28724 29288
rect 28675 29257 28687 29260
rect 28629 29251 28687 29257
rect 28718 29248 28724 29260
rect 28776 29248 28782 29300
rect 32582 29288 32588 29300
rect 32543 29260 32588 29288
rect 32582 29248 32588 29260
rect 32640 29248 32646 29300
rect 34057 29291 34115 29297
rect 34057 29257 34069 29291
rect 34103 29288 34115 29291
rect 34146 29288 34152 29300
rect 34103 29260 34152 29288
rect 34103 29257 34115 29260
rect 34057 29251 34115 29257
rect 34146 29248 34152 29260
rect 34204 29288 34210 29300
rect 34609 29291 34667 29297
rect 34609 29288 34621 29291
rect 34204 29260 34621 29288
rect 34204 29248 34210 29260
rect 34609 29257 34621 29260
rect 34655 29257 34667 29291
rect 34609 29251 34667 29257
rect 36722 29248 36728 29300
rect 36780 29288 36786 29300
rect 40221 29291 40279 29297
rect 40221 29288 40233 29291
rect 36780 29260 40233 29288
rect 36780 29248 36786 29260
rect 40221 29257 40233 29260
rect 40267 29257 40279 29291
rect 44818 29288 44824 29300
rect 44779 29260 44824 29288
rect 40221 29251 40279 29257
rect 11330 29220 11336 29232
rect 11243 29192 11336 29220
rect 11330 29180 11336 29192
rect 11388 29220 11394 29232
rect 13464 29220 13492 29248
rect 11388 29192 13492 29220
rect 11388 29180 11394 29192
rect 18782 29180 18788 29232
rect 18840 29220 18846 29232
rect 19245 29223 19303 29229
rect 19245 29220 19257 29223
rect 18840 29192 19257 29220
rect 18840 29180 18846 29192
rect 19245 29189 19257 29192
rect 19291 29189 19303 29223
rect 20438 29220 20444 29232
rect 20399 29192 20444 29220
rect 19245 29183 19303 29189
rect 20438 29180 20444 29192
rect 20496 29220 20502 29232
rect 20496 29192 27108 29220
rect 20496 29180 20502 29192
rect 10870 29112 10876 29164
rect 10928 29152 10934 29164
rect 10965 29155 11023 29161
rect 10965 29152 10977 29155
rect 10928 29124 10977 29152
rect 10928 29112 10934 29124
rect 10965 29121 10977 29124
rect 11011 29152 11023 29155
rect 11609 29155 11667 29161
rect 11609 29152 11621 29155
rect 11011 29124 11621 29152
rect 11011 29121 11023 29124
rect 10965 29115 11023 29121
rect 11609 29121 11621 29124
rect 11655 29121 11667 29155
rect 12986 29152 12992 29164
rect 12947 29124 12992 29152
rect 11609 29115 11667 29121
rect 12986 29112 12992 29124
rect 13044 29152 13050 29164
rect 13817 29155 13875 29161
rect 13817 29152 13829 29155
rect 13044 29124 13829 29152
rect 13044 29112 13050 29124
rect 13817 29121 13829 29124
rect 13863 29121 13875 29155
rect 13817 29115 13875 29121
rect 16942 29112 16948 29164
rect 17000 29152 17006 29164
rect 17129 29155 17187 29161
rect 17129 29152 17141 29155
rect 17000 29124 17141 29152
rect 17000 29112 17006 29124
rect 17129 29121 17141 29124
rect 17175 29152 17187 29155
rect 17773 29155 17831 29161
rect 17773 29152 17785 29155
rect 17175 29124 17785 29152
rect 17175 29121 17187 29124
rect 17129 29115 17187 29121
rect 17773 29121 17785 29124
rect 17819 29121 17831 29155
rect 17773 29115 17831 29121
rect 18690 29112 18696 29164
rect 18748 29152 18754 29164
rect 19978 29152 19984 29164
rect 18748 29124 19984 29152
rect 18748 29112 18754 29124
rect 19978 29112 19984 29124
rect 20036 29152 20042 29164
rect 20533 29155 20591 29161
rect 20533 29152 20545 29155
rect 20036 29124 20545 29152
rect 20036 29112 20042 29124
rect 20533 29121 20545 29124
rect 20579 29152 20591 29155
rect 20898 29152 20904 29164
rect 20579 29124 20904 29152
rect 20579 29121 20591 29124
rect 20533 29115 20591 29121
rect 20898 29112 20904 29124
rect 20956 29112 20962 29164
rect 21082 29112 21088 29164
rect 21140 29152 21146 29164
rect 21177 29155 21235 29161
rect 21177 29152 21189 29155
rect 21140 29124 21189 29152
rect 21140 29112 21146 29124
rect 21177 29121 21189 29124
rect 21223 29121 21235 29155
rect 21177 29115 21235 29121
rect 22462 29112 22468 29164
rect 22520 29152 22526 29164
rect 22741 29155 22799 29161
rect 22741 29152 22753 29155
rect 22520 29124 22753 29152
rect 22520 29112 22526 29124
rect 22741 29121 22753 29124
rect 22787 29121 22799 29155
rect 22741 29115 22799 29121
rect 24029 29155 24087 29161
rect 24029 29121 24041 29155
rect 24075 29152 24087 29155
rect 24118 29152 24124 29164
rect 24075 29124 24124 29152
rect 24075 29121 24087 29124
rect 24029 29115 24087 29121
rect 24118 29112 24124 29124
rect 24176 29112 24182 29164
rect 26050 29152 26056 29164
rect 26011 29124 26056 29152
rect 26050 29112 26056 29124
rect 26108 29112 26114 29164
rect 27080 29161 27108 29192
rect 32766 29180 32772 29232
rect 32824 29220 32830 29232
rect 33502 29220 33508 29232
rect 32824 29192 33508 29220
rect 32824 29180 32830 29192
rect 33502 29180 33508 29192
rect 33560 29180 33566 29232
rect 39853 29223 39911 29229
rect 39853 29220 39865 29223
rect 37108 29192 39865 29220
rect 27065 29155 27123 29161
rect 27065 29121 27077 29155
rect 27111 29152 27123 29155
rect 27614 29152 27620 29164
rect 27111 29124 27620 29152
rect 27111 29121 27123 29124
rect 27065 29115 27123 29121
rect 27614 29112 27620 29124
rect 27672 29112 27678 29164
rect 30558 29112 30564 29164
rect 30616 29152 30622 29164
rect 31113 29155 31171 29161
rect 31113 29152 31125 29155
rect 30616 29124 31125 29152
rect 30616 29112 30622 29124
rect 31113 29121 31125 29124
rect 31159 29152 31171 29155
rect 31294 29152 31300 29164
rect 31159 29124 31300 29152
rect 31159 29121 31171 29124
rect 31113 29115 31171 29121
rect 31294 29112 31300 29124
rect 31352 29112 31358 29164
rect 31386 29112 31392 29164
rect 31444 29152 31450 29164
rect 31444 29124 31892 29152
rect 31444 29112 31450 29124
rect 10226 29084 10232 29096
rect 10187 29056 10232 29084
rect 10226 29044 10232 29056
rect 10284 29044 10290 29096
rect 10781 29087 10839 29093
rect 10781 29053 10793 29087
rect 10827 29053 10839 29087
rect 12434 29084 12440 29096
rect 12395 29056 12440 29084
rect 10781 29047 10839 29053
rect 9490 28976 9496 29028
rect 9548 29016 9554 29028
rect 9769 29019 9827 29025
rect 9769 29016 9781 29019
rect 9548 28988 9781 29016
rect 9548 28976 9554 28988
rect 9769 28985 9781 28988
rect 9815 29016 9827 29019
rect 10686 29016 10692 29028
rect 9815 28988 10692 29016
rect 9815 28985 9827 28988
rect 9769 28979 9827 28985
rect 10686 28976 10692 28988
rect 10744 29016 10750 29028
rect 10796 29016 10824 29047
rect 12434 29044 12440 29056
rect 12492 29044 12498 29096
rect 12526 29044 12532 29096
rect 12584 29084 12590 29096
rect 12897 29087 12955 29093
rect 12897 29084 12909 29087
rect 12584 29056 12909 29084
rect 12584 29044 12590 29056
rect 12897 29053 12909 29056
rect 12943 29084 12955 29087
rect 12943 29056 13814 29084
rect 12943 29053 12955 29056
rect 12897 29047 12955 29053
rect 12544 29016 12572 29044
rect 10744 28988 12572 29016
rect 13786 29016 13814 29056
rect 14458 29044 14464 29096
rect 14516 29084 14522 29096
rect 14772 29087 14830 29093
rect 14772 29084 14784 29087
rect 14516 29056 14784 29084
rect 14516 29044 14522 29056
rect 14772 29053 14784 29056
rect 14818 29084 14830 29087
rect 14918 29084 14924 29096
rect 14818 29056 14924 29084
rect 14818 29053 14830 29056
rect 14772 29047 14830 29053
rect 14918 29044 14924 29056
rect 14976 29084 14982 29096
rect 15197 29087 15255 29093
rect 15197 29084 15209 29087
rect 14976 29056 15209 29084
rect 14976 29044 14982 29056
rect 15197 29053 15209 29056
rect 15243 29053 15255 29087
rect 16206 29084 16212 29096
rect 16167 29056 16212 29084
rect 15197 29047 15255 29053
rect 16206 29044 16212 29056
rect 16264 29084 16270 29096
rect 16393 29087 16451 29093
rect 16393 29084 16405 29087
rect 16264 29056 16405 29084
rect 16264 29044 16270 29056
rect 16393 29053 16405 29056
rect 16439 29084 16451 29087
rect 16574 29084 16580 29096
rect 16439 29056 16580 29084
rect 16439 29053 16451 29056
rect 16393 29047 16451 29053
rect 16574 29044 16580 29056
rect 16632 29044 16638 29096
rect 16853 29087 16911 29093
rect 16853 29053 16865 29087
rect 16899 29053 16911 29087
rect 16853 29047 16911 29053
rect 18116 29087 18174 29093
rect 18116 29053 18128 29087
rect 18162 29084 18174 29087
rect 18414 29084 18420 29096
rect 18162 29056 18420 29084
rect 18162 29053 18174 29056
rect 18116 29047 18174 29053
rect 16298 29016 16304 29028
rect 13786 28988 16304 29016
rect 10744 28976 10750 28988
rect 16298 28976 16304 28988
rect 16356 29016 16362 29028
rect 16868 29016 16896 29047
rect 18414 29044 18420 29056
rect 18472 29044 18478 29096
rect 21542 29044 21548 29096
rect 21600 29084 21606 29096
rect 21729 29087 21787 29093
rect 21729 29084 21741 29087
rect 21600 29056 21741 29084
rect 21600 29044 21606 29056
rect 21729 29053 21741 29056
rect 21775 29053 21787 29087
rect 21729 29047 21787 29053
rect 22189 29087 22247 29093
rect 22189 29053 22201 29087
rect 22235 29053 22247 29087
rect 22189 29047 22247 29053
rect 16356 28988 16896 29016
rect 16356 28976 16362 28988
rect 17310 28976 17316 29028
rect 17368 29016 17374 29028
rect 17405 29019 17463 29025
rect 17405 29016 17417 29019
rect 17368 28988 17417 29016
rect 17368 28976 17374 28988
rect 17405 28985 17417 28988
rect 17451 29016 17463 29019
rect 18506 29016 18512 29028
rect 17451 28988 18512 29016
rect 17451 28985 17463 28988
rect 17405 28979 17463 28985
rect 18506 28976 18512 28988
rect 18564 28976 18570 29028
rect 20165 29019 20223 29025
rect 20165 28985 20177 29019
rect 20211 29016 20223 29019
rect 20346 29016 20352 29028
rect 20211 28988 20352 29016
rect 20211 28985 20223 28988
rect 20165 28979 20223 28985
rect 20346 28976 20352 28988
rect 20404 28976 20410 29028
rect 20898 29016 20904 29028
rect 20859 28988 20904 29016
rect 20898 28976 20904 28988
rect 20956 29016 20962 29028
rect 21634 29016 21640 29028
rect 20956 28988 21640 29016
rect 20956 28976 20962 28988
rect 21634 28976 21640 28988
rect 21692 29016 21698 29028
rect 22204 29016 22232 29047
rect 26234 29044 26240 29096
rect 26292 29084 26298 29096
rect 26973 29087 27031 29093
rect 26973 29084 26985 29087
rect 26292 29056 26985 29084
rect 26292 29044 26298 29056
rect 26973 29053 26985 29056
rect 27019 29084 27031 29087
rect 27709 29087 27767 29093
rect 27709 29084 27721 29087
rect 27019 29056 27721 29084
rect 27019 29053 27031 29056
rect 26973 29047 27031 29053
rect 27709 29053 27721 29056
rect 27755 29084 27767 29087
rect 27798 29084 27804 29096
rect 27755 29056 27804 29084
rect 27755 29053 27767 29056
rect 27709 29047 27767 29053
rect 27798 29044 27804 29056
rect 27856 29044 27862 29096
rect 28902 29044 28908 29096
rect 28960 29084 28966 29096
rect 29270 29084 29276 29096
rect 28960 29056 29276 29084
rect 28960 29044 28966 29056
rect 29270 29044 29276 29056
rect 29328 29044 29334 29096
rect 30193 29087 30251 29093
rect 30193 29053 30205 29087
rect 30239 29084 30251 29087
rect 30837 29087 30895 29093
rect 30837 29084 30849 29087
rect 30239 29056 30849 29084
rect 30239 29053 30251 29056
rect 30193 29047 30251 29053
rect 30837 29053 30849 29056
rect 30883 29053 30895 29087
rect 30837 29047 30895 29053
rect 21692 28988 22232 29016
rect 22557 29019 22615 29025
rect 21692 28976 21698 28988
rect 22557 28985 22569 29019
rect 22603 29016 22615 29019
rect 25222 29016 25228 29028
rect 22603 28988 25228 29016
rect 22603 28985 22615 28988
rect 22557 28979 22615 28985
rect 25222 28976 25228 28988
rect 25280 28976 25286 29028
rect 25593 29019 25651 29025
rect 25593 29016 25605 29019
rect 25332 28988 25605 29016
rect 14875 28951 14933 28957
rect 14875 28917 14887 28951
rect 14921 28948 14933 28951
rect 15010 28948 15016 28960
rect 14921 28920 15016 28948
rect 14921 28917 14933 28920
rect 14875 28911 14933 28917
rect 15010 28908 15016 28920
rect 15068 28908 15074 28960
rect 17494 28908 17500 28960
rect 17552 28948 17558 28960
rect 18187 28951 18245 28957
rect 18187 28948 18199 28951
rect 17552 28920 18199 28948
rect 17552 28908 17558 28920
rect 18187 28917 18199 28920
rect 18233 28917 18245 28951
rect 21542 28948 21548 28960
rect 21503 28920 21548 28948
rect 18187 28911 18245 28917
rect 21542 28908 21548 28920
rect 21600 28908 21606 28960
rect 21818 28948 21824 28960
rect 21779 28920 21824 28948
rect 21818 28908 21824 28920
rect 21876 28908 21882 28960
rect 25332 28957 25360 28988
rect 25593 28985 25605 28988
rect 25639 28985 25651 29019
rect 25593 28979 25651 28985
rect 25685 29019 25743 29025
rect 25685 28985 25697 29019
rect 25731 28985 25743 29019
rect 26602 29016 26608 29028
rect 26563 28988 26608 29016
rect 25685 28979 25743 28985
rect 24489 28951 24547 28957
rect 24489 28917 24501 28951
rect 24535 28948 24547 28951
rect 25317 28951 25375 28957
rect 25317 28948 25329 28951
rect 24535 28920 25329 28948
rect 24535 28917 24547 28920
rect 24489 28911 24547 28917
rect 25317 28917 25329 28920
rect 25363 28917 25375 28951
rect 25317 28911 25375 28917
rect 25406 28908 25412 28960
rect 25464 28948 25470 28960
rect 25700 28948 25728 28979
rect 26602 28976 26608 28988
rect 26660 28976 26666 29028
rect 29594 29019 29652 29025
rect 29594 29016 29606 29019
rect 29012 28988 29606 29016
rect 29012 28960 29040 28988
rect 29594 28985 29606 28988
rect 29640 28985 29652 29019
rect 29594 28979 29652 28985
rect 28994 28948 29000 28960
rect 25464 28920 25728 28948
rect 28955 28920 29000 28948
rect 25464 28908 25470 28920
rect 28994 28908 29000 28920
rect 29052 28908 29058 28960
rect 30190 28908 30196 28960
rect 30248 28948 30254 28960
rect 30374 28948 30380 28960
rect 30248 28920 30380 28948
rect 30248 28908 30254 28920
rect 30374 28908 30380 28920
rect 30432 28948 30438 28960
rect 30469 28951 30527 28957
rect 30469 28948 30481 28951
rect 30432 28920 30481 28948
rect 30432 28908 30438 28920
rect 30469 28917 30481 28920
rect 30515 28917 30527 28951
rect 30852 28948 30880 29047
rect 31205 29019 31263 29025
rect 31205 28985 31217 29019
rect 31251 28985 31263 29019
rect 31864 29016 31892 29124
rect 31938 29112 31944 29164
rect 31996 29152 32002 29164
rect 32861 29155 32919 29161
rect 32861 29152 32873 29155
rect 31996 29124 32873 29152
rect 31996 29112 32002 29124
rect 32861 29121 32873 29124
rect 32907 29152 32919 29155
rect 32950 29152 32956 29164
rect 32907 29124 32956 29152
rect 32907 29121 32919 29124
rect 32861 29115 32919 29121
rect 32950 29112 32956 29124
rect 33008 29112 33014 29164
rect 34977 29155 35035 29161
rect 34977 29121 34989 29155
rect 35023 29152 35035 29155
rect 35342 29152 35348 29164
rect 35023 29124 35348 29152
rect 35023 29121 35035 29124
rect 34977 29115 35035 29121
rect 35342 29112 35348 29124
rect 35400 29112 35406 29164
rect 35434 29112 35440 29164
rect 35492 29152 35498 29164
rect 35492 29124 35537 29152
rect 35492 29112 35498 29124
rect 36630 29084 36636 29096
rect 36591 29056 36636 29084
rect 36630 29044 36636 29056
rect 36688 29044 36694 29096
rect 36814 29044 36820 29096
rect 36872 29084 36878 29096
rect 37108 29093 37136 29192
rect 39853 29189 39865 29192
rect 39899 29189 39911 29223
rect 39853 29183 39911 29189
rect 37369 29155 37427 29161
rect 37369 29121 37381 29155
rect 37415 29152 37427 29155
rect 37734 29152 37740 29164
rect 37415 29124 37740 29152
rect 37415 29121 37427 29124
rect 37369 29115 37427 29121
rect 37734 29112 37740 29124
rect 37792 29112 37798 29164
rect 37826 29112 37832 29164
rect 37884 29152 37890 29164
rect 38562 29152 38568 29164
rect 37884 29124 37929 29152
rect 38523 29124 38568 29152
rect 37884 29112 37890 29124
rect 38562 29112 38568 29124
rect 38620 29112 38626 29164
rect 39390 29112 39396 29164
rect 39448 29152 39454 29164
rect 39485 29155 39543 29161
rect 39485 29152 39497 29155
rect 39448 29124 39497 29152
rect 39448 29112 39454 29124
rect 39485 29121 39497 29124
rect 39531 29121 39543 29155
rect 39485 29115 39543 29121
rect 37093 29087 37151 29093
rect 37093 29084 37105 29087
rect 36872 29056 37105 29084
rect 36872 29044 36878 29056
rect 37093 29053 37105 29056
rect 37139 29053 37151 29087
rect 37093 29047 37151 29053
rect 31864 28988 32628 29016
rect 31205 28979 31263 28985
rect 31220 28948 31248 28979
rect 32122 28948 32128 28960
rect 30852 28920 31248 28948
rect 32083 28920 32128 28948
rect 30469 28911 30527 28917
rect 32122 28908 32128 28920
rect 32180 28908 32186 28960
rect 32600 28948 32628 28988
rect 32950 28976 32956 29028
rect 33008 29016 33014 29028
rect 33505 29019 33563 29025
rect 33505 29016 33517 29019
rect 33008 28988 33053 29016
rect 33106 28988 33517 29016
rect 33008 28976 33014 28988
rect 33106 28948 33134 28988
rect 33505 28985 33517 28988
rect 33551 28985 33563 29019
rect 33505 28979 33563 28985
rect 35066 28976 35072 29028
rect 35124 29016 35130 29028
rect 35124 28988 35169 29016
rect 35124 28976 35130 28988
rect 35434 28976 35440 29028
rect 35492 29016 35498 29028
rect 36446 29016 36452 29028
rect 35492 28988 36452 29016
rect 35492 28976 35498 28988
rect 36446 28976 36452 28988
rect 36504 28976 36510 29028
rect 38286 29016 38292 29028
rect 38247 28988 38292 29016
rect 38286 28976 38292 28988
rect 38344 28976 38350 29028
rect 38381 29019 38439 29025
rect 38381 28985 38393 29019
rect 38427 29016 38439 29019
rect 38654 29016 38660 29028
rect 38427 28988 38660 29016
rect 38427 28985 38439 28988
rect 38381 28979 38439 28985
rect 38654 28976 38660 28988
rect 38712 28976 38718 29028
rect 35526 28948 35532 28960
rect 32600 28920 33134 28948
rect 35439 28920 35532 28948
rect 35526 28908 35532 28920
rect 35584 28948 35590 28960
rect 35897 28951 35955 28957
rect 35897 28948 35909 28951
rect 35584 28920 35909 28948
rect 35584 28908 35590 28920
rect 35897 28917 35909 28920
rect 35943 28917 35955 28951
rect 39500 28948 39528 29115
rect 39868 29016 39896 29183
rect 40236 29084 40264 29251
rect 44818 29248 44824 29260
rect 44876 29248 44882 29300
rect 42978 29180 42984 29232
rect 43036 29220 43042 29232
rect 44361 29223 44419 29229
rect 44361 29220 44373 29223
rect 43036 29192 44373 29220
rect 43036 29180 43042 29192
rect 44361 29189 44373 29192
rect 44407 29189 44419 29223
rect 44361 29183 44419 29189
rect 42426 29152 42432 29164
rect 40972 29124 42432 29152
rect 40972 29093 41000 29124
rect 42426 29112 42432 29124
rect 42484 29152 42490 29164
rect 42702 29152 42708 29164
rect 42484 29124 42564 29152
rect 42663 29124 42708 29152
rect 42484 29112 42490 29124
rect 40497 29087 40555 29093
rect 40497 29084 40509 29087
rect 40236 29056 40509 29084
rect 40497 29053 40509 29056
rect 40543 29053 40555 29087
rect 40497 29047 40555 29053
rect 40957 29087 41015 29093
rect 40957 29053 40969 29087
rect 41003 29053 41015 29087
rect 40957 29047 41015 29053
rect 40972 29016 41000 29047
rect 41046 29044 41052 29096
rect 41104 29084 41110 29096
rect 42536 29093 42564 29124
rect 42702 29112 42708 29124
rect 42760 29112 42766 29164
rect 42797 29155 42855 29161
rect 42797 29121 42809 29155
rect 42843 29152 42855 29155
rect 43346 29152 43352 29164
rect 42843 29124 43352 29152
rect 42843 29121 42855 29124
rect 42797 29115 42855 29121
rect 43346 29112 43352 29124
rect 43404 29112 43410 29164
rect 43809 29155 43867 29161
rect 43809 29121 43821 29155
rect 43855 29152 43867 29155
rect 44836 29152 44864 29248
rect 43855 29124 44864 29152
rect 43855 29121 43867 29124
rect 43809 29115 43867 29121
rect 41969 29087 42027 29093
rect 41969 29084 41981 29087
rect 41104 29056 41981 29084
rect 41104 29044 41110 29056
rect 41969 29053 41981 29056
rect 42015 29084 42027 29087
rect 42061 29087 42119 29093
rect 42061 29084 42073 29087
rect 42015 29056 42073 29084
rect 42015 29053 42027 29056
rect 41969 29047 42027 29053
rect 42061 29053 42073 29056
rect 42107 29053 42119 29087
rect 42061 29047 42119 29053
rect 42521 29087 42579 29093
rect 42521 29053 42533 29087
rect 42567 29053 42579 29087
rect 42521 29047 42579 29053
rect 41230 29016 41236 29028
rect 39868 28988 41000 29016
rect 41191 28988 41236 29016
rect 41230 28976 41236 28988
rect 41288 28976 41294 29028
rect 43898 29016 43904 29028
rect 43859 28988 43904 29016
rect 43898 28976 43904 28988
rect 43956 28976 43962 29028
rect 41138 28948 41144 28960
rect 39500 28920 41144 28948
rect 35897 28911 35955 28917
rect 41138 28908 41144 28920
rect 41196 28948 41202 28960
rect 41509 28951 41567 28957
rect 41509 28948 41521 28951
rect 41196 28920 41521 28948
rect 41196 28908 41202 28920
rect 41509 28917 41521 28920
rect 41555 28917 41567 28951
rect 43346 28948 43352 28960
rect 43307 28920 43352 28948
rect 41509 28911 41567 28917
rect 43346 28908 43352 28920
rect 43404 28908 43410 28960
rect 44358 28908 44364 28960
rect 44416 28948 44422 28960
rect 45094 28948 45100 28960
rect 44416 28920 45100 28948
rect 44416 28908 44422 28920
rect 45094 28908 45100 28920
rect 45152 28908 45158 28960
rect 1104 28858 48852 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 48852 28858
rect 1104 28784 48852 28806
rect 9858 28744 9864 28756
rect 9819 28716 9864 28744
rect 9858 28704 9864 28716
rect 9916 28704 9922 28756
rect 15010 28744 15016 28756
rect 14971 28716 15016 28744
rect 15010 28704 15016 28716
rect 15068 28744 15074 28756
rect 15068 28716 15424 28744
rect 15068 28704 15074 28716
rect 12158 28676 12164 28688
rect 12119 28648 12164 28676
rect 12158 28636 12164 28648
rect 12216 28636 12222 28688
rect 15396 28685 15424 28716
rect 16298 28704 16304 28756
rect 16356 28744 16362 28756
rect 16393 28747 16451 28753
rect 16393 28744 16405 28747
rect 16356 28716 16405 28744
rect 16356 28704 16362 28716
rect 16393 28713 16405 28716
rect 16439 28713 16451 28747
rect 16393 28707 16451 28713
rect 21450 28704 21456 28756
rect 21508 28744 21514 28756
rect 21545 28747 21603 28753
rect 21545 28744 21557 28747
rect 21508 28716 21557 28744
rect 21508 28704 21514 28716
rect 21545 28713 21557 28716
rect 21591 28713 21603 28747
rect 21545 28707 21603 28713
rect 15381 28679 15439 28685
rect 15381 28645 15393 28679
rect 15427 28645 15439 28679
rect 15381 28639 15439 28645
rect 15470 28636 15476 28688
rect 15528 28676 15534 28688
rect 15528 28648 15573 28676
rect 15528 28636 15534 28648
rect 17218 28636 17224 28688
rect 17276 28676 17282 28688
rect 17313 28679 17371 28685
rect 17313 28676 17325 28679
rect 17276 28648 17325 28676
rect 17276 28636 17282 28648
rect 17313 28645 17325 28648
rect 17359 28645 17371 28679
rect 21560 28676 21588 28707
rect 22186 28704 22192 28756
rect 22244 28744 22250 28756
rect 22373 28747 22431 28753
rect 22373 28744 22385 28747
rect 22244 28716 22385 28744
rect 22244 28704 22250 28716
rect 22373 28713 22385 28716
rect 22419 28713 22431 28747
rect 22373 28707 22431 28713
rect 29178 28704 29184 28756
rect 29236 28744 29242 28756
rect 29273 28747 29331 28753
rect 29273 28744 29285 28747
rect 29236 28716 29285 28744
rect 29236 28704 29242 28716
rect 29273 28713 29285 28716
rect 29319 28713 29331 28747
rect 30098 28744 30104 28756
rect 30059 28716 30104 28744
rect 29273 28707 29331 28713
rect 30098 28704 30104 28716
rect 30156 28704 30162 28756
rect 30653 28747 30711 28753
rect 30653 28713 30665 28747
rect 30699 28744 30711 28747
rect 30926 28744 30932 28756
rect 30699 28716 30932 28744
rect 30699 28713 30711 28716
rect 30653 28707 30711 28713
rect 30926 28704 30932 28716
rect 30984 28704 30990 28756
rect 31294 28744 31300 28756
rect 31255 28716 31300 28744
rect 31294 28704 31300 28716
rect 31352 28704 31358 28756
rect 31938 28744 31944 28756
rect 31899 28716 31944 28744
rect 31938 28704 31944 28716
rect 31996 28704 32002 28756
rect 33410 28744 33416 28756
rect 33371 28716 33416 28744
rect 33410 28704 33416 28716
rect 33468 28704 33474 28756
rect 33965 28747 34023 28753
rect 33965 28713 33977 28747
rect 34011 28744 34023 28747
rect 34146 28744 34152 28756
rect 34011 28716 34152 28744
rect 34011 28713 34023 28716
rect 33965 28707 34023 28713
rect 34146 28704 34152 28716
rect 34204 28744 34210 28756
rect 35066 28744 35072 28756
rect 34204 28716 35072 28744
rect 34204 28704 34210 28716
rect 22462 28676 22468 28688
rect 21560 28648 22468 28676
rect 17313 28639 17371 28645
rect 22462 28636 22468 28648
rect 22520 28636 22526 28688
rect 23106 28676 23112 28688
rect 22566 28648 23112 28676
rect 10318 28608 10324 28620
rect 10279 28580 10324 28608
rect 10318 28568 10324 28580
rect 10376 28568 10382 28620
rect 10594 28568 10600 28620
rect 10652 28608 10658 28620
rect 10781 28611 10839 28617
rect 10781 28608 10793 28611
rect 10652 28580 10793 28608
rect 10652 28568 10658 28580
rect 10781 28577 10793 28580
rect 10827 28577 10839 28611
rect 10781 28571 10839 28577
rect 14185 28611 14243 28617
rect 14185 28577 14197 28611
rect 14231 28608 14243 28611
rect 14274 28608 14280 28620
rect 14231 28580 14280 28608
rect 14231 28577 14243 28580
rect 14185 28571 14243 28577
rect 14274 28568 14280 28580
rect 14332 28568 14338 28620
rect 17954 28568 17960 28620
rect 18012 28608 18018 28620
rect 18598 28608 18604 28620
rect 18012 28580 18604 28608
rect 18012 28568 18018 28580
rect 18598 28568 18604 28580
rect 18656 28608 18662 28620
rect 18728 28611 18786 28617
rect 18728 28608 18740 28611
rect 18656 28580 18740 28608
rect 18656 28568 18662 28580
rect 18728 28577 18740 28580
rect 18774 28577 18786 28611
rect 18728 28571 18786 28577
rect 22097 28611 22155 28617
rect 22097 28577 22109 28611
rect 22143 28608 22155 28611
rect 22566 28608 22594 28648
rect 23106 28636 23112 28648
rect 23164 28636 23170 28688
rect 25038 28676 25044 28688
rect 24999 28648 25044 28676
rect 25038 28636 25044 28648
rect 25096 28636 25102 28688
rect 25590 28676 25596 28688
rect 25551 28648 25596 28676
rect 25590 28636 25596 28648
rect 25648 28636 25654 28688
rect 26694 28676 26700 28688
rect 26655 28648 26700 28676
rect 26694 28636 26700 28648
rect 26752 28636 26758 28688
rect 28902 28676 28908 28688
rect 28863 28648 28908 28676
rect 28902 28636 28908 28648
rect 28960 28636 28966 28688
rect 32490 28636 32496 28688
rect 32548 28676 32554 28688
rect 34992 28685 35020 28716
rect 35066 28704 35072 28716
rect 35124 28704 35130 28756
rect 36814 28704 36820 28756
rect 36872 28744 36878 28756
rect 37093 28747 37151 28753
rect 37093 28744 37105 28747
rect 36872 28716 37105 28744
rect 36872 28704 36878 28716
rect 37093 28713 37105 28716
rect 37139 28713 37151 28747
rect 37093 28707 37151 28713
rect 37553 28747 37611 28753
rect 37553 28713 37565 28747
rect 37599 28744 37611 28747
rect 37734 28744 37740 28756
rect 37599 28716 37740 28744
rect 37599 28713 37611 28716
rect 37553 28707 37611 28713
rect 37734 28704 37740 28716
rect 37792 28704 37798 28756
rect 38473 28747 38531 28753
rect 38473 28713 38485 28747
rect 38519 28744 38531 28747
rect 38654 28744 38660 28756
rect 38519 28716 38660 28744
rect 38519 28713 38531 28716
rect 38473 28707 38531 28713
rect 38654 28704 38660 28716
rect 38712 28704 38718 28756
rect 39574 28744 39580 28756
rect 39535 28716 39580 28744
rect 39574 28704 39580 28716
rect 39632 28704 39638 28756
rect 41230 28704 41236 28756
rect 41288 28744 41294 28756
rect 41325 28747 41383 28753
rect 41325 28744 41337 28747
rect 41288 28716 41337 28744
rect 41288 28704 41294 28716
rect 41325 28713 41337 28716
rect 41371 28713 41383 28747
rect 42426 28744 42432 28756
rect 42387 28716 42432 28744
rect 41325 28707 41383 28713
rect 42426 28704 42432 28716
rect 42484 28704 42490 28756
rect 43898 28744 43904 28756
rect 43859 28716 43904 28744
rect 43898 28704 43904 28716
rect 43956 28704 43962 28756
rect 34241 28679 34299 28685
rect 34241 28676 34253 28679
rect 32548 28648 34253 28676
rect 32548 28636 32554 28648
rect 34241 28645 34253 28648
rect 34287 28645 34299 28679
rect 34241 28639 34299 28645
rect 34977 28679 35035 28685
rect 34977 28645 34989 28679
rect 35023 28645 35035 28679
rect 34977 28639 35035 28645
rect 35250 28636 35256 28688
rect 35308 28676 35314 28688
rect 35529 28679 35587 28685
rect 35529 28676 35541 28679
rect 35308 28648 35541 28676
rect 35308 28636 35314 28648
rect 35529 28645 35541 28648
rect 35575 28645 35587 28679
rect 35529 28639 35587 28645
rect 38286 28636 38292 28688
rect 38344 28676 38350 28688
rect 38749 28679 38807 28685
rect 38749 28676 38761 28679
rect 38344 28648 38761 28676
rect 38344 28636 38350 28648
rect 38749 28645 38761 28648
rect 38795 28645 38807 28679
rect 40678 28676 40684 28688
rect 40591 28648 40684 28676
rect 38749 28639 38807 28645
rect 22143 28580 22594 28608
rect 22143 28577 22155 28580
rect 22097 28571 22155 28577
rect 27890 28568 27896 28620
rect 27948 28608 27954 28620
rect 28169 28611 28227 28617
rect 28169 28608 28181 28611
rect 27948 28580 28181 28608
rect 27948 28568 27954 28580
rect 28169 28577 28181 28580
rect 28215 28577 28227 28611
rect 28718 28608 28724 28620
rect 28631 28580 28724 28608
rect 28169 28571 28227 28577
rect 28718 28568 28724 28580
rect 28776 28608 28782 28620
rect 29362 28608 29368 28620
rect 28776 28580 29368 28608
rect 28776 28568 28782 28580
rect 29362 28568 29368 28580
rect 29420 28568 29426 28620
rect 30282 28568 30288 28620
rect 30340 28608 30346 28620
rect 30929 28611 30987 28617
rect 30929 28608 30941 28611
rect 30340 28580 30941 28608
rect 30340 28568 30346 28580
rect 30929 28577 30941 28580
rect 30975 28577 30987 28611
rect 33042 28608 33048 28620
rect 32955 28580 33048 28608
rect 30929 28571 30987 28577
rect 33042 28568 33048 28580
rect 33100 28608 33106 28620
rect 33686 28608 33692 28620
rect 33100 28580 33692 28608
rect 33100 28568 33106 28580
rect 33686 28568 33692 28580
rect 33744 28568 33750 28620
rect 35618 28568 35624 28620
rect 35676 28608 35682 28620
rect 36700 28611 36758 28617
rect 36700 28608 36712 28611
rect 35676 28580 36712 28608
rect 35676 28568 35682 28580
rect 36700 28577 36712 28580
rect 36746 28608 36758 28611
rect 36814 28608 36820 28620
rect 36746 28580 36820 28608
rect 36746 28577 36758 28580
rect 36700 28571 36758 28577
rect 36814 28568 36820 28580
rect 36872 28568 36878 28620
rect 37182 28568 37188 28620
rect 37240 28608 37246 28620
rect 37956 28611 38014 28617
rect 37956 28608 37968 28611
rect 37240 28580 37968 28608
rect 37240 28568 37246 28580
rect 37956 28577 37968 28580
rect 38002 28608 38014 28611
rect 38562 28608 38568 28620
rect 38002 28580 38568 28608
rect 38002 28577 38014 28580
rect 37956 28571 38014 28577
rect 38562 28568 38568 28580
rect 38620 28568 38626 28620
rect 40604 28617 40632 28648
rect 40678 28636 40684 28648
rect 40736 28676 40742 28688
rect 41046 28676 41052 28688
rect 40736 28648 41052 28676
rect 40736 28636 40742 28648
rect 41046 28636 41052 28648
rect 41104 28636 41110 28688
rect 42702 28636 42708 28688
rect 42760 28676 42766 28688
rect 44177 28679 44235 28685
rect 44177 28676 44189 28679
rect 42760 28648 44189 28676
rect 42760 28636 42766 28648
rect 44177 28645 44189 28648
rect 44223 28645 44235 28679
rect 44177 28639 44235 28645
rect 38984 28611 39042 28617
rect 38984 28577 38996 28611
rect 39030 28577 39042 28611
rect 38984 28571 39042 28577
rect 40589 28611 40647 28617
rect 40589 28577 40601 28611
rect 40635 28577 40647 28611
rect 40589 28571 40647 28577
rect 40773 28611 40831 28617
rect 40773 28577 40785 28611
rect 40819 28577 40831 28611
rect 40773 28571 40831 28577
rect 41944 28611 42002 28617
rect 41944 28577 41956 28611
rect 41990 28577 42002 28611
rect 41944 28571 42002 28577
rect 10870 28540 10876 28552
rect 10831 28512 10876 28540
rect 10870 28500 10876 28512
rect 10928 28500 10934 28552
rect 12066 28540 12072 28552
rect 12027 28512 12072 28540
rect 12066 28500 12072 28512
rect 12124 28500 12130 28552
rect 12713 28543 12771 28549
rect 12713 28509 12725 28543
rect 12759 28540 12771 28543
rect 12802 28540 12808 28552
rect 12759 28512 12808 28540
rect 12759 28509 12771 28512
rect 12713 28503 12771 28509
rect 12802 28500 12808 28512
rect 12860 28500 12866 28552
rect 15654 28540 15660 28552
rect 15615 28512 15660 28540
rect 15654 28500 15660 28512
rect 15712 28500 15718 28552
rect 17221 28543 17279 28549
rect 17221 28509 17233 28543
rect 17267 28540 17279 28543
rect 17494 28540 17500 28552
rect 17267 28512 17500 28540
rect 17267 28509 17279 28512
rect 17221 28503 17279 28509
rect 17494 28500 17500 28512
rect 17552 28500 17558 28552
rect 17586 28500 17592 28552
rect 17644 28540 17650 28552
rect 21174 28540 21180 28552
rect 17644 28512 17689 28540
rect 21135 28512 21180 28540
rect 17644 28500 17650 28512
rect 21174 28500 21180 28512
rect 21232 28500 21238 28552
rect 23017 28543 23075 28549
rect 23017 28509 23029 28543
rect 23063 28509 23075 28543
rect 23290 28540 23296 28552
rect 23251 28512 23296 28540
rect 23017 28503 23075 28509
rect 19935 28475 19993 28481
rect 19935 28441 19947 28475
rect 19981 28472 19993 28475
rect 23032 28472 23060 28503
rect 23290 28500 23296 28512
rect 23348 28500 23354 28552
rect 24762 28540 24768 28552
rect 24675 28512 24768 28540
rect 24762 28500 24768 28512
rect 24820 28540 24826 28552
rect 24949 28543 25007 28549
rect 24949 28540 24961 28543
rect 24820 28512 24961 28540
rect 24820 28500 24826 28512
rect 24949 28509 24961 28512
rect 24995 28509 25007 28543
rect 26602 28540 26608 28552
rect 26563 28512 26608 28540
rect 24949 28503 25007 28509
rect 26602 28500 26608 28512
rect 26660 28500 26666 28552
rect 26881 28543 26939 28549
rect 26881 28509 26893 28543
rect 26927 28509 26939 28543
rect 29730 28540 29736 28552
rect 29691 28512 29736 28540
rect 26881 28503 26939 28509
rect 23658 28472 23664 28484
rect 19981 28444 23664 28472
rect 19981 28441 19993 28444
rect 19935 28435 19993 28441
rect 23658 28432 23664 28444
rect 23716 28432 23722 28484
rect 25958 28432 25964 28484
rect 26016 28472 26022 28484
rect 26896 28472 26924 28503
rect 29730 28500 29736 28512
rect 29788 28500 29794 28552
rect 34885 28543 34943 28549
rect 34885 28509 34897 28543
rect 34931 28540 34943 28543
rect 35250 28540 35256 28552
rect 34931 28512 35256 28540
rect 34931 28509 34943 28512
rect 34885 28503 34943 28509
rect 35250 28500 35256 28512
rect 35308 28540 35314 28552
rect 35986 28540 35992 28552
rect 35308 28512 35992 28540
rect 35308 28500 35314 28512
rect 35986 28500 35992 28512
rect 36044 28500 36050 28552
rect 37642 28500 37648 28552
rect 37700 28540 37706 28552
rect 38999 28540 39027 28571
rect 39298 28540 39304 28552
rect 37700 28512 39304 28540
rect 37700 28500 37706 28512
rect 39298 28500 39304 28512
rect 39356 28500 39362 28552
rect 40218 28500 40224 28552
rect 40276 28540 40282 28552
rect 40788 28540 40816 28571
rect 41046 28540 41052 28552
rect 40276 28512 40816 28540
rect 41007 28512 41052 28540
rect 40276 28500 40282 28512
rect 41046 28500 41052 28512
rect 41104 28500 41110 28552
rect 41959 28540 41987 28571
rect 42334 28568 42340 28620
rect 42392 28608 42398 28620
rect 43254 28608 43260 28620
rect 42392 28580 43260 28608
rect 42392 28568 42398 28580
rect 43254 28568 43260 28580
rect 43312 28568 43318 28620
rect 43622 28568 43628 28620
rect 43680 28608 43686 28620
rect 44396 28611 44454 28617
rect 44396 28608 44408 28611
rect 43680 28580 44408 28608
rect 43680 28568 43686 28580
rect 44396 28577 44408 28580
rect 44442 28608 44454 28611
rect 44634 28608 44640 28620
rect 44442 28580 44640 28608
rect 44442 28577 44454 28580
rect 44396 28571 44454 28577
rect 44634 28568 44640 28580
rect 44692 28568 44698 28620
rect 42518 28540 42524 28552
rect 41959 28512 42524 28540
rect 42518 28500 42524 28512
rect 42576 28540 42582 28552
rect 42794 28540 42800 28552
rect 42576 28512 42800 28540
rect 42576 28500 42582 28512
rect 42794 28500 42800 28512
rect 42852 28500 42858 28552
rect 26016 28444 26924 28472
rect 36771 28475 36829 28481
rect 26016 28432 26022 28444
rect 36771 28441 36783 28475
rect 36817 28472 36829 28475
rect 39574 28472 39580 28484
rect 36817 28444 39580 28472
rect 36817 28441 36829 28444
rect 36771 28435 36829 28441
rect 39574 28432 39580 28444
rect 39632 28432 39638 28484
rect 41138 28432 41144 28484
rect 41196 28472 41202 28484
rect 43346 28472 43352 28484
rect 41196 28444 43352 28472
rect 41196 28432 41202 28444
rect 43346 28432 43352 28444
rect 43404 28432 43410 28484
rect 10502 28364 10508 28416
rect 10560 28404 10566 28416
rect 11333 28407 11391 28413
rect 11333 28404 11345 28407
rect 10560 28376 11345 28404
rect 10560 28364 10566 28376
rect 11333 28373 11345 28376
rect 11379 28373 11391 28407
rect 11333 28367 11391 28373
rect 14323 28407 14381 28413
rect 14323 28373 14335 28407
rect 14369 28404 14381 28407
rect 15010 28404 15016 28416
rect 14369 28376 15016 28404
rect 14369 28373 14381 28376
rect 14323 28367 14381 28373
rect 15010 28364 15016 28376
rect 15068 28364 15074 28416
rect 18138 28404 18144 28416
rect 18099 28376 18144 28404
rect 18138 28364 18144 28376
rect 18196 28364 18202 28416
rect 18690 28364 18696 28416
rect 18748 28404 18754 28416
rect 18831 28407 18889 28413
rect 18831 28404 18843 28407
rect 18748 28376 18843 28404
rect 18748 28364 18754 28376
rect 18831 28373 18843 28376
rect 18877 28373 18889 28407
rect 19702 28404 19708 28416
rect 19663 28376 19708 28404
rect 18831 28367 18889 28373
rect 19702 28364 19708 28376
rect 19760 28364 19766 28416
rect 20346 28404 20352 28416
rect 20307 28376 20352 28404
rect 20346 28364 20352 28376
rect 20404 28364 20410 28416
rect 23014 28364 23020 28416
rect 23072 28404 23078 28416
rect 27706 28404 27712 28416
rect 23072 28376 27712 28404
rect 23072 28364 23078 28376
rect 27706 28364 27712 28376
rect 27764 28364 27770 28416
rect 32214 28364 32220 28416
rect 32272 28404 32278 28416
rect 32309 28407 32367 28413
rect 32309 28404 32321 28407
rect 32272 28376 32321 28404
rect 32272 28364 32278 28376
rect 32309 28373 32321 28376
rect 32355 28373 32367 28407
rect 32858 28404 32864 28416
rect 32819 28376 32864 28404
rect 32309 28367 32367 28373
rect 32858 28364 32864 28376
rect 32916 28364 32922 28416
rect 37826 28364 37832 28416
rect 37884 28404 37890 28416
rect 38059 28407 38117 28413
rect 38059 28404 38071 28407
rect 37884 28376 38071 28404
rect 37884 28364 37890 28376
rect 38059 28373 38071 28376
rect 38105 28373 38117 28407
rect 38059 28367 38117 28373
rect 38930 28364 38936 28416
rect 38988 28404 38994 28416
rect 39071 28407 39129 28413
rect 39071 28404 39083 28407
rect 38988 28376 39083 28404
rect 38988 28364 38994 28376
rect 39071 28373 39083 28376
rect 39117 28373 39129 28407
rect 39071 28367 39129 28373
rect 41322 28364 41328 28416
rect 41380 28404 41386 28416
rect 41693 28407 41751 28413
rect 41693 28404 41705 28407
rect 41380 28376 41705 28404
rect 41380 28364 41386 28376
rect 41693 28373 41705 28376
rect 41739 28373 41751 28407
rect 41693 28367 41751 28373
rect 42015 28407 42073 28413
rect 42015 28373 42027 28407
rect 42061 28404 42073 28407
rect 42242 28404 42248 28416
rect 42061 28376 42248 28404
rect 42061 28373 42073 28376
rect 42015 28367 42073 28373
rect 42242 28364 42248 28376
rect 42300 28364 42306 28416
rect 43487 28407 43545 28413
rect 43487 28373 43499 28407
rect 43533 28404 43545 28407
rect 43714 28404 43720 28416
rect 43533 28376 43720 28404
rect 43533 28373 43545 28376
rect 43487 28367 43545 28373
rect 43714 28364 43720 28376
rect 43772 28364 43778 28416
rect 44499 28407 44557 28413
rect 44499 28373 44511 28407
rect 44545 28404 44557 28407
rect 45462 28404 45468 28416
rect 44545 28376 45468 28404
rect 44545 28373 44557 28376
rect 44499 28367 44557 28373
rect 45462 28364 45468 28376
rect 45520 28364 45526 28416
rect 1104 28314 48852 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 48852 28314
rect 1104 28240 48852 28262
rect 12526 28160 12532 28212
rect 12584 28200 12590 28212
rect 16485 28203 16543 28209
rect 12584 28172 13814 28200
rect 12584 28160 12590 28172
rect 13786 28132 13814 28172
rect 16485 28169 16497 28203
rect 16531 28200 16543 28203
rect 17494 28200 17500 28212
rect 16531 28172 17500 28200
rect 16531 28169 16543 28172
rect 16485 28163 16543 28169
rect 17494 28160 17500 28172
rect 17552 28160 17558 28212
rect 22554 28160 22560 28212
rect 22612 28200 22618 28212
rect 22741 28203 22799 28209
rect 22741 28200 22753 28203
rect 22612 28172 22753 28200
rect 22612 28160 22618 28172
rect 22741 28169 22753 28172
rect 22787 28169 22799 28203
rect 23106 28200 23112 28212
rect 23067 28172 23112 28200
rect 22741 28163 22799 28169
rect 23106 28160 23112 28172
rect 23164 28200 23170 28212
rect 24443 28203 24501 28209
rect 23164 28172 23474 28200
rect 23164 28160 23170 28172
rect 19702 28132 19708 28144
rect 13786 28104 19708 28132
rect 19702 28092 19708 28104
rect 19760 28132 19766 28144
rect 19797 28135 19855 28141
rect 19797 28132 19809 28135
rect 19760 28104 19809 28132
rect 19760 28092 19766 28104
rect 19797 28101 19809 28104
rect 19843 28101 19855 28135
rect 23446 28132 23474 28172
rect 24443 28169 24455 28203
rect 24489 28200 24501 28203
rect 24762 28200 24768 28212
rect 24489 28172 24768 28200
rect 24489 28169 24501 28172
rect 24443 28163 24501 28169
rect 24762 28160 24768 28172
rect 24820 28160 24826 28212
rect 26602 28160 26608 28212
rect 26660 28200 26666 28212
rect 27019 28203 27077 28209
rect 27019 28200 27031 28203
rect 26660 28172 27031 28200
rect 26660 28160 26666 28172
rect 27019 28169 27031 28172
rect 27065 28169 27077 28203
rect 27019 28163 27077 28169
rect 27338 28160 27344 28212
rect 27396 28200 27402 28212
rect 28626 28200 28632 28212
rect 27396 28172 28632 28200
rect 27396 28160 27402 28172
rect 28626 28160 28632 28172
rect 28684 28200 28690 28212
rect 29086 28200 29092 28212
rect 28684 28172 29092 28200
rect 28684 28160 28690 28172
rect 29086 28160 29092 28172
rect 29144 28160 29150 28212
rect 30190 28200 30196 28212
rect 30151 28172 30196 28200
rect 30190 28160 30196 28172
rect 30248 28160 30254 28212
rect 31251 28203 31309 28209
rect 31251 28169 31263 28203
rect 31297 28200 31309 28203
rect 32490 28200 32496 28212
rect 31297 28172 32496 28200
rect 31297 28169 31309 28172
rect 31251 28163 31309 28169
rect 32490 28160 32496 28172
rect 32548 28160 32554 28212
rect 33686 28200 33692 28212
rect 33647 28172 33692 28200
rect 33686 28160 33692 28172
rect 33744 28160 33750 28212
rect 34146 28160 34152 28212
rect 34204 28200 34210 28212
rect 34241 28203 34299 28209
rect 34241 28200 34253 28203
rect 34204 28172 34253 28200
rect 34204 28160 34210 28172
rect 34241 28169 34253 28172
rect 34287 28200 34299 28203
rect 34609 28203 34667 28209
rect 34609 28200 34621 28203
rect 34287 28172 34621 28200
rect 34287 28169 34299 28172
rect 34241 28163 34299 28169
rect 34609 28169 34621 28172
rect 34655 28169 34667 28203
rect 35894 28200 35900 28212
rect 35855 28172 35900 28200
rect 34609 28163 34667 28169
rect 24213 28135 24271 28141
rect 24213 28132 24225 28135
rect 23446 28104 24225 28132
rect 19797 28095 19855 28101
rect 24213 28101 24225 28104
rect 24259 28132 24271 28135
rect 25038 28132 25044 28144
rect 24259 28104 25044 28132
rect 24259 28101 24271 28104
rect 24213 28095 24271 28101
rect 25038 28092 25044 28104
rect 25096 28132 25102 28144
rect 25225 28135 25283 28141
rect 25225 28132 25237 28135
rect 25096 28104 25237 28132
rect 25096 28092 25102 28104
rect 25225 28101 25237 28104
rect 25271 28132 25283 28135
rect 26513 28135 26571 28141
rect 26513 28132 26525 28135
rect 25271 28104 26525 28132
rect 25271 28101 25283 28104
rect 25225 28095 25283 28101
rect 26513 28101 26525 28104
rect 26559 28132 26571 28135
rect 26694 28132 26700 28144
rect 26559 28104 26700 28132
rect 26559 28101 26571 28104
rect 26513 28095 26571 28101
rect 10502 28064 10508 28076
rect 10463 28036 10508 28064
rect 10502 28024 10508 28036
rect 10560 28024 10566 28076
rect 11790 28024 11796 28076
rect 11848 28064 11854 28076
rect 12069 28067 12127 28073
rect 12069 28064 12081 28067
rect 11848 28036 12081 28064
rect 11848 28024 11854 28036
rect 12069 28033 12081 28036
rect 12115 28064 12127 28067
rect 12158 28064 12164 28076
rect 12115 28036 12164 28064
rect 12115 28033 12127 28036
rect 12069 28027 12127 28033
rect 12158 28024 12164 28036
rect 12216 28064 12222 28076
rect 12989 28067 13047 28073
rect 12989 28064 13001 28067
rect 12216 28036 13001 28064
rect 12216 28024 12222 28036
rect 12989 28033 13001 28036
rect 13035 28064 13047 28067
rect 13262 28064 13268 28076
rect 13035 28036 13268 28064
rect 13035 28033 13047 28036
rect 12989 28027 13047 28033
rect 13262 28024 13268 28036
rect 13320 28024 13326 28076
rect 13817 28067 13875 28073
rect 13817 28033 13829 28067
rect 13863 28064 13875 28067
rect 14182 28064 14188 28076
rect 13863 28036 14188 28064
rect 13863 28033 13875 28036
rect 13817 28027 13875 28033
rect 14182 28024 14188 28036
rect 14240 28064 14246 28076
rect 15286 28064 15292 28076
rect 14240 28036 15292 28064
rect 14240 28024 14246 28036
rect 15286 28024 15292 28036
rect 15344 28064 15350 28076
rect 17586 28064 17592 28076
rect 15344 28036 17592 28064
rect 15344 28024 15350 28036
rect 17586 28024 17592 28036
rect 17644 28024 17650 28076
rect 21174 28064 21180 28076
rect 21087 28036 21180 28064
rect 21174 28024 21180 28036
rect 21232 28064 21238 28076
rect 21821 28067 21879 28073
rect 21821 28064 21833 28067
rect 21232 28036 21833 28064
rect 21232 28024 21238 28036
rect 21821 28033 21833 28036
rect 21867 28033 21879 28067
rect 21821 28027 21879 28033
rect 9560 27999 9618 28005
rect 9560 27965 9572 27999
rect 9606 27996 9618 27999
rect 11330 27996 11336 28008
rect 9606 27968 10088 27996
rect 9606 27965 9618 27968
rect 9560 27959 9618 27965
rect 9631 27863 9689 27869
rect 9631 27829 9643 27863
rect 9677 27860 9689 27863
rect 9858 27860 9864 27872
rect 9677 27832 9864 27860
rect 9677 27829 9689 27832
rect 9631 27823 9689 27829
rect 9858 27820 9864 27832
rect 9916 27820 9922 27872
rect 10060 27869 10088 27968
rect 10882 27968 11336 27996
rect 10882 27937 10910 27968
rect 11330 27956 11336 27968
rect 11388 27956 11394 28008
rect 14274 27996 14280 28008
rect 14235 27968 14280 27996
rect 14274 27956 14280 27968
rect 14332 27956 14338 28008
rect 17012 27999 17070 28005
rect 17012 27965 17024 27999
rect 17058 27996 17070 27999
rect 17497 27999 17555 28005
rect 17497 27996 17509 27999
rect 17058 27968 17509 27996
rect 17058 27965 17070 27968
rect 17012 27959 17070 27965
rect 17497 27965 17509 27968
rect 17543 27996 17555 27999
rect 17678 27996 17684 28008
rect 17543 27968 17684 27996
rect 17543 27965 17555 27968
rect 17497 27959 17555 27965
rect 17678 27956 17684 27968
rect 17736 27956 17742 28008
rect 18138 27996 18144 28008
rect 18099 27968 18144 27996
rect 18138 27956 18144 27968
rect 18196 27956 18202 28008
rect 20441 27999 20499 28005
rect 20441 27996 20453 27999
rect 20272 27968 20453 27996
rect 10413 27931 10471 27937
rect 10413 27897 10425 27931
rect 10459 27928 10471 27931
rect 10867 27931 10925 27937
rect 10867 27928 10879 27931
rect 10459 27900 10879 27928
rect 10459 27897 10471 27900
rect 10413 27891 10471 27897
rect 10867 27897 10879 27900
rect 10913 27897 10925 27931
rect 11698 27928 11704 27940
rect 10867 27891 10925 27897
rect 11164 27900 11704 27928
rect 10045 27863 10103 27869
rect 10045 27829 10057 27863
rect 10091 27860 10103 27863
rect 11164 27860 11192 27900
rect 11698 27888 11704 27900
rect 11756 27928 11762 27940
rect 12526 27928 12532 27940
rect 11756 27900 12532 27928
rect 11756 27888 11762 27900
rect 12526 27888 12532 27900
rect 12584 27888 12590 27940
rect 13173 27931 13231 27937
rect 13173 27897 13185 27931
rect 13219 27897 13231 27931
rect 13173 27891 13231 27897
rect 11422 27860 11428 27872
rect 10091 27832 11192 27860
rect 11383 27832 11428 27860
rect 10091 27829 10103 27832
rect 10045 27823 10103 27829
rect 11422 27820 11428 27832
rect 11480 27820 11486 27872
rect 13078 27820 13084 27872
rect 13136 27860 13142 27872
rect 13188 27860 13216 27891
rect 13262 27888 13268 27940
rect 13320 27928 13326 27940
rect 15102 27928 15108 27940
rect 13320 27900 13365 27928
rect 15063 27900 15108 27928
rect 13320 27888 13326 27900
rect 15102 27888 15108 27900
rect 15160 27888 15166 27940
rect 15197 27931 15255 27937
rect 15197 27897 15209 27931
rect 15243 27928 15255 27931
rect 15470 27928 15476 27940
rect 15243 27900 15476 27928
rect 15243 27897 15255 27900
rect 15197 27891 15255 27897
rect 13136 27832 13216 27860
rect 13136 27820 13142 27832
rect 13722 27820 13728 27872
rect 13780 27860 13786 27872
rect 14829 27863 14887 27869
rect 14829 27860 14841 27863
rect 13780 27832 14841 27860
rect 13780 27820 13786 27832
rect 14829 27829 14841 27832
rect 14875 27860 14887 27863
rect 15212 27860 15240 27891
rect 15470 27888 15476 27900
rect 15528 27888 15534 27940
rect 15746 27928 15752 27940
rect 15707 27900 15752 27928
rect 15746 27888 15752 27900
rect 15804 27888 15810 27940
rect 16853 27931 16911 27937
rect 16853 27897 16865 27931
rect 16899 27928 16911 27931
rect 17218 27928 17224 27940
rect 16899 27900 17224 27928
rect 16899 27897 16911 27900
rect 16853 27891 16911 27897
rect 17218 27888 17224 27900
rect 17276 27888 17282 27940
rect 18598 27888 18604 27940
rect 18656 27928 18662 27940
rect 19337 27931 19395 27937
rect 19337 27928 19349 27931
rect 18656 27900 19349 27928
rect 18656 27888 18662 27900
rect 19337 27897 19349 27900
rect 19383 27897 19395 27931
rect 19337 27891 19395 27897
rect 14875 27832 15240 27860
rect 15488 27860 15516 27888
rect 20272 27872 20300 27968
rect 20441 27965 20453 27968
rect 20487 27965 20499 27999
rect 20441 27959 20499 27965
rect 20898 27956 20904 28008
rect 20956 27996 20962 28008
rect 20993 27999 21051 28005
rect 20993 27996 21005 27999
rect 20956 27968 21005 27996
rect 20956 27956 20962 27968
rect 20993 27965 21005 27968
rect 21039 27996 21051 27999
rect 21634 27996 21640 28008
rect 21039 27968 21640 27996
rect 21039 27965 21051 27968
rect 20993 27959 21051 27965
rect 21634 27956 21640 27968
rect 21692 27956 21698 28008
rect 21726 27956 21732 28008
rect 21784 27996 21790 28008
rect 22348 27999 22406 28005
rect 22348 27996 22360 27999
rect 21784 27968 22360 27996
rect 21784 27956 21790 27968
rect 22348 27965 22360 27968
rect 22394 27996 22406 27999
rect 22554 27996 22560 28008
rect 22394 27968 22560 27996
rect 22394 27965 22406 27968
rect 22348 27959 22406 27965
rect 22554 27956 22560 27968
rect 22612 27956 22618 28008
rect 24372 27999 24430 28005
rect 24372 27965 24384 27999
rect 24418 27996 24430 27999
rect 24418 27968 24900 27996
rect 24418 27965 24430 27968
rect 24372 27959 24430 27965
rect 16025 27863 16083 27869
rect 16025 27860 16037 27863
rect 15488 27832 16037 27860
rect 14875 27829 14887 27832
rect 14829 27823 14887 27829
rect 16025 27829 16037 27832
rect 16071 27829 16083 27863
rect 16025 27823 16083 27829
rect 16942 27820 16948 27872
rect 17000 27860 17006 27872
rect 17083 27863 17141 27869
rect 17083 27860 17095 27863
rect 17000 27832 17095 27860
rect 17000 27820 17006 27832
rect 17083 27829 17095 27832
rect 17129 27829 17141 27863
rect 17083 27823 17141 27829
rect 17865 27863 17923 27869
rect 17865 27829 17877 27863
rect 17911 27860 17923 27863
rect 18506 27860 18512 27872
rect 17911 27832 18512 27860
rect 17911 27829 17923 27832
rect 17865 27823 17923 27829
rect 18506 27820 18512 27832
rect 18564 27820 18570 27872
rect 18782 27820 18788 27872
rect 18840 27860 18846 27872
rect 19061 27863 19119 27869
rect 19061 27860 19073 27863
rect 18840 27832 19073 27860
rect 18840 27820 18846 27832
rect 19061 27829 19073 27832
rect 19107 27829 19119 27863
rect 20254 27860 20260 27872
rect 20215 27832 20260 27860
rect 19061 27823 19119 27829
rect 20254 27820 20260 27832
rect 20312 27820 20318 27872
rect 21450 27860 21456 27872
rect 21411 27832 21456 27860
rect 21450 27820 21456 27832
rect 21508 27820 21514 27872
rect 22419 27863 22477 27869
rect 22419 27829 22431 27863
rect 22465 27860 22477 27863
rect 22554 27860 22560 27872
rect 22465 27832 22560 27860
rect 22465 27829 22477 27832
rect 22419 27823 22477 27829
rect 22554 27820 22560 27832
rect 22612 27820 22618 27872
rect 24872 27869 24900 27968
rect 25240 27928 25268 28095
rect 26694 28092 26700 28104
rect 26752 28092 26758 28144
rect 32858 28092 32864 28144
rect 32916 28132 32922 28144
rect 33045 28135 33103 28141
rect 33045 28132 33057 28135
rect 32916 28104 33057 28132
rect 32916 28092 32922 28104
rect 33045 28101 33057 28104
rect 33091 28101 33103 28135
rect 33410 28132 33416 28144
rect 33371 28104 33416 28132
rect 33045 28095 33103 28101
rect 33410 28092 33416 28104
rect 33468 28092 33474 28144
rect 25409 28067 25467 28073
rect 25409 28033 25421 28067
rect 25455 28064 25467 28067
rect 25590 28064 25596 28076
rect 25455 28036 25596 28064
rect 25455 28033 25467 28036
rect 25409 28027 25467 28033
rect 25590 28024 25596 28036
rect 25648 28064 25654 28076
rect 28031 28067 28089 28073
rect 28031 28064 28043 28067
rect 25648 28036 28043 28064
rect 25648 28024 25654 28036
rect 28031 28033 28043 28036
rect 28077 28033 28089 28067
rect 28031 28027 28089 28033
rect 29178 28024 29184 28076
rect 29236 28064 29242 28076
rect 29273 28067 29331 28073
rect 29273 28064 29285 28067
rect 29236 28036 29285 28064
rect 29236 28024 29242 28036
rect 29273 28033 29285 28036
rect 29319 28033 29331 28067
rect 31941 28067 31999 28073
rect 31941 28064 31953 28067
rect 29273 28027 29331 28033
rect 30944 28036 31953 28064
rect 26050 27956 26056 28008
rect 26108 27996 26114 28008
rect 27338 27996 27344 28008
rect 26108 27968 26153 27996
rect 27299 27968 27344 27996
rect 26108 27956 26114 27968
rect 27338 27956 27344 27968
rect 27396 27956 27402 28008
rect 27944 27999 28002 28005
rect 27944 27965 27956 27999
rect 27990 27996 28002 27999
rect 27990 27968 28304 27996
rect 27990 27965 28002 27968
rect 27944 27959 28002 27965
rect 25501 27931 25559 27937
rect 25501 27928 25513 27931
rect 25240 27900 25513 27928
rect 25501 27897 25513 27900
rect 25547 27897 25559 27931
rect 25501 27891 25559 27897
rect 26789 27931 26847 27937
rect 26789 27897 26801 27931
rect 26835 27928 26847 27931
rect 27356 27928 27384 27956
rect 26835 27900 27384 27928
rect 26835 27897 26847 27900
rect 26789 27891 26847 27897
rect 28276 27872 28304 27968
rect 29635 27931 29693 27937
rect 29635 27897 29647 27931
rect 29681 27897 29693 27931
rect 29635 27891 29693 27897
rect 24857 27863 24915 27869
rect 24857 27829 24869 27863
rect 24903 27860 24915 27863
rect 25314 27860 25320 27872
rect 24903 27832 25320 27860
rect 24903 27829 24915 27832
rect 24857 27823 24915 27829
rect 25314 27820 25320 27832
rect 25372 27820 25378 27872
rect 27801 27863 27859 27869
rect 27801 27829 27813 27863
rect 27847 27860 27859 27863
rect 27890 27860 27896 27872
rect 27847 27832 27896 27860
rect 27847 27829 27859 27832
rect 27801 27823 27859 27829
rect 27890 27820 27896 27832
rect 27948 27820 27954 27872
rect 28258 27820 28264 27872
rect 28316 27860 28322 27872
rect 28353 27863 28411 27869
rect 28353 27860 28365 27863
rect 28316 27832 28365 27860
rect 28316 27820 28322 27832
rect 28353 27829 28365 27832
rect 28399 27829 28411 27863
rect 28994 27860 29000 27872
rect 28955 27832 29000 27860
rect 28353 27823 28411 27829
rect 28994 27820 29000 27832
rect 29052 27860 29058 27872
rect 29650 27860 29678 27891
rect 29730 27888 29736 27940
rect 29788 27928 29794 27940
rect 30837 27931 30895 27937
rect 30837 27928 30849 27931
rect 29788 27900 30849 27928
rect 29788 27888 29794 27900
rect 30837 27897 30849 27900
rect 30883 27897 30895 27931
rect 30837 27891 30895 27897
rect 30098 27860 30104 27872
rect 29052 27832 30104 27860
rect 29052 27820 29058 27832
rect 30098 27820 30104 27832
rect 30156 27860 30162 27872
rect 30469 27863 30527 27869
rect 30469 27860 30481 27863
rect 30156 27832 30481 27860
rect 30156 27820 30162 27832
rect 30469 27829 30481 27832
rect 30515 27860 30527 27863
rect 30944 27860 30972 28036
rect 31941 28033 31953 28036
rect 31987 28064 31999 28067
rect 31987 28036 32489 28064
rect 31987 28033 31999 28036
rect 31941 28027 31999 28033
rect 31180 27999 31238 28005
rect 31180 27965 31192 27999
rect 31226 27996 31238 27999
rect 32125 27999 32183 28005
rect 31226 27968 31708 27996
rect 31226 27965 31238 27968
rect 31180 27959 31238 27965
rect 31680 27872 31708 27968
rect 32125 27965 32137 27999
rect 32171 27996 32183 27999
rect 32214 27996 32220 28008
rect 32171 27968 32220 27996
rect 32171 27965 32183 27968
rect 32125 27959 32183 27965
rect 32214 27956 32220 27968
rect 32272 27956 32278 28008
rect 32461 27937 32489 28036
rect 32446 27931 32504 27937
rect 32446 27897 32458 27931
rect 32492 27928 32504 27931
rect 33410 27928 33416 27940
rect 32492 27900 33416 27928
rect 32492 27897 32504 27900
rect 32446 27891 32504 27897
rect 33410 27888 33416 27900
rect 33468 27888 33474 27940
rect 34624 27928 34652 28163
rect 35894 28160 35900 28172
rect 35952 28160 35958 28212
rect 37182 28200 37188 28212
rect 37143 28172 37188 28200
rect 37182 28160 37188 28172
rect 37240 28160 37246 28212
rect 39298 28200 39304 28212
rect 39259 28172 39304 28200
rect 39298 28160 39304 28172
rect 39356 28160 39362 28212
rect 40678 28200 40684 28212
rect 40639 28172 40684 28200
rect 40678 28160 40684 28172
rect 40736 28160 40742 28212
rect 41138 28200 41144 28212
rect 41099 28172 41144 28200
rect 41138 28160 41144 28172
rect 41196 28160 41202 28212
rect 43254 28160 43260 28212
rect 43312 28200 43318 28212
rect 43349 28203 43407 28209
rect 43349 28200 43361 28203
rect 43312 28172 43361 28200
rect 43312 28160 43318 28172
rect 43349 28169 43361 28172
rect 43395 28169 43407 28203
rect 44634 28200 44640 28212
rect 44595 28172 44640 28200
rect 43349 28163 43407 28169
rect 44634 28160 44640 28172
rect 44692 28160 44698 28212
rect 34977 28067 35035 28073
rect 34977 28033 34989 28067
rect 35023 28064 35035 28067
rect 35912 28064 35940 28160
rect 38562 28092 38568 28144
rect 38620 28132 38626 28144
rect 40696 28132 40724 28160
rect 38620 28104 40724 28132
rect 38620 28092 38626 28104
rect 35023 28036 35940 28064
rect 37415 28067 37473 28073
rect 35023 28033 35035 28036
rect 34977 28027 35035 28033
rect 37415 28033 37427 28067
rect 37461 28064 37473 28067
rect 38381 28067 38439 28073
rect 38381 28064 38393 28067
rect 37461 28036 38393 28064
rect 37461 28033 37473 28036
rect 37415 28027 37473 28033
rect 38381 28033 38393 28036
rect 38427 28064 38439 28067
rect 39669 28067 39727 28073
rect 39669 28064 39681 28067
rect 38427 28036 39681 28064
rect 38427 28033 38439 28036
rect 38381 28027 38439 28033
rect 39669 28033 39681 28036
rect 39715 28033 39727 28067
rect 41322 28064 41328 28076
rect 41283 28036 41328 28064
rect 39669 28027 39727 28033
rect 41322 28024 41328 28036
rect 41380 28024 41386 28076
rect 43073 28067 43131 28073
rect 43073 28033 43085 28067
rect 43119 28064 43131 28067
rect 43714 28064 43720 28076
rect 43119 28036 43720 28064
rect 43119 28033 43131 28036
rect 43073 28027 43131 28033
rect 43714 28024 43720 28036
rect 43772 28024 43778 28076
rect 43806 28024 43812 28076
rect 43864 28064 43870 28076
rect 43993 28067 44051 28073
rect 43993 28064 44005 28067
rect 43864 28036 44005 28064
rect 43864 28024 43870 28036
rect 43993 28033 44005 28036
rect 44039 28033 44051 28067
rect 43993 28027 44051 28033
rect 37328 27999 37386 28005
rect 37328 27965 37340 27999
rect 37374 27996 37386 27999
rect 37374 27968 37872 27996
rect 37374 27965 37386 27968
rect 37328 27959 37386 27965
rect 35069 27931 35127 27937
rect 35069 27928 35081 27931
rect 34624 27900 35081 27928
rect 35069 27897 35081 27900
rect 35115 27897 35127 27931
rect 35069 27891 35127 27897
rect 35621 27931 35679 27937
rect 35621 27897 35633 27931
rect 35667 27897 35679 27931
rect 35621 27891 35679 27897
rect 31662 27860 31668 27872
rect 30515 27832 30972 27860
rect 31623 27832 31668 27860
rect 30515 27829 30527 27832
rect 30469 27823 30527 27829
rect 31662 27820 31668 27832
rect 31720 27820 31726 27872
rect 33226 27820 33232 27872
rect 33284 27860 33290 27872
rect 35636 27860 35664 27891
rect 33284 27832 35664 27860
rect 36725 27863 36783 27869
rect 33284 27820 33290 27832
rect 36725 27829 36737 27863
rect 36771 27860 36783 27863
rect 36814 27860 36820 27872
rect 36771 27832 36820 27860
rect 36771 27829 36783 27832
rect 36725 27823 36783 27829
rect 36814 27820 36820 27832
rect 36872 27820 36878 27872
rect 37844 27869 37872 27968
rect 41874 27956 41880 28008
rect 41932 27996 41938 28008
rect 42245 27999 42303 28005
rect 42245 27996 42257 27999
rect 41932 27968 42257 27996
rect 41932 27956 41938 27968
rect 42245 27965 42257 27968
rect 42291 27996 42303 27999
rect 42291 27968 42794 27996
rect 42291 27965 42303 27968
rect 42245 27959 42303 27965
rect 38197 27931 38255 27937
rect 38197 27897 38209 27931
rect 38243 27928 38255 27931
rect 38473 27931 38531 27937
rect 38473 27928 38485 27931
rect 38243 27900 38485 27928
rect 38243 27897 38255 27900
rect 38197 27891 38255 27897
rect 38473 27897 38485 27900
rect 38519 27928 38531 27931
rect 38654 27928 38660 27940
rect 38519 27900 38660 27928
rect 38519 27897 38531 27900
rect 38473 27891 38531 27897
rect 38654 27888 38660 27900
rect 38712 27888 38718 27940
rect 38838 27888 38844 27940
rect 38896 27928 38902 27940
rect 39025 27931 39083 27937
rect 39025 27928 39037 27931
rect 38896 27900 39037 27928
rect 38896 27888 38902 27900
rect 39025 27897 39037 27900
rect 39071 27897 39083 27931
rect 39025 27891 39083 27897
rect 41138 27888 41144 27940
rect 41196 27928 41202 27940
rect 41506 27928 41512 27940
rect 41196 27900 41512 27928
rect 41196 27888 41202 27900
rect 41506 27888 41512 27900
rect 41564 27928 41570 27940
rect 41646 27931 41704 27937
rect 41646 27928 41658 27931
rect 41564 27900 41658 27928
rect 41564 27888 41570 27900
rect 41646 27897 41658 27900
rect 41692 27897 41704 27931
rect 42766 27928 42794 27968
rect 43809 27931 43867 27937
rect 43809 27928 43821 27931
rect 42766 27900 43821 27928
rect 41646 27891 41704 27897
rect 43809 27897 43821 27900
rect 43855 27897 43867 27931
rect 43809 27891 43867 27897
rect 37829 27863 37887 27869
rect 37829 27829 37841 27863
rect 37875 27860 37887 27863
rect 38010 27860 38016 27872
rect 37875 27832 38016 27860
rect 37875 27829 37887 27832
rect 37829 27823 37887 27829
rect 38010 27820 38016 27832
rect 38068 27860 38074 27872
rect 38746 27860 38752 27872
rect 38068 27832 38752 27860
rect 38068 27820 38074 27832
rect 38746 27820 38752 27832
rect 38804 27820 38810 27872
rect 40218 27860 40224 27872
rect 40179 27832 40224 27860
rect 40218 27820 40224 27832
rect 40276 27820 40282 27872
rect 42518 27860 42524 27872
rect 42479 27832 42524 27860
rect 42518 27820 42524 27832
rect 42576 27820 42582 27872
rect 43622 27820 43628 27872
rect 43680 27860 43686 27872
rect 43824 27860 43852 27891
rect 43680 27832 43852 27860
rect 43680 27820 43686 27832
rect 1104 27770 48852 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 48852 27770
rect 1104 27696 48852 27718
rect 11422 27616 11428 27668
rect 11480 27656 11486 27668
rect 12437 27659 12495 27665
rect 12437 27656 12449 27659
rect 11480 27628 12449 27656
rect 11480 27616 11486 27628
rect 12437 27625 12449 27628
rect 12483 27656 12495 27659
rect 12618 27656 12624 27668
rect 12483 27628 12624 27656
rect 12483 27625 12495 27628
rect 12437 27619 12495 27625
rect 12618 27616 12624 27628
rect 12676 27656 12682 27668
rect 13722 27656 13728 27668
rect 12676 27628 13728 27656
rect 12676 27616 12682 27628
rect 10318 27548 10324 27600
rect 10376 27588 10382 27600
rect 10413 27591 10471 27597
rect 10413 27588 10425 27591
rect 10376 27560 10425 27588
rect 10376 27548 10382 27560
rect 10413 27557 10425 27560
rect 10459 27588 10471 27591
rect 11235 27591 11293 27597
rect 10459 27560 11192 27588
rect 10459 27557 10471 27560
rect 10413 27551 10471 27557
rect 10870 27520 10876 27532
rect 10831 27492 10876 27520
rect 10870 27480 10876 27492
rect 10928 27480 10934 27532
rect 11164 27520 11192 27560
rect 11235 27557 11247 27591
rect 11281 27588 11293 27591
rect 11330 27588 11336 27600
rect 11281 27560 11336 27588
rect 11281 27557 11293 27560
rect 11235 27551 11293 27557
rect 11330 27548 11336 27560
rect 11388 27548 11394 27600
rect 13648 27597 13676 27628
rect 13722 27616 13728 27628
rect 13780 27616 13786 27668
rect 20254 27656 20260 27668
rect 14292 27628 20260 27656
rect 12253 27591 12311 27597
rect 12253 27588 12265 27591
rect 11486 27560 12265 27588
rect 11486 27520 11514 27560
rect 12253 27557 12265 27560
rect 12299 27557 12311 27591
rect 12253 27551 12311 27557
rect 13633 27591 13691 27597
rect 13633 27557 13645 27591
rect 13679 27557 13691 27591
rect 14182 27588 14188 27600
rect 14143 27560 14188 27588
rect 13633 27551 13691 27557
rect 14182 27548 14188 27560
rect 14240 27548 14246 27600
rect 11790 27520 11796 27532
rect 11164 27492 11514 27520
rect 11751 27492 11796 27520
rect 11790 27480 11796 27492
rect 11848 27480 11854 27532
rect 8573 27455 8631 27461
rect 8573 27421 8585 27455
rect 8619 27452 8631 27455
rect 9999 27455 10057 27461
rect 8619 27424 9674 27452
rect 8619 27421 8631 27424
rect 8573 27415 8631 27421
rect 9646 27384 9674 27424
rect 9999 27421 10011 27455
rect 10045 27452 10057 27455
rect 13541 27455 13599 27461
rect 13541 27452 13553 27455
rect 10045 27424 13553 27452
rect 10045 27421 10057 27424
rect 9999 27415 10057 27421
rect 13541 27421 13553 27424
rect 13587 27452 13599 27455
rect 13814 27452 13820 27464
rect 13587 27424 13820 27452
rect 13587 27421 13599 27424
rect 13541 27415 13599 27421
rect 13814 27412 13820 27424
rect 13872 27412 13878 27464
rect 12158 27384 12164 27396
rect 9646 27356 12164 27384
rect 12158 27344 12164 27356
rect 12216 27344 12222 27396
rect 12250 27344 12256 27396
rect 12308 27384 12314 27396
rect 14292 27384 14320 27628
rect 20254 27616 20260 27628
rect 20312 27616 20318 27668
rect 23658 27656 23664 27668
rect 23619 27628 23664 27656
rect 23658 27616 23664 27628
rect 23716 27616 23722 27668
rect 25590 27656 25596 27668
rect 25551 27628 25596 27656
rect 25590 27616 25596 27628
rect 25648 27616 25654 27668
rect 26602 27616 26608 27668
rect 26660 27656 26666 27668
rect 26697 27659 26755 27665
rect 26697 27656 26709 27659
rect 26660 27628 26709 27656
rect 26660 27616 26666 27628
rect 26697 27625 26709 27628
rect 26743 27625 26755 27659
rect 32214 27656 32220 27668
rect 32175 27628 32220 27656
rect 26697 27619 26755 27625
rect 32214 27616 32220 27628
rect 32272 27616 32278 27668
rect 35161 27659 35219 27665
rect 35161 27625 35173 27659
rect 35207 27656 35219 27659
rect 35250 27656 35256 27668
rect 35207 27628 35256 27656
rect 35207 27625 35219 27628
rect 35161 27619 35219 27625
rect 35250 27616 35256 27628
rect 35308 27616 35314 27668
rect 38102 27656 38108 27668
rect 38063 27628 38108 27656
rect 38102 27616 38108 27628
rect 38160 27616 38166 27668
rect 38654 27656 38660 27668
rect 38615 27628 38660 27656
rect 38654 27616 38660 27628
rect 38712 27656 38718 27668
rect 38933 27659 38991 27665
rect 38933 27656 38945 27659
rect 38712 27628 38945 27656
rect 38712 27616 38718 27628
rect 38933 27625 38945 27628
rect 38979 27656 38991 27659
rect 39482 27656 39488 27668
rect 38979 27628 39488 27656
rect 38979 27625 38991 27628
rect 38933 27619 38991 27625
rect 39482 27616 39488 27628
rect 39540 27656 39546 27668
rect 41506 27656 41512 27668
rect 39540 27628 39712 27656
rect 41467 27628 41512 27656
rect 39540 27616 39546 27628
rect 15470 27588 15476 27600
rect 15431 27560 15476 27588
rect 15470 27548 15476 27560
rect 15528 27548 15534 27600
rect 16942 27548 16948 27600
rect 17000 27588 17006 27600
rect 17129 27591 17187 27597
rect 17129 27588 17141 27591
rect 17000 27560 17141 27588
rect 17000 27548 17006 27560
rect 17129 27557 17141 27560
rect 17175 27557 17187 27591
rect 17129 27551 17187 27557
rect 17218 27548 17224 27600
rect 17276 27588 17282 27600
rect 18509 27591 18567 27597
rect 17276 27560 17321 27588
rect 17276 27548 17282 27560
rect 18509 27557 18521 27591
rect 18555 27588 18567 27591
rect 18690 27588 18696 27600
rect 18555 27560 18696 27588
rect 18555 27557 18567 27560
rect 18509 27551 18567 27557
rect 18690 27548 18696 27560
rect 18748 27548 18754 27600
rect 18782 27548 18788 27600
rect 18840 27588 18846 27600
rect 19981 27591 20039 27597
rect 18840 27560 18885 27588
rect 18840 27548 18846 27560
rect 19981 27557 19993 27591
rect 20027 27588 20039 27591
rect 20438 27588 20444 27600
rect 20027 27560 20444 27588
rect 20027 27557 20039 27560
rect 19981 27551 20039 27557
rect 20438 27548 20444 27560
rect 20496 27548 20502 27600
rect 22554 27548 22560 27600
rect 22612 27588 22618 27600
rect 22741 27591 22799 27597
rect 22741 27588 22753 27591
rect 22612 27560 22753 27588
rect 22612 27548 22618 27560
rect 22741 27557 22753 27560
rect 22787 27557 22799 27591
rect 22741 27551 22799 27557
rect 22833 27591 22891 27597
rect 22833 27557 22845 27591
rect 22879 27588 22891 27591
rect 23014 27588 23020 27600
rect 22879 27560 23020 27588
rect 22879 27557 22891 27560
rect 22833 27551 22891 27557
rect 23014 27548 23020 27560
rect 23072 27588 23078 27600
rect 25130 27588 25136 27600
rect 23072 27560 25136 27588
rect 23072 27548 23078 27560
rect 25130 27548 25136 27560
rect 25188 27548 25194 27600
rect 27985 27591 28043 27597
rect 27985 27557 27997 27591
rect 28031 27588 28043 27591
rect 30374 27588 30380 27600
rect 28031 27560 30380 27588
rect 28031 27557 28043 27560
rect 27985 27551 28043 27557
rect 30374 27548 30380 27560
rect 30432 27548 30438 27600
rect 31159 27591 31217 27597
rect 31159 27557 31171 27591
rect 31205 27588 31217 27591
rect 34790 27588 34796 27600
rect 31205 27560 34796 27588
rect 31205 27557 31217 27560
rect 31159 27551 31217 27557
rect 34790 27548 34796 27560
rect 34848 27548 34854 27600
rect 39574 27588 39580 27600
rect 39535 27560 39580 27588
rect 39574 27548 39580 27560
rect 39632 27548 39638 27600
rect 39684 27597 39712 27628
rect 41506 27616 41512 27628
rect 41564 27616 41570 27668
rect 42242 27616 42248 27668
rect 42300 27656 42306 27668
rect 42337 27659 42395 27665
rect 42337 27656 42349 27659
rect 42300 27628 42349 27656
rect 42300 27616 42306 27628
rect 42337 27625 42349 27628
rect 42383 27625 42395 27659
rect 42337 27619 42395 27625
rect 39669 27591 39727 27597
rect 39669 27557 39681 27591
rect 39715 27557 39727 27591
rect 39669 27551 39727 27557
rect 43622 27548 43628 27600
rect 43680 27588 43686 27600
rect 43993 27591 44051 27597
rect 43993 27588 44005 27591
rect 43680 27560 44005 27588
rect 43680 27548 43686 27560
rect 43993 27557 44005 27560
rect 44039 27557 44051 27591
rect 45462 27588 45468 27600
rect 45423 27560 45468 27588
rect 43993 27551 44051 27557
rect 45462 27548 45468 27560
rect 45520 27548 45526 27600
rect 45554 27548 45560 27600
rect 45612 27588 45618 27600
rect 45612 27560 45657 27588
rect 45612 27548 45618 27560
rect 21082 27520 21088 27532
rect 21043 27492 21088 27520
rect 21082 27480 21088 27492
rect 21140 27480 21146 27532
rect 21634 27520 21640 27532
rect 21595 27492 21640 27520
rect 21634 27480 21640 27492
rect 21692 27480 21698 27532
rect 24740 27523 24798 27529
rect 24740 27489 24752 27523
rect 24786 27520 24798 27523
rect 24854 27520 24860 27532
rect 24786 27492 24860 27520
rect 24786 27489 24798 27492
rect 24740 27483 24798 27489
rect 24854 27480 24860 27492
rect 24912 27480 24918 27532
rect 27246 27520 27252 27532
rect 27207 27492 27252 27520
rect 27246 27480 27252 27492
rect 27304 27480 27310 27532
rect 28718 27480 28724 27532
rect 28776 27520 28782 27532
rect 28813 27523 28871 27529
rect 28813 27520 28825 27523
rect 28776 27492 28825 27520
rect 28776 27480 28782 27492
rect 28813 27489 28825 27492
rect 28859 27489 28871 27523
rect 29362 27520 29368 27532
rect 29323 27492 29368 27520
rect 28813 27483 28871 27489
rect 29362 27480 29368 27492
rect 29420 27480 29426 27532
rect 29549 27523 29607 27529
rect 29549 27489 29561 27523
rect 29595 27520 29607 27523
rect 29730 27520 29736 27532
rect 29595 27492 29736 27520
rect 29595 27489 29607 27492
rect 29549 27483 29607 27489
rect 29730 27480 29736 27492
rect 29788 27480 29794 27532
rect 31072 27523 31130 27529
rect 31072 27489 31084 27523
rect 31118 27489 31130 27523
rect 31072 27483 31130 27489
rect 15378 27452 15384 27464
rect 15339 27424 15384 27452
rect 15378 27412 15384 27424
rect 15436 27412 15442 27464
rect 15746 27452 15752 27464
rect 15707 27424 15752 27452
rect 15746 27412 15752 27424
rect 15804 27452 15810 27464
rect 17126 27452 17132 27464
rect 15804 27424 17132 27452
rect 15804 27412 15810 27424
rect 17126 27412 17132 27424
rect 17184 27452 17190 27464
rect 17405 27455 17463 27461
rect 17405 27452 17417 27455
rect 17184 27424 17417 27452
rect 17184 27412 17190 27424
rect 17405 27421 17417 27424
rect 17451 27421 17463 27455
rect 17405 27415 17463 27421
rect 18874 27412 18880 27464
rect 18932 27452 18938 27464
rect 18969 27455 19027 27461
rect 18969 27452 18981 27455
rect 18932 27424 18981 27452
rect 18932 27412 18938 27424
rect 18969 27421 18981 27424
rect 19015 27421 19027 27455
rect 18969 27415 19027 27421
rect 20533 27455 20591 27461
rect 20533 27421 20545 27455
rect 20579 27452 20591 27455
rect 21652 27452 21680 27480
rect 21818 27452 21824 27464
rect 20579 27424 21680 27452
rect 21779 27424 21824 27452
rect 20579 27421 20591 27424
rect 20533 27415 20591 27421
rect 21818 27412 21824 27424
rect 21876 27412 21882 27464
rect 27522 27412 27528 27464
rect 27580 27452 27586 27464
rect 27617 27455 27675 27461
rect 27617 27452 27629 27455
rect 27580 27424 27629 27452
rect 27580 27412 27586 27424
rect 27617 27421 27629 27424
rect 27663 27421 27675 27455
rect 27617 27415 27675 27421
rect 28353 27455 28411 27461
rect 28353 27421 28365 27455
rect 28399 27452 28411 27455
rect 29380 27452 29408 27480
rect 28399 27424 29408 27452
rect 31087 27452 31115 27483
rect 32306 27480 32312 27532
rect 32364 27520 32370 27532
rect 32401 27523 32459 27529
rect 32401 27520 32413 27523
rect 32364 27492 32413 27520
rect 32364 27480 32370 27492
rect 32401 27489 32413 27492
rect 32447 27489 32459 27523
rect 32582 27520 32588 27532
rect 32543 27492 32588 27520
rect 32401 27483 32459 27489
rect 31202 27452 31208 27464
rect 31087 27424 31208 27452
rect 28399 27421 28411 27424
rect 28353 27415 28411 27421
rect 31202 27412 31208 27424
rect 31260 27412 31266 27464
rect 32416 27452 32444 27483
rect 32582 27480 32588 27492
rect 32640 27480 32646 27532
rect 34054 27480 34060 27532
rect 34112 27520 34118 27532
rect 34698 27529 34704 27532
rect 34644 27523 34704 27529
rect 34644 27520 34656 27523
rect 34112 27492 34656 27520
rect 34112 27480 34118 27492
rect 34644 27489 34656 27492
rect 34690 27489 34704 27523
rect 34644 27483 34704 27489
rect 34698 27480 34704 27483
rect 34756 27480 34762 27532
rect 36170 27520 36176 27532
rect 36131 27492 36176 27520
rect 36170 27480 36176 27492
rect 36228 27480 36234 27532
rect 36541 27523 36599 27529
rect 36541 27489 36553 27523
rect 36587 27520 36599 27523
rect 37090 27520 37096 27532
rect 36587 27492 37096 27520
rect 36587 27489 36599 27492
rect 36541 27483 36599 27489
rect 32858 27452 32864 27464
rect 32416 27424 32864 27452
rect 32858 27412 32864 27424
rect 32916 27412 32922 27464
rect 35710 27412 35716 27464
rect 35768 27452 35774 27464
rect 36556 27452 36584 27483
rect 37090 27480 37096 27492
rect 37148 27480 37154 27532
rect 37553 27523 37611 27529
rect 37553 27489 37565 27523
rect 37599 27520 37611 27523
rect 38930 27520 38936 27532
rect 37599 27492 38936 27520
rect 37599 27489 37611 27492
rect 37553 27483 37611 27489
rect 38930 27480 38936 27492
rect 38988 27480 38994 27532
rect 41046 27480 41052 27532
rect 41104 27520 41110 27532
rect 41141 27523 41199 27529
rect 41141 27520 41153 27523
rect 41104 27492 41153 27520
rect 41104 27480 41110 27492
rect 41141 27489 41153 27492
rect 41187 27489 41199 27523
rect 41141 27483 41199 27489
rect 35768 27424 36584 27452
rect 36817 27455 36875 27461
rect 35768 27412 35774 27424
rect 36817 27421 36829 27455
rect 36863 27452 36875 27455
rect 37458 27452 37464 27464
rect 36863 27424 37464 27452
rect 36863 27421 36875 27424
rect 36817 27415 36875 27421
rect 37458 27412 37464 27424
rect 37516 27452 37522 27464
rect 37737 27455 37795 27461
rect 37737 27452 37749 27455
rect 37516 27424 37749 27452
rect 37516 27412 37522 27424
rect 37737 27421 37749 27424
rect 37783 27421 37795 27455
rect 37737 27415 37795 27421
rect 39853 27455 39911 27461
rect 39853 27421 39865 27455
rect 39899 27421 39911 27455
rect 43898 27452 43904 27464
rect 43859 27424 43904 27452
rect 39853 27415 39911 27421
rect 23290 27384 23296 27396
rect 12308 27356 14320 27384
rect 23251 27356 23296 27384
rect 12308 27344 12314 27356
rect 23290 27344 23296 27356
rect 23348 27344 23354 27396
rect 28718 27344 28724 27396
rect 28776 27384 28782 27396
rect 36630 27384 36636 27396
rect 28776 27356 36636 27384
rect 28776 27344 28782 27356
rect 36630 27344 36636 27356
rect 36688 27344 36694 27396
rect 39206 27344 39212 27396
rect 39264 27384 39270 27396
rect 39868 27384 39896 27415
rect 43898 27412 43904 27424
rect 43956 27412 43962 27464
rect 44545 27455 44603 27461
rect 44545 27421 44557 27455
rect 44591 27452 44603 27455
rect 44818 27452 44824 27464
rect 44591 27424 44824 27452
rect 44591 27421 44603 27424
rect 44545 27415 44603 27421
rect 44818 27412 44824 27424
rect 44876 27412 44882 27464
rect 45741 27455 45799 27461
rect 45741 27421 45753 27455
rect 45787 27421 45799 27455
rect 45741 27415 45799 27421
rect 39264 27356 39896 27384
rect 39264 27344 39270 27356
rect 43806 27344 43812 27396
rect 43864 27384 43870 27396
rect 45756 27384 45784 27415
rect 43864 27356 45784 27384
rect 43864 27344 43870 27356
rect 9769 27319 9827 27325
rect 9769 27285 9781 27319
rect 9815 27316 9827 27319
rect 9950 27316 9956 27328
rect 9815 27288 9956 27316
rect 9815 27285 9827 27288
rect 9769 27279 9827 27285
rect 9950 27276 9956 27288
rect 10008 27276 10014 27328
rect 10594 27276 10600 27328
rect 10652 27316 10658 27328
rect 10689 27319 10747 27325
rect 10689 27316 10701 27319
rect 10652 27288 10701 27316
rect 10652 27276 10658 27288
rect 10689 27285 10701 27288
rect 10735 27285 10747 27319
rect 12066 27316 12072 27328
rect 12027 27288 12072 27316
rect 10689 27279 10747 27285
rect 12066 27276 12072 27288
rect 12124 27276 12130 27328
rect 13078 27316 13084 27328
rect 13039 27288 13084 27316
rect 13078 27276 13084 27288
rect 13136 27276 13142 27328
rect 15102 27316 15108 27328
rect 15063 27288 15108 27316
rect 15102 27276 15108 27288
rect 15160 27276 15166 27328
rect 18141 27319 18199 27325
rect 18141 27285 18153 27319
rect 18187 27316 18199 27319
rect 18230 27316 18236 27328
rect 18187 27288 18236 27316
rect 18187 27285 18199 27288
rect 18141 27279 18199 27285
rect 18230 27276 18236 27288
rect 18288 27276 18294 27328
rect 24811 27319 24869 27325
rect 24811 27285 24823 27319
rect 24857 27316 24869 27319
rect 24946 27316 24952 27328
rect 24857 27288 24952 27316
rect 24857 27285 24869 27288
rect 24811 27279 24869 27285
rect 24946 27276 24952 27288
rect 25004 27276 25010 27328
rect 27154 27276 27160 27328
rect 27212 27316 27218 27328
rect 27387 27319 27445 27325
rect 27387 27316 27399 27319
rect 27212 27288 27399 27316
rect 27212 27276 27218 27288
rect 27387 27285 27399 27288
rect 27433 27285 27445 27319
rect 27387 27279 27445 27285
rect 27525 27319 27583 27325
rect 27525 27285 27537 27319
rect 27571 27316 27583 27319
rect 27614 27316 27620 27328
rect 27571 27288 27620 27316
rect 27571 27285 27583 27288
rect 27525 27279 27583 27285
rect 27614 27276 27620 27288
rect 27672 27276 27678 27328
rect 30190 27316 30196 27328
rect 30151 27288 30196 27316
rect 30190 27276 30196 27288
rect 30248 27276 30254 27328
rect 34747 27319 34805 27325
rect 34747 27285 34759 27319
rect 34793 27316 34805 27319
rect 36722 27316 36728 27328
rect 34793 27288 36728 27316
rect 34793 27285 34805 27288
rect 34747 27279 34805 27285
rect 36722 27276 36728 27288
rect 36780 27276 36786 27328
rect 40218 27276 40224 27328
rect 40276 27316 40282 27328
rect 40497 27319 40555 27325
rect 40497 27316 40509 27319
rect 40276 27288 40509 27316
rect 40276 27276 40282 27288
rect 40497 27285 40509 27288
rect 40543 27285 40555 27319
rect 42058 27316 42064 27328
rect 42019 27288 42064 27316
rect 40497 27279 40555 27285
rect 42058 27276 42064 27288
rect 42116 27276 42122 27328
rect 43622 27316 43628 27328
rect 43583 27288 43628 27316
rect 43622 27276 43628 27288
rect 43680 27276 43686 27328
rect 1104 27226 48852 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 48852 27226
rect 1104 27152 48852 27174
rect 10870 27072 10876 27124
rect 10928 27112 10934 27124
rect 11425 27115 11483 27121
rect 11425 27112 11437 27115
rect 10928 27084 11437 27112
rect 10928 27072 10934 27084
rect 11425 27081 11437 27084
rect 11471 27081 11483 27115
rect 12158 27112 12164 27124
rect 12119 27084 12164 27112
rect 11425 27075 11483 27081
rect 12158 27072 12164 27084
rect 12216 27112 12222 27124
rect 12216 27084 12572 27112
rect 12216 27072 12222 27084
rect 10502 27004 10508 27056
rect 10560 27044 10566 27056
rect 11146 27044 11152 27056
rect 10560 27016 10640 27044
rect 11059 27016 11152 27044
rect 10560 27004 10566 27016
rect 10612 26985 10640 27016
rect 11146 27004 11152 27016
rect 11204 27044 11210 27056
rect 11330 27044 11336 27056
rect 11204 27016 11336 27044
rect 11204 27004 11210 27016
rect 11330 27004 11336 27016
rect 11388 27004 11394 27056
rect 12544 26985 12572 27084
rect 13814 27072 13820 27124
rect 13872 27112 13878 27124
rect 13872 27084 13917 27112
rect 13872 27072 13878 27084
rect 15102 27072 15108 27124
rect 15160 27112 15166 27124
rect 16623 27115 16681 27121
rect 16623 27112 16635 27115
rect 15160 27084 16635 27112
rect 15160 27072 15166 27084
rect 16623 27081 16635 27084
rect 16669 27081 16681 27115
rect 16623 27075 16681 27081
rect 17218 27072 17224 27124
rect 17276 27112 17282 27124
rect 17405 27115 17463 27121
rect 17405 27112 17417 27115
rect 17276 27084 17417 27112
rect 17276 27072 17282 27084
rect 17405 27081 17417 27084
rect 17451 27112 17463 27115
rect 18782 27112 18788 27124
rect 17451 27084 18788 27112
rect 17451 27081 17463 27084
rect 17405 27075 17463 27081
rect 18782 27072 18788 27084
rect 18840 27072 18846 27124
rect 19150 27072 19156 27124
rect 19208 27112 19214 27124
rect 19337 27115 19395 27121
rect 19337 27112 19349 27115
rect 19208 27084 19349 27112
rect 19208 27072 19214 27084
rect 19337 27081 19349 27084
rect 19383 27112 19395 27115
rect 20027 27115 20085 27121
rect 20027 27112 20039 27115
rect 19383 27084 20039 27112
rect 19383 27081 19395 27084
rect 19337 27075 19395 27081
rect 20027 27081 20039 27084
rect 20073 27081 20085 27115
rect 20027 27075 20085 27081
rect 20165 27115 20223 27121
rect 20165 27081 20177 27115
rect 20211 27112 20223 27115
rect 20438 27112 20444 27124
rect 20211 27084 20444 27112
rect 20211 27081 20223 27084
rect 20165 27075 20223 27081
rect 20438 27072 20444 27084
rect 20496 27072 20502 27124
rect 22741 27115 22799 27121
rect 22741 27081 22753 27115
rect 22787 27112 22799 27115
rect 23014 27112 23020 27124
rect 22787 27084 23020 27112
rect 22787 27081 22799 27084
rect 22741 27075 22799 27081
rect 23014 27072 23020 27084
rect 23072 27072 23078 27124
rect 24486 27072 24492 27124
rect 24544 27112 24550 27124
rect 24854 27112 24860 27124
rect 24544 27084 24860 27112
rect 24544 27072 24550 27084
rect 24854 27072 24860 27084
rect 24912 27072 24918 27124
rect 27614 27072 27620 27124
rect 27672 27112 27678 27124
rect 27893 27115 27951 27121
rect 27893 27112 27905 27115
rect 27672 27084 27905 27112
rect 27672 27072 27678 27084
rect 27893 27081 27905 27084
rect 27939 27081 27951 27115
rect 27893 27075 27951 27081
rect 28718 27072 28724 27124
rect 28776 27112 28782 27124
rect 28813 27115 28871 27121
rect 28813 27112 28825 27115
rect 28776 27084 28825 27112
rect 28776 27072 28782 27084
rect 28813 27081 28825 27084
rect 28859 27081 28871 27115
rect 28813 27075 28871 27081
rect 29362 27072 29368 27124
rect 29420 27112 29426 27124
rect 29549 27115 29607 27121
rect 29549 27112 29561 27115
rect 29420 27084 29561 27112
rect 29420 27072 29426 27084
rect 29549 27081 29561 27084
rect 29595 27112 29607 27115
rect 31757 27115 31815 27121
rect 31757 27112 31769 27115
rect 29595 27084 31769 27112
rect 29595 27081 29607 27084
rect 29549 27075 29607 27081
rect 31757 27081 31769 27084
rect 31803 27112 31815 27115
rect 32582 27112 32588 27124
rect 31803 27084 32588 27112
rect 31803 27081 31815 27084
rect 31757 27075 31815 27081
rect 32582 27072 32588 27084
rect 32640 27072 32646 27124
rect 34698 27112 34704 27124
rect 34659 27084 34704 27112
rect 34698 27072 34704 27084
rect 34756 27072 34762 27124
rect 35710 27112 35716 27124
rect 35671 27084 35716 27112
rect 35710 27072 35716 27084
rect 35768 27072 35774 27124
rect 37829 27115 37887 27121
rect 37829 27081 37841 27115
rect 37875 27112 37887 27115
rect 38102 27112 38108 27124
rect 37875 27084 38108 27112
rect 37875 27081 37887 27084
rect 37829 27075 37887 27081
rect 38102 27072 38108 27084
rect 38160 27072 38166 27124
rect 39482 27112 39488 27124
rect 39443 27084 39488 27112
rect 39482 27072 39488 27084
rect 39540 27072 39546 27124
rect 39574 27072 39580 27124
rect 39632 27112 39638 27124
rect 39853 27115 39911 27121
rect 39853 27112 39865 27115
rect 39632 27084 39865 27112
rect 39632 27072 39638 27084
rect 39853 27081 39865 27084
rect 39899 27081 39911 27115
rect 41506 27112 41512 27124
rect 41467 27084 41512 27112
rect 39853 27075 39911 27081
rect 41506 27072 41512 27084
rect 41564 27072 41570 27124
rect 41969 27115 42027 27121
rect 41969 27081 41981 27115
rect 42015 27112 42027 27115
rect 42058 27112 42064 27124
rect 42015 27084 42064 27112
rect 42015 27081 42027 27084
rect 41969 27075 42027 27081
rect 42058 27072 42064 27084
rect 42116 27072 42122 27124
rect 45462 27072 45468 27124
rect 45520 27112 45526 27124
rect 45741 27115 45799 27121
rect 45741 27112 45753 27115
rect 45520 27084 45753 27112
rect 45520 27072 45526 27084
rect 45741 27081 45753 27084
rect 45787 27081 45799 27115
rect 45741 27075 45799 27081
rect 12710 27004 12716 27056
rect 12768 27044 12774 27056
rect 17037 27047 17095 27053
rect 12768 27016 16563 27044
rect 12768 27004 12774 27016
rect 10597 26979 10655 26985
rect 10597 26945 10609 26979
rect 10643 26945 10655 26979
rect 10597 26939 10655 26945
rect 12529 26979 12587 26985
rect 12529 26945 12541 26979
rect 12575 26945 12587 26979
rect 12802 26976 12808 26988
rect 12763 26948 12808 26976
rect 12529 26939 12587 26945
rect 12802 26936 12808 26948
rect 12860 26936 12866 26988
rect 15010 26976 15016 26988
rect 14971 26948 15016 26976
rect 15010 26936 15016 26948
rect 15068 26936 15074 26988
rect 15654 26976 15660 26988
rect 15615 26948 15660 26976
rect 15654 26936 15660 26948
rect 15712 26936 15718 26988
rect 9858 26868 9864 26920
rect 9916 26908 9922 26920
rect 10045 26911 10103 26917
rect 10045 26908 10057 26911
rect 9916 26880 10057 26908
rect 9916 26868 9922 26880
rect 10045 26877 10057 26880
rect 10091 26908 10103 26911
rect 10410 26908 10416 26920
rect 10091 26880 10416 26908
rect 10091 26877 10103 26880
rect 10045 26871 10103 26877
rect 10410 26868 10416 26880
rect 10468 26868 10474 26920
rect 16535 26917 16563 27016
rect 17037 27013 17049 27047
rect 17083 27044 17095 27047
rect 20990 27044 20996 27056
rect 17083 27016 20996 27044
rect 17083 27013 17095 27016
rect 17037 27007 17095 27013
rect 10505 26911 10563 26917
rect 10505 26877 10517 26911
rect 10551 26877 10563 26911
rect 16535 26911 16610 26917
rect 16535 26880 16564 26911
rect 10505 26871 10563 26877
rect 16552 26877 16564 26880
rect 16598 26908 16610 26911
rect 17052 26908 17080 27007
rect 20990 27004 20996 27016
rect 21048 27004 21054 27056
rect 22554 27004 22560 27056
rect 22612 27044 22618 27056
rect 23385 27047 23443 27053
rect 23385 27044 23397 27047
rect 22612 27016 23397 27044
rect 22612 27004 22618 27016
rect 23385 27013 23397 27016
rect 23431 27013 23443 27047
rect 23385 27007 23443 27013
rect 25222 27004 25228 27056
rect 25280 27044 25286 27056
rect 25593 27047 25651 27053
rect 25593 27044 25605 27047
rect 25280 27016 25605 27044
rect 25280 27004 25286 27016
rect 25593 27013 25605 27016
rect 25639 27044 25651 27047
rect 25958 27044 25964 27056
rect 25639 27016 25964 27044
rect 25639 27013 25651 27016
rect 25593 27007 25651 27013
rect 25958 27004 25964 27016
rect 26016 27004 26022 27056
rect 26050 27004 26056 27056
rect 26108 27044 26114 27056
rect 26786 27044 26792 27056
rect 26108 27016 26792 27044
rect 26108 27004 26114 27016
rect 26786 27004 26792 27016
rect 26844 27044 26850 27056
rect 30009 27047 30067 27053
rect 26844 27016 26924 27044
rect 26844 27004 26850 27016
rect 19797 26979 19855 26985
rect 19797 26945 19809 26979
rect 19843 26976 19855 26979
rect 20257 26979 20315 26985
rect 20257 26976 20269 26979
rect 19843 26948 20269 26976
rect 19843 26945 19855 26948
rect 19797 26939 19855 26945
rect 20257 26945 20269 26948
rect 20303 26976 20315 26979
rect 20898 26976 20904 26988
rect 20303 26948 20904 26976
rect 20303 26945 20315 26948
rect 20257 26939 20315 26945
rect 20898 26936 20904 26948
rect 20956 26936 20962 26988
rect 21818 26976 21824 26988
rect 21779 26948 21824 26976
rect 21818 26936 21824 26948
rect 21876 26936 21882 26988
rect 24213 26979 24271 26985
rect 24213 26945 24225 26979
rect 24259 26976 24271 26979
rect 26605 26979 26663 26985
rect 26605 26976 26617 26979
rect 24259 26948 26617 26976
rect 24259 26945 24271 26948
rect 24213 26939 24271 26945
rect 26605 26945 26617 26948
rect 26651 26976 26663 26979
rect 26694 26976 26700 26988
rect 26651 26948 26700 26976
rect 26651 26945 26663 26948
rect 26605 26939 26663 26945
rect 26694 26936 26700 26948
rect 26752 26936 26758 26988
rect 26896 26985 26924 27016
rect 30009 27013 30021 27047
rect 30055 27044 30067 27047
rect 32122 27044 32128 27056
rect 30055 27016 32128 27044
rect 30055 27013 30067 27016
rect 30009 27007 30067 27013
rect 26881 26979 26939 26985
rect 26881 26945 26893 26979
rect 26927 26945 26939 26979
rect 26881 26939 26939 26945
rect 18049 26911 18107 26917
rect 18049 26908 18061 26911
rect 16598 26880 17080 26908
rect 17880 26880 18061 26908
rect 16598 26877 16610 26880
rect 16552 26871 16610 26877
rect 9585 26843 9643 26849
rect 9585 26809 9597 26843
rect 9631 26840 9643 26843
rect 10520 26840 10548 26871
rect 10594 26840 10600 26852
rect 9631 26812 10600 26840
rect 9631 26809 9643 26812
rect 9585 26803 9643 26809
rect 10594 26800 10600 26812
rect 10652 26800 10658 26852
rect 12618 26840 12624 26852
rect 12579 26812 12624 26840
rect 12618 26800 12624 26812
rect 12676 26800 12682 26852
rect 13262 26800 13268 26852
rect 13320 26840 13326 26852
rect 14737 26843 14795 26849
rect 14737 26840 14749 26843
rect 13320 26812 14749 26840
rect 13320 26800 13326 26812
rect 14737 26809 14749 26812
rect 14783 26840 14795 26843
rect 15105 26843 15163 26849
rect 15105 26840 15117 26843
rect 14783 26812 15117 26840
rect 14783 26809 14795 26812
rect 14737 26803 14795 26809
rect 15105 26809 15117 26812
rect 15151 26809 15163 26843
rect 15105 26803 15163 26809
rect 9950 26772 9956 26784
rect 9911 26744 9956 26772
rect 9950 26732 9956 26744
rect 10008 26732 10014 26784
rect 12636 26772 12664 26800
rect 13449 26775 13507 26781
rect 13449 26772 13461 26775
rect 12636 26744 13461 26772
rect 13449 26741 13461 26744
rect 13495 26741 13507 26775
rect 15120 26772 15148 26803
rect 17880 26784 17908 26880
rect 18049 26877 18061 26880
rect 18095 26877 18107 26911
rect 18049 26871 18107 26877
rect 18230 26868 18236 26920
rect 18288 26908 18294 26920
rect 18509 26911 18567 26917
rect 18509 26908 18521 26911
rect 18288 26880 18521 26908
rect 18288 26868 18294 26880
rect 18509 26877 18521 26880
rect 18555 26877 18567 26911
rect 18509 26871 18567 26877
rect 19889 26911 19947 26917
rect 19889 26877 19901 26911
rect 19935 26908 19947 26911
rect 20070 26908 20076 26920
rect 19935 26880 20076 26908
rect 19935 26877 19947 26880
rect 19889 26871 19947 26877
rect 20070 26868 20076 26880
rect 20128 26868 20134 26920
rect 24004 26911 24062 26917
rect 24004 26877 24016 26911
rect 24050 26908 24062 26911
rect 24394 26908 24400 26920
rect 24050 26880 24400 26908
rect 24050 26877 24062 26880
rect 24004 26871 24062 26877
rect 24394 26868 24400 26880
rect 24452 26868 24458 26920
rect 28128 26911 28186 26917
rect 28128 26877 28140 26911
rect 28174 26908 28186 26911
rect 28350 26908 28356 26920
rect 28174 26880 28356 26908
rect 28174 26877 28186 26880
rect 28128 26871 28186 26877
rect 28350 26868 28356 26880
rect 28408 26868 28414 26920
rect 29086 26868 29092 26920
rect 29144 26908 29150 26920
rect 30116 26917 30144 27016
rect 32122 27004 32128 27016
rect 32180 27044 32186 27056
rect 39758 27044 39764 27056
rect 32180 27016 32530 27044
rect 32180 27004 32186 27016
rect 32398 26976 32404 26988
rect 32359 26948 32404 26976
rect 32398 26936 32404 26948
rect 32456 26936 32462 26988
rect 32502 26976 32530 27016
rect 33152 27016 39764 27044
rect 33152 26976 33180 27016
rect 39758 27004 39764 27016
rect 39816 27004 39822 27056
rect 33502 26976 33508 26988
rect 32502 26948 33180 26976
rect 33244 26948 33508 26976
rect 30101 26911 30159 26917
rect 30101 26908 30113 26911
rect 29144 26880 30113 26908
rect 29144 26868 29150 26880
rect 30101 26877 30113 26880
rect 30147 26877 30159 26911
rect 30101 26871 30159 26877
rect 30190 26868 30196 26920
rect 30248 26908 30254 26920
rect 30653 26911 30711 26917
rect 30653 26908 30665 26911
rect 30248 26880 30665 26908
rect 30248 26868 30254 26880
rect 30653 26877 30665 26880
rect 30699 26908 30711 26911
rect 30699 26880 30972 26908
rect 30699 26877 30711 26880
rect 30653 26871 30711 26877
rect 22142 26843 22200 26849
rect 22142 26809 22154 26843
rect 22188 26809 22200 26843
rect 22142 26803 22200 26809
rect 15470 26772 15476 26784
rect 15120 26744 15476 26772
rect 13449 26735 13507 26741
rect 15470 26732 15476 26744
rect 15528 26772 15534 26784
rect 15933 26775 15991 26781
rect 15933 26772 15945 26775
rect 15528 26744 15945 26772
rect 15528 26732 15534 26744
rect 15933 26741 15945 26744
rect 15979 26741 15991 26775
rect 17862 26772 17868 26784
rect 17823 26744 17868 26772
rect 15933 26735 15991 26741
rect 17862 26732 17868 26744
rect 17920 26732 17926 26784
rect 18138 26772 18144 26784
rect 18099 26744 18144 26772
rect 18138 26732 18144 26744
rect 18196 26732 18202 26784
rect 20530 26772 20536 26784
rect 20491 26744 20536 26772
rect 20530 26732 20536 26744
rect 20588 26732 20594 26784
rect 21082 26772 21088 26784
rect 21043 26744 21088 26772
rect 21082 26732 21088 26744
rect 21140 26732 21146 26784
rect 21450 26732 21456 26784
rect 21508 26772 21514 26784
rect 21729 26775 21787 26781
rect 21729 26772 21741 26775
rect 21508 26744 21741 26772
rect 21508 26732 21514 26744
rect 21729 26741 21741 26744
rect 21775 26772 21787 26775
rect 22157 26772 22185 26803
rect 24854 26800 24860 26852
rect 24912 26840 24918 26852
rect 25041 26843 25099 26849
rect 25041 26840 25053 26843
rect 24912 26812 25053 26840
rect 24912 26800 24918 26812
rect 25041 26809 25053 26812
rect 25087 26809 25099 26843
rect 25041 26803 25099 26809
rect 25130 26800 25136 26852
rect 25188 26840 25194 26852
rect 26697 26843 26755 26849
rect 26697 26840 26709 26843
rect 25188 26812 25233 26840
rect 25976 26812 26709 26840
rect 25188 26800 25194 26812
rect 22738 26772 22744 26784
rect 21775 26744 22744 26772
rect 21775 26741 21787 26744
rect 21729 26735 21787 26741
rect 22738 26732 22744 26744
rect 22796 26732 22802 26784
rect 25148 26772 25176 26800
rect 25976 26781 26004 26812
rect 26697 26809 26709 26812
rect 26743 26809 26755 26843
rect 26697 26803 26755 26809
rect 26970 26800 26976 26852
rect 27028 26840 27034 26852
rect 28215 26843 28273 26849
rect 28215 26840 28227 26843
rect 27028 26812 28227 26840
rect 27028 26800 27034 26812
rect 28215 26809 28227 26812
rect 28261 26809 28273 26843
rect 30834 26840 30840 26852
rect 30795 26812 30840 26840
rect 28215 26803 28273 26809
rect 30834 26800 30840 26812
rect 30892 26800 30898 26852
rect 30944 26840 30972 26880
rect 31662 26868 31668 26920
rect 31720 26908 31726 26920
rect 31916 26911 31974 26917
rect 31916 26908 31928 26911
rect 31720 26880 31928 26908
rect 31720 26868 31726 26880
rect 31916 26877 31928 26880
rect 31962 26908 31974 26911
rect 32416 26908 32444 26936
rect 33244 26917 33272 26948
rect 33502 26936 33508 26948
rect 33560 26976 33566 26988
rect 33870 26976 33876 26988
rect 33560 26948 33876 26976
rect 33560 26936 33566 26948
rect 33870 26936 33876 26948
rect 33928 26976 33934 26988
rect 38289 26979 38347 26985
rect 33928 26948 37872 26976
rect 33928 26936 33934 26948
rect 31962 26880 32444 26908
rect 33137 26911 33195 26917
rect 31962 26877 31974 26880
rect 31916 26871 31974 26877
rect 33137 26877 33149 26911
rect 33183 26908 33195 26911
rect 33229 26911 33287 26917
rect 33229 26908 33241 26911
rect 33183 26880 33241 26908
rect 33183 26877 33195 26880
rect 33137 26871 33195 26877
rect 33229 26877 33241 26880
rect 33275 26877 33287 26911
rect 33229 26871 33287 26877
rect 33318 26868 33324 26920
rect 33376 26908 33382 26920
rect 33689 26911 33747 26917
rect 33689 26908 33701 26911
rect 33376 26880 33701 26908
rect 33376 26868 33382 26880
rect 33689 26877 33701 26880
rect 33735 26877 33747 26911
rect 33689 26871 33747 26877
rect 36633 26911 36691 26917
rect 36633 26877 36645 26911
rect 36679 26877 36691 26911
rect 37090 26908 37096 26920
rect 37051 26880 37096 26908
rect 36633 26871 36691 26877
rect 33336 26840 33364 26868
rect 33962 26840 33968 26852
rect 30944 26812 33364 26840
rect 33923 26812 33968 26840
rect 33962 26800 33968 26812
rect 34020 26800 34026 26852
rect 36446 26840 36452 26852
rect 36407 26812 36452 26840
rect 36446 26800 36452 26812
rect 36504 26840 36510 26852
rect 36648 26840 36676 26871
rect 37090 26868 37096 26880
rect 37148 26868 37154 26920
rect 37366 26840 37372 26852
rect 36504 26812 36676 26840
rect 37327 26812 37372 26840
rect 36504 26800 36510 26812
rect 37366 26800 37372 26812
rect 37424 26800 37430 26852
rect 25961 26775 26019 26781
rect 25961 26772 25973 26775
rect 25148 26744 25973 26772
rect 25961 26741 25973 26744
rect 26007 26741 26019 26775
rect 25961 26735 26019 26741
rect 26421 26775 26479 26781
rect 26421 26741 26433 26775
rect 26467 26772 26479 26775
rect 27246 26772 27252 26784
rect 26467 26744 27252 26772
rect 26467 26741 26479 26744
rect 26421 26735 26479 26741
rect 27246 26732 27252 26744
rect 27304 26732 27310 26784
rect 27522 26772 27528 26784
rect 27483 26744 27528 26772
rect 27522 26732 27528 26744
rect 27580 26732 27586 26784
rect 31202 26772 31208 26784
rect 31163 26744 31208 26772
rect 31202 26732 31208 26744
rect 31260 26732 31266 26784
rect 31987 26775 32045 26781
rect 31987 26741 31999 26775
rect 32033 26772 32045 26775
rect 32214 26772 32220 26784
rect 32033 26744 32220 26772
rect 32033 26741 32045 26744
rect 31987 26735 32045 26741
rect 32214 26732 32220 26744
rect 32272 26732 32278 26784
rect 32769 26775 32827 26781
rect 32769 26741 32781 26775
rect 32815 26772 32827 26775
rect 32858 26772 32864 26784
rect 32815 26744 32864 26772
rect 32815 26741 32827 26744
rect 32769 26735 32827 26741
rect 32858 26732 32864 26744
rect 32916 26732 32922 26784
rect 34882 26772 34888 26784
rect 34843 26744 34888 26772
rect 34882 26732 34888 26744
rect 34940 26732 34946 26784
rect 36170 26772 36176 26784
rect 36131 26744 36176 26772
rect 36170 26732 36176 26744
rect 36228 26732 36234 26784
rect 37844 26772 37872 26948
rect 38289 26945 38301 26979
rect 38335 26976 38347 26979
rect 38930 26976 38936 26988
rect 38335 26948 38936 26976
rect 38335 26945 38347 26948
rect 38289 26939 38347 26945
rect 38930 26936 38936 26948
rect 38988 26936 38994 26988
rect 40218 26936 40224 26988
rect 40276 26976 40282 26988
rect 41233 26979 41291 26985
rect 40276 26948 41000 26976
rect 40276 26936 40282 26948
rect 40972 26917 41000 26948
rect 41233 26945 41245 26979
rect 41279 26976 41291 26979
rect 41322 26976 41328 26988
rect 41279 26948 41328 26976
rect 41279 26945 41291 26948
rect 41233 26939 41291 26945
rect 41322 26936 41328 26948
rect 41380 26936 41386 26988
rect 42153 26979 42211 26985
rect 42153 26945 42165 26979
rect 42199 26976 42211 26979
rect 42242 26976 42248 26988
rect 42199 26948 42248 26976
rect 42199 26945 42211 26948
rect 42153 26939 42211 26945
rect 42242 26936 42248 26948
rect 42300 26936 42306 26988
rect 42426 26976 42432 26988
rect 42387 26948 42432 26976
rect 42426 26936 42432 26948
rect 42484 26936 42490 26988
rect 43993 26979 44051 26985
rect 43993 26976 44005 26979
rect 42812 26948 44005 26976
rect 40313 26911 40371 26917
rect 40313 26877 40325 26911
rect 40359 26908 40371 26911
rect 40497 26911 40555 26917
rect 40497 26908 40509 26911
rect 40359 26880 40509 26908
rect 40359 26877 40371 26880
rect 40313 26871 40371 26877
rect 40497 26877 40509 26880
rect 40543 26877 40555 26911
rect 40497 26871 40555 26877
rect 40957 26911 41015 26917
rect 40957 26877 40969 26911
rect 41003 26877 41015 26911
rect 40957 26871 41015 26877
rect 38381 26843 38439 26849
rect 38381 26809 38393 26843
rect 38427 26840 38439 26843
rect 38654 26840 38660 26852
rect 38427 26812 38660 26840
rect 38427 26809 38439 26812
rect 38381 26803 38439 26809
rect 38654 26800 38660 26812
rect 38712 26800 38718 26852
rect 38933 26843 38991 26849
rect 38933 26809 38945 26843
rect 38979 26840 38991 26843
rect 39114 26840 39120 26852
rect 38979 26812 39120 26840
rect 38979 26809 38991 26812
rect 38933 26803 38991 26809
rect 39114 26800 39120 26812
rect 39172 26800 39178 26852
rect 40328 26772 40356 26871
rect 42245 26843 42303 26849
rect 42245 26809 42257 26843
rect 42291 26840 42303 26843
rect 42812 26840 42840 26948
rect 43993 26945 44005 26948
rect 44039 26976 44051 26979
rect 44266 26976 44272 26988
rect 44039 26948 44272 26976
rect 44039 26945 44051 26948
rect 43993 26939 44051 26945
rect 44266 26936 44272 26948
rect 44324 26976 44330 26988
rect 45465 26979 45523 26985
rect 45465 26976 45477 26979
rect 44324 26948 45477 26976
rect 44324 26936 44330 26948
rect 45465 26945 45477 26948
rect 45511 26976 45523 26979
rect 45554 26976 45560 26988
rect 45511 26948 45560 26976
rect 45511 26945 45523 26948
rect 45465 26939 45523 26945
rect 45554 26936 45560 26948
rect 45612 26936 45618 26988
rect 42291 26812 42840 26840
rect 43257 26843 43315 26849
rect 42291 26809 42303 26812
rect 42245 26803 42303 26809
rect 43257 26809 43269 26843
rect 43303 26840 43315 26843
rect 44174 26840 44180 26852
rect 43303 26812 44180 26840
rect 43303 26809 43315 26812
rect 43257 26803 43315 26809
rect 37844 26744 40356 26772
rect 42058 26732 42064 26784
rect 42116 26772 42122 26784
rect 42260 26772 42288 26803
rect 44174 26800 44180 26812
rect 44232 26800 44238 26852
rect 44266 26800 44272 26852
rect 44324 26840 44330 26852
rect 44818 26840 44824 26852
rect 44324 26812 44369 26840
rect 44779 26812 44824 26840
rect 44324 26800 44330 26812
rect 44818 26800 44824 26812
rect 44876 26800 44882 26852
rect 43622 26772 43628 26784
rect 42116 26744 42288 26772
rect 43583 26744 43628 26772
rect 42116 26732 42122 26744
rect 43622 26732 43628 26744
rect 43680 26732 43686 26784
rect 1104 26682 48852 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 48852 26682
rect 1104 26608 48852 26630
rect 13078 26528 13084 26580
rect 13136 26568 13142 26580
rect 13219 26571 13277 26577
rect 13219 26568 13231 26571
rect 13136 26540 13231 26568
rect 13136 26528 13142 26540
rect 13219 26537 13231 26540
rect 13265 26537 13277 26571
rect 15010 26568 15016 26580
rect 14971 26540 15016 26568
rect 13219 26531 13277 26537
rect 15010 26528 15016 26540
rect 15068 26528 15074 26580
rect 15378 26528 15384 26580
rect 15436 26568 15442 26580
rect 15473 26571 15531 26577
rect 15473 26568 15485 26571
rect 15436 26540 15485 26568
rect 15436 26528 15442 26540
rect 15473 26537 15485 26540
rect 15519 26537 15531 26571
rect 15473 26531 15531 26537
rect 16942 26528 16948 26580
rect 17000 26568 17006 26580
rect 17037 26571 17095 26577
rect 17037 26568 17049 26571
rect 17000 26540 17049 26568
rect 17000 26528 17006 26540
rect 17037 26537 17049 26540
rect 17083 26537 17095 26571
rect 17037 26531 17095 26537
rect 18693 26571 18751 26577
rect 18693 26537 18705 26571
rect 18739 26568 18751 26571
rect 18782 26568 18788 26580
rect 18739 26540 18788 26568
rect 18739 26537 18751 26540
rect 18693 26531 18751 26537
rect 18782 26528 18788 26540
rect 18840 26528 18846 26580
rect 20070 26528 20076 26580
rect 20128 26568 20134 26580
rect 20257 26571 20315 26577
rect 20257 26568 20269 26571
rect 20128 26540 20269 26568
rect 20128 26528 20134 26540
rect 20257 26537 20269 26540
rect 20303 26537 20315 26571
rect 21818 26568 21824 26580
rect 21779 26540 21824 26568
rect 20257 26531 20315 26537
rect 21818 26528 21824 26540
rect 21876 26528 21882 26580
rect 23983 26571 24041 26577
rect 23983 26537 23995 26571
rect 24029 26568 24041 26571
rect 24765 26571 24823 26577
rect 24765 26568 24777 26571
rect 24029 26540 24777 26568
rect 24029 26537 24041 26540
rect 23983 26531 24041 26537
rect 24765 26537 24777 26540
rect 24811 26568 24823 26571
rect 24854 26568 24860 26580
rect 24811 26540 24860 26568
rect 24811 26537 24823 26540
rect 24765 26531 24823 26537
rect 24854 26528 24860 26540
rect 24912 26528 24918 26580
rect 26694 26568 26700 26580
rect 26655 26540 26700 26568
rect 26694 26528 26700 26540
rect 26752 26528 26758 26580
rect 28350 26568 28356 26580
rect 28311 26540 28356 26568
rect 28350 26528 28356 26540
rect 28408 26528 28414 26580
rect 30190 26568 30196 26580
rect 28460 26540 30196 26568
rect 11330 26460 11336 26512
rect 11388 26500 11394 26512
rect 11701 26503 11759 26509
rect 11701 26500 11713 26503
rect 11388 26472 11713 26500
rect 11388 26460 11394 26472
rect 11701 26469 11713 26472
rect 11747 26469 11759 26503
rect 11701 26463 11759 26469
rect 12066 26460 12072 26512
rect 12124 26500 12130 26512
rect 14231 26503 14289 26509
rect 14231 26500 14243 26503
rect 12124 26472 14243 26500
rect 12124 26460 12130 26472
rect 14231 26469 14243 26472
rect 14277 26469 14289 26503
rect 16022 26500 16028 26512
rect 15983 26472 16028 26500
rect 14231 26463 14289 26469
rect 16022 26460 16028 26472
rect 16080 26460 16086 26512
rect 16206 26460 16212 26512
rect 16264 26500 16270 26512
rect 19981 26503 20039 26509
rect 19981 26500 19993 26503
rect 16264 26472 17540 26500
rect 16264 26460 16270 26472
rect 17512 26444 17540 26472
rect 18248 26472 19993 26500
rect 18248 26444 18276 26472
rect 19981 26469 19993 26472
rect 20027 26469 20039 26503
rect 19981 26463 20039 26469
rect 10042 26392 10048 26444
rect 10100 26432 10106 26444
rect 10502 26432 10508 26444
rect 10100 26404 10508 26432
rect 10100 26392 10106 26404
rect 10502 26392 10508 26404
rect 10560 26392 10566 26444
rect 12253 26435 12311 26441
rect 12253 26401 12265 26435
rect 12299 26432 12311 26435
rect 12802 26432 12808 26444
rect 12299 26404 12808 26432
rect 12299 26401 12311 26404
rect 12253 26395 12311 26401
rect 12802 26392 12808 26404
rect 12860 26392 12866 26444
rect 13081 26435 13139 26441
rect 13081 26401 13093 26435
rect 13127 26432 13139 26435
rect 13170 26432 13176 26444
rect 13127 26404 13176 26432
rect 13127 26401 13139 26404
rect 13081 26395 13139 26401
rect 13170 26392 13176 26404
rect 13228 26392 13234 26444
rect 14144 26435 14202 26441
rect 14144 26401 14156 26435
rect 14190 26432 14202 26435
rect 14366 26432 14372 26444
rect 14190 26404 14372 26432
rect 14190 26401 14202 26404
rect 14144 26395 14202 26401
rect 14366 26392 14372 26404
rect 14424 26392 14430 26444
rect 17494 26432 17500 26444
rect 17407 26404 17500 26432
rect 17494 26392 17500 26404
rect 17552 26392 17558 26444
rect 17957 26435 18015 26441
rect 17957 26401 17969 26435
rect 18003 26432 18015 26435
rect 18230 26432 18236 26444
rect 18003 26404 18236 26432
rect 18003 26401 18015 26404
rect 17957 26395 18015 26401
rect 18230 26392 18236 26404
rect 18288 26392 18294 26444
rect 19245 26435 19303 26441
rect 19245 26401 19257 26435
rect 19291 26432 19303 26435
rect 19518 26432 19524 26444
rect 19291 26404 19524 26432
rect 19291 26401 19303 26404
rect 19245 26395 19303 26401
rect 19518 26392 19524 26404
rect 19576 26432 19582 26444
rect 20088 26432 20116 26528
rect 22459 26503 22517 26509
rect 22459 26469 22471 26503
rect 22505 26500 22517 26503
rect 22738 26500 22744 26512
rect 22505 26472 22744 26500
rect 22505 26469 22517 26472
rect 22459 26463 22517 26469
rect 22738 26460 22744 26472
rect 22796 26460 22802 26512
rect 24946 26500 24952 26512
rect 24907 26472 24952 26500
rect 24946 26460 24952 26472
rect 25004 26460 25010 26512
rect 25041 26503 25099 26509
rect 25041 26469 25053 26503
rect 25087 26500 25099 26503
rect 25130 26500 25136 26512
rect 25087 26472 25136 26500
rect 25087 26469 25099 26472
rect 25041 26463 25099 26469
rect 25130 26460 25136 26472
rect 25188 26460 25194 26512
rect 25593 26503 25651 26509
rect 25593 26469 25605 26503
rect 25639 26500 25651 26503
rect 25682 26500 25688 26512
rect 25639 26472 25688 26500
rect 25639 26469 25651 26472
rect 25593 26463 25651 26469
rect 25682 26460 25688 26472
rect 25740 26460 25746 26512
rect 27982 26500 27988 26512
rect 27895 26472 27988 26500
rect 27982 26460 27988 26472
rect 28040 26500 28046 26512
rect 28460 26500 28488 26540
rect 30190 26528 30196 26540
rect 30248 26528 30254 26580
rect 30834 26568 30840 26580
rect 30795 26540 30840 26568
rect 30834 26528 30840 26540
rect 30892 26528 30898 26580
rect 33962 26528 33968 26580
rect 34020 26568 34026 26580
rect 34790 26568 34796 26580
rect 34020 26540 34796 26568
rect 34020 26528 34026 26540
rect 34790 26528 34796 26540
rect 34848 26528 34854 26580
rect 35342 26528 35348 26580
rect 35400 26568 35406 26580
rect 36679 26571 36737 26577
rect 36679 26568 36691 26571
rect 35400 26540 36691 26568
rect 35400 26528 35406 26540
rect 36679 26537 36691 26540
rect 36725 26537 36737 26571
rect 37090 26568 37096 26580
rect 37051 26540 37096 26568
rect 36679 26531 36737 26537
rect 37090 26528 37096 26540
rect 37148 26528 37154 26580
rect 37458 26568 37464 26580
rect 37419 26540 37464 26568
rect 37458 26528 37464 26540
rect 37516 26528 37522 26580
rect 41046 26528 41052 26580
rect 41104 26568 41110 26580
rect 41141 26571 41199 26577
rect 41141 26568 41153 26571
rect 41104 26540 41153 26568
rect 41104 26528 41110 26540
rect 41141 26537 41153 26540
rect 41187 26537 41199 26571
rect 41141 26531 41199 26537
rect 43165 26571 43223 26577
rect 43165 26537 43177 26571
rect 43211 26568 43223 26571
rect 43487 26571 43545 26577
rect 43487 26568 43499 26571
rect 43211 26540 43499 26568
rect 43211 26537 43223 26540
rect 43165 26531 43223 26537
rect 43487 26537 43499 26540
rect 43533 26568 43545 26571
rect 43898 26568 43904 26580
rect 43533 26540 43904 26568
rect 43533 26537 43545 26540
rect 43487 26531 43545 26537
rect 43898 26528 43904 26540
rect 43956 26528 43962 26580
rect 44174 26528 44180 26580
rect 44232 26568 44238 26580
rect 44499 26571 44557 26577
rect 44499 26568 44511 26571
rect 44232 26540 44511 26568
rect 44232 26528 44238 26540
rect 44499 26537 44511 26540
rect 44545 26537 44557 26571
rect 44499 26531 44557 26537
rect 28040 26472 28488 26500
rect 28040 26460 28046 26472
rect 28902 26460 28908 26512
rect 28960 26500 28966 26512
rect 29365 26503 29423 26509
rect 29365 26500 29377 26503
rect 28960 26472 29377 26500
rect 28960 26460 28966 26472
rect 29365 26469 29377 26472
rect 29411 26469 29423 26503
rect 32306 26500 32312 26512
rect 32267 26472 32312 26500
rect 29365 26463 29423 26469
rect 32306 26460 32312 26472
rect 32364 26460 32370 26512
rect 32490 26460 32496 26512
rect 32548 26500 32554 26512
rect 35161 26503 35219 26509
rect 32548 26472 34008 26500
rect 32548 26460 32554 26472
rect 33980 26444 34008 26472
rect 35161 26469 35173 26503
rect 35207 26500 35219 26503
rect 35802 26500 35808 26512
rect 35207 26472 35808 26500
rect 35207 26469 35219 26472
rect 35161 26463 35219 26469
rect 35802 26460 35808 26472
rect 35860 26460 35866 26512
rect 38102 26460 38108 26512
rect 38160 26500 38166 26512
rect 38334 26503 38392 26509
rect 38334 26500 38346 26503
rect 38160 26472 38346 26500
rect 38160 26460 38166 26472
rect 38334 26469 38346 26472
rect 38380 26469 38392 26503
rect 41874 26500 41880 26512
rect 41835 26472 41880 26500
rect 38334 26463 38392 26469
rect 41874 26460 41880 26472
rect 41932 26460 41938 26512
rect 42150 26460 42156 26512
rect 42208 26500 42214 26512
rect 43993 26503 44051 26509
rect 42208 26472 42794 26500
rect 42208 26460 42214 26472
rect 19576 26404 20116 26432
rect 19576 26392 19582 26404
rect 21082 26392 21088 26444
rect 21140 26432 21146 26444
rect 23845 26435 23903 26441
rect 21140 26404 23474 26432
rect 21140 26392 21146 26404
rect 10643 26367 10701 26373
rect 10643 26333 10655 26367
rect 10689 26364 10701 26367
rect 11609 26367 11667 26373
rect 11609 26364 11621 26367
rect 10689 26336 11621 26364
rect 10689 26333 10701 26336
rect 10643 26327 10701 26333
rect 11609 26333 11621 26336
rect 11655 26364 11667 26367
rect 11882 26364 11888 26376
rect 11655 26336 11888 26364
rect 11655 26333 11667 26336
rect 11609 26327 11667 26333
rect 11882 26324 11888 26336
rect 11940 26324 11946 26376
rect 15194 26324 15200 26376
rect 15252 26364 15258 26376
rect 15933 26367 15991 26373
rect 15933 26364 15945 26367
rect 15252 26336 15945 26364
rect 15252 26324 15258 26336
rect 15933 26333 15945 26336
rect 15979 26333 15991 26367
rect 15933 26327 15991 26333
rect 16209 26367 16267 26373
rect 16209 26333 16221 26367
rect 16255 26333 16267 26367
rect 18046 26364 18052 26376
rect 18007 26336 18052 26364
rect 16209 26327 16267 26333
rect 15654 26256 15660 26308
rect 15712 26296 15718 26308
rect 16224 26296 16252 26327
rect 18046 26324 18052 26336
rect 18104 26324 18110 26376
rect 19150 26324 19156 26376
rect 19208 26364 19214 26376
rect 19392 26367 19450 26373
rect 19392 26364 19404 26367
rect 19208 26336 19404 26364
rect 19208 26324 19214 26336
rect 19392 26333 19404 26336
rect 19438 26333 19450 26367
rect 19610 26364 19616 26376
rect 19523 26336 19616 26364
rect 19392 26327 19450 26333
rect 19610 26324 19616 26336
rect 19668 26364 19674 26376
rect 19978 26364 19984 26376
rect 19668 26336 19984 26364
rect 19668 26324 19674 26336
rect 19978 26324 19984 26336
rect 20036 26324 20042 26376
rect 22097 26367 22155 26373
rect 22097 26333 22109 26367
rect 22143 26364 22155 26367
rect 22186 26364 22192 26376
rect 22143 26336 22192 26364
rect 22143 26333 22155 26336
rect 22097 26327 22155 26333
rect 22186 26324 22192 26336
rect 22244 26324 22250 26376
rect 23446 26364 23474 26404
rect 23845 26401 23857 26435
rect 23891 26432 23903 26435
rect 23934 26432 23940 26444
rect 23891 26404 23940 26432
rect 23891 26401 23903 26404
rect 23845 26395 23903 26401
rect 23934 26392 23940 26404
rect 23992 26392 23998 26444
rect 27246 26432 27252 26444
rect 27207 26404 27252 26432
rect 27246 26392 27252 26404
rect 27304 26392 27310 26444
rect 29086 26432 29092 26444
rect 27448 26404 29092 26432
rect 27448 26364 27476 26404
rect 29086 26392 29092 26404
rect 29144 26392 29150 26444
rect 30926 26432 30932 26444
rect 30887 26404 30932 26432
rect 30926 26392 30932 26404
rect 30984 26392 30990 26444
rect 33962 26432 33968 26444
rect 33923 26404 33968 26432
rect 33962 26392 33968 26404
rect 34020 26392 34026 26444
rect 36538 26432 36544 26444
rect 36499 26404 36544 26432
rect 36538 26392 36544 26404
rect 36596 26392 36602 26444
rect 37366 26392 37372 26444
rect 37424 26432 37430 26444
rect 38013 26435 38071 26441
rect 38013 26432 38025 26435
rect 37424 26404 38025 26432
rect 37424 26392 37430 26404
rect 38013 26401 38025 26404
rect 38059 26401 38071 26435
rect 39758 26432 39764 26444
rect 39719 26404 39764 26432
rect 38013 26395 38071 26401
rect 39758 26392 39764 26404
rect 39816 26392 39822 26444
rect 40218 26432 40224 26444
rect 40179 26404 40224 26432
rect 40218 26392 40224 26404
rect 40276 26392 40282 26444
rect 42766 26432 42794 26472
rect 43993 26469 44005 26503
rect 44039 26500 44051 26503
rect 44266 26500 44272 26512
rect 44039 26472 44272 26500
rect 44039 26469 44051 26472
rect 43993 26463 44051 26469
rect 44266 26460 44272 26472
rect 44324 26460 44330 26512
rect 43416 26435 43474 26441
rect 43416 26432 43428 26435
rect 42766 26404 43428 26432
rect 43416 26401 43428 26404
rect 43462 26432 43474 26435
rect 43714 26432 43720 26444
rect 43462 26404 43720 26432
rect 43462 26401 43474 26404
rect 43416 26395 43474 26401
rect 43714 26392 43720 26404
rect 43772 26392 43778 26444
rect 44358 26432 44364 26444
rect 44319 26404 44364 26432
rect 44358 26392 44364 26404
rect 44416 26392 44422 26444
rect 27614 26364 27620 26376
rect 23446 26336 27476 26364
rect 27575 26336 27620 26364
rect 27614 26324 27620 26336
rect 27672 26324 27678 26376
rect 29270 26364 29276 26376
rect 29231 26336 29276 26364
rect 29270 26324 29276 26336
rect 29328 26324 29334 26376
rect 29917 26367 29975 26373
rect 29917 26333 29929 26367
rect 29963 26364 29975 26367
rect 30006 26364 30012 26376
rect 29963 26336 30012 26364
rect 29963 26333 29975 26336
rect 29917 26327 29975 26333
rect 30006 26324 30012 26336
rect 30064 26324 30070 26376
rect 31159 26367 31217 26373
rect 31159 26333 31171 26367
rect 31205 26364 31217 26367
rect 31846 26364 31852 26376
rect 31205 26336 31852 26364
rect 31205 26333 31217 26336
rect 31159 26327 31217 26333
rect 31846 26324 31852 26336
rect 31904 26364 31910 26376
rect 32217 26367 32275 26373
rect 32217 26364 32229 26367
rect 31904 26336 32229 26364
rect 31904 26324 31910 26336
rect 32217 26333 32229 26336
rect 32263 26333 32275 26367
rect 32217 26327 32275 26333
rect 32493 26367 32551 26373
rect 32493 26333 32505 26367
rect 32539 26333 32551 26367
rect 32493 26327 32551 26333
rect 17770 26296 17776 26308
rect 15712 26268 17776 26296
rect 15712 26256 15718 26268
rect 17770 26256 17776 26268
rect 17828 26256 17834 26308
rect 19521 26299 19579 26305
rect 19521 26265 19533 26299
rect 19567 26296 19579 26299
rect 20438 26296 20444 26308
rect 19567 26268 20444 26296
rect 19567 26265 19579 26268
rect 19521 26259 19579 26265
rect 20438 26256 20444 26268
rect 20496 26256 20502 26308
rect 30024 26296 30052 26324
rect 32508 26296 32536 26327
rect 34882 26324 34888 26376
rect 34940 26364 34946 26376
rect 35069 26367 35127 26373
rect 35069 26364 35081 26367
rect 34940 26336 35081 26364
rect 34940 26324 34946 26336
rect 35069 26333 35081 26336
rect 35115 26364 35127 26367
rect 36078 26364 36084 26376
rect 35115 26336 36084 26364
rect 35115 26333 35127 26336
rect 35069 26327 35127 26333
rect 36078 26324 36084 26336
rect 36136 26324 36142 26376
rect 40494 26364 40500 26376
rect 40455 26336 40500 26364
rect 40494 26324 40500 26336
rect 40552 26324 40558 26376
rect 41782 26364 41788 26376
rect 41743 26336 41788 26364
rect 41782 26324 41788 26336
rect 41840 26324 41846 26376
rect 42058 26364 42064 26376
rect 42019 26336 42064 26364
rect 42058 26324 42064 26336
rect 42116 26364 42122 26376
rect 42426 26364 42432 26376
rect 42116 26336 42432 26364
rect 42116 26324 42122 26336
rect 42426 26324 42432 26336
rect 42484 26324 42490 26376
rect 35250 26296 35256 26308
rect 30024 26268 35256 26296
rect 35250 26256 35256 26268
rect 35308 26256 35314 26308
rect 35618 26296 35624 26308
rect 35579 26268 35624 26296
rect 35618 26256 35624 26268
rect 35676 26256 35682 26308
rect 9858 26188 9864 26240
rect 9916 26228 9922 26240
rect 10045 26231 10103 26237
rect 10045 26228 10057 26231
rect 9916 26200 10057 26228
rect 9916 26188 9922 26200
rect 10045 26197 10057 26200
rect 10091 26197 10103 26231
rect 18966 26228 18972 26240
rect 18927 26200 18972 26228
rect 10045 26191 10103 26197
rect 18966 26188 18972 26200
rect 19024 26188 19030 26240
rect 21177 26231 21235 26237
rect 21177 26197 21189 26231
rect 21223 26228 21235 26231
rect 21634 26228 21640 26240
rect 21223 26200 21640 26228
rect 21223 26197 21235 26200
rect 21177 26191 21235 26197
rect 21634 26188 21640 26200
rect 21692 26228 21698 26240
rect 22094 26228 22100 26240
rect 21692 26200 22100 26228
rect 21692 26188 21698 26200
rect 22094 26188 22100 26200
rect 22152 26188 22158 26240
rect 23014 26228 23020 26240
rect 22975 26200 23020 26228
rect 23014 26188 23020 26200
rect 23072 26188 23078 26240
rect 26510 26188 26516 26240
rect 26568 26228 26574 26240
rect 27154 26228 27160 26240
rect 26568 26200 27160 26228
rect 26568 26188 26574 26200
rect 27154 26188 27160 26200
rect 27212 26228 27218 26240
rect 27387 26231 27445 26237
rect 27387 26228 27399 26231
rect 27212 26200 27399 26228
rect 27212 26188 27218 26200
rect 27387 26197 27399 26200
rect 27433 26197 27445 26231
rect 27387 26191 27445 26197
rect 27525 26231 27583 26237
rect 27525 26197 27537 26231
rect 27571 26228 27583 26231
rect 27798 26228 27804 26240
rect 27571 26200 27804 26228
rect 27571 26197 27583 26200
rect 27525 26191 27583 26197
rect 27798 26188 27804 26200
rect 27856 26188 27862 26240
rect 33318 26228 33324 26240
rect 33279 26200 33324 26228
rect 33318 26188 33324 26200
rect 33376 26188 33382 26240
rect 34103 26231 34161 26237
rect 34103 26197 34115 26231
rect 34149 26228 34161 26231
rect 34698 26228 34704 26240
rect 34149 26200 34704 26228
rect 34149 26197 34161 26200
rect 34103 26191 34161 26197
rect 34698 26188 34704 26200
rect 34756 26188 34762 26240
rect 38930 26228 38936 26240
rect 38891 26200 38936 26228
rect 38930 26188 38936 26200
rect 38988 26188 38994 26240
rect 39206 26228 39212 26240
rect 39167 26200 39212 26228
rect 39206 26188 39212 26200
rect 39264 26188 39270 26240
rect 1104 26138 48852 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 48852 26138
rect 1104 26064 48852 26086
rect 9953 26027 10011 26033
rect 9953 25993 9965 26027
rect 9999 26024 10011 26027
rect 10226 26024 10232 26036
rect 9999 25996 10232 26024
rect 9999 25993 10011 25996
rect 9953 25987 10011 25993
rect 10226 25984 10232 25996
rect 10284 25984 10290 26036
rect 11882 26024 11888 26036
rect 11843 25996 11888 26024
rect 11882 25984 11888 25996
rect 11940 25984 11946 26036
rect 14277 26027 14335 26033
rect 14277 25993 14289 26027
rect 14323 26024 14335 26027
rect 14366 26024 14372 26036
rect 14323 25996 14372 26024
rect 14323 25993 14335 25996
rect 14277 25987 14335 25993
rect 14366 25984 14372 25996
rect 14424 26024 14430 26036
rect 17678 26024 17684 26036
rect 14424 25996 17684 26024
rect 14424 25984 14430 25996
rect 17678 25984 17684 25996
rect 17736 25984 17742 26036
rect 19610 26024 19616 26036
rect 19571 25996 19616 26024
rect 19610 25984 19616 25996
rect 19668 25984 19674 26036
rect 19981 26027 20039 26033
rect 19981 25993 19993 26027
rect 20027 26024 20039 26027
rect 20438 26024 20444 26036
rect 20027 25996 20444 26024
rect 20027 25993 20039 25996
rect 19981 25987 20039 25993
rect 20438 25984 20444 25996
rect 20496 25984 20502 26036
rect 24949 26027 25007 26033
rect 24949 25993 24961 26027
rect 24995 26024 25007 26027
rect 25130 26024 25136 26036
rect 24995 25996 25136 26024
rect 24995 25993 25007 25996
rect 24949 25987 25007 25993
rect 25130 25984 25136 25996
rect 25188 25984 25194 26036
rect 25332 25996 27108 26024
rect 11330 25916 11336 25968
rect 11388 25956 11394 25968
rect 14553 25959 14611 25965
rect 14553 25956 14565 25959
rect 11388 25928 14565 25956
rect 11388 25916 11394 25928
rect 14553 25925 14565 25928
rect 14599 25956 14611 25959
rect 14918 25956 14924 25968
rect 14599 25928 14924 25956
rect 14599 25925 14611 25928
rect 14553 25919 14611 25925
rect 14918 25916 14924 25928
rect 14976 25956 14982 25968
rect 15841 25959 15899 25965
rect 15841 25956 15853 25959
rect 14976 25928 15853 25956
rect 14976 25916 14982 25928
rect 15841 25925 15853 25928
rect 15887 25956 15899 25959
rect 16022 25956 16028 25968
rect 15887 25928 16028 25956
rect 15887 25925 15899 25928
rect 15841 25919 15899 25925
rect 16022 25916 16028 25928
rect 16080 25916 16086 25968
rect 17494 25956 17500 25968
rect 17455 25928 17500 25956
rect 17494 25916 17500 25928
rect 17552 25956 17558 25968
rect 19242 25956 19248 25968
rect 17552 25928 19248 25956
rect 17552 25916 17558 25928
rect 19242 25916 19248 25928
rect 19300 25956 19306 25968
rect 23934 25956 23940 25968
rect 19300 25928 20116 25956
rect 23847 25928 23940 25956
rect 19300 25916 19306 25928
rect 13262 25848 13268 25900
rect 13320 25888 13326 25900
rect 15286 25888 15292 25900
rect 13320 25860 13365 25888
rect 15247 25860 15292 25888
rect 13320 25848 13326 25860
rect 15286 25848 15292 25860
rect 15344 25848 15350 25900
rect 16393 25891 16451 25897
rect 16393 25857 16405 25891
rect 16439 25888 16451 25891
rect 16850 25888 16856 25900
rect 16439 25860 16856 25888
rect 16439 25857 16451 25860
rect 16393 25851 16451 25857
rect 16850 25848 16856 25860
rect 16908 25848 16914 25900
rect 17037 25891 17095 25897
rect 17037 25857 17049 25891
rect 17083 25888 17095 25891
rect 17126 25888 17132 25900
rect 17083 25860 17132 25888
rect 17083 25857 17095 25860
rect 17037 25851 17095 25857
rect 17126 25848 17132 25860
rect 17184 25848 17190 25900
rect 17770 25848 17776 25900
rect 17828 25888 17834 25900
rect 18601 25891 18659 25897
rect 18601 25888 18613 25891
rect 17828 25860 18613 25888
rect 17828 25848 17834 25860
rect 18601 25857 18613 25860
rect 18647 25888 18659 25891
rect 18874 25888 18880 25900
rect 18647 25860 18880 25888
rect 18647 25857 18659 25860
rect 18601 25851 18659 25857
rect 18874 25848 18880 25860
rect 18932 25848 18938 25900
rect 20088 25832 20116 25928
rect 23934 25916 23940 25928
rect 23992 25956 23998 25968
rect 25332 25956 25360 25996
rect 27080 25956 27108 25996
rect 28534 25984 28540 26036
rect 28592 26024 28598 26036
rect 28629 26027 28687 26033
rect 28629 26024 28641 26027
rect 28592 25996 28641 26024
rect 28592 25984 28598 25996
rect 28629 25993 28641 25996
rect 28675 25993 28687 26027
rect 28629 25987 28687 25993
rect 29270 25984 29276 26036
rect 29328 26024 29334 26036
rect 29411 26027 29469 26033
rect 29411 26024 29423 26027
rect 29328 25996 29423 26024
rect 29328 25984 29334 25996
rect 29411 25993 29423 25996
rect 29457 26024 29469 26027
rect 30101 26027 30159 26033
rect 30101 26024 30113 26027
rect 29457 25996 30113 26024
rect 29457 25993 29469 25996
rect 29411 25987 29469 25993
rect 30101 25993 30113 25996
rect 30147 25993 30159 26027
rect 36078 26024 36084 26036
rect 36039 25996 36084 26024
rect 30101 25987 30159 25993
rect 36078 25984 36084 25996
rect 36136 25984 36142 26036
rect 37366 25984 37372 26036
rect 37424 26024 37430 26036
rect 37645 26027 37703 26033
rect 37645 26024 37657 26027
rect 37424 25996 37657 26024
rect 37424 25984 37430 25996
rect 37645 25993 37657 25996
rect 37691 25993 37703 26027
rect 37645 25987 37703 25993
rect 38749 26027 38807 26033
rect 38749 25993 38761 26027
rect 38795 26024 38807 26027
rect 38930 26024 38936 26036
rect 38795 25996 38936 26024
rect 38795 25993 38807 25996
rect 38749 25987 38807 25993
rect 38930 25984 38936 25996
rect 38988 25984 38994 26036
rect 39758 25984 39764 26036
rect 39816 26024 39822 26036
rect 39853 26027 39911 26033
rect 39853 26024 39865 26027
rect 39816 25996 39865 26024
rect 39816 25984 39822 25996
rect 39853 25993 39865 25996
rect 39899 25993 39911 26027
rect 39853 25987 39911 25993
rect 40865 26027 40923 26033
rect 40865 25993 40877 26027
rect 40911 26024 40923 26027
rect 41782 26024 41788 26036
rect 40911 25996 41788 26024
rect 40911 25993 40923 25996
rect 40865 25987 40923 25993
rect 41782 25984 41788 25996
rect 41840 26024 41846 26036
rect 43027 26027 43085 26033
rect 43027 26024 43039 26027
rect 41840 25996 43039 26024
rect 41840 25984 41846 25996
rect 43027 25993 43039 25996
rect 43073 25993 43085 26027
rect 43714 26024 43720 26036
rect 43675 25996 43720 26024
rect 43027 25987 43085 25993
rect 43714 25984 43720 25996
rect 43772 25984 43778 26036
rect 44726 26024 44732 26036
rect 43824 25996 44732 26024
rect 30926 25956 30932 25968
rect 23992 25928 25360 25956
rect 25424 25928 27016 25956
rect 27080 25928 30932 25956
rect 23992 25916 23998 25928
rect 25424 25900 25452 25928
rect 22186 25888 22192 25900
rect 22147 25860 22192 25888
rect 22186 25848 22192 25860
rect 22244 25848 22250 25900
rect 25133 25891 25191 25897
rect 25133 25857 25145 25891
rect 25179 25888 25191 25891
rect 25222 25888 25228 25900
rect 25179 25860 25228 25888
rect 25179 25857 25191 25860
rect 25133 25851 25191 25857
rect 25222 25848 25228 25860
rect 25280 25848 25286 25900
rect 25406 25888 25412 25900
rect 25367 25860 25412 25888
rect 25406 25848 25412 25860
rect 25464 25848 25470 25900
rect 26510 25888 26516 25900
rect 26471 25860 26516 25888
rect 26510 25848 26516 25860
rect 26568 25848 26574 25900
rect 26697 25891 26755 25897
rect 26697 25857 26709 25891
rect 26743 25888 26755 25891
rect 26786 25888 26792 25900
rect 26743 25860 26792 25888
rect 26743 25857 26755 25860
rect 26697 25851 26755 25857
rect 26786 25848 26792 25860
rect 26844 25848 26850 25900
rect 26988 25897 27016 25928
rect 30926 25916 30932 25928
rect 30984 25916 30990 25968
rect 31202 25916 31208 25968
rect 31260 25956 31266 25968
rect 36446 25956 36452 25968
rect 31260 25928 36452 25956
rect 31260 25916 31266 25928
rect 36446 25916 36452 25928
rect 36504 25916 36510 25968
rect 36538 25916 36544 25968
rect 36596 25956 36602 25968
rect 40034 25956 40040 25968
rect 36596 25928 40040 25956
rect 36596 25916 36602 25928
rect 40034 25916 40040 25928
rect 40092 25916 40098 25968
rect 41874 25916 41880 25968
rect 41932 25956 41938 25968
rect 42337 25959 42395 25965
rect 42337 25956 42349 25959
rect 41932 25928 42349 25956
rect 41932 25916 41938 25928
rect 42337 25925 42349 25928
rect 42383 25925 42395 25959
rect 42337 25919 42395 25925
rect 43441 25959 43499 25965
rect 43441 25925 43453 25959
rect 43487 25956 43499 25959
rect 43824 25956 43852 25996
rect 44726 25984 44732 25996
rect 44784 25984 44790 26036
rect 45281 25959 45339 25965
rect 45281 25956 45293 25959
rect 43487 25928 43852 25956
rect 44008 25928 45293 25956
rect 43487 25925 43499 25928
rect 43441 25919 43499 25925
rect 26973 25891 27031 25897
rect 26973 25857 26985 25891
rect 27019 25857 27031 25891
rect 26973 25851 27031 25857
rect 28350 25848 28356 25900
rect 28408 25888 28414 25900
rect 28994 25888 29000 25900
rect 28408 25860 29000 25888
rect 28408 25848 28414 25860
rect 28994 25848 29000 25860
rect 29052 25888 29058 25900
rect 30561 25891 30619 25897
rect 30561 25888 30573 25891
rect 29052 25860 30573 25888
rect 29052 25848 29058 25860
rect 30561 25857 30573 25860
rect 30607 25888 30619 25891
rect 30650 25888 30656 25900
rect 30607 25860 30656 25888
rect 30607 25857 30619 25860
rect 30561 25851 30619 25857
rect 30650 25848 30656 25860
rect 30708 25848 30714 25900
rect 30745 25891 30803 25897
rect 30745 25857 30757 25891
rect 30791 25888 30803 25891
rect 30834 25888 30840 25900
rect 30791 25860 30840 25888
rect 30791 25857 30803 25860
rect 30745 25851 30803 25857
rect 30834 25848 30840 25860
rect 30892 25848 30898 25900
rect 32214 25848 32220 25900
rect 32272 25888 32278 25900
rect 32585 25891 32643 25897
rect 32585 25888 32597 25891
rect 32272 25860 32597 25888
rect 32272 25848 32278 25860
rect 32585 25857 32597 25860
rect 32631 25888 32643 25891
rect 33505 25891 33563 25897
rect 33505 25888 33517 25891
rect 32631 25860 33517 25888
rect 32631 25857 32643 25860
rect 32585 25851 32643 25857
rect 33505 25857 33517 25860
rect 33551 25857 33563 25891
rect 33505 25851 33563 25857
rect 34790 25848 34796 25900
rect 34848 25888 34854 25900
rect 34885 25891 34943 25897
rect 34885 25888 34897 25891
rect 34848 25860 34897 25888
rect 34848 25848 34854 25860
rect 34885 25857 34897 25860
rect 34931 25857 34943 25891
rect 34885 25851 34943 25857
rect 35342 25848 35348 25900
rect 35400 25888 35406 25900
rect 36556 25888 36584 25916
rect 36722 25888 36728 25900
rect 35400 25860 36584 25888
rect 36683 25860 36728 25888
rect 35400 25848 35406 25860
rect 36722 25848 36728 25860
rect 36780 25848 36786 25900
rect 36906 25848 36912 25900
rect 36964 25888 36970 25900
rect 37001 25891 37059 25897
rect 37001 25888 37013 25891
rect 36964 25860 37013 25888
rect 36964 25848 36970 25860
rect 37001 25857 37013 25860
rect 37047 25857 37059 25891
rect 37001 25851 37059 25857
rect 38933 25891 38991 25897
rect 38933 25857 38945 25891
rect 38979 25888 38991 25891
rect 39206 25888 39212 25900
rect 38979 25860 39212 25888
rect 38979 25857 38991 25860
rect 38933 25851 38991 25857
rect 39206 25848 39212 25860
rect 39264 25888 39270 25900
rect 41693 25891 41751 25897
rect 41693 25888 41705 25891
rect 39264 25860 41705 25888
rect 39264 25848 39270 25860
rect 41693 25857 41705 25860
rect 41739 25888 41751 25891
rect 42058 25888 42064 25900
rect 41739 25860 42064 25888
rect 41739 25857 41751 25860
rect 41693 25851 41751 25857
rect 42058 25848 42064 25860
rect 42116 25848 42122 25900
rect 10226 25820 10232 25832
rect 10187 25792 10232 25820
rect 10226 25780 10232 25792
rect 10284 25780 10290 25832
rect 10594 25820 10600 25832
rect 10555 25792 10600 25820
rect 10594 25780 10600 25792
rect 10652 25780 10658 25832
rect 20070 25820 20076 25832
rect 19983 25792 20076 25820
rect 20070 25780 20076 25792
rect 20128 25780 20134 25832
rect 20530 25820 20536 25832
rect 20491 25792 20536 25820
rect 20530 25780 20536 25792
rect 20588 25780 20594 25832
rect 21634 25820 21640 25832
rect 21595 25792 21640 25820
rect 21634 25780 21640 25792
rect 21692 25780 21698 25832
rect 22094 25820 22100 25832
rect 22055 25792 22100 25820
rect 22094 25780 22100 25792
rect 22152 25780 22158 25832
rect 28236 25823 28294 25829
rect 28236 25789 28248 25823
rect 28282 25820 28294 25823
rect 28534 25820 28540 25832
rect 28282 25792 28540 25820
rect 28282 25789 28294 25792
rect 28236 25783 28294 25789
rect 28534 25780 28540 25792
rect 28592 25780 28598 25832
rect 28810 25780 28816 25832
rect 28868 25820 28874 25832
rect 29340 25823 29398 25829
rect 29340 25820 29352 25823
rect 28868 25792 29352 25820
rect 28868 25780 28874 25792
rect 29340 25789 29352 25792
rect 29386 25820 29398 25823
rect 29825 25823 29883 25829
rect 29825 25820 29837 25823
rect 29386 25792 29837 25820
rect 29386 25789 29398 25792
rect 29340 25783 29398 25789
rect 29825 25789 29837 25792
rect 29871 25820 29883 25823
rect 31478 25820 31484 25832
rect 29871 25792 31484 25820
rect 29871 25789 29883 25792
rect 29825 25783 29883 25789
rect 31478 25780 31484 25792
rect 31536 25780 31542 25832
rect 33226 25780 33232 25832
rect 33284 25820 33290 25832
rect 35618 25820 35624 25832
rect 33284 25792 35624 25820
rect 33284 25780 33290 25792
rect 35618 25780 35624 25792
rect 35676 25780 35682 25832
rect 42956 25823 43014 25829
rect 42956 25789 42968 25823
rect 43002 25820 43014 25823
rect 43346 25820 43352 25832
rect 43002 25792 43352 25820
rect 43002 25789 43014 25792
rect 42956 25783 43014 25789
rect 43346 25780 43352 25792
rect 43404 25820 43410 25832
rect 43456 25820 43484 25919
rect 44008 25900 44036 25928
rect 45281 25925 45293 25928
rect 45327 25925 45339 25959
rect 45281 25919 45339 25925
rect 43990 25888 43996 25900
rect 43903 25860 43996 25888
rect 43990 25848 43996 25860
rect 44048 25848 44054 25900
rect 44082 25848 44088 25900
rect 44140 25888 44146 25900
rect 44269 25891 44327 25897
rect 44269 25888 44281 25891
rect 44140 25860 44281 25888
rect 44140 25848 44146 25860
rect 44269 25857 44281 25860
rect 44315 25857 44327 25891
rect 44269 25851 44327 25857
rect 43404 25792 43484 25820
rect 43404 25780 43410 25792
rect 10778 25752 10784 25764
rect 10739 25724 10784 25752
rect 10778 25712 10784 25724
rect 10836 25712 10842 25764
rect 12713 25755 12771 25761
rect 12713 25721 12725 25755
rect 12759 25752 12771 25755
rect 13357 25755 13415 25761
rect 13357 25752 13369 25755
rect 12759 25724 13369 25752
rect 12759 25721 12771 25724
rect 12713 25715 12771 25721
rect 13357 25721 13369 25724
rect 13403 25752 13415 25755
rect 13538 25752 13544 25764
rect 13403 25724 13544 25752
rect 13403 25721 13415 25724
rect 13357 25715 13415 25721
rect 13538 25712 13544 25724
rect 13596 25712 13602 25764
rect 13906 25752 13912 25764
rect 13867 25724 13912 25752
rect 13906 25712 13912 25724
rect 13964 25712 13970 25764
rect 14826 25752 14832 25764
rect 14787 25724 14832 25752
rect 14826 25712 14832 25724
rect 14884 25712 14890 25764
rect 14918 25712 14924 25764
rect 14976 25752 14982 25764
rect 14976 25724 15021 25752
rect 14976 25712 14982 25724
rect 16022 25712 16028 25764
rect 16080 25752 16086 25764
rect 16482 25752 16488 25764
rect 16080 25724 16488 25752
rect 16080 25712 16086 25724
rect 16482 25712 16488 25724
rect 16540 25712 16546 25764
rect 18693 25755 18751 25761
rect 18693 25721 18705 25755
rect 18739 25752 18751 25755
rect 18966 25752 18972 25764
rect 18739 25724 18972 25752
rect 18739 25721 18751 25724
rect 18693 25715 18751 25721
rect 18966 25712 18972 25724
rect 19024 25712 19030 25764
rect 19058 25712 19064 25764
rect 19116 25752 19122 25764
rect 19245 25755 19303 25761
rect 19245 25752 19257 25755
rect 19116 25724 19257 25752
rect 19116 25712 19122 25724
rect 19245 25721 19257 25724
rect 19291 25752 19303 25755
rect 22278 25752 22284 25764
rect 19291 25724 22284 25752
rect 19291 25721 19303 25724
rect 19245 25715 19303 25721
rect 22278 25712 22284 25724
rect 22336 25712 22342 25764
rect 24581 25755 24639 25761
rect 24581 25721 24593 25755
rect 24627 25752 24639 25755
rect 24762 25752 24768 25764
rect 24627 25724 24768 25752
rect 24627 25721 24639 25724
rect 24581 25715 24639 25721
rect 24762 25712 24768 25724
rect 24820 25752 24826 25764
rect 25225 25755 25283 25761
rect 24820 25724 25084 25752
rect 24820 25712 24826 25724
rect 9398 25644 9404 25696
rect 9456 25684 9462 25696
rect 10502 25684 10508 25696
rect 9456 25656 10508 25684
rect 9456 25644 9462 25656
rect 10502 25644 10508 25656
rect 10560 25684 10566 25696
rect 11054 25684 11060 25696
rect 10560 25656 11060 25684
rect 10560 25644 10566 25656
rect 11054 25644 11060 25656
rect 11112 25644 11118 25696
rect 11330 25644 11336 25696
rect 11388 25684 11394 25696
rect 11517 25687 11575 25693
rect 11517 25684 11529 25687
rect 11388 25656 11529 25684
rect 11388 25644 11394 25656
rect 11517 25653 11529 25656
rect 11563 25653 11575 25687
rect 11517 25647 11575 25653
rect 13081 25687 13139 25693
rect 13081 25653 13093 25687
rect 13127 25684 13139 25687
rect 13170 25684 13176 25696
rect 13127 25656 13176 25684
rect 13127 25653 13139 25656
rect 13081 25647 13139 25653
rect 13170 25644 13176 25656
rect 13228 25644 13234 25696
rect 18230 25684 18236 25696
rect 18191 25656 18236 25684
rect 18230 25644 18236 25656
rect 18288 25644 18294 25696
rect 20162 25684 20168 25696
rect 20123 25656 20168 25684
rect 20162 25644 20168 25656
rect 20220 25644 20226 25696
rect 20622 25644 20628 25696
rect 20680 25684 20686 25696
rect 21453 25687 21511 25693
rect 21453 25684 21465 25687
rect 20680 25656 21465 25684
rect 20680 25644 20686 25656
rect 21453 25653 21465 25656
rect 21499 25684 21511 25687
rect 21634 25684 21640 25696
rect 21499 25656 21640 25684
rect 21499 25653 21511 25656
rect 21453 25647 21511 25653
rect 21634 25644 21640 25656
rect 21692 25644 21698 25696
rect 22738 25684 22744 25696
rect 22699 25656 22744 25684
rect 22738 25644 22744 25656
rect 22796 25644 22802 25696
rect 25056 25684 25084 25724
rect 25225 25721 25237 25755
rect 25271 25721 25283 25755
rect 25225 25715 25283 25721
rect 26145 25755 26203 25761
rect 26145 25721 26157 25755
rect 26191 25752 26203 25755
rect 26510 25752 26516 25764
rect 26191 25724 26516 25752
rect 26191 25721 26203 25724
rect 26145 25715 26203 25721
rect 25240 25684 25268 25715
rect 26510 25712 26516 25724
rect 26568 25712 26574 25764
rect 26694 25712 26700 25764
rect 26752 25752 26758 25764
rect 26789 25755 26847 25761
rect 26789 25752 26801 25755
rect 26752 25724 26801 25752
rect 26752 25712 26758 25724
rect 26789 25721 26801 25724
rect 26835 25721 26847 25755
rect 26789 25715 26847 25721
rect 30650 25712 30656 25764
rect 30708 25752 30714 25764
rect 31066 25755 31124 25761
rect 31066 25752 31078 25755
rect 30708 25724 31078 25752
rect 30708 25712 30714 25724
rect 31066 25721 31078 25724
rect 31112 25721 31124 25755
rect 32677 25755 32735 25761
rect 32677 25752 32689 25755
rect 31066 25715 31124 25721
rect 32324 25724 32689 25752
rect 32324 25696 32352 25724
rect 32677 25721 32689 25724
rect 32723 25721 32735 25755
rect 35206 25755 35264 25761
rect 35206 25752 35218 25755
rect 32677 25715 32735 25721
rect 34624 25724 35218 25752
rect 25056 25656 25268 25684
rect 26878 25644 26884 25696
rect 26936 25684 26942 25696
rect 27614 25684 27620 25696
rect 26936 25656 27620 25684
rect 26936 25644 26942 25656
rect 27614 25644 27620 25656
rect 27672 25644 27678 25696
rect 27798 25644 27804 25696
rect 27856 25684 27862 25696
rect 27985 25687 28043 25693
rect 27985 25684 27997 25687
rect 27856 25656 27997 25684
rect 27856 25644 27862 25656
rect 27985 25653 27997 25656
rect 28031 25653 28043 25687
rect 27985 25647 28043 25653
rect 28307 25687 28365 25693
rect 28307 25653 28319 25687
rect 28353 25684 28365 25687
rect 28534 25684 28540 25696
rect 28353 25656 28540 25684
rect 28353 25653 28365 25656
rect 28307 25647 28365 25653
rect 28534 25644 28540 25656
rect 28592 25644 28598 25696
rect 28902 25644 28908 25696
rect 28960 25684 28966 25696
rect 28997 25687 29055 25693
rect 28997 25684 29009 25687
rect 28960 25656 29009 25684
rect 28960 25644 28966 25656
rect 28997 25653 29009 25656
rect 29043 25653 29055 25687
rect 31662 25684 31668 25696
rect 31623 25656 31668 25684
rect 28997 25647 29055 25653
rect 31662 25644 31668 25656
rect 31720 25684 31726 25696
rect 31941 25687 31999 25693
rect 31941 25684 31953 25687
rect 31720 25656 31953 25684
rect 31720 25644 31726 25656
rect 31941 25653 31953 25656
rect 31987 25684 31999 25687
rect 32306 25684 32312 25696
rect 31987 25656 32312 25684
rect 31987 25653 31999 25656
rect 31941 25647 31999 25653
rect 32306 25644 32312 25656
rect 32364 25644 32370 25696
rect 33410 25644 33416 25696
rect 33468 25684 33474 25696
rect 33962 25684 33968 25696
rect 33468 25656 33968 25684
rect 33468 25644 33474 25656
rect 33962 25644 33968 25656
rect 34020 25644 34026 25696
rect 34422 25644 34428 25696
rect 34480 25684 34486 25696
rect 34624 25693 34652 25724
rect 35206 25721 35218 25724
rect 35252 25721 35264 25755
rect 36817 25755 36875 25761
rect 36817 25752 36829 25755
rect 35206 25715 35264 25721
rect 35820 25724 36829 25752
rect 35820 25696 35848 25724
rect 36817 25721 36829 25724
rect 36863 25752 36875 25755
rect 36998 25752 37004 25764
rect 36863 25724 37004 25752
rect 36863 25721 36875 25724
rect 36817 25715 36875 25721
rect 36998 25712 37004 25724
rect 37056 25712 37062 25764
rect 39022 25712 39028 25764
rect 39080 25752 39086 25764
rect 39574 25752 39580 25764
rect 39080 25724 39125 25752
rect 39535 25724 39580 25752
rect 39080 25712 39086 25724
rect 39574 25712 39580 25724
rect 39632 25712 39638 25764
rect 39758 25712 39764 25764
rect 39816 25752 39822 25764
rect 40218 25752 40224 25764
rect 39816 25724 40224 25752
rect 39816 25712 39822 25724
rect 40218 25712 40224 25724
rect 40276 25712 40282 25764
rect 41414 25752 41420 25764
rect 41375 25724 41420 25752
rect 41414 25712 41420 25724
rect 41472 25712 41478 25764
rect 41509 25755 41567 25761
rect 41509 25721 41521 25755
rect 41555 25721 41567 25755
rect 41509 25715 41567 25721
rect 44085 25755 44143 25761
rect 44085 25721 44097 25755
rect 44131 25752 44143 25755
rect 44266 25752 44272 25764
rect 44131 25724 44272 25752
rect 44131 25721 44143 25724
rect 44085 25715 44143 25721
rect 34609 25687 34667 25693
rect 34609 25684 34621 25687
rect 34480 25656 34621 25684
rect 34480 25644 34486 25656
rect 34609 25653 34621 25656
rect 34655 25653 34667 25687
rect 35802 25684 35808 25696
rect 35715 25656 35808 25684
rect 34609 25647 34667 25653
rect 35802 25644 35808 25656
rect 35860 25644 35866 25696
rect 38102 25684 38108 25696
rect 38063 25656 38108 25684
rect 38102 25644 38108 25656
rect 38160 25644 38166 25696
rect 41233 25687 41291 25693
rect 41233 25653 41245 25687
rect 41279 25684 41291 25687
rect 41524 25684 41552 25715
rect 44266 25712 44272 25724
rect 44324 25712 44330 25764
rect 41690 25684 41696 25696
rect 41279 25656 41696 25684
rect 41279 25653 41291 25656
rect 41233 25647 41291 25653
rect 41690 25644 41696 25656
rect 41748 25644 41754 25696
rect 43806 25644 43812 25696
rect 43864 25684 43870 25696
rect 44358 25684 44364 25696
rect 43864 25656 44364 25684
rect 43864 25644 43870 25656
rect 44358 25644 44364 25656
rect 44416 25684 44422 25696
rect 44913 25687 44971 25693
rect 44913 25684 44925 25687
rect 44416 25656 44925 25684
rect 44416 25644 44422 25656
rect 44913 25653 44925 25656
rect 44959 25653 44971 25687
rect 44913 25647 44971 25653
rect 1104 25594 48852 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 48852 25594
rect 1104 25520 48852 25542
rect 11330 25480 11336 25492
rect 11291 25452 11336 25480
rect 11330 25440 11336 25452
rect 11388 25440 11394 25492
rect 14323 25483 14381 25489
rect 14323 25449 14335 25483
rect 14369 25480 14381 25483
rect 14737 25483 14795 25489
rect 14737 25480 14749 25483
rect 14369 25452 14749 25480
rect 14369 25449 14381 25452
rect 14323 25443 14381 25449
rect 14737 25449 14749 25452
rect 14783 25480 14795 25483
rect 14826 25480 14832 25492
rect 14783 25452 14832 25480
rect 14783 25449 14795 25452
rect 14737 25443 14795 25449
rect 14826 25440 14832 25452
rect 14884 25440 14890 25492
rect 16482 25480 16488 25492
rect 16443 25452 16488 25480
rect 16482 25440 16488 25452
rect 16540 25440 16546 25492
rect 17770 25480 17776 25492
rect 17731 25452 17776 25480
rect 17770 25440 17776 25452
rect 17828 25440 17834 25492
rect 18877 25483 18935 25489
rect 18877 25449 18889 25483
rect 18923 25480 18935 25483
rect 18966 25480 18972 25492
rect 18923 25452 18972 25480
rect 18923 25449 18935 25452
rect 18877 25443 18935 25449
rect 18966 25440 18972 25452
rect 19024 25440 19030 25492
rect 19150 25440 19156 25492
rect 19208 25480 19214 25492
rect 19245 25483 19303 25489
rect 19245 25480 19257 25483
rect 19208 25452 19257 25480
rect 19208 25440 19214 25452
rect 19245 25449 19257 25452
rect 19291 25480 19303 25483
rect 20070 25480 20076 25492
rect 19291 25452 19380 25480
rect 20031 25452 20076 25480
rect 19291 25449 19303 25452
rect 19245 25443 19303 25449
rect 10318 25372 10324 25424
rect 10376 25412 10382 25424
rect 10775 25415 10833 25421
rect 10775 25412 10787 25415
rect 10376 25384 10787 25412
rect 10376 25372 10382 25384
rect 10775 25381 10787 25384
rect 10821 25412 10833 25415
rect 11146 25412 11152 25424
rect 10821 25384 11152 25412
rect 10821 25381 10833 25384
rect 10775 25375 10833 25381
rect 11146 25372 11152 25384
rect 11204 25372 11210 25424
rect 12621 25415 12679 25421
rect 12621 25412 12633 25415
rect 12268 25384 12633 25412
rect 10226 25304 10232 25356
rect 10284 25344 10290 25356
rect 11882 25344 11888 25356
rect 10284 25316 11888 25344
rect 10284 25304 10290 25316
rect 11882 25304 11888 25316
rect 11940 25304 11946 25356
rect 10413 25279 10471 25285
rect 10413 25245 10425 25279
rect 10459 25276 10471 25279
rect 10778 25276 10784 25288
rect 10459 25248 10784 25276
rect 10459 25245 10471 25248
rect 10413 25239 10471 25245
rect 10778 25236 10784 25248
rect 10836 25236 10842 25288
rect 10042 25140 10048 25152
rect 10003 25112 10048 25140
rect 10042 25100 10048 25112
rect 10100 25100 10106 25152
rect 12066 25100 12072 25152
rect 12124 25140 12130 25152
rect 12268 25149 12296 25384
rect 12621 25381 12633 25384
rect 12667 25381 12679 25415
rect 12621 25375 12679 25381
rect 13262 25372 13268 25424
rect 13320 25412 13326 25424
rect 13541 25415 13599 25421
rect 13541 25412 13553 25415
rect 13320 25384 13553 25412
rect 13320 25372 13326 25384
rect 13541 25381 13553 25384
rect 13587 25412 13599 25415
rect 15286 25412 15292 25424
rect 13587 25384 15292 25412
rect 13587 25381 13599 25384
rect 13541 25375 13599 25381
rect 15286 25372 15292 25384
rect 15344 25372 15350 25424
rect 15470 25372 15476 25424
rect 15528 25412 15534 25424
rect 15651 25415 15709 25421
rect 15651 25412 15663 25415
rect 15528 25384 15663 25412
rect 15528 25372 15534 25384
rect 15651 25381 15663 25384
rect 15697 25412 15709 25415
rect 18319 25415 18377 25421
rect 18319 25412 18331 25415
rect 15697 25384 18331 25412
rect 15697 25381 15709 25384
rect 15651 25375 15709 25381
rect 18319 25381 18331 25384
rect 18365 25412 18377 25415
rect 18506 25412 18512 25424
rect 18365 25384 18512 25412
rect 18365 25381 18377 25384
rect 18319 25375 18377 25381
rect 18506 25372 18512 25384
rect 18564 25372 18570 25424
rect 13630 25304 13636 25356
rect 13688 25344 13694 25356
rect 14182 25344 14188 25356
rect 14240 25353 14246 25356
rect 14240 25347 14278 25353
rect 13688 25316 14188 25344
rect 13688 25304 13694 25316
rect 14182 25304 14188 25316
rect 14266 25313 14278 25347
rect 14240 25307 14278 25313
rect 17957 25347 18015 25353
rect 17957 25313 17969 25347
rect 18003 25344 18015 25347
rect 18046 25344 18052 25356
rect 18003 25316 18052 25344
rect 18003 25313 18015 25316
rect 17957 25307 18015 25313
rect 14240 25304 14246 25307
rect 18046 25304 18052 25316
rect 18104 25304 18110 25356
rect 19352 25344 19380 25452
rect 20070 25440 20076 25452
rect 20128 25440 20134 25492
rect 22186 25480 22192 25492
rect 22147 25452 22192 25480
rect 22186 25440 22192 25452
rect 22244 25440 22250 25492
rect 24765 25483 24823 25489
rect 24765 25449 24777 25483
rect 24811 25480 24823 25483
rect 24946 25480 24952 25492
rect 24811 25452 24952 25480
rect 24811 25449 24823 25452
rect 24765 25443 24823 25449
rect 24946 25440 24952 25452
rect 25004 25440 25010 25492
rect 25222 25440 25228 25492
rect 25280 25480 25286 25492
rect 25869 25483 25927 25489
rect 25869 25480 25881 25483
rect 25280 25452 25881 25480
rect 25280 25440 25286 25452
rect 25869 25449 25881 25452
rect 25915 25449 25927 25483
rect 26786 25480 26792 25492
rect 26747 25452 26792 25480
rect 25869 25443 25927 25449
rect 26786 25440 26792 25452
rect 26844 25440 26850 25492
rect 28350 25480 28356 25492
rect 28311 25452 28356 25480
rect 28350 25440 28356 25452
rect 28408 25440 28414 25492
rect 31846 25480 31852 25492
rect 31807 25452 31852 25480
rect 31846 25440 31852 25452
rect 31904 25440 31910 25492
rect 34514 25440 34520 25492
rect 34572 25480 34578 25492
rect 34885 25483 34943 25489
rect 34885 25480 34897 25483
rect 34572 25452 34897 25480
rect 34572 25440 34578 25452
rect 34885 25449 34897 25452
rect 34931 25480 34943 25483
rect 34931 25452 35204 25480
rect 34931 25449 34943 25452
rect 34885 25443 34943 25449
rect 19426 25372 19432 25424
rect 19484 25412 19490 25424
rect 19613 25415 19671 25421
rect 19613 25412 19625 25415
rect 19484 25384 19625 25412
rect 19484 25372 19490 25384
rect 19613 25381 19625 25384
rect 19659 25381 19671 25415
rect 19613 25375 19671 25381
rect 19628 25344 19656 25375
rect 23014 25372 23020 25424
rect 23072 25412 23078 25424
rect 23385 25415 23443 25421
rect 23385 25412 23397 25415
rect 23072 25384 23397 25412
rect 23072 25372 23078 25384
rect 23385 25381 23397 25384
rect 23431 25381 23443 25415
rect 25038 25412 25044 25424
rect 24999 25384 25044 25412
rect 23385 25375 23443 25381
rect 25038 25372 25044 25384
rect 25096 25372 25102 25424
rect 25130 25372 25136 25424
rect 25188 25412 25194 25424
rect 25682 25412 25688 25424
rect 25188 25384 25688 25412
rect 25188 25372 25194 25384
rect 25682 25372 25688 25384
rect 25740 25372 25746 25424
rect 29914 25412 29920 25424
rect 29875 25384 29920 25412
rect 29914 25372 29920 25384
rect 29972 25372 29978 25424
rect 32306 25412 32312 25424
rect 32267 25384 32312 25412
rect 32306 25372 32312 25384
rect 32364 25372 32370 25424
rect 34698 25372 34704 25424
rect 34756 25412 34762 25424
rect 35176 25421 35204 25452
rect 36722 25440 36728 25492
rect 36780 25480 36786 25492
rect 37369 25483 37427 25489
rect 37369 25480 37381 25483
rect 36780 25452 37381 25480
rect 36780 25440 36786 25452
rect 37369 25449 37381 25452
rect 37415 25449 37427 25483
rect 37369 25443 37427 25449
rect 40635 25483 40693 25489
rect 40635 25449 40647 25483
rect 40681 25480 40693 25483
rect 41414 25480 41420 25492
rect 40681 25452 41420 25480
rect 40681 25449 40693 25452
rect 40635 25443 40693 25449
rect 41414 25440 41420 25452
rect 41472 25440 41478 25492
rect 35069 25415 35127 25421
rect 35069 25412 35081 25415
rect 34756 25384 35081 25412
rect 34756 25372 34762 25384
rect 35069 25381 35081 25384
rect 35115 25381 35127 25415
rect 35069 25375 35127 25381
rect 35161 25415 35219 25421
rect 35161 25381 35173 25415
rect 35207 25412 35219 25415
rect 35802 25412 35808 25424
rect 35207 25384 35808 25412
rect 35207 25381 35219 25384
rect 35161 25375 35219 25381
rect 35802 25372 35808 25384
rect 35860 25372 35866 25424
rect 36998 25412 37004 25424
rect 36959 25384 37004 25412
rect 36998 25372 37004 25384
rect 37056 25372 37062 25424
rect 38930 25412 38936 25424
rect 38891 25384 38936 25412
rect 38930 25372 38936 25384
rect 38988 25372 38994 25424
rect 41690 25412 41696 25424
rect 41651 25384 41696 25412
rect 41690 25372 41696 25384
rect 41748 25372 41754 25424
rect 43622 25372 43628 25424
rect 43680 25412 43686 25424
rect 43993 25415 44051 25421
rect 43993 25412 44005 25415
rect 43680 25384 44005 25412
rect 43680 25372 43686 25384
rect 43993 25381 44005 25384
rect 44039 25381 44051 25415
rect 43993 25375 44051 25381
rect 20346 25344 20352 25356
rect 19352 25316 19564 25344
rect 19628 25316 20352 25344
rect 12529 25279 12587 25285
rect 12529 25245 12541 25279
rect 12575 25276 12587 25279
rect 12802 25276 12808 25288
rect 12575 25248 12808 25276
rect 12575 25245 12587 25248
rect 12529 25239 12587 25245
rect 12802 25236 12808 25248
rect 12860 25236 12866 25288
rect 13173 25279 13231 25285
rect 13173 25245 13185 25279
rect 13219 25276 13231 25279
rect 13219 25248 13814 25276
rect 13219 25245 13231 25248
rect 13173 25239 13231 25245
rect 13786 25208 13814 25248
rect 15102 25236 15108 25288
rect 15160 25276 15166 25288
rect 15289 25279 15347 25285
rect 15289 25276 15301 25279
rect 15160 25248 15301 25276
rect 15160 25236 15166 25248
rect 15289 25245 15301 25248
rect 15335 25245 15347 25279
rect 19536 25276 19564 25316
rect 20346 25304 20352 25316
rect 20404 25304 20410 25356
rect 26418 25304 26424 25356
rect 26476 25344 26482 25356
rect 27062 25353 27068 25356
rect 27008 25347 27068 25353
rect 27008 25344 27020 25347
rect 26476 25316 27020 25344
rect 26476 25304 26482 25316
rect 27008 25313 27020 25316
rect 27054 25313 27068 25347
rect 27008 25307 27068 25313
rect 27062 25304 27068 25307
rect 27120 25304 27126 25356
rect 33594 25304 33600 25356
rect 33652 25344 33658 25356
rect 34000 25347 34058 25353
rect 34000 25344 34012 25347
rect 33652 25316 34012 25344
rect 33652 25304 33658 25316
rect 34000 25313 34012 25316
rect 34046 25313 34058 25347
rect 34000 25307 34058 25313
rect 36446 25304 36452 25356
rect 36504 25344 36510 25356
rect 36576 25347 36634 25353
rect 36576 25344 36588 25347
rect 36504 25316 36588 25344
rect 36504 25304 36510 25316
rect 36576 25313 36588 25316
rect 36622 25313 36634 25347
rect 36576 25307 36634 25313
rect 37642 25304 37648 25356
rect 37700 25344 37706 25356
rect 37772 25347 37830 25353
rect 37772 25344 37784 25347
rect 37700 25316 37784 25344
rect 37700 25304 37706 25316
rect 37772 25313 37784 25316
rect 37818 25313 37830 25347
rect 37772 25307 37830 25313
rect 40310 25304 40316 25356
rect 40368 25344 40374 25356
rect 40532 25347 40590 25353
rect 40532 25344 40544 25347
rect 40368 25316 40544 25344
rect 40368 25304 40374 25316
rect 40532 25313 40544 25316
rect 40578 25313 40590 25347
rect 40532 25307 40590 25313
rect 20070 25276 20076 25288
rect 19536 25248 20076 25276
rect 15289 25239 15347 25245
rect 20070 25236 20076 25248
rect 20128 25236 20134 25288
rect 23290 25276 23296 25288
rect 23251 25248 23296 25276
rect 23290 25236 23296 25248
rect 23348 25236 23354 25288
rect 24949 25279 25007 25285
rect 24949 25245 24961 25279
rect 24995 25276 25007 25279
rect 25130 25276 25136 25288
rect 24995 25248 25136 25276
rect 24995 25245 25007 25248
rect 24949 25239 25007 25245
rect 25130 25236 25136 25248
rect 25188 25236 25194 25288
rect 25225 25279 25283 25285
rect 25225 25245 25237 25279
rect 25271 25276 25283 25279
rect 25406 25276 25412 25288
rect 25271 25248 25412 25276
rect 25271 25245 25283 25248
rect 25225 25239 25283 25245
rect 13906 25208 13912 25220
rect 13786 25180 13912 25208
rect 13906 25168 13912 25180
rect 13964 25208 13970 25220
rect 16298 25208 16304 25220
rect 13964 25180 16304 25208
rect 13964 25168 13970 25180
rect 16298 25168 16304 25180
rect 16356 25168 16362 25220
rect 23845 25211 23903 25217
rect 23845 25177 23857 25211
rect 23891 25208 23903 25211
rect 25240 25208 25268 25239
rect 25406 25236 25412 25248
rect 25464 25236 25470 25288
rect 27985 25279 28043 25285
rect 27985 25245 27997 25279
rect 28031 25276 28043 25279
rect 28166 25276 28172 25288
rect 28031 25248 28172 25276
rect 28031 25245 28043 25248
rect 27985 25239 28043 25245
rect 28166 25236 28172 25248
rect 28224 25236 28230 25288
rect 28534 25236 28540 25288
rect 28592 25276 28598 25288
rect 29825 25279 29883 25285
rect 29825 25276 29837 25279
rect 28592 25248 29837 25276
rect 28592 25236 28598 25248
rect 29825 25245 29837 25248
rect 29871 25276 29883 25279
rect 30098 25276 30104 25288
rect 29871 25248 30104 25276
rect 29871 25245 29883 25248
rect 29825 25239 29883 25245
rect 30098 25236 30104 25248
rect 30156 25236 30162 25288
rect 32217 25279 32275 25285
rect 32217 25245 32229 25279
rect 32263 25276 32275 25279
rect 32582 25276 32588 25288
rect 32263 25248 32588 25276
rect 32263 25245 32275 25248
rect 32217 25239 32275 25245
rect 32582 25236 32588 25248
rect 32640 25236 32646 25288
rect 35345 25279 35403 25285
rect 35345 25276 35357 25279
rect 32784 25248 35357 25276
rect 23891 25180 25268 25208
rect 27111 25211 27169 25217
rect 23891 25177 23903 25180
rect 23845 25171 23903 25177
rect 27111 25177 27123 25211
rect 27157 25208 27169 25211
rect 29273 25211 29331 25217
rect 29273 25208 29285 25211
rect 27157 25180 29285 25208
rect 27157 25177 27169 25180
rect 27111 25171 27169 25177
rect 29273 25177 29285 25180
rect 29319 25208 29331 25211
rect 29362 25208 29368 25220
rect 29319 25180 29368 25208
rect 29319 25177 29331 25180
rect 29273 25171 29331 25177
rect 29362 25168 29368 25180
rect 29420 25168 29426 25220
rect 30374 25208 30380 25220
rect 30335 25180 30380 25208
rect 30374 25168 30380 25180
rect 30432 25208 30438 25220
rect 32784 25217 32812 25248
rect 35345 25245 35357 25248
rect 35391 25276 35403 25279
rect 35802 25276 35808 25288
rect 35391 25248 35808 25276
rect 35391 25245 35403 25248
rect 35345 25239 35403 25245
rect 35802 25236 35808 25248
rect 35860 25236 35866 25288
rect 38838 25276 38844 25288
rect 38799 25248 38844 25276
rect 38838 25236 38844 25248
rect 38896 25236 38902 25288
rect 39022 25236 39028 25288
rect 39080 25276 39086 25288
rect 39117 25279 39175 25285
rect 39117 25276 39129 25279
rect 39080 25248 39129 25276
rect 39080 25236 39086 25248
rect 39117 25245 39129 25248
rect 39163 25276 39175 25279
rect 39574 25276 39580 25288
rect 39163 25248 39580 25276
rect 39163 25245 39175 25248
rect 39117 25239 39175 25245
rect 39574 25236 39580 25248
rect 39632 25236 39638 25288
rect 41598 25276 41604 25288
rect 41559 25248 41604 25276
rect 41598 25236 41604 25248
rect 41656 25236 41662 25288
rect 41877 25279 41935 25285
rect 41877 25245 41889 25279
rect 41923 25276 41935 25279
rect 43714 25276 43720 25288
rect 41923 25248 43720 25276
rect 41923 25245 41935 25248
rect 41877 25239 41935 25245
rect 32769 25211 32827 25217
rect 32769 25208 32781 25211
rect 30432 25180 32781 25208
rect 30432 25168 30438 25180
rect 32769 25177 32781 25180
rect 32815 25177 32827 25211
rect 35434 25208 35440 25220
rect 32769 25171 32827 25177
rect 33106 25180 35440 25208
rect 12253 25143 12311 25149
rect 12253 25140 12265 25143
rect 12124 25112 12265 25140
rect 12124 25100 12130 25112
rect 12253 25109 12265 25112
rect 12299 25109 12311 25143
rect 12253 25103 12311 25109
rect 15105 25143 15163 25149
rect 15105 25109 15117 25143
rect 15151 25140 15163 25143
rect 15194 25140 15200 25152
rect 15151 25112 15200 25140
rect 15151 25109 15163 25112
rect 15105 25103 15163 25109
rect 15194 25100 15200 25112
rect 15252 25100 15258 25152
rect 16206 25140 16212 25152
rect 16167 25112 16212 25140
rect 16206 25100 16212 25112
rect 16264 25100 16270 25152
rect 16850 25140 16856 25152
rect 16811 25112 16856 25140
rect 16850 25100 16856 25112
rect 16908 25100 16914 25152
rect 19334 25100 19340 25152
rect 19392 25140 19398 25152
rect 20441 25143 20499 25149
rect 20441 25140 20453 25143
rect 19392 25112 20453 25140
rect 19392 25100 19398 25112
rect 20441 25109 20453 25112
rect 20487 25140 20499 25143
rect 20530 25140 20536 25152
rect 20487 25112 20536 25140
rect 20487 25109 20499 25112
rect 20441 25103 20499 25109
rect 20530 25100 20536 25112
rect 20588 25100 20594 25152
rect 21729 25143 21787 25149
rect 21729 25109 21741 25143
rect 21775 25140 21787 25143
rect 22094 25140 22100 25152
rect 21775 25112 22100 25140
rect 21775 25109 21787 25112
rect 21729 25103 21787 25109
rect 22094 25100 22100 25112
rect 22152 25140 22158 25152
rect 22646 25140 22652 25152
rect 22152 25112 22652 25140
rect 22152 25100 22158 25112
rect 22646 25100 22652 25112
rect 22704 25100 22710 25152
rect 23934 25100 23940 25152
rect 23992 25140 23998 25152
rect 24213 25143 24271 25149
rect 24213 25140 24225 25143
rect 23992 25112 24225 25140
rect 23992 25100 23998 25112
rect 24213 25109 24225 25112
rect 24259 25109 24271 25143
rect 24213 25103 24271 25109
rect 26510 25100 26516 25152
rect 26568 25140 26574 25152
rect 27246 25140 27252 25152
rect 26568 25112 27252 25140
rect 26568 25100 26574 25112
rect 27246 25100 27252 25112
rect 27304 25140 27310 25152
rect 27433 25143 27491 25149
rect 27433 25140 27445 25143
rect 27304 25112 27445 25140
rect 27304 25100 27310 25112
rect 27433 25109 27445 25112
rect 27479 25109 27491 25143
rect 28902 25140 28908 25152
rect 28863 25112 28908 25140
rect 27433 25103 27491 25109
rect 28902 25100 28908 25112
rect 28960 25100 28966 25152
rect 30926 25100 30932 25152
rect 30984 25140 30990 25152
rect 31113 25143 31171 25149
rect 31113 25140 31125 25143
rect 30984 25112 31125 25140
rect 30984 25100 30990 25112
rect 31113 25109 31125 25112
rect 31159 25140 31171 25143
rect 33106 25140 33134 25180
rect 35434 25168 35440 25180
rect 35492 25168 35498 25220
rect 35986 25168 35992 25220
rect 36044 25208 36050 25220
rect 37875 25211 37933 25217
rect 37875 25208 37887 25211
rect 36044 25180 37887 25208
rect 36044 25168 36050 25180
rect 37875 25177 37887 25180
rect 37921 25177 37933 25211
rect 37875 25171 37933 25177
rect 39206 25168 39212 25220
rect 39264 25208 39270 25220
rect 41892 25208 41920 25239
rect 43714 25236 43720 25248
rect 43772 25236 43778 25288
rect 43901 25279 43959 25285
rect 43901 25245 43913 25279
rect 43947 25276 43959 25279
rect 44634 25276 44640 25288
rect 43947 25248 44640 25276
rect 43947 25245 43959 25248
rect 43901 25239 43959 25245
rect 44634 25236 44640 25248
rect 44692 25276 44698 25288
rect 45373 25279 45431 25285
rect 45373 25276 45385 25279
rect 44692 25248 45385 25276
rect 44692 25236 44698 25248
rect 45373 25245 45385 25248
rect 45419 25245 45431 25279
rect 45373 25239 45431 25245
rect 39264 25180 41920 25208
rect 39264 25168 39270 25180
rect 44082 25168 44088 25220
rect 44140 25208 44146 25220
rect 44453 25211 44511 25217
rect 44453 25208 44465 25211
rect 44140 25180 44465 25208
rect 44140 25168 44146 25180
rect 44453 25177 44465 25180
rect 44499 25177 44511 25211
rect 44453 25171 44511 25177
rect 31159 25112 33134 25140
rect 34103 25143 34161 25149
rect 31159 25109 31171 25112
rect 31113 25103 31171 25109
rect 34103 25109 34115 25143
rect 34149 25140 34161 25143
rect 34425 25143 34483 25149
rect 34425 25140 34437 25143
rect 34149 25112 34437 25140
rect 34149 25109 34161 25112
rect 34103 25103 34161 25109
rect 34425 25109 34437 25112
rect 34471 25140 34483 25143
rect 34698 25140 34704 25152
rect 34471 25112 34704 25140
rect 34471 25109 34483 25112
rect 34425 25103 34483 25109
rect 34698 25100 34704 25112
rect 34756 25100 34762 25152
rect 36538 25100 36544 25152
rect 36596 25140 36602 25152
rect 36679 25143 36737 25149
rect 36679 25140 36691 25143
rect 36596 25112 36691 25140
rect 36596 25100 36602 25112
rect 36679 25109 36691 25112
rect 36725 25109 36737 25143
rect 38194 25140 38200 25152
rect 38155 25112 38200 25140
rect 36679 25103 36737 25109
rect 38194 25100 38200 25112
rect 38252 25100 38258 25152
rect 1104 25050 48852 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 48852 25050
rect 1104 24976 48852 24998
rect 10318 24936 10324 24948
rect 10279 24908 10324 24936
rect 10318 24896 10324 24908
rect 10376 24896 10382 24948
rect 11517 24939 11575 24945
rect 11517 24905 11529 24939
rect 11563 24936 11575 24939
rect 12802 24936 12808 24948
rect 11563 24908 12808 24936
rect 11563 24905 11575 24908
rect 11517 24899 11575 24905
rect 12802 24896 12808 24908
rect 12860 24896 12866 24948
rect 13538 24936 13544 24948
rect 13499 24908 13544 24936
rect 13538 24896 13544 24908
rect 13596 24896 13602 24948
rect 14550 24896 14556 24948
rect 14608 24936 14614 24948
rect 15470 24936 15476 24948
rect 14608 24908 15476 24936
rect 14608 24896 14614 24908
rect 15470 24896 15476 24908
rect 15528 24896 15534 24948
rect 17129 24939 17187 24945
rect 17129 24905 17141 24939
rect 17175 24936 17187 24939
rect 18046 24936 18052 24948
rect 17175 24908 18052 24936
rect 17175 24905 17187 24908
rect 17129 24899 17187 24905
rect 18046 24896 18052 24908
rect 18104 24896 18110 24948
rect 23014 24936 23020 24948
rect 22975 24908 23020 24936
rect 23014 24896 23020 24908
rect 23072 24896 23078 24948
rect 24857 24939 24915 24945
rect 24857 24905 24869 24939
rect 24903 24936 24915 24939
rect 25038 24936 25044 24948
rect 24903 24908 25044 24936
rect 24903 24905 24915 24908
rect 24857 24899 24915 24905
rect 25038 24896 25044 24908
rect 25096 24936 25102 24948
rect 25133 24939 25191 24945
rect 25133 24936 25145 24939
rect 25096 24908 25145 24936
rect 25096 24896 25102 24908
rect 25133 24905 25145 24908
rect 25179 24905 25191 24939
rect 26602 24936 26608 24948
rect 26563 24908 26608 24936
rect 25133 24899 25191 24905
rect 26602 24896 26608 24908
rect 26660 24896 26666 24948
rect 27062 24936 27068 24948
rect 27023 24908 27068 24936
rect 27062 24896 27068 24908
rect 27120 24896 27126 24948
rect 34514 24896 34520 24948
rect 34572 24936 34578 24948
rect 34609 24939 34667 24945
rect 34609 24936 34621 24939
rect 34572 24908 34621 24936
rect 34572 24896 34578 24908
rect 34609 24905 34621 24908
rect 34655 24905 34667 24939
rect 34609 24899 34667 24905
rect 34790 24896 34796 24948
rect 34848 24936 34854 24948
rect 35897 24939 35955 24945
rect 35897 24936 35909 24939
rect 34848 24908 35909 24936
rect 34848 24896 34854 24908
rect 35897 24905 35909 24908
rect 35943 24905 35955 24939
rect 35897 24899 35955 24905
rect 36357 24939 36415 24945
rect 36357 24905 36369 24939
rect 36403 24936 36415 24939
rect 36446 24936 36452 24948
rect 36403 24908 36452 24936
rect 36403 24905 36415 24908
rect 36357 24899 36415 24905
rect 36446 24896 36452 24908
rect 36504 24896 36510 24948
rect 36998 24896 37004 24948
rect 37056 24936 37062 24948
rect 37277 24939 37335 24945
rect 37277 24936 37289 24939
rect 37056 24908 37289 24936
rect 37056 24896 37062 24908
rect 37277 24905 37289 24908
rect 37323 24936 37335 24939
rect 37642 24936 37648 24948
rect 37323 24908 37648 24936
rect 37323 24905 37335 24908
rect 37277 24899 37335 24905
rect 37642 24896 37648 24908
rect 37700 24896 37706 24948
rect 38930 24936 38936 24948
rect 38891 24908 38936 24936
rect 38930 24896 38936 24908
rect 38988 24896 38994 24948
rect 39482 24896 39488 24948
rect 39540 24936 39546 24948
rect 40310 24936 40316 24948
rect 39540 24908 40316 24936
rect 39540 24896 39546 24908
rect 40310 24896 40316 24908
rect 40368 24936 40374 24948
rect 40681 24939 40739 24945
rect 40681 24936 40693 24939
rect 40368 24908 40693 24936
rect 40368 24896 40374 24908
rect 40681 24905 40693 24908
rect 40727 24905 40739 24939
rect 41690 24936 41696 24948
rect 41651 24908 41696 24936
rect 40681 24899 40739 24905
rect 41690 24896 41696 24908
rect 41748 24896 41754 24948
rect 43622 24936 43628 24948
rect 43583 24908 43628 24936
rect 43622 24896 43628 24908
rect 43680 24896 43686 24948
rect 43855 24939 43913 24945
rect 43855 24905 43867 24939
rect 43901 24936 43913 24939
rect 43990 24936 43996 24948
rect 43901 24908 43996 24936
rect 43901 24905 43913 24908
rect 43855 24899 43913 24905
rect 43990 24896 43996 24908
rect 44048 24896 44054 24948
rect 44085 24939 44143 24945
rect 44085 24905 44097 24939
rect 44131 24936 44143 24939
rect 44269 24939 44327 24945
rect 44269 24936 44281 24939
rect 44131 24908 44281 24936
rect 44131 24905 44143 24908
rect 44085 24899 44143 24905
rect 44269 24905 44281 24908
rect 44315 24936 44327 24939
rect 44450 24936 44456 24948
rect 44315 24908 44456 24936
rect 44315 24905 44327 24908
rect 44269 24899 44327 24905
rect 44450 24896 44456 24908
rect 44508 24896 44514 24948
rect 44634 24936 44640 24948
rect 44595 24908 44640 24936
rect 44634 24896 44640 24908
rect 44692 24896 44698 24948
rect 11238 24828 11244 24880
rect 11296 24868 11302 24880
rect 12161 24871 12219 24877
rect 12161 24868 12173 24871
rect 11296 24840 12173 24868
rect 11296 24828 11302 24840
rect 12161 24837 12173 24840
rect 12207 24868 12219 24871
rect 12529 24871 12587 24877
rect 12529 24868 12541 24871
rect 12207 24840 12541 24868
rect 12207 24837 12219 24840
rect 12161 24831 12219 24837
rect 12529 24837 12541 24840
rect 12575 24837 12587 24871
rect 18230 24868 18236 24880
rect 12529 24831 12587 24837
rect 14844 24840 18236 24868
rect 9953 24803 10011 24809
rect 9953 24769 9965 24803
rect 9999 24800 10011 24803
rect 10042 24800 10048 24812
rect 9999 24772 10048 24800
rect 9999 24769 10011 24772
rect 9953 24763 10011 24769
rect 10042 24760 10048 24772
rect 10100 24800 10106 24812
rect 10594 24800 10600 24812
rect 10100 24772 10600 24800
rect 10100 24760 10106 24772
rect 10594 24760 10600 24772
rect 10652 24800 10658 24812
rect 10652 24772 13492 24800
rect 10652 24760 10658 24772
rect 10410 24732 10416 24744
rect 10371 24704 10416 24732
rect 10410 24692 10416 24704
rect 10468 24692 10474 24744
rect 10980 24741 11008 24772
rect 10965 24735 11023 24741
rect 10965 24701 10977 24735
rect 11011 24701 11023 24735
rect 10965 24695 11023 24701
rect 11885 24735 11943 24741
rect 11885 24701 11897 24735
rect 11931 24732 11943 24735
rect 12618 24732 12624 24744
rect 11931 24704 12624 24732
rect 11931 24701 11943 24704
rect 11885 24695 11943 24701
rect 12618 24692 12624 24704
rect 12676 24692 12682 24744
rect 13464 24676 13492 24772
rect 14366 24732 14372 24744
rect 14327 24704 14372 24732
rect 14366 24692 14372 24704
rect 14424 24692 14430 24744
rect 14844 24741 14872 24840
rect 18230 24828 18236 24840
rect 18288 24828 18294 24880
rect 27890 24868 27896 24880
rect 22296 24840 27896 24868
rect 16025 24803 16083 24809
rect 16025 24769 16037 24803
rect 16071 24800 16083 24803
rect 16114 24800 16120 24812
rect 16071 24772 16120 24800
rect 16071 24769 16083 24772
rect 16025 24763 16083 24769
rect 16114 24760 16120 24772
rect 16172 24800 16178 24812
rect 17126 24800 17132 24812
rect 16172 24772 17132 24800
rect 16172 24760 16178 24772
rect 17126 24760 17132 24772
rect 17184 24760 17190 24812
rect 17773 24803 17831 24809
rect 17773 24769 17785 24803
rect 17819 24800 17831 24803
rect 18506 24800 18512 24812
rect 17819 24772 18512 24800
rect 17819 24769 17831 24772
rect 17773 24763 17831 24769
rect 18506 24760 18512 24772
rect 18564 24800 18570 24812
rect 20162 24800 20168 24812
rect 18564 24772 19288 24800
rect 20123 24772 20168 24800
rect 18564 24760 18570 24772
rect 14829 24735 14887 24741
rect 14829 24701 14841 24735
rect 14875 24701 14887 24735
rect 14829 24695 14887 24701
rect 17497 24735 17555 24741
rect 17497 24701 17509 24735
rect 17543 24732 17555 24735
rect 17862 24732 17868 24744
rect 17543 24704 17868 24732
rect 17543 24701 17555 24704
rect 17497 24695 17555 24701
rect 11146 24664 11152 24676
rect 11107 24636 11152 24664
rect 11146 24624 11152 24636
rect 11204 24624 11210 24676
rect 12529 24667 12587 24673
rect 12529 24633 12541 24667
rect 12575 24664 12587 24667
rect 12943 24667 13001 24673
rect 12943 24664 12955 24667
rect 12575 24636 12955 24664
rect 12575 24633 12587 24636
rect 12529 24627 12587 24633
rect 12943 24633 12955 24636
rect 12989 24633 13001 24667
rect 12943 24627 13001 24633
rect 13446 24624 13452 24676
rect 13504 24664 13510 24676
rect 13817 24667 13875 24673
rect 13817 24664 13829 24667
rect 13504 24636 13829 24664
rect 13504 24624 13510 24636
rect 13817 24633 13829 24636
rect 13863 24664 13875 24667
rect 14844 24664 14872 24695
rect 17862 24692 17868 24704
rect 17920 24732 17926 24744
rect 18046 24732 18052 24744
rect 17920 24704 18052 24732
rect 17920 24692 17926 24704
rect 18046 24692 18052 24704
rect 18104 24692 18110 24744
rect 18601 24735 18659 24741
rect 18601 24701 18613 24735
rect 18647 24732 18659 24735
rect 19260 24732 19288 24772
rect 20162 24760 20168 24772
rect 20220 24760 20226 24812
rect 18647 24704 19196 24732
rect 19260 24704 20116 24732
rect 18647 24701 18659 24704
rect 18601 24695 18659 24701
rect 15102 24664 15108 24676
rect 13863 24636 14872 24664
rect 15063 24636 15108 24664
rect 13863 24633 13875 24636
rect 13817 24627 13875 24633
rect 15102 24624 15108 24636
rect 15160 24624 15166 24676
rect 16117 24667 16175 24673
rect 16117 24633 16129 24667
rect 16163 24664 16175 24667
rect 16206 24664 16212 24676
rect 16163 24636 16212 24664
rect 16163 24633 16175 24636
rect 16117 24627 16175 24633
rect 14182 24596 14188 24608
rect 14143 24568 14188 24596
rect 14182 24556 14188 24568
rect 14240 24556 14246 24608
rect 15841 24599 15899 24605
rect 15841 24565 15853 24599
rect 15887 24596 15899 24599
rect 16132 24596 16160 24627
rect 16206 24624 16212 24636
rect 16264 24624 16270 24676
rect 16298 24624 16304 24676
rect 16356 24664 16362 24676
rect 16669 24667 16727 24673
rect 16669 24664 16681 24667
rect 16356 24636 16681 24664
rect 16356 24624 16362 24636
rect 16669 24633 16681 24636
rect 16715 24664 16727 24667
rect 19058 24664 19064 24676
rect 16715 24636 19064 24664
rect 16715 24633 16727 24636
rect 16669 24627 16727 24633
rect 19058 24624 19064 24636
rect 19116 24624 19122 24676
rect 18138 24596 18144 24608
rect 15887 24568 16160 24596
rect 18099 24568 18144 24596
rect 15887 24565 15899 24568
rect 15841 24559 15899 24565
rect 18138 24556 18144 24568
rect 18196 24556 18202 24608
rect 19168 24605 19196 24704
rect 19153 24599 19211 24605
rect 19153 24565 19165 24599
rect 19199 24596 19211 24599
rect 19334 24596 19340 24608
rect 19199 24568 19340 24596
rect 19199 24565 19211 24568
rect 19153 24559 19211 24565
rect 19334 24556 19340 24568
rect 19392 24556 19398 24608
rect 20088 24605 20116 24704
rect 21266 24692 21272 24744
rect 21324 24732 21330 24744
rect 22296 24741 22324 24840
rect 27890 24828 27896 24840
rect 27948 24828 27954 24880
rect 33137 24871 33195 24877
rect 33137 24837 33149 24871
rect 33183 24868 33195 24871
rect 35342 24868 35348 24880
rect 33183 24840 35348 24868
rect 33183 24837 33195 24840
rect 33137 24831 33195 24837
rect 22741 24803 22799 24809
rect 22741 24769 22753 24803
rect 22787 24800 22799 24803
rect 23934 24800 23940 24812
rect 22787 24772 23940 24800
rect 22787 24769 22799 24772
rect 22741 24763 22799 24769
rect 23934 24760 23940 24772
rect 23992 24760 23998 24812
rect 29362 24800 29368 24812
rect 29323 24772 29368 24800
rect 29362 24760 29368 24772
rect 29420 24760 29426 24812
rect 29822 24760 29828 24812
rect 29880 24800 29886 24812
rect 30009 24803 30067 24809
rect 30009 24800 30021 24803
rect 29880 24772 30021 24800
rect 29880 24760 29886 24772
rect 30009 24769 30021 24772
rect 30055 24800 30067 24803
rect 30055 24772 32444 24800
rect 30055 24769 30067 24772
rect 30009 24763 30067 24769
rect 21913 24735 21971 24741
rect 21913 24732 21925 24735
rect 21324 24704 21925 24732
rect 21324 24692 21330 24704
rect 21913 24701 21925 24704
rect 21959 24732 21971 24735
rect 22281 24735 22339 24741
rect 22281 24732 22293 24735
rect 21959 24704 22293 24732
rect 21959 24701 21971 24704
rect 21913 24695 21971 24701
rect 22281 24701 22293 24704
rect 22327 24701 22339 24735
rect 22281 24695 22339 24701
rect 22557 24735 22615 24741
rect 22557 24701 22569 24735
rect 22603 24732 22615 24735
rect 22646 24732 22652 24744
rect 22603 24704 22652 24732
rect 22603 24701 22615 24704
rect 22557 24695 22615 24701
rect 22646 24692 22652 24704
rect 22704 24692 22710 24744
rect 25682 24732 25688 24744
rect 25643 24704 25688 24732
rect 25682 24692 25688 24704
rect 25740 24692 25746 24744
rect 27430 24732 27436 24744
rect 27391 24704 27436 24732
rect 27430 24692 27436 24704
rect 27488 24692 27494 24744
rect 27982 24732 27988 24744
rect 27943 24704 27988 24732
rect 27982 24692 27988 24704
rect 28040 24692 28046 24744
rect 32416 24676 32444 24772
rect 33279 24741 33307 24840
rect 35342 24828 35348 24840
rect 35400 24828 35406 24880
rect 38838 24828 38844 24880
rect 38896 24868 38902 24880
rect 39301 24871 39359 24877
rect 39301 24868 39313 24871
rect 38896 24840 39313 24868
rect 38896 24828 38902 24840
rect 39301 24837 39313 24840
rect 39347 24868 39359 24871
rect 42521 24871 42579 24877
rect 42521 24868 42533 24871
rect 39347 24840 42533 24868
rect 39347 24837 39359 24840
rect 39301 24831 39359 24837
rect 42521 24837 42533 24840
rect 42567 24868 42579 24871
rect 44818 24868 44824 24880
rect 42567 24840 44824 24868
rect 42567 24837 42579 24840
rect 42521 24831 42579 24837
rect 44818 24828 44824 24840
rect 44876 24828 44882 24880
rect 34698 24760 34704 24812
rect 34756 24800 34762 24812
rect 34977 24803 35035 24809
rect 34977 24800 34989 24803
rect 34756 24772 34989 24800
rect 34756 24760 34762 24772
rect 34977 24769 34989 24772
rect 35023 24769 35035 24803
rect 35250 24800 35256 24812
rect 35211 24772 35256 24800
rect 34977 24763 35035 24769
rect 35250 24760 35256 24772
rect 35308 24760 35314 24812
rect 37734 24800 37740 24812
rect 37647 24772 37740 24800
rect 37734 24760 37740 24772
rect 37792 24800 37798 24812
rect 38194 24800 38200 24812
rect 37792 24772 38200 24800
rect 37792 24760 37798 24772
rect 38194 24760 38200 24772
rect 38252 24760 38258 24812
rect 42889 24803 42947 24809
rect 42889 24800 42901 24803
rect 41800 24772 42901 24800
rect 33264 24735 33322 24741
rect 33264 24701 33276 24735
rect 33310 24701 33322 24735
rect 33264 24695 33322 24701
rect 36354 24692 36360 24744
rect 36412 24732 36418 24744
rect 36484 24735 36542 24741
rect 36484 24732 36496 24735
rect 36412 24704 36496 24732
rect 36412 24692 36418 24704
rect 36484 24701 36496 24704
rect 36530 24701 36542 24735
rect 36484 24695 36542 24701
rect 39850 24692 39856 24744
rect 39908 24732 39914 24744
rect 40862 24732 40868 24744
rect 40920 24741 40926 24744
rect 40920 24735 40958 24741
rect 39908 24704 40868 24732
rect 39908 24692 39914 24704
rect 40862 24692 40868 24704
rect 40946 24732 40958 24735
rect 41325 24735 41383 24741
rect 41325 24732 41337 24735
rect 40946 24704 41337 24732
rect 40946 24701 40958 24704
rect 40920 24695 40958 24701
rect 41325 24701 41337 24704
rect 41371 24701 41383 24735
rect 41325 24695 41383 24701
rect 40920 24692 40926 24695
rect 20527 24667 20585 24673
rect 20527 24633 20539 24667
rect 20573 24664 20585 24667
rect 22738 24664 22744 24676
rect 20573 24636 22744 24664
rect 20573 24633 20585 24636
rect 20527 24627 20585 24633
rect 20073 24599 20131 24605
rect 20073 24565 20085 24599
rect 20119 24596 20131 24599
rect 20542 24596 20570 24627
rect 22738 24624 22744 24636
rect 22796 24664 22802 24676
rect 23385 24667 23443 24673
rect 23385 24664 23397 24667
rect 22796 24636 23397 24664
rect 22796 24624 22802 24636
rect 23385 24633 23397 24636
rect 23431 24664 23443 24667
rect 24210 24664 24216 24676
rect 23431 24636 24216 24664
rect 23431 24633 23443 24636
rect 23385 24627 23443 24633
rect 24210 24624 24216 24636
rect 24268 24673 24274 24676
rect 24268 24667 24316 24673
rect 24268 24633 24270 24667
rect 24304 24664 24316 24667
rect 25501 24667 25559 24673
rect 25501 24664 25513 24667
rect 24304 24636 25513 24664
rect 24304 24633 24316 24636
rect 24268 24627 24316 24633
rect 25501 24633 25513 24636
rect 25547 24664 25559 24667
rect 26006 24667 26064 24673
rect 26006 24664 26018 24667
rect 25547 24636 26018 24664
rect 25547 24633 25559 24636
rect 25501 24627 25559 24633
rect 26006 24633 26018 24636
rect 26052 24633 26064 24667
rect 28166 24664 28172 24676
rect 28127 24636 28172 24664
rect 26006 24627 26064 24633
rect 24268 24624 24274 24627
rect 20714 24596 20720 24608
rect 20119 24568 20720 24596
rect 20119 24565 20131 24568
rect 20073 24559 20131 24565
rect 20714 24556 20720 24568
rect 20772 24556 20778 24608
rect 20990 24556 20996 24608
rect 21048 24596 21054 24608
rect 21085 24599 21143 24605
rect 21085 24596 21097 24599
rect 21048 24568 21097 24596
rect 21048 24556 21054 24568
rect 21085 24565 21097 24568
rect 21131 24565 21143 24599
rect 26021 24596 26049 24627
rect 28166 24624 28172 24636
rect 28224 24624 28230 24676
rect 28902 24624 28908 24676
rect 28960 24664 28966 24676
rect 29089 24667 29147 24673
rect 29089 24664 29101 24667
rect 28960 24636 29101 24664
rect 28960 24624 28966 24636
rect 29089 24633 29101 24636
rect 29135 24664 29147 24667
rect 29457 24667 29515 24673
rect 29457 24664 29469 24667
rect 29135 24636 29469 24664
rect 29135 24633 29147 24636
rect 29089 24627 29147 24633
rect 29457 24633 29469 24636
rect 29503 24633 29515 24667
rect 31754 24664 31760 24676
rect 31715 24636 31760 24664
rect 29457 24627 29515 24633
rect 28258 24596 28264 24608
rect 26021 24568 28264 24596
rect 21085 24559 21143 24565
rect 28258 24556 28264 24568
rect 28316 24596 28322 24608
rect 28445 24599 28503 24605
rect 28445 24596 28457 24599
rect 28316 24568 28457 24596
rect 28316 24556 28322 24568
rect 28445 24565 28457 24568
rect 28491 24565 28503 24599
rect 29472 24596 29500 24627
rect 31754 24624 31760 24636
rect 31812 24624 31818 24676
rect 31849 24667 31907 24673
rect 31849 24633 31861 24667
rect 31895 24633 31907 24667
rect 32398 24664 32404 24676
rect 32359 24636 32404 24664
rect 31849 24627 31907 24633
rect 29914 24596 29920 24608
rect 29472 24568 29920 24596
rect 28445 24559 28503 24565
rect 29914 24556 29920 24568
rect 29972 24596 29978 24608
rect 30285 24599 30343 24605
rect 30285 24596 30297 24599
rect 29972 24568 30297 24596
rect 29972 24556 29978 24568
rect 30285 24565 30297 24568
rect 30331 24565 30343 24599
rect 30285 24559 30343 24565
rect 31573 24599 31631 24605
rect 31573 24565 31585 24599
rect 31619 24596 31631 24599
rect 31662 24596 31668 24608
rect 31619 24568 31668 24596
rect 31619 24565 31631 24568
rect 31573 24559 31631 24565
rect 31662 24556 31668 24568
rect 31720 24596 31726 24608
rect 31864 24596 31892 24627
rect 32398 24624 32404 24636
rect 32456 24624 32462 24676
rect 32582 24624 32588 24676
rect 32640 24664 32646 24676
rect 33367 24667 33425 24673
rect 33367 24664 33379 24667
rect 32640 24636 33379 24664
rect 32640 24624 32646 24636
rect 33367 24633 33379 24636
rect 33413 24633 33425 24667
rect 33367 24627 33425 24633
rect 34514 24624 34520 24676
rect 34572 24664 34578 24676
rect 35066 24664 35072 24676
rect 34572 24636 35072 24664
rect 34572 24624 34578 24636
rect 35066 24624 35072 24636
rect 35124 24624 35130 24676
rect 37645 24667 37703 24673
rect 37645 24633 37657 24667
rect 37691 24664 37703 24667
rect 38010 24664 38016 24676
rect 37691 24636 38016 24664
rect 37691 24633 37703 24636
rect 37645 24627 37703 24633
rect 38010 24624 38016 24636
rect 38068 24624 38074 24676
rect 41003 24667 41061 24673
rect 41003 24633 41015 24667
rect 41049 24664 41061 24667
rect 41800 24664 41828 24772
rect 42889 24769 42901 24772
rect 42935 24769 42947 24803
rect 42889 24763 42947 24769
rect 43784 24735 43842 24741
rect 43784 24701 43796 24735
rect 43830 24732 43842 24735
rect 44085 24735 44143 24741
rect 44085 24732 44097 24735
rect 43830 24704 44097 24732
rect 43830 24701 43842 24704
rect 43784 24695 43842 24701
rect 44085 24701 44097 24704
rect 44131 24732 44143 24735
rect 44266 24732 44272 24744
rect 44131 24704 44272 24732
rect 44131 24701 44143 24704
rect 44085 24695 44143 24701
rect 44266 24692 44272 24704
rect 44324 24692 44330 24744
rect 41969 24667 42027 24673
rect 41969 24664 41981 24667
rect 41049 24636 41981 24664
rect 41049 24633 41061 24636
rect 41003 24627 41061 24633
rect 41969 24633 41981 24636
rect 42015 24633 42027 24667
rect 41969 24627 42027 24633
rect 42061 24667 42119 24673
rect 42061 24633 42073 24667
rect 42107 24633 42119 24667
rect 42061 24627 42119 24633
rect 32677 24599 32735 24605
rect 32677 24596 32689 24599
rect 31720 24568 32689 24596
rect 31720 24556 31726 24568
rect 32677 24565 32689 24568
rect 32723 24565 32735 24599
rect 32677 24559 32735 24565
rect 33594 24556 33600 24608
rect 33652 24596 33658 24608
rect 33965 24599 34023 24605
rect 33965 24596 33977 24599
rect 33652 24568 33977 24596
rect 33652 24556 33658 24568
rect 33965 24565 33977 24568
rect 34011 24565 34023 24599
rect 33965 24559 34023 24565
rect 36354 24556 36360 24608
rect 36412 24596 36418 24608
rect 36587 24599 36645 24605
rect 36587 24596 36599 24599
rect 36412 24568 36599 24596
rect 36412 24556 36418 24568
rect 36587 24565 36599 24568
rect 36633 24565 36645 24599
rect 38654 24596 38660 24608
rect 38615 24568 38660 24596
rect 36587 24559 36645 24565
rect 38654 24556 38660 24568
rect 38712 24556 38718 24608
rect 41690 24556 41696 24608
rect 41748 24596 41754 24608
rect 42076 24596 42104 24627
rect 41748 24568 42104 24596
rect 41748 24556 41754 24568
rect 1104 24506 48852 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 48852 24506
rect 1104 24432 48852 24454
rect 10410 24392 10416 24404
rect 10371 24364 10416 24392
rect 10410 24352 10416 24364
rect 10468 24352 10474 24404
rect 10778 24392 10784 24404
rect 10739 24364 10784 24392
rect 10778 24352 10784 24364
rect 10836 24352 10842 24404
rect 12066 24392 12072 24404
rect 12027 24364 12072 24392
rect 12066 24352 12072 24364
rect 12124 24352 12130 24404
rect 12618 24352 12624 24404
rect 12676 24392 12682 24404
rect 12989 24395 13047 24401
rect 12989 24392 13001 24395
rect 12676 24364 13001 24392
rect 12676 24352 12682 24364
rect 12989 24361 13001 24364
rect 13035 24361 13047 24395
rect 12989 24355 13047 24361
rect 13354 24352 13360 24404
rect 13412 24392 13418 24404
rect 14366 24392 14372 24404
rect 13412 24364 13814 24392
rect 14327 24364 14372 24392
rect 13412 24352 13418 24364
rect 11238 24284 11244 24336
rect 11296 24324 11302 24336
rect 11470 24327 11528 24333
rect 11470 24324 11482 24327
rect 11296 24296 11482 24324
rect 11296 24284 11302 24296
rect 11470 24293 11482 24296
rect 11516 24293 11528 24327
rect 11470 24287 11528 24293
rect 12434 24216 12440 24268
rect 12492 24256 12498 24268
rect 12897 24259 12955 24265
rect 12897 24256 12909 24259
rect 12492 24228 12909 24256
rect 12492 24216 12498 24228
rect 12897 24225 12909 24228
rect 12943 24256 12955 24259
rect 13262 24256 13268 24268
rect 12943 24228 13268 24256
rect 12943 24225 12955 24228
rect 12897 24219 12955 24225
rect 13262 24216 13268 24228
rect 13320 24216 13326 24268
rect 13446 24256 13452 24268
rect 13407 24228 13452 24256
rect 13446 24216 13452 24228
rect 13504 24216 13510 24268
rect 13786 24256 13814 24364
rect 14366 24352 14372 24364
rect 14424 24352 14430 24404
rect 15102 24352 15108 24404
rect 15160 24392 15166 24404
rect 15473 24395 15531 24401
rect 15473 24392 15485 24395
rect 15160 24364 15485 24392
rect 15160 24352 15166 24364
rect 15473 24361 15485 24364
rect 15519 24361 15531 24395
rect 15473 24355 15531 24361
rect 15795 24395 15853 24401
rect 15795 24361 15807 24395
rect 15841 24392 15853 24395
rect 16850 24392 16856 24404
rect 15841 24364 16856 24392
rect 15841 24361 15853 24364
rect 15795 24355 15853 24361
rect 16850 24352 16856 24364
rect 16908 24352 16914 24404
rect 20162 24392 20168 24404
rect 20123 24364 20168 24392
rect 20162 24352 20168 24364
rect 20220 24352 20226 24404
rect 21174 24392 21180 24404
rect 21135 24364 21180 24392
rect 21174 24352 21180 24364
rect 21232 24352 21238 24404
rect 23290 24392 23296 24404
rect 23251 24364 23296 24392
rect 23290 24352 23296 24364
rect 23348 24352 23354 24404
rect 24210 24392 24216 24404
rect 24171 24364 24216 24392
rect 24210 24352 24216 24364
rect 24268 24352 24274 24404
rect 24762 24392 24768 24404
rect 24723 24364 24768 24392
rect 24762 24352 24768 24364
rect 24820 24352 24826 24404
rect 25130 24392 25136 24404
rect 25091 24364 25136 24392
rect 25130 24352 25136 24364
rect 25188 24352 25194 24404
rect 27893 24395 27951 24401
rect 27893 24361 27905 24395
rect 27939 24392 27951 24395
rect 27982 24392 27988 24404
rect 27939 24364 27988 24392
rect 27939 24361 27951 24364
rect 27893 24355 27951 24361
rect 27982 24352 27988 24364
rect 28040 24352 28046 24404
rect 28166 24392 28172 24404
rect 28127 24364 28172 24392
rect 28166 24352 28172 24364
rect 28224 24352 28230 24404
rect 28810 24392 28816 24404
rect 28771 24364 28816 24392
rect 28810 24352 28816 24364
rect 28868 24352 28874 24404
rect 30098 24392 30104 24404
rect 30059 24364 30104 24392
rect 30098 24352 30104 24364
rect 30156 24352 30162 24404
rect 31754 24392 31760 24404
rect 31715 24364 31760 24392
rect 31754 24352 31760 24364
rect 31812 24392 31818 24404
rect 32263 24395 32321 24401
rect 32263 24392 32275 24395
rect 31812 24364 32275 24392
rect 31812 24352 31818 24364
rect 32263 24361 32275 24364
rect 32309 24361 32321 24395
rect 32582 24392 32588 24404
rect 32543 24364 32588 24392
rect 32263 24355 32321 24361
rect 32582 24352 32588 24364
rect 32640 24352 32646 24404
rect 35066 24392 35072 24404
rect 35027 24364 35072 24392
rect 35066 24352 35072 24364
rect 35124 24352 35130 24404
rect 36446 24392 36452 24404
rect 36407 24364 36452 24392
rect 36446 24352 36452 24364
rect 36504 24392 36510 24404
rect 37366 24392 37372 24404
rect 36504 24364 37372 24392
rect 36504 24352 36510 24364
rect 37366 24352 37372 24364
rect 37424 24352 37430 24404
rect 38841 24395 38899 24401
rect 38841 24361 38853 24395
rect 38887 24392 38899 24395
rect 38930 24392 38936 24404
rect 38887 24364 38936 24392
rect 38887 24361 38899 24364
rect 38841 24355 38899 24361
rect 38930 24352 38936 24364
rect 38988 24352 38994 24404
rect 41417 24395 41475 24401
rect 41417 24361 41429 24395
rect 41463 24361 41475 24395
rect 41417 24355 41475 24361
rect 16114 24324 16120 24336
rect 16075 24296 16120 24324
rect 16114 24284 16120 24296
rect 16172 24284 16178 24336
rect 18319 24327 18377 24333
rect 18319 24293 18331 24327
rect 18365 24324 18377 24327
rect 18506 24324 18512 24336
rect 18365 24296 18512 24324
rect 18365 24293 18377 24296
rect 18319 24287 18377 24293
rect 18506 24284 18512 24296
rect 18564 24284 18570 24336
rect 20530 24284 20536 24336
rect 20588 24324 20594 24336
rect 22097 24327 22155 24333
rect 20588 24296 21404 24324
rect 20588 24284 20594 24296
rect 15724 24259 15782 24265
rect 15724 24256 15736 24259
rect 13786 24228 15736 24256
rect 15724 24225 15736 24228
rect 15770 24256 15782 24259
rect 16022 24256 16028 24268
rect 15770 24228 16028 24256
rect 15770 24225 15782 24228
rect 15724 24219 15782 24225
rect 16022 24216 16028 24228
rect 16080 24216 16086 24268
rect 16720 24259 16778 24265
rect 16720 24225 16732 24259
rect 16766 24256 16778 24259
rect 17402 24256 17408 24268
rect 16766 24228 17408 24256
rect 16766 24225 16778 24228
rect 16720 24219 16778 24225
rect 17402 24216 17408 24228
rect 17460 24216 17466 24268
rect 17957 24259 18015 24265
rect 17957 24225 17969 24259
rect 18003 24256 18015 24259
rect 18138 24256 18144 24268
rect 18003 24228 18144 24256
rect 18003 24225 18015 24228
rect 17957 24219 18015 24225
rect 18138 24216 18144 24228
rect 18196 24216 18202 24268
rect 19772 24259 19830 24265
rect 19772 24225 19784 24259
rect 19818 24256 19830 24259
rect 19886 24256 19892 24268
rect 19818 24228 19892 24256
rect 19818 24225 19830 24228
rect 19772 24219 19830 24225
rect 19886 24216 19892 24228
rect 19944 24216 19950 24268
rect 21177 24259 21235 24265
rect 21177 24225 21189 24259
rect 21223 24256 21235 24259
rect 21266 24256 21272 24268
rect 21223 24228 21272 24256
rect 21223 24225 21235 24228
rect 21177 24219 21235 24225
rect 21266 24216 21272 24228
rect 21324 24216 21330 24268
rect 21376 24265 21404 24296
rect 22097 24293 22109 24327
rect 22143 24324 22155 24327
rect 22646 24324 22652 24336
rect 22143 24296 22652 24324
rect 22143 24293 22155 24296
rect 22097 24287 22155 24293
rect 22646 24284 22652 24296
rect 22704 24324 22710 24336
rect 28000 24324 28028 24352
rect 30466 24324 30472 24336
rect 22704 24296 23474 24324
rect 28000 24296 29224 24324
rect 30427 24296 30472 24324
rect 22704 24284 22710 24296
rect 21361 24259 21419 24265
rect 21361 24225 21373 24259
rect 21407 24256 21419 24259
rect 22186 24256 22192 24268
rect 21407 24228 22192 24256
rect 21407 24225 21419 24228
rect 21361 24219 21419 24225
rect 22186 24216 22192 24228
rect 22244 24216 22250 24268
rect 22278 24216 22284 24268
rect 22336 24256 22342 24268
rect 22532 24259 22590 24265
rect 22532 24256 22544 24259
rect 22336 24228 22544 24256
rect 22336 24216 22342 24228
rect 22532 24225 22544 24228
rect 22578 24256 22590 24259
rect 22922 24256 22928 24268
rect 22578 24228 22928 24256
rect 22578 24225 22590 24228
rect 22532 24219 22590 24225
rect 22922 24216 22928 24228
rect 22980 24216 22986 24268
rect 11146 24188 11152 24200
rect 11107 24160 11152 24188
rect 11146 24148 11152 24160
rect 11204 24148 11210 24200
rect 15194 24148 15200 24200
rect 15252 24188 15258 24200
rect 16807 24191 16865 24197
rect 16807 24188 16819 24191
rect 15252 24160 16819 24188
rect 15252 24148 15258 24160
rect 16807 24157 16819 24160
rect 16853 24157 16865 24191
rect 16807 24151 16865 24157
rect 14366 24080 14372 24132
rect 14424 24120 14430 24132
rect 18414 24120 18420 24132
rect 14424 24092 18420 24120
rect 14424 24080 14430 24092
rect 18414 24080 18420 24092
rect 18472 24080 18478 24132
rect 18782 24080 18788 24132
rect 18840 24120 18846 24132
rect 19843 24123 19901 24129
rect 19843 24120 19855 24123
rect 18840 24092 19855 24120
rect 18840 24080 18846 24092
rect 19843 24089 19855 24092
rect 19889 24089 19901 24123
rect 22603 24123 22661 24129
rect 22603 24120 22615 24123
rect 19843 24083 19901 24089
rect 21652 24092 22615 24120
rect 21652 24064 21680 24092
rect 22603 24089 22615 24092
rect 22649 24089 22661 24123
rect 22603 24083 22661 24089
rect 12342 24012 12348 24064
rect 12400 24052 12406 24064
rect 12437 24055 12495 24061
rect 12437 24052 12449 24055
rect 12400 24024 12449 24052
rect 12400 24012 12406 24024
rect 12437 24021 12449 24024
rect 12483 24021 12495 24055
rect 18874 24052 18880 24064
rect 18835 24024 18880 24052
rect 12437 24015 12495 24021
rect 18874 24012 18880 24024
rect 18932 24012 18938 24064
rect 19150 24052 19156 24064
rect 19111 24024 19156 24052
rect 19150 24012 19156 24024
rect 19208 24012 19214 24064
rect 21634 24012 21640 24064
rect 21692 24012 21698 24064
rect 23446 24052 23474 24296
rect 25406 24216 25412 24268
rect 25464 24256 25470 24268
rect 26418 24256 26424 24268
rect 25464 24228 26424 24256
rect 25464 24216 25470 24228
rect 26418 24216 26424 24228
rect 26476 24256 26482 24268
rect 26548 24259 26606 24265
rect 26548 24256 26560 24259
rect 26476 24228 26560 24256
rect 26476 24216 26482 24228
rect 26548 24225 26560 24228
rect 26594 24225 26606 24259
rect 28718 24256 28724 24268
rect 28679 24228 28724 24256
rect 26548 24219 26606 24225
rect 28718 24216 28724 24228
rect 28776 24216 28782 24268
rect 29196 24265 29224 24296
rect 30466 24284 30472 24296
rect 30524 24284 30530 24336
rect 35342 24324 35348 24336
rect 35303 24296 35348 24324
rect 35342 24284 35348 24296
rect 35400 24284 35406 24336
rect 35618 24284 35624 24336
rect 35676 24324 35682 24336
rect 35897 24327 35955 24333
rect 35897 24324 35909 24327
rect 35676 24296 35909 24324
rect 35676 24284 35682 24296
rect 35897 24293 35909 24296
rect 35943 24293 35955 24327
rect 35897 24287 35955 24293
rect 38102 24284 38108 24336
rect 38160 24324 38166 24336
rect 38242 24327 38300 24333
rect 38242 24324 38254 24327
rect 38160 24296 38254 24324
rect 38160 24284 38166 24296
rect 38242 24293 38254 24296
rect 38288 24324 38300 24327
rect 40818 24327 40876 24333
rect 40818 24324 40830 24327
rect 38288 24296 40830 24324
rect 38288 24293 38300 24296
rect 38242 24287 38300 24293
rect 40818 24293 40830 24296
rect 40864 24324 40876 24327
rect 41230 24324 41236 24336
rect 40864 24296 41236 24324
rect 40864 24293 40876 24296
rect 40818 24287 40876 24293
rect 41230 24284 41236 24296
rect 41288 24284 41294 24336
rect 41432 24324 41460 24355
rect 41598 24352 41604 24404
rect 41656 24392 41662 24404
rect 42061 24395 42119 24401
rect 42061 24392 42073 24395
rect 41656 24364 42073 24392
rect 41656 24352 41662 24364
rect 42061 24361 42073 24364
rect 42107 24392 42119 24395
rect 42383 24395 42441 24401
rect 42383 24392 42395 24395
rect 42107 24364 42395 24392
rect 42107 24361 42119 24364
rect 42061 24355 42119 24361
rect 42383 24361 42395 24364
rect 42429 24361 42441 24395
rect 42383 24355 42441 24361
rect 41690 24324 41696 24336
rect 41432 24296 41696 24324
rect 41690 24284 41696 24296
rect 41748 24324 41754 24336
rect 43254 24324 43260 24336
rect 41748 24296 43260 24324
rect 41748 24284 41754 24296
rect 43254 24284 43260 24296
rect 43312 24324 43318 24336
rect 43533 24327 43591 24333
rect 43533 24324 43545 24327
rect 43312 24296 43545 24324
rect 43312 24284 43318 24296
rect 43533 24293 43545 24296
rect 43579 24293 43591 24327
rect 43533 24287 43591 24293
rect 29181 24259 29239 24265
rect 29181 24225 29193 24259
rect 29227 24256 29239 24259
rect 29454 24256 29460 24268
rect 29227 24228 29460 24256
rect 29227 24225 29239 24228
rect 29181 24219 29239 24225
rect 29454 24216 29460 24228
rect 29512 24216 29518 24268
rect 31754 24216 31760 24268
rect 31812 24256 31818 24268
rect 32160 24259 32218 24265
rect 32160 24256 32172 24259
rect 31812 24228 32172 24256
rect 31812 24216 31818 24228
rect 32160 24225 32172 24228
rect 32206 24225 32218 24259
rect 33778 24256 33784 24268
rect 32160 24219 32218 24225
rect 33106 24228 33784 24256
rect 23842 24188 23848 24200
rect 23803 24160 23848 24188
rect 23842 24148 23848 24160
rect 23900 24148 23906 24200
rect 27430 24188 27436 24200
rect 27391 24160 27436 24188
rect 27430 24148 27436 24160
rect 27488 24148 27494 24200
rect 30374 24188 30380 24200
rect 30335 24160 30380 24188
rect 30374 24148 30380 24160
rect 30432 24148 30438 24200
rect 31018 24188 31024 24200
rect 30979 24160 31024 24188
rect 31018 24148 31024 24160
rect 31076 24148 31082 24200
rect 32674 24148 32680 24200
rect 32732 24188 32738 24200
rect 33106 24188 33134 24228
rect 33778 24216 33784 24228
rect 33836 24216 33842 24268
rect 34054 24256 34060 24268
rect 34015 24228 34060 24256
rect 34054 24216 34060 24228
rect 34112 24216 34118 24268
rect 40494 24256 40500 24268
rect 40455 24228 40500 24256
rect 40494 24216 40500 24228
rect 40552 24216 40558 24268
rect 42312 24259 42370 24265
rect 42312 24225 42324 24259
rect 42358 24256 42370 24259
rect 42794 24256 42800 24268
rect 42358 24228 42800 24256
rect 42358 24225 42370 24228
rect 42312 24219 42370 24225
rect 42794 24216 42800 24228
rect 42852 24216 42858 24268
rect 34330 24188 34336 24200
rect 32732 24160 33134 24188
rect 34291 24160 34336 24188
rect 32732 24148 32738 24160
rect 34330 24148 34336 24160
rect 34388 24148 34394 24200
rect 34701 24191 34759 24197
rect 34701 24157 34713 24191
rect 34747 24188 34759 24191
rect 35253 24191 35311 24197
rect 35253 24188 35265 24191
rect 34747 24160 35265 24188
rect 34747 24157 34759 24160
rect 34701 24151 34759 24157
rect 35253 24157 35265 24160
rect 35299 24188 35311 24191
rect 36354 24188 36360 24200
rect 35299 24160 36360 24188
rect 35299 24157 35311 24160
rect 35253 24151 35311 24157
rect 36354 24148 36360 24160
rect 36412 24148 36418 24200
rect 37918 24188 37924 24200
rect 37879 24160 37924 24188
rect 37918 24148 37924 24160
rect 37976 24148 37982 24200
rect 43438 24188 43444 24200
rect 43399 24160 43444 24188
rect 43438 24148 43444 24160
rect 43496 24148 43502 24200
rect 44082 24188 44088 24200
rect 44043 24160 44088 24188
rect 44082 24148 44088 24160
rect 44140 24148 44146 24200
rect 23753 24055 23811 24061
rect 23753 24052 23765 24055
rect 23446 24024 23765 24052
rect 23753 24021 23765 24024
rect 23799 24052 23811 24055
rect 24026 24052 24032 24064
rect 23799 24024 24032 24052
rect 23799 24021 23811 24024
rect 23753 24015 23811 24021
rect 24026 24012 24032 24024
rect 24084 24012 24090 24064
rect 25682 24052 25688 24064
rect 25643 24024 25688 24052
rect 25682 24012 25688 24024
rect 25740 24012 25746 24064
rect 26651 24055 26709 24061
rect 26651 24021 26663 24055
rect 26697 24052 26709 24055
rect 27338 24052 27344 24064
rect 26697 24024 27344 24052
rect 26697 24021 26709 24024
rect 26651 24015 26709 24021
rect 27338 24012 27344 24024
rect 27396 24012 27402 24064
rect 29730 24052 29736 24064
rect 29691 24024 29736 24052
rect 29730 24012 29736 24024
rect 29788 24012 29794 24064
rect 1104 23962 48852 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 48852 23962
rect 1104 23888 48852 23910
rect 11146 23808 11152 23860
rect 11204 23848 11210 23860
rect 11517 23851 11575 23857
rect 11517 23848 11529 23851
rect 11204 23820 11529 23848
rect 11204 23808 11210 23820
rect 11517 23817 11529 23820
rect 11563 23817 11575 23851
rect 12250 23848 12256 23860
rect 12211 23820 12256 23848
rect 11517 23811 11575 23817
rect 12250 23808 12256 23820
rect 12308 23808 12314 23860
rect 13262 23808 13268 23860
rect 13320 23848 13326 23860
rect 13449 23851 13507 23857
rect 13449 23848 13461 23851
rect 13320 23820 13461 23848
rect 13320 23808 13326 23820
rect 13449 23817 13461 23820
rect 13495 23848 13507 23851
rect 17402 23848 17408 23860
rect 13495 23820 17126 23848
rect 17363 23820 17408 23848
rect 13495 23817 13507 23820
rect 13449 23811 13507 23817
rect 11238 23780 11244 23792
rect 11199 23752 11244 23780
rect 11238 23740 11244 23752
rect 11296 23740 11302 23792
rect 14921 23783 14979 23789
rect 14921 23749 14933 23783
rect 14967 23780 14979 23783
rect 15562 23780 15568 23792
rect 14967 23752 15568 23780
rect 14967 23749 14979 23752
rect 14921 23743 14979 23749
rect 15562 23740 15568 23752
rect 15620 23740 15626 23792
rect 12342 23672 12348 23724
rect 12400 23712 12406 23724
rect 12986 23712 12992 23724
rect 12400 23684 12801 23712
rect 12947 23684 12992 23712
rect 12400 23672 12406 23684
rect 10410 23604 10416 23656
rect 10468 23644 10474 23656
rect 12250 23644 12256 23656
rect 10468 23616 12256 23644
rect 10468 23604 10474 23616
rect 12250 23604 12256 23616
rect 12308 23644 12314 23656
rect 12437 23647 12495 23653
rect 12437 23644 12449 23647
rect 12308 23616 12449 23644
rect 12308 23604 12314 23616
rect 12437 23613 12449 23616
rect 12483 23613 12495 23647
rect 12773 23644 12801 23684
rect 12986 23672 12992 23684
rect 13044 23672 13050 23724
rect 14366 23712 14372 23724
rect 13786 23684 14372 23712
rect 12897 23647 12955 23653
rect 12897 23644 12909 23647
rect 12773 23616 12909 23644
rect 12437 23607 12495 23613
rect 12897 23613 12909 23616
rect 12943 23613 12955 23647
rect 12897 23607 12955 23613
rect 9950 23536 9956 23588
rect 10008 23576 10014 23588
rect 13786 23576 13814 23684
rect 14366 23672 14372 23684
rect 14424 23712 14430 23724
rect 17098 23712 17126 23820
rect 17402 23808 17408 23820
rect 17460 23808 17466 23860
rect 17865 23851 17923 23857
rect 17865 23817 17877 23851
rect 17911 23848 17923 23851
rect 18138 23848 18144 23860
rect 17911 23820 18144 23848
rect 17911 23817 17923 23820
rect 17865 23811 17923 23817
rect 18138 23808 18144 23820
rect 18196 23808 18202 23860
rect 18325 23851 18383 23857
rect 18325 23817 18337 23851
rect 18371 23848 18383 23851
rect 18506 23848 18512 23860
rect 18371 23820 18512 23848
rect 18371 23817 18383 23820
rect 18325 23811 18383 23817
rect 18506 23808 18512 23820
rect 18564 23808 18570 23860
rect 18693 23851 18751 23857
rect 18693 23817 18705 23851
rect 18739 23848 18751 23851
rect 18874 23848 18880 23860
rect 18739 23820 18880 23848
rect 18739 23817 18751 23820
rect 18693 23811 18751 23817
rect 18874 23808 18880 23820
rect 18932 23808 18938 23860
rect 19886 23848 19892 23860
rect 19847 23820 19892 23848
rect 19886 23808 19892 23820
rect 19944 23808 19950 23860
rect 20530 23848 20536 23860
rect 20443 23820 20536 23848
rect 20530 23808 20536 23820
rect 20588 23848 20594 23860
rect 21266 23848 21272 23860
rect 20588 23820 21272 23848
rect 20588 23808 20594 23820
rect 21266 23808 21272 23820
rect 21324 23808 21330 23860
rect 22186 23848 22192 23860
rect 22147 23820 22192 23848
rect 22186 23808 22192 23820
rect 22244 23808 22250 23860
rect 22922 23848 22928 23860
rect 22883 23820 22928 23848
rect 22922 23808 22928 23820
rect 22980 23808 22986 23860
rect 24210 23808 24216 23860
rect 24268 23848 24274 23860
rect 24673 23851 24731 23857
rect 24673 23848 24685 23851
rect 24268 23820 24685 23848
rect 24268 23808 24274 23820
rect 24673 23817 24685 23820
rect 24719 23817 24731 23851
rect 26418 23848 26424 23860
rect 26379 23820 26424 23848
rect 24673 23811 24731 23817
rect 26418 23808 26424 23820
rect 26476 23808 26482 23860
rect 27249 23851 27307 23857
rect 27249 23817 27261 23851
rect 27295 23848 27307 23851
rect 27614 23848 27620 23860
rect 27295 23820 27620 23848
rect 27295 23817 27307 23820
rect 27249 23811 27307 23817
rect 27614 23808 27620 23820
rect 27672 23848 27678 23860
rect 27890 23848 27896 23860
rect 27672 23820 27896 23848
rect 27672 23808 27678 23820
rect 27890 23808 27896 23820
rect 27948 23808 27954 23860
rect 28718 23848 28724 23860
rect 28679 23820 28724 23848
rect 28718 23808 28724 23820
rect 28776 23808 28782 23860
rect 29454 23848 29460 23860
rect 29415 23820 29460 23848
rect 29454 23808 29460 23820
rect 29512 23808 29518 23860
rect 30466 23808 30472 23860
rect 30524 23848 30530 23860
rect 30745 23851 30803 23857
rect 30745 23848 30757 23851
rect 30524 23820 30757 23848
rect 30524 23808 30530 23820
rect 30745 23817 30757 23820
rect 30791 23817 30803 23851
rect 30745 23811 30803 23817
rect 33689 23851 33747 23857
rect 33689 23817 33701 23851
rect 33735 23848 33747 23851
rect 33778 23848 33784 23860
rect 33735 23820 33784 23848
rect 33735 23817 33747 23820
rect 33689 23811 33747 23817
rect 33778 23808 33784 23820
rect 33836 23848 33842 23860
rect 34238 23848 34244 23860
rect 33836 23820 34244 23848
rect 33836 23808 33842 23820
rect 34238 23808 34244 23820
rect 34296 23808 34302 23860
rect 36538 23848 36544 23860
rect 36499 23820 36544 23848
rect 36538 23808 36544 23820
rect 36596 23808 36602 23860
rect 36630 23808 36636 23860
rect 36688 23848 36694 23860
rect 36909 23851 36967 23857
rect 36909 23848 36921 23851
rect 36688 23820 36921 23848
rect 36688 23808 36694 23820
rect 36909 23817 36921 23820
rect 36955 23817 36967 23851
rect 36909 23811 36967 23817
rect 38565 23851 38623 23857
rect 38565 23817 38577 23851
rect 38611 23848 38623 23851
rect 38654 23848 38660 23860
rect 38611 23820 38660 23848
rect 38611 23817 38623 23820
rect 38565 23811 38623 23817
rect 19426 23780 19432 23792
rect 19387 23752 19432 23780
rect 19426 23740 19432 23752
rect 19484 23740 19490 23792
rect 20070 23740 20076 23792
rect 20128 23780 20134 23792
rect 21726 23780 21732 23792
rect 20128 23752 21732 23780
rect 20128 23740 20134 23752
rect 21726 23740 21732 23752
rect 21784 23740 21790 23792
rect 30377 23783 30435 23789
rect 30377 23749 30389 23783
rect 30423 23780 30435 23783
rect 31018 23780 31024 23792
rect 30423 23752 31024 23780
rect 30423 23749 30435 23752
rect 30377 23743 30435 23749
rect 31018 23740 31024 23752
rect 31076 23780 31082 23792
rect 32953 23783 33011 23789
rect 32953 23780 32965 23783
rect 31076 23752 32965 23780
rect 31076 23740 31082 23752
rect 32953 23749 32965 23752
rect 32999 23749 33011 23783
rect 35802 23780 35808 23792
rect 35763 23752 35808 23780
rect 32953 23743 33011 23749
rect 35802 23740 35808 23752
rect 35860 23740 35866 23792
rect 18138 23712 18144 23724
rect 14424 23684 15792 23712
rect 17098 23684 18144 23712
rect 14424 23672 14430 23684
rect 14052 23647 14110 23653
rect 14052 23613 14064 23647
rect 14098 23644 14110 23647
rect 14458 23644 14464 23656
rect 14098 23616 14464 23644
rect 14098 23613 14110 23616
rect 14052 23607 14110 23613
rect 14458 23604 14464 23616
rect 14516 23604 14522 23656
rect 15764 23644 15792 23684
rect 18138 23672 18144 23684
rect 18196 23672 18202 23724
rect 18877 23715 18935 23721
rect 18877 23681 18889 23715
rect 18923 23712 18935 23715
rect 19150 23712 19156 23724
rect 18923 23684 19156 23712
rect 18923 23681 18935 23684
rect 18877 23675 18935 23681
rect 19150 23672 19156 23684
rect 19208 23672 19214 23724
rect 20993 23715 21051 23721
rect 20993 23681 21005 23715
rect 21039 23712 21051 23715
rect 21174 23712 21180 23724
rect 21039 23684 21180 23712
rect 21039 23681 21051 23684
rect 20993 23675 21051 23681
rect 21174 23672 21180 23684
rect 21232 23712 21238 23724
rect 22557 23715 22615 23721
rect 22557 23712 22569 23715
rect 21232 23684 22569 23712
rect 21232 23672 21238 23684
rect 22557 23681 22569 23684
rect 22603 23681 22615 23715
rect 22557 23675 22615 23681
rect 24397 23715 24455 23721
rect 24397 23681 24409 23715
rect 24443 23712 24455 23715
rect 25682 23712 25688 23724
rect 24443 23684 25688 23712
rect 24443 23681 24455 23684
rect 24397 23675 24455 23681
rect 25682 23672 25688 23684
rect 25740 23672 25746 23724
rect 26881 23715 26939 23721
rect 26881 23681 26893 23715
rect 26927 23712 26939 23715
rect 29822 23712 29828 23724
rect 26927 23684 27936 23712
rect 29783 23684 29828 23712
rect 26927 23681 26939 23684
rect 26881 23675 26939 23681
rect 16644 23647 16702 23653
rect 16644 23644 16656 23647
rect 15764 23616 16656 23644
rect 16644 23613 16656 23616
rect 16690 23644 16702 23647
rect 17037 23647 17095 23653
rect 17037 23644 17049 23647
rect 16690 23616 17049 23644
rect 16690 23613 16702 23616
rect 16644 23607 16702 23613
rect 17037 23613 17049 23616
rect 17083 23613 17095 23647
rect 17037 23607 17095 23613
rect 23477 23647 23535 23653
rect 23477 23613 23489 23647
rect 23523 23644 23535 23647
rect 23934 23644 23940 23656
rect 23523 23616 23940 23644
rect 23523 23613 23535 23616
rect 23477 23607 23535 23613
rect 23934 23604 23940 23616
rect 23992 23604 23998 23656
rect 24026 23604 24032 23656
rect 24084 23644 24090 23656
rect 24121 23647 24179 23653
rect 24121 23644 24133 23647
rect 24084 23616 24133 23644
rect 24084 23604 24090 23616
rect 24121 23613 24133 23616
rect 24167 23613 24179 23647
rect 27614 23644 27620 23656
rect 27575 23616 27620 23644
rect 24121 23607 24179 23613
rect 27614 23604 27620 23616
rect 27672 23604 27678 23656
rect 27908 23653 27936 23684
rect 29822 23672 29828 23684
rect 29880 23712 29886 23724
rect 30098 23712 30104 23724
rect 29880 23684 30104 23712
rect 29880 23672 29886 23684
rect 30098 23672 30104 23684
rect 30156 23672 30162 23724
rect 31481 23715 31539 23721
rect 31481 23681 31493 23715
rect 31527 23712 31539 23715
rect 32401 23715 32459 23721
rect 32401 23712 32413 23715
rect 31527 23684 32413 23712
rect 31527 23681 31539 23684
rect 31481 23675 31539 23681
rect 32401 23681 32413 23684
rect 32447 23712 32459 23715
rect 33226 23712 33232 23724
rect 32447 23684 33232 23712
rect 32447 23681 32459 23684
rect 32401 23675 32459 23681
rect 33226 23672 33232 23684
rect 33284 23672 33290 23724
rect 35253 23715 35311 23721
rect 35253 23681 35265 23715
rect 35299 23712 35311 23715
rect 36556 23712 36584 23808
rect 35299 23684 36584 23712
rect 35299 23681 35311 23684
rect 35253 23675 35311 23681
rect 27893 23647 27951 23653
rect 27893 23613 27905 23647
rect 27939 23644 27951 23647
rect 27982 23644 27988 23656
rect 27939 23616 27988 23644
rect 27939 23613 27951 23616
rect 27893 23607 27951 23613
rect 27982 23604 27988 23616
rect 28040 23604 28046 23656
rect 36354 23604 36360 23656
rect 36412 23644 36418 23656
rect 36924 23644 36952 23811
rect 38654 23808 38660 23820
rect 38712 23808 38718 23860
rect 40313 23851 40371 23857
rect 40313 23817 40325 23851
rect 40359 23848 40371 23851
rect 40494 23848 40500 23860
rect 40359 23820 40500 23848
rect 40359 23817 40371 23820
rect 40313 23811 40371 23817
rect 40494 23808 40500 23820
rect 40552 23808 40558 23860
rect 41230 23848 41236 23860
rect 41191 23820 41236 23848
rect 41230 23808 41236 23820
rect 41288 23808 41294 23860
rect 43438 23848 43444 23860
rect 42766 23820 43444 23848
rect 40911 23783 40969 23789
rect 40911 23749 40923 23783
rect 40957 23780 40969 23783
rect 42766 23780 42794 23820
rect 43438 23808 43444 23820
rect 43496 23848 43502 23860
rect 43717 23851 43775 23857
rect 43717 23848 43729 23851
rect 43496 23820 43729 23848
rect 43496 23808 43502 23820
rect 43717 23817 43729 23820
rect 43763 23817 43775 23851
rect 43717 23811 43775 23817
rect 40957 23752 42794 23780
rect 40957 23749 40969 23752
rect 40911 23743 40969 23749
rect 43254 23740 43260 23792
rect 43312 23780 43318 23792
rect 43349 23783 43407 23789
rect 43349 23780 43361 23783
rect 43312 23752 43361 23780
rect 43312 23740 43318 23752
rect 43349 23749 43361 23752
rect 43395 23749 43407 23783
rect 43349 23743 43407 23749
rect 37734 23712 37740 23724
rect 37695 23684 37740 23712
rect 37734 23672 37740 23684
rect 37792 23672 37798 23724
rect 38749 23715 38807 23721
rect 38749 23681 38761 23715
rect 38795 23712 38807 23715
rect 39114 23712 39120 23724
rect 38795 23684 39120 23712
rect 38795 23681 38807 23684
rect 38749 23675 38807 23681
rect 39114 23672 39120 23684
rect 39172 23672 39178 23724
rect 41877 23715 41935 23721
rect 41877 23681 41889 23715
rect 41923 23712 41935 23715
rect 42150 23712 42156 23724
rect 41923 23684 42156 23712
rect 41923 23681 41935 23684
rect 41877 23675 41935 23681
rect 42150 23672 42156 23684
rect 42208 23672 42214 23724
rect 37093 23647 37151 23653
rect 37093 23644 37105 23647
rect 36412 23616 37105 23644
rect 36412 23604 36418 23616
rect 37093 23613 37105 23616
rect 37139 23613 37151 23647
rect 37093 23607 37151 23613
rect 37182 23604 37188 23656
rect 37240 23644 37246 23656
rect 37553 23647 37611 23653
rect 37553 23644 37565 23647
rect 37240 23616 37565 23644
rect 37240 23604 37246 23616
rect 37553 23613 37565 23616
rect 37599 23644 37611 23647
rect 38194 23644 38200 23656
rect 37599 23616 38200 23644
rect 37599 23613 37611 23616
rect 37553 23607 37611 23613
rect 38194 23604 38200 23616
rect 38252 23604 38258 23656
rect 40770 23644 40776 23656
rect 40828 23653 40834 23656
rect 40828 23647 40866 23653
rect 40718 23616 40776 23644
rect 40770 23604 40776 23616
rect 40854 23644 40866 23647
rect 41601 23647 41659 23653
rect 41601 23644 41613 23647
rect 40854 23616 41613 23644
rect 40854 23613 40866 23616
rect 40828 23607 40866 23613
rect 41601 23613 41613 23616
rect 41647 23613 41659 23647
rect 41601 23607 41659 23613
rect 40828 23604 40834 23607
rect 10008 23548 13814 23576
rect 14139 23579 14197 23585
rect 10008 23536 10014 23548
rect 14139 23545 14151 23579
rect 14185 23576 14197 23579
rect 14734 23576 14740 23588
rect 14185 23548 14740 23576
rect 14185 23545 14197 23548
rect 14139 23539 14197 23545
rect 14734 23536 14740 23548
rect 14792 23536 14798 23588
rect 15102 23576 15108 23588
rect 15063 23548 15108 23576
rect 15102 23536 15108 23548
rect 15160 23536 15166 23588
rect 15206 23579 15264 23585
rect 15206 23545 15218 23579
rect 15252 23576 15264 23579
rect 15562 23576 15568 23588
rect 15252 23548 15568 23576
rect 15252 23545 15264 23548
rect 15206 23539 15264 23545
rect 15562 23536 15568 23548
rect 15620 23536 15626 23588
rect 15749 23579 15807 23585
rect 15749 23545 15761 23579
rect 15795 23576 15807 23579
rect 15838 23576 15844 23588
rect 15795 23548 15844 23576
rect 15795 23545 15807 23548
rect 15749 23539 15807 23545
rect 15838 23536 15844 23548
rect 15896 23536 15902 23588
rect 16022 23576 16028 23588
rect 15935 23548 16028 23576
rect 16022 23536 16028 23548
rect 16080 23536 16086 23588
rect 18874 23536 18880 23588
rect 18932 23576 18938 23588
rect 18969 23579 19027 23585
rect 18969 23576 18981 23579
rect 18932 23548 18981 23576
rect 18932 23536 18938 23548
rect 18969 23545 18981 23548
rect 19015 23545 19027 23579
rect 21314 23579 21372 23585
rect 21314 23576 21326 23579
rect 18969 23539 19027 23545
rect 20824 23548 21326 23576
rect 16114 23468 16120 23520
rect 16172 23508 16178 23520
rect 16715 23511 16773 23517
rect 16715 23508 16727 23511
rect 16172 23480 16727 23508
rect 16172 23468 16178 23480
rect 16715 23477 16727 23480
rect 16761 23477 16773 23511
rect 16715 23471 16773 23477
rect 20714 23468 20720 23520
rect 20772 23508 20778 23520
rect 20824 23517 20852 23548
rect 21314 23545 21326 23548
rect 21360 23545 21372 23579
rect 28074 23576 28080 23588
rect 28035 23548 28080 23576
rect 21314 23539 21372 23545
rect 28074 23536 28080 23548
rect 28132 23536 28138 23588
rect 28994 23536 29000 23588
rect 29052 23576 29058 23588
rect 29917 23579 29975 23585
rect 29052 23548 29776 23576
rect 29052 23536 29058 23548
rect 29748 23520 29776 23548
rect 29917 23545 29929 23579
rect 29963 23545 29975 23579
rect 29917 23539 29975 23545
rect 31849 23579 31907 23585
rect 31849 23545 31861 23579
rect 31895 23576 31907 23579
rect 32493 23579 32551 23585
rect 31895 23548 32327 23576
rect 31895 23545 31907 23548
rect 31849 23539 31907 23545
rect 20809 23511 20867 23517
rect 20809 23508 20821 23511
rect 20772 23480 20821 23508
rect 20772 23468 20778 23480
rect 20809 23477 20821 23480
rect 20855 23477 20867 23511
rect 20809 23471 20867 23477
rect 21450 23468 21456 23520
rect 21508 23508 21514 23520
rect 21913 23511 21971 23517
rect 21913 23508 21925 23511
rect 21508 23480 21925 23508
rect 21508 23468 21514 23480
rect 21913 23477 21925 23480
rect 21959 23477 21971 23511
rect 29730 23508 29736 23520
rect 29643 23480 29736 23508
rect 21913 23471 21971 23477
rect 29730 23468 29736 23480
rect 29788 23508 29794 23520
rect 29932 23508 29960 23539
rect 29788 23480 29960 23508
rect 29788 23468 29794 23480
rect 31754 23468 31760 23520
rect 31812 23508 31818 23520
rect 32125 23511 32183 23517
rect 32125 23508 32137 23511
rect 31812 23480 32137 23508
rect 31812 23468 31818 23480
rect 32125 23477 32137 23480
rect 32171 23477 32183 23511
rect 32299 23508 32327 23548
rect 32493 23545 32505 23579
rect 32539 23545 32551 23579
rect 32493 23539 32551 23545
rect 32508 23508 32536 23539
rect 33318 23536 33324 23588
rect 33376 23576 33382 23588
rect 33965 23579 34023 23585
rect 33965 23576 33977 23579
rect 33376 23548 33977 23576
rect 33376 23536 33382 23548
rect 33965 23545 33977 23548
rect 34011 23576 34023 23579
rect 34054 23576 34060 23588
rect 34011 23548 34060 23576
rect 34011 23545 34023 23548
rect 33965 23539 34023 23545
rect 34054 23536 34060 23548
rect 34112 23536 34118 23588
rect 35342 23585 35348 23588
rect 34701 23579 34759 23585
rect 34701 23545 34713 23579
rect 34747 23576 34759 23579
rect 35338 23576 35348 23585
rect 34747 23548 35348 23576
rect 34747 23545 34759 23548
rect 34701 23539 34759 23545
rect 35338 23539 35348 23548
rect 35400 23576 35406 23588
rect 36173 23579 36231 23585
rect 36173 23576 36185 23579
rect 35400 23548 36185 23576
rect 35342 23536 35348 23539
rect 35400 23536 35406 23548
rect 36173 23545 36185 23548
rect 36219 23545 36231 23579
rect 36173 23539 36231 23545
rect 38838 23536 38844 23588
rect 38896 23576 38902 23588
rect 38896 23548 38941 23576
rect 38896 23536 38902 23548
rect 39022 23536 39028 23588
rect 39080 23576 39086 23588
rect 39393 23579 39451 23585
rect 39393 23576 39405 23579
rect 39080 23548 39405 23576
rect 39080 23536 39086 23548
rect 39393 23545 39405 23548
rect 39439 23576 39451 23579
rect 39439 23548 41736 23576
rect 39439 23545 39451 23548
rect 39393 23539 39451 23545
rect 32950 23508 32956 23520
rect 32299 23480 32956 23508
rect 32125 23471 32183 23477
rect 32950 23468 32956 23480
rect 33008 23468 33014 23520
rect 38102 23508 38108 23520
rect 38063 23480 38108 23508
rect 38102 23468 38108 23480
rect 38160 23468 38166 23520
rect 41708 23508 41736 23548
rect 41966 23536 41972 23588
rect 42024 23576 42030 23588
rect 42521 23579 42579 23585
rect 42521 23576 42533 23579
rect 42024 23548 42069 23576
rect 42260 23548 42533 23576
rect 42024 23536 42030 23548
rect 42260 23508 42288 23548
rect 42521 23545 42533 23548
rect 42567 23545 42579 23579
rect 42521 23539 42579 23545
rect 41708 23480 42288 23508
rect 42794 23468 42800 23520
rect 42852 23508 42858 23520
rect 42852 23480 42897 23508
rect 42852 23468 42858 23480
rect 1104 23418 48852 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 48852 23418
rect 1104 23344 48852 23366
rect 12989 23307 13047 23313
rect 12989 23273 13001 23307
rect 13035 23304 13047 23307
rect 13446 23304 13452 23316
rect 13035 23276 13452 23304
rect 13035 23273 13047 23276
rect 12989 23267 13047 23273
rect 13446 23264 13452 23276
rect 13504 23264 13510 23316
rect 14323 23307 14381 23313
rect 14323 23273 14335 23307
rect 14369 23304 14381 23307
rect 15102 23304 15108 23316
rect 14369 23276 15108 23304
rect 14369 23273 14381 23276
rect 14323 23267 14381 23273
rect 15102 23264 15108 23276
rect 15160 23264 15166 23316
rect 15562 23304 15568 23316
rect 15475 23276 15568 23304
rect 15488 23245 15516 23276
rect 15562 23264 15568 23276
rect 15620 23304 15626 23316
rect 15930 23304 15936 23316
rect 15620 23276 15936 23304
rect 15620 23264 15626 23276
rect 15930 23264 15936 23276
rect 15988 23264 15994 23316
rect 18782 23304 18788 23316
rect 18743 23276 18788 23304
rect 18782 23264 18788 23276
rect 18840 23264 18846 23316
rect 19242 23264 19248 23316
rect 19300 23304 19306 23316
rect 19978 23304 19984 23316
rect 19300 23276 19984 23304
rect 19300 23264 19306 23276
rect 19978 23264 19984 23276
rect 20036 23264 20042 23316
rect 20346 23264 20352 23316
rect 20404 23304 20410 23316
rect 20806 23304 20812 23316
rect 20404 23276 20812 23304
rect 20404 23264 20410 23276
rect 20806 23264 20812 23276
rect 20864 23304 20870 23316
rect 23842 23304 23848 23316
rect 20864 23276 21680 23304
rect 20864 23264 20870 23276
rect 15473 23239 15531 23245
rect 15473 23205 15485 23239
rect 15519 23205 15531 23239
rect 15473 23199 15531 23205
rect 17129 23239 17187 23245
rect 17129 23205 17141 23239
rect 17175 23236 17187 23239
rect 17218 23236 17224 23248
rect 17175 23208 17224 23236
rect 17175 23205 17187 23208
rect 17129 23199 17187 23205
rect 17218 23196 17224 23208
rect 17276 23196 17282 23248
rect 19058 23196 19064 23248
rect 19116 23236 19122 23248
rect 19116 23208 19161 23236
rect 19116 23196 19122 23208
rect 20990 23196 20996 23248
rect 21048 23236 21054 23248
rect 21085 23239 21143 23245
rect 21085 23236 21097 23239
rect 21048 23208 21097 23236
rect 21048 23196 21054 23208
rect 21085 23205 21097 23208
rect 21131 23205 21143 23239
rect 21085 23199 21143 23205
rect 11882 23168 11888 23180
rect 11843 23140 11888 23168
rect 11882 23128 11888 23140
rect 11940 23128 11946 23180
rect 12342 23168 12348 23180
rect 12303 23140 12348 23168
rect 12342 23128 12348 23140
rect 12400 23128 12406 23180
rect 14185 23171 14243 23177
rect 14185 23137 14197 23171
rect 14231 23168 14243 23171
rect 14274 23168 14280 23180
rect 14231 23140 14280 23168
rect 14231 23137 14243 23140
rect 14185 23131 14243 23137
rect 14274 23128 14280 23140
rect 14332 23128 14338 23180
rect 12434 23100 12440 23112
rect 12395 23072 12440 23100
rect 12434 23060 12440 23072
rect 12492 23060 12498 23112
rect 15378 23100 15384 23112
rect 15339 23072 15384 23100
rect 15378 23060 15384 23072
rect 15436 23060 15442 23112
rect 15838 23060 15844 23112
rect 15896 23100 15902 23112
rect 17034 23100 17040 23112
rect 15896 23072 16942 23100
rect 16995 23072 17040 23100
rect 15896 23060 15902 23072
rect 15933 23035 15991 23041
rect 15933 23001 15945 23035
rect 15979 23001 15991 23035
rect 16914 23032 16942 23072
rect 17034 23060 17040 23072
rect 17092 23060 17098 23112
rect 17313 23103 17371 23109
rect 17313 23069 17325 23103
rect 17359 23069 17371 23103
rect 18966 23100 18972 23112
rect 18927 23072 18972 23100
rect 17313 23063 17371 23069
rect 17328 23032 17356 23063
rect 18966 23060 18972 23072
rect 19024 23060 19030 23112
rect 19610 23100 19616 23112
rect 19571 23072 19616 23100
rect 19610 23060 19616 23072
rect 19668 23060 19674 23112
rect 20993 23103 21051 23109
rect 20993 23069 21005 23103
rect 21039 23069 21051 23103
rect 21652 23100 21680 23276
rect 23676 23276 23848 23304
rect 23676 23245 23704 23276
rect 23842 23264 23848 23276
rect 23900 23304 23906 23316
rect 23937 23307 23995 23313
rect 23937 23304 23949 23307
rect 23900 23276 23949 23304
rect 23900 23264 23906 23276
rect 23937 23273 23949 23276
rect 23983 23273 23995 23307
rect 23937 23267 23995 23273
rect 27433 23307 27491 23313
rect 27433 23273 27445 23307
rect 27479 23304 27491 23307
rect 27890 23304 27896 23316
rect 27479 23276 27896 23304
rect 27479 23273 27491 23276
rect 27433 23267 27491 23273
rect 27890 23264 27896 23276
rect 27948 23264 27954 23316
rect 29365 23307 29423 23313
rect 29365 23273 29377 23307
rect 29411 23304 29423 23307
rect 30098 23304 30104 23316
rect 29411 23276 30104 23304
rect 29411 23273 29423 23276
rect 29365 23267 29423 23273
rect 30098 23264 30104 23276
rect 30156 23264 30162 23316
rect 30377 23307 30435 23313
rect 30377 23273 30389 23307
rect 30423 23304 30435 23307
rect 30466 23304 30472 23316
rect 30423 23276 30472 23304
rect 30423 23273 30435 23276
rect 30377 23267 30435 23273
rect 30466 23264 30472 23276
rect 30524 23264 30530 23316
rect 32950 23264 32956 23316
rect 33008 23304 33014 23316
rect 33045 23307 33103 23313
rect 33045 23304 33057 23307
rect 33008 23276 33057 23304
rect 33008 23264 33014 23276
rect 33045 23273 33057 23276
rect 33091 23273 33103 23307
rect 37090 23304 37096 23316
rect 37051 23276 37096 23304
rect 33045 23267 33103 23273
rect 37090 23264 37096 23276
rect 37148 23264 37154 23316
rect 37918 23264 37924 23316
rect 37976 23304 37982 23316
rect 38013 23307 38071 23313
rect 38013 23304 38025 23307
rect 37976 23276 38025 23304
rect 37976 23264 37982 23276
rect 38013 23273 38025 23276
rect 38059 23304 38071 23307
rect 38749 23307 38807 23313
rect 38749 23304 38761 23307
rect 38059 23276 38761 23304
rect 38059 23273 38071 23276
rect 38013 23267 38071 23273
rect 38749 23273 38761 23276
rect 38795 23273 38807 23307
rect 39206 23304 39212 23316
rect 39167 23276 39212 23304
rect 38749 23267 38807 23273
rect 39206 23264 39212 23276
rect 39264 23264 39270 23316
rect 41230 23304 41236 23316
rect 41191 23276 41236 23304
rect 41230 23264 41236 23276
rect 41288 23264 41294 23316
rect 41785 23307 41843 23313
rect 41785 23273 41797 23307
rect 41831 23304 41843 23307
rect 41966 23304 41972 23316
rect 41831 23276 41972 23304
rect 41831 23273 41843 23276
rect 41785 23267 41843 23273
rect 41966 23264 41972 23276
rect 42024 23304 42030 23316
rect 42061 23307 42119 23313
rect 42061 23304 42073 23307
rect 42024 23276 42073 23304
rect 42024 23264 42030 23276
rect 42061 23273 42073 23276
rect 42107 23273 42119 23307
rect 42061 23267 42119 23273
rect 42150 23264 42156 23316
rect 42208 23304 42214 23316
rect 42429 23307 42487 23313
rect 42429 23304 42441 23307
rect 42208 23276 42441 23304
rect 42208 23264 42214 23276
rect 42429 23273 42441 23276
rect 42475 23304 42487 23307
rect 44082 23304 44088 23316
rect 42475 23276 44088 23304
rect 42475 23273 42487 23276
rect 42429 23267 42487 23273
rect 44082 23264 44088 23276
rect 44140 23264 44146 23316
rect 23661 23239 23719 23245
rect 23661 23205 23673 23239
rect 23707 23205 23719 23239
rect 23661 23199 23719 23205
rect 28071 23239 28129 23245
rect 28071 23205 28083 23239
rect 28117 23236 28129 23239
rect 28258 23236 28264 23248
rect 28117 23208 28264 23236
rect 28117 23205 28129 23208
rect 28071 23199 28129 23205
rect 28258 23196 28264 23208
rect 28316 23236 28322 23248
rect 29778 23239 29836 23245
rect 29778 23236 29790 23239
rect 28316 23208 29790 23236
rect 28316 23196 28322 23208
rect 29778 23205 29790 23208
rect 29824 23205 29836 23239
rect 29778 23199 29836 23205
rect 32487 23239 32545 23245
rect 32487 23205 32499 23239
rect 32533 23236 32545 23239
rect 32582 23236 32588 23248
rect 32533 23208 32588 23236
rect 32533 23205 32545 23208
rect 32487 23199 32545 23205
rect 32582 23196 32588 23208
rect 32640 23196 32646 23248
rect 34422 23196 34428 23248
rect 34480 23236 34486 23248
rect 34698 23236 34704 23248
rect 34480 23208 34704 23236
rect 34480 23196 34486 23208
rect 34698 23196 34704 23208
rect 34756 23236 34762 23248
rect 34838 23239 34896 23245
rect 34838 23236 34850 23239
rect 34756 23208 34850 23236
rect 34756 23196 34762 23208
rect 34838 23205 34850 23208
rect 34884 23205 34896 23239
rect 34838 23199 34896 23205
rect 22922 23168 22928 23180
rect 22883 23140 22928 23168
rect 22922 23128 22928 23140
rect 22980 23128 22986 23180
rect 23382 23128 23388 23180
rect 23440 23168 23446 23180
rect 23477 23171 23535 23177
rect 23477 23168 23489 23171
rect 23440 23140 23489 23168
rect 23440 23128 23446 23140
rect 23477 23137 23489 23140
rect 23523 23168 23535 23171
rect 24026 23168 24032 23180
rect 23523 23140 24032 23168
rect 23523 23137 23535 23140
rect 23477 23131 23535 23137
rect 24026 23128 24032 23140
rect 24084 23128 24090 23180
rect 24486 23168 24492 23180
rect 24447 23140 24492 23168
rect 24486 23128 24492 23140
rect 24544 23128 24550 23180
rect 25222 23168 25228 23180
rect 25183 23140 25228 23168
rect 25222 23128 25228 23140
rect 25280 23128 25286 23180
rect 26326 23128 26332 23180
rect 26384 23168 26390 23180
rect 26513 23171 26571 23177
rect 26513 23168 26525 23171
rect 26384 23140 26525 23168
rect 26384 23128 26390 23140
rect 26513 23137 26525 23140
rect 26559 23168 26571 23171
rect 26970 23168 26976 23180
rect 26559 23140 26976 23168
rect 26559 23137 26571 23140
rect 26513 23131 26571 23137
rect 26970 23128 26976 23140
rect 27028 23128 27034 23180
rect 30374 23128 30380 23180
rect 30432 23168 30438 23180
rect 30653 23171 30711 23177
rect 30653 23168 30665 23171
rect 30432 23140 30665 23168
rect 30432 23128 30438 23140
rect 30653 23137 30665 23140
rect 30699 23137 30711 23171
rect 36262 23168 36268 23180
rect 36223 23140 36268 23168
rect 30653 23131 30711 23137
rect 36262 23128 36268 23140
rect 36320 23128 36326 23180
rect 37918 23168 37924 23180
rect 37879 23140 37924 23168
rect 37918 23128 37924 23140
rect 37976 23128 37982 23180
rect 38286 23168 38292 23180
rect 38247 23140 38292 23168
rect 38286 23128 38292 23140
rect 38344 23128 38350 23180
rect 39298 23168 39304 23180
rect 39259 23140 39304 23168
rect 39298 23128 39304 23140
rect 39356 23128 39362 23180
rect 39758 23168 39764 23180
rect 39719 23140 39764 23168
rect 39758 23128 39764 23140
rect 39816 23128 39822 23180
rect 40218 23128 40224 23180
rect 40276 23168 40282 23180
rect 42794 23168 42800 23180
rect 40276 23140 42800 23168
rect 40276 23128 40282 23140
rect 42794 23128 42800 23140
rect 42852 23128 42858 23180
rect 24857 23103 24915 23109
rect 24857 23100 24869 23103
rect 21652 23072 24869 23100
rect 20993 23063 21051 23069
rect 24857 23069 24869 23072
rect 24903 23100 24915 23103
rect 26418 23100 26424 23112
rect 24903 23072 26424 23100
rect 24903 23069 24915 23072
rect 24857 23063 24915 23069
rect 19426 23032 19432 23044
rect 16914 23004 19432 23032
rect 15933 22995 15991 23001
rect 15654 22924 15660 22976
rect 15712 22964 15718 22976
rect 15948 22964 15976 22995
rect 19426 22992 19432 23004
rect 19484 23032 19490 23044
rect 21008 23032 21036 23063
rect 26418 23060 26424 23072
rect 26476 23060 26482 23112
rect 27065 23103 27123 23109
rect 27065 23069 27077 23103
rect 27111 23100 27123 23103
rect 27706 23100 27712 23112
rect 27111 23072 27712 23100
rect 27111 23069 27123 23072
rect 27065 23063 27123 23069
rect 27706 23060 27712 23072
rect 27764 23060 27770 23112
rect 28810 23060 28816 23112
rect 28868 23100 28874 23112
rect 29457 23103 29515 23109
rect 29457 23100 29469 23103
rect 28868 23072 29469 23100
rect 28868 23060 28874 23072
rect 29457 23069 29469 23072
rect 29503 23069 29515 23103
rect 32122 23100 32128 23112
rect 32083 23072 32128 23100
rect 29457 23063 29515 23069
rect 32122 23060 32128 23072
rect 32180 23060 32186 23112
rect 34514 23100 34520 23112
rect 34475 23072 34520 23100
rect 34514 23060 34520 23072
rect 34572 23060 34578 23112
rect 40037 23103 40095 23109
rect 40037 23069 40049 23103
rect 40083 23100 40095 23103
rect 40865 23103 40923 23109
rect 40865 23100 40877 23103
rect 40083 23072 40877 23100
rect 40083 23069 40095 23072
rect 40037 23063 40095 23069
rect 40865 23069 40877 23072
rect 40911 23100 40923 23103
rect 41690 23100 41696 23112
rect 40911 23072 41696 23100
rect 40911 23069 40923 23072
rect 40865 23063 40923 23069
rect 41690 23060 41696 23072
rect 41748 23060 41754 23112
rect 21542 23032 21548 23044
rect 19484 23004 21036 23032
rect 21503 23004 21548 23032
rect 19484 22992 19490 23004
rect 21542 22992 21548 23004
rect 21600 22992 21606 23044
rect 25314 22992 25320 23044
rect 25372 23032 25378 23044
rect 31018 23032 31024 23044
rect 25372 23004 31024 23032
rect 25372 22992 25378 23004
rect 31018 22992 31024 23004
rect 31076 22992 31082 23044
rect 17770 22964 17776 22976
rect 15712 22936 17776 22964
rect 15712 22924 15718 22936
rect 17770 22924 17776 22936
rect 17828 22924 17834 22976
rect 26694 22964 26700 22976
rect 26655 22936 26700 22964
rect 26694 22924 26700 22936
rect 26752 22924 26758 22976
rect 28626 22964 28632 22976
rect 28587 22936 28632 22964
rect 28626 22924 28632 22936
rect 28684 22924 28690 22976
rect 35342 22924 35348 22976
rect 35400 22964 35406 22976
rect 35437 22967 35495 22973
rect 35437 22964 35449 22967
rect 35400 22936 35449 22964
rect 35400 22924 35406 22936
rect 35437 22933 35449 22936
rect 35483 22964 35495 22967
rect 35713 22967 35771 22973
rect 35713 22964 35725 22967
rect 35483 22936 35725 22964
rect 35483 22933 35495 22936
rect 35437 22927 35495 22933
rect 35713 22933 35725 22936
rect 35759 22933 35771 22967
rect 35713 22927 35771 22933
rect 35802 22924 35808 22976
rect 35860 22964 35866 22976
rect 36403 22967 36461 22973
rect 36403 22964 36415 22967
rect 35860 22936 36415 22964
rect 35860 22924 35866 22936
rect 36403 22933 36415 22936
rect 36449 22933 36461 22967
rect 36403 22927 36461 22933
rect 1104 22874 48852 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 48852 22874
rect 1104 22800 48852 22822
rect 13357 22763 13415 22769
rect 13357 22729 13369 22763
rect 13403 22760 13415 22763
rect 14274 22760 14280 22772
rect 13403 22732 13814 22760
rect 14235 22732 14280 22760
rect 13403 22729 13415 22732
rect 13357 22723 13415 22729
rect 13786 22692 13814 22732
rect 14274 22720 14280 22732
rect 14332 22720 14338 22772
rect 16577 22763 16635 22769
rect 16577 22729 16589 22763
rect 16623 22760 16635 22763
rect 16807 22763 16865 22769
rect 16807 22760 16819 22763
rect 16623 22732 16819 22760
rect 16623 22729 16635 22732
rect 16577 22723 16635 22729
rect 16807 22729 16819 22732
rect 16853 22760 16865 22763
rect 17034 22760 17040 22772
rect 16853 22732 17040 22760
rect 16853 22729 16865 22732
rect 16807 22723 16865 22729
rect 17034 22720 17040 22732
rect 17092 22720 17098 22772
rect 17221 22763 17279 22769
rect 17221 22729 17233 22763
rect 17267 22760 17279 22763
rect 17310 22760 17316 22772
rect 17267 22732 17316 22760
rect 17267 22729 17279 22732
rect 17221 22723 17279 22729
rect 15470 22692 15476 22704
rect 13786 22664 15476 22692
rect 15470 22652 15476 22664
rect 15528 22652 15534 22704
rect 15654 22692 15660 22704
rect 15615 22664 15660 22692
rect 15654 22652 15660 22664
rect 15712 22652 15718 22704
rect 12434 22624 12440 22636
rect 12395 22596 12440 22624
rect 12434 22584 12440 22596
rect 12492 22584 12498 22636
rect 15102 22624 15108 22636
rect 15015 22596 15108 22624
rect 15102 22584 15108 22596
rect 15160 22624 15166 22636
rect 16114 22624 16120 22636
rect 15160 22596 16120 22624
rect 15160 22584 15166 22596
rect 16114 22584 16120 22596
rect 16172 22584 16178 22636
rect 16736 22559 16794 22565
rect 16736 22525 16748 22559
rect 16782 22556 16794 22559
rect 17236 22556 17264 22723
rect 17310 22720 17316 22732
rect 17368 22720 17374 22772
rect 19426 22720 19432 22772
rect 19484 22760 19490 22772
rect 20165 22763 20223 22769
rect 20165 22760 20177 22763
rect 19484 22732 20177 22760
rect 19484 22720 19490 22732
rect 20165 22729 20177 22732
rect 20211 22729 20223 22763
rect 20990 22760 20996 22772
rect 20951 22732 20996 22760
rect 20165 22723 20223 22729
rect 20990 22720 20996 22732
rect 21048 22720 21054 22772
rect 21085 22763 21143 22769
rect 21085 22729 21097 22763
rect 21131 22760 21143 22763
rect 22922 22760 22928 22772
rect 21131 22732 22928 22760
rect 21131 22729 21143 22732
rect 21085 22723 21143 22729
rect 22922 22720 22928 22732
rect 22980 22720 22986 22772
rect 23382 22760 23388 22772
rect 23343 22732 23388 22760
rect 23382 22720 23388 22732
rect 23440 22720 23446 22772
rect 24486 22760 24492 22772
rect 24447 22732 24492 22760
rect 24486 22720 24492 22732
rect 24544 22720 24550 22772
rect 28258 22720 28264 22772
rect 28316 22760 28322 22772
rect 28353 22763 28411 22769
rect 28353 22760 28365 22763
rect 28316 22732 28365 22760
rect 28316 22720 28322 22732
rect 28353 22729 28365 22732
rect 28399 22729 28411 22763
rect 28353 22723 28411 22729
rect 28810 22720 28816 22772
rect 28868 22760 28874 22772
rect 28997 22763 29055 22769
rect 28997 22760 29009 22763
rect 28868 22732 29009 22760
rect 28868 22720 28874 22732
rect 28997 22729 29009 22732
rect 29043 22729 29055 22763
rect 28997 22723 29055 22729
rect 31018 22720 31024 22772
rect 31076 22760 31082 22772
rect 32674 22760 32680 22772
rect 31076 22732 32680 22760
rect 31076 22720 31082 22732
rect 32674 22720 32680 22732
rect 32732 22760 32738 22772
rect 36262 22760 36268 22772
rect 32732 22732 36268 22760
rect 32732 22720 32738 22732
rect 36262 22720 36268 22732
rect 36320 22720 36326 22772
rect 38286 22720 38292 22772
rect 38344 22760 38350 22772
rect 38381 22763 38439 22769
rect 38381 22760 38393 22763
rect 38344 22732 38393 22760
rect 38344 22720 38350 22732
rect 38381 22729 38393 22732
rect 38427 22760 38439 22763
rect 39758 22760 39764 22772
rect 38427 22732 39764 22760
rect 38427 22729 38439 22732
rect 38381 22723 38439 22729
rect 39758 22720 39764 22732
rect 39816 22720 39822 22772
rect 41049 22763 41107 22769
rect 41049 22729 41061 22763
rect 41095 22760 41107 22763
rect 41230 22760 41236 22772
rect 41095 22732 41236 22760
rect 41095 22729 41107 22732
rect 41049 22723 41107 22729
rect 41230 22720 41236 22732
rect 41288 22720 41294 22772
rect 41690 22760 41696 22772
rect 41651 22732 41696 22760
rect 41690 22720 41696 22732
rect 41748 22720 41754 22772
rect 17770 22652 17776 22704
rect 17828 22692 17834 22704
rect 19610 22692 19616 22704
rect 17828 22664 19616 22692
rect 17828 22652 17834 22664
rect 19610 22652 19616 22664
rect 19668 22692 19674 22704
rect 22189 22695 22247 22701
rect 22189 22692 22201 22695
rect 19668 22664 22201 22692
rect 19668 22652 19674 22664
rect 18782 22624 18788 22636
rect 18743 22596 18788 22624
rect 18782 22584 18788 22596
rect 18840 22584 18846 22636
rect 19058 22624 19064 22636
rect 19019 22596 19064 22624
rect 19058 22584 19064 22596
rect 19116 22584 19122 22636
rect 19978 22584 19984 22636
rect 20036 22624 20042 22636
rect 21284 22633 21312 22664
rect 22189 22661 22201 22664
rect 22235 22661 22247 22695
rect 22189 22655 22247 22661
rect 21085 22627 21143 22633
rect 21085 22624 21097 22627
rect 20036 22596 21097 22624
rect 20036 22584 20042 22596
rect 21085 22593 21097 22596
rect 21131 22593 21143 22627
rect 21085 22587 21143 22593
rect 21269 22627 21327 22633
rect 21269 22593 21281 22627
rect 21315 22593 21327 22627
rect 21542 22624 21548 22636
rect 21503 22596 21548 22624
rect 21269 22587 21327 22593
rect 21542 22584 21548 22596
rect 21600 22584 21606 22636
rect 22940 22624 22968 22720
rect 23934 22652 23940 22704
rect 23992 22692 23998 22704
rect 23992 22664 28298 22692
rect 23992 22652 23998 22664
rect 27614 22624 27620 22636
rect 22940 22596 27292 22624
rect 23566 22556 23572 22568
rect 16782 22528 17264 22556
rect 23527 22528 23572 22556
rect 16782 22525 16794 22528
rect 16736 22519 16794 22525
rect 23566 22516 23572 22528
rect 23624 22516 23630 22568
rect 24213 22559 24271 22565
rect 24213 22525 24225 22559
rect 24259 22556 24271 22559
rect 25222 22556 25228 22568
rect 24259 22528 25228 22556
rect 24259 22525 24271 22528
rect 24213 22519 24271 22525
rect 25222 22516 25228 22528
rect 25280 22556 25286 22568
rect 25317 22559 25375 22565
rect 25317 22556 25329 22559
rect 25280 22528 25329 22556
rect 25280 22516 25286 22528
rect 25317 22525 25329 22528
rect 25363 22556 25375 22559
rect 26142 22556 26148 22568
rect 25363 22528 25820 22556
rect 26055 22528 26148 22556
rect 25363 22525 25375 22528
rect 25317 22519 25375 22525
rect 10502 22448 10508 22500
rect 10560 22488 10566 22500
rect 11793 22491 11851 22497
rect 11793 22488 11805 22491
rect 10560 22460 11805 22488
rect 10560 22448 10566 22460
rect 11793 22457 11805 22460
rect 11839 22488 11851 22491
rect 11882 22488 11888 22500
rect 11839 22460 11888 22488
rect 11839 22457 11851 22460
rect 11793 22451 11851 22457
rect 11882 22448 11888 22460
rect 11940 22448 11946 22500
rect 12802 22497 12808 22500
rect 12253 22491 12311 22497
rect 12253 22457 12265 22491
rect 12299 22488 12311 22491
rect 12758 22491 12808 22497
rect 12758 22488 12770 22491
rect 12299 22460 12770 22488
rect 12299 22457 12311 22460
rect 12253 22451 12311 22457
rect 12758 22457 12770 22460
rect 12804 22457 12808 22491
rect 12758 22451 12808 22457
rect 12802 22448 12808 22451
rect 12860 22448 12866 22500
rect 15197 22491 15255 22497
rect 15197 22457 15209 22491
rect 15243 22457 15255 22491
rect 15197 22451 15255 22457
rect 11238 22380 11244 22432
rect 11296 22420 11302 22432
rect 11425 22423 11483 22429
rect 11425 22420 11437 22423
rect 11296 22392 11437 22420
rect 11296 22380 11302 22392
rect 11425 22389 11437 22392
rect 11471 22389 11483 22423
rect 11425 22383 11483 22389
rect 14921 22423 14979 22429
rect 14921 22389 14933 22423
rect 14967 22420 14979 22423
rect 15212 22420 15240 22451
rect 15470 22448 15476 22500
rect 15528 22488 15534 22500
rect 17218 22488 17224 22500
rect 15528 22460 17224 22488
rect 15528 22448 15534 22460
rect 17218 22448 17224 22460
rect 17276 22488 17282 22500
rect 17497 22491 17555 22497
rect 17497 22488 17509 22491
rect 17276 22460 17509 22488
rect 17276 22448 17282 22460
rect 17497 22457 17509 22460
rect 17543 22457 17555 22491
rect 17497 22451 17555 22457
rect 18601 22491 18659 22497
rect 18601 22457 18613 22491
rect 18647 22488 18659 22491
rect 18874 22488 18880 22500
rect 18647 22460 18880 22488
rect 18647 22457 18659 22460
rect 18601 22451 18659 22457
rect 18874 22448 18880 22460
rect 18932 22448 18938 22500
rect 21361 22491 21419 22497
rect 21361 22457 21373 22491
rect 21407 22488 21419 22491
rect 21450 22488 21456 22500
rect 21407 22460 21456 22488
rect 21407 22457 21419 22460
rect 21361 22451 21419 22457
rect 15746 22420 15752 22432
rect 14967 22392 15752 22420
rect 14967 22389 14979 22392
rect 14921 22383 14979 22389
rect 15746 22380 15752 22392
rect 15804 22380 15810 22432
rect 15930 22380 15936 22432
rect 15988 22420 15994 22432
rect 16025 22423 16083 22429
rect 16025 22420 16037 22423
rect 15988 22392 16037 22420
rect 15988 22380 15994 22392
rect 16025 22389 16037 22392
rect 16071 22389 16083 22423
rect 18892 22420 18920 22448
rect 19705 22423 19763 22429
rect 19705 22420 19717 22423
rect 18892 22392 19717 22420
rect 16025 22383 16083 22389
rect 19705 22389 19717 22392
rect 19751 22389 19763 22423
rect 19705 22383 19763 22389
rect 20625 22423 20683 22429
rect 20625 22389 20637 22423
rect 20671 22420 20683 22423
rect 21376 22420 21404 22451
rect 21450 22448 21456 22460
rect 21508 22448 21514 22500
rect 24670 22488 24676 22500
rect 24631 22460 24676 22488
rect 24670 22448 24676 22460
rect 24728 22448 24734 22500
rect 25792 22432 25820 22528
rect 26142 22516 26148 22528
rect 26200 22556 26206 22568
rect 27264 22565 27292 22596
rect 27540 22596 27620 22624
rect 27540 22565 27568 22596
rect 27614 22584 27620 22596
rect 27672 22584 27678 22636
rect 27706 22584 27712 22636
rect 27764 22624 27770 22636
rect 27893 22627 27951 22633
rect 27893 22624 27905 22627
rect 27764 22596 27905 22624
rect 27764 22584 27770 22596
rect 27893 22593 27905 22596
rect 27939 22593 27951 22627
rect 28270 22624 28298 22664
rect 28718 22652 28724 22704
rect 28776 22692 28782 22704
rect 30098 22692 30104 22704
rect 28776 22664 30104 22692
rect 28776 22652 28782 22664
rect 30098 22652 30104 22664
rect 30156 22652 30162 22704
rect 32766 22692 32772 22704
rect 31588 22664 32772 22692
rect 29641 22627 29699 22633
rect 29641 22624 29653 22627
rect 28270 22596 29653 22624
rect 27893 22587 27951 22593
rect 29641 22593 29653 22596
rect 29687 22593 29699 22627
rect 29641 22587 29699 22593
rect 29825 22627 29883 22633
rect 29825 22593 29837 22627
rect 29871 22624 29883 22627
rect 30006 22624 30012 22636
rect 29871 22596 30012 22624
rect 29871 22593 29883 22596
rect 29825 22587 29883 22593
rect 30006 22584 30012 22596
rect 30064 22584 30070 22636
rect 30469 22627 30527 22633
rect 30469 22593 30481 22627
rect 30515 22624 30527 22627
rect 30926 22624 30932 22636
rect 30515 22596 30932 22624
rect 30515 22593 30527 22596
rect 30469 22587 30527 22593
rect 30926 22584 30932 22596
rect 30984 22584 30990 22636
rect 26237 22559 26295 22565
rect 26237 22556 26249 22559
rect 26200 22528 26249 22556
rect 26200 22516 26206 22528
rect 26237 22525 26249 22528
rect 26283 22525 26295 22559
rect 26237 22519 26295 22525
rect 27249 22559 27307 22565
rect 27249 22525 27261 22559
rect 27295 22556 27307 22559
rect 27525 22559 27583 22565
rect 27525 22556 27537 22559
rect 27295 22528 27537 22556
rect 27295 22525 27307 22528
rect 27249 22519 27307 22525
rect 27525 22525 27537 22528
rect 27571 22525 27583 22559
rect 27525 22519 27583 22525
rect 27801 22559 27859 22565
rect 27801 22525 27813 22559
rect 27847 22556 27859 22559
rect 27982 22556 27988 22568
rect 27847 22528 27988 22556
rect 27847 22525 27859 22528
rect 27801 22519 27859 22525
rect 27982 22516 27988 22528
rect 28040 22516 28046 22568
rect 31588 22565 31616 22664
rect 32766 22652 32772 22664
rect 32824 22652 32830 22704
rect 33594 22652 33600 22704
rect 33652 22692 33658 22704
rect 33962 22692 33968 22704
rect 33652 22664 33968 22692
rect 33652 22652 33658 22664
rect 33962 22652 33968 22664
rect 34020 22652 34026 22704
rect 32122 22584 32128 22636
rect 32180 22624 32186 22636
rect 32309 22627 32367 22633
rect 32309 22624 32321 22627
rect 32180 22596 32321 22624
rect 32180 22584 32186 22596
rect 32309 22593 32321 22596
rect 32355 22624 32367 22627
rect 32953 22627 33011 22633
rect 32953 22624 32965 22627
rect 32355 22596 32965 22624
rect 32355 22593 32367 22596
rect 32309 22587 32367 22593
rect 32953 22593 32965 22596
rect 32999 22593 33011 22627
rect 32953 22587 33011 22593
rect 35250 22584 35256 22636
rect 35308 22624 35314 22636
rect 35529 22627 35587 22633
rect 35529 22624 35541 22627
rect 35308 22596 35541 22624
rect 35308 22584 35314 22596
rect 35529 22593 35541 22596
rect 35575 22593 35587 22627
rect 36280 22624 36308 22720
rect 38562 22652 38568 22704
rect 38620 22692 38626 22704
rect 38746 22692 38752 22704
rect 38620 22664 38752 22692
rect 38620 22652 38626 22664
rect 38746 22652 38752 22664
rect 38804 22652 38810 22704
rect 39298 22692 39304 22704
rect 39259 22664 39304 22692
rect 39298 22652 39304 22664
rect 39356 22652 39362 22704
rect 42475 22695 42533 22701
rect 42475 22661 42487 22695
rect 42521 22692 42533 22695
rect 43438 22692 43444 22704
rect 42521 22664 43444 22692
rect 42521 22661 42533 22664
rect 42475 22655 42533 22661
rect 43438 22652 43444 22664
rect 43496 22652 43502 22704
rect 41325 22627 41383 22633
rect 41325 22624 41337 22627
rect 36280 22596 41337 22624
rect 35529 22587 35587 22593
rect 31297 22559 31355 22565
rect 31297 22525 31309 22559
rect 31343 22556 31355 22559
rect 31573 22559 31631 22565
rect 31573 22556 31585 22559
rect 31343 22528 31585 22556
rect 31343 22525 31355 22528
rect 31297 22519 31355 22525
rect 31573 22525 31585 22528
rect 31619 22525 31631 22559
rect 31573 22519 31631 22525
rect 31662 22516 31668 22568
rect 31720 22556 31726 22568
rect 32033 22559 32091 22565
rect 32033 22556 32045 22559
rect 31720 22528 32045 22556
rect 31720 22516 31726 22528
rect 32033 22525 32045 22528
rect 32079 22556 32091 22559
rect 33318 22556 33324 22568
rect 32079 22528 33324 22556
rect 32079 22525 32091 22528
rect 32033 22519 32091 22525
rect 33318 22516 33324 22528
rect 33376 22516 33382 22568
rect 33689 22559 33747 22565
rect 33689 22525 33701 22559
rect 33735 22556 33747 22559
rect 33778 22556 33784 22568
rect 33836 22565 33842 22568
rect 33836 22559 33874 22565
rect 33735 22528 33784 22556
rect 33735 22525 33747 22528
rect 33689 22519 33747 22525
rect 26326 22448 26332 22500
rect 26384 22488 26390 22500
rect 26697 22491 26755 22497
rect 26697 22488 26709 22491
rect 26384 22460 26709 22488
rect 26384 22448 26390 22460
rect 26697 22457 26709 22460
rect 26743 22457 26755 22491
rect 26697 22451 26755 22457
rect 28626 22448 28632 22500
rect 28684 22488 28690 22500
rect 29822 22488 29828 22500
rect 28684 22460 29828 22488
rect 28684 22448 28690 22460
rect 29822 22448 29828 22460
rect 29880 22488 29886 22500
rect 29917 22491 29975 22497
rect 29917 22488 29929 22491
rect 29880 22460 29929 22488
rect 29880 22448 29886 22460
rect 29917 22457 29929 22460
rect 29963 22457 29975 22491
rect 29917 22451 29975 22457
rect 30098 22448 30104 22500
rect 30156 22488 30162 22500
rect 33704 22488 33732 22519
rect 33778 22516 33784 22528
rect 33862 22525 33874 22559
rect 36909 22559 36967 22565
rect 36909 22556 36921 22559
rect 33836 22519 33874 22525
rect 36740 22528 36921 22556
rect 33836 22516 33842 22519
rect 30156 22460 33732 22488
rect 33919 22491 33977 22497
rect 30156 22448 30162 22460
rect 33919 22457 33931 22491
rect 33965 22488 33977 22491
rect 34882 22488 34888 22500
rect 33965 22460 34888 22488
rect 33965 22457 33977 22460
rect 33919 22451 33977 22457
rect 34882 22448 34888 22460
rect 34940 22488 34946 22500
rect 35253 22491 35311 22497
rect 35253 22488 35265 22491
rect 34940 22460 35265 22488
rect 34940 22448 34946 22460
rect 35253 22457 35265 22460
rect 35299 22457 35311 22491
rect 35253 22451 35311 22457
rect 35342 22448 35348 22500
rect 35400 22488 35406 22500
rect 35400 22460 35445 22488
rect 35400 22448 35406 22460
rect 20671 22392 21404 22420
rect 20671 22389 20683 22392
rect 20625 22383 20683 22389
rect 23658 22380 23664 22432
rect 23716 22420 23722 22432
rect 23799 22423 23857 22429
rect 23799 22420 23811 22423
rect 23716 22392 23811 22420
rect 23716 22380 23722 22392
rect 23799 22389 23811 22392
rect 23845 22389 23857 22423
rect 25774 22420 25780 22432
rect 25735 22392 25780 22420
rect 23799 22383 23857 22389
rect 25774 22380 25780 22392
rect 25832 22380 25838 22432
rect 26418 22420 26424 22432
rect 26379 22392 26424 22420
rect 26418 22380 26424 22392
rect 26476 22380 26482 22432
rect 28258 22380 28264 22432
rect 28316 22420 28322 22432
rect 29457 22423 29515 22429
rect 29457 22420 29469 22423
rect 28316 22392 29469 22420
rect 28316 22380 28322 22392
rect 29457 22389 29469 22392
rect 29503 22389 29515 22423
rect 29457 22383 29515 22389
rect 29638 22380 29644 22432
rect 29696 22420 29702 22432
rect 31297 22423 31355 22429
rect 31297 22420 31309 22423
rect 29696 22392 31309 22420
rect 29696 22380 29702 22392
rect 31297 22389 31309 22392
rect 31343 22420 31355 22423
rect 31389 22423 31447 22429
rect 31389 22420 31401 22423
rect 31343 22392 31401 22420
rect 31343 22389 31355 22392
rect 31297 22383 31355 22389
rect 31389 22389 31401 22392
rect 31435 22389 31447 22423
rect 32582 22420 32588 22432
rect 32543 22392 32588 22420
rect 31389 22383 31447 22389
rect 32582 22380 32588 22392
rect 32640 22420 32646 22432
rect 34517 22423 34575 22429
rect 34517 22420 34529 22423
rect 32640 22392 34529 22420
rect 32640 22380 32646 22392
rect 34517 22389 34529 22392
rect 34563 22420 34575 22423
rect 34698 22420 34704 22432
rect 34563 22392 34704 22420
rect 34563 22389 34575 22392
rect 34517 22383 34575 22389
rect 34698 22380 34704 22392
rect 34756 22380 34762 22432
rect 35710 22380 35716 22432
rect 35768 22420 35774 22432
rect 36170 22420 36176 22432
rect 35768 22392 36176 22420
rect 35768 22380 35774 22392
rect 36170 22380 36176 22392
rect 36228 22420 36234 22432
rect 36740 22429 36768 22528
rect 36909 22525 36921 22528
rect 36955 22525 36967 22559
rect 36909 22519 36967 22525
rect 37090 22516 37096 22568
rect 37148 22556 37154 22568
rect 37369 22559 37427 22565
rect 37369 22556 37381 22559
rect 37148 22528 37381 22556
rect 37148 22516 37154 22528
rect 37369 22525 37381 22528
rect 37415 22525 37427 22559
rect 37369 22519 37427 22525
rect 38524 22559 38582 22565
rect 38524 22525 38536 22559
rect 38570 22556 38582 22559
rect 38933 22559 38991 22565
rect 38933 22556 38945 22559
rect 38570 22528 38945 22556
rect 38570 22525 38582 22528
rect 38524 22519 38582 22525
rect 38933 22525 38945 22528
rect 38979 22556 38991 22559
rect 39022 22556 39028 22568
rect 38979 22528 39028 22556
rect 38979 22525 38991 22528
rect 38933 22519 38991 22525
rect 39022 22516 39028 22528
rect 39080 22516 39086 22568
rect 40547 22565 40575 22596
rect 41325 22593 41337 22596
rect 41371 22593 41383 22627
rect 41325 22587 41383 22593
rect 40532 22559 40590 22565
rect 40532 22525 40544 22559
rect 40578 22525 40590 22559
rect 41340 22556 41368 22587
rect 42372 22559 42430 22565
rect 42372 22556 42384 22559
rect 41340 22528 42384 22556
rect 40532 22519 40590 22525
rect 42372 22525 42384 22528
rect 42418 22556 42430 22559
rect 42518 22556 42524 22568
rect 42418 22528 42524 22556
rect 42418 22525 42430 22528
rect 42372 22519 42430 22525
rect 42518 22516 42524 22528
rect 42576 22556 42582 22568
rect 42797 22559 42855 22565
rect 42797 22556 42809 22559
rect 42576 22528 42809 22556
rect 42576 22516 42582 22528
rect 42797 22525 42809 22528
rect 42843 22525 42855 22559
rect 42797 22519 42855 22525
rect 43416 22559 43474 22565
rect 43416 22525 43428 22559
rect 43462 22556 43474 22559
rect 43806 22556 43812 22568
rect 43462 22528 43812 22556
rect 43462 22525 43474 22528
rect 43416 22519 43474 22525
rect 43806 22516 43812 22528
rect 43864 22516 43870 22568
rect 37642 22488 37648 22500
rect 37603 22460 37648 22488
rect 37642 22448 37648 22460
rect 37700 22448 37706 22500
rect 38378 22488 38384 22500
rect 37936 22460 38384 22488
rect 37936 22432 37964 22460
rect 38378 22448 38384 22460
rect 38436 22448 38442 22500
rect 36725 22423 36783 22429
rect 36725 22420 36737 22423
rect 36228 22392 36737 22420
rect 36228 22380 36234 22392
rect 36725 22389 36737 22392
rect 36771 22389 36783 22423
rect 37918 22420 37924 22432
rect 37879 22392 37924 22420
rect 36725 22383 36783 22389
rect 37918 22380 37924 22392
rect 37976 22380 37982 22432
rect 38010 22380 38016 22432
rect 38068 22420 38074 22432
rect 38611 22423 38669 22429
rect 38611 22420 38623 22423
rect 38068 22392 38623 22420
rect 38068 22380 38074 22392
rect 38611 22389 38623 22392
rect 38657 22389 38669 22423
rect 38611 22383 38669 22389
rect 38746 22380 38752 22432
rect 38804 22420 38810 22432
rect 40635 22423 40693 22429
rect 40635 22420 40647 22423
rect 38804 22392 40647 22420
rect 38804 22380 38810 22392
rect 40635 22389 40647 22392
rect 40681 22389 40693 22423
rect 40635 22383 40693 22389
rect 43487 22423 43545 22429
rect 43487 22389 43499 22423
rect 43533 22420 43545 22423
rect 43714 22420 43720 22432
rect 43533 22392 43720 22420
rect 43533 22389 43545 22392
rect 43487 22383 43545 22389
rect 43714 22380 43720 22392
rect 43772 22380 43778 22432
rect 1104 22330 48852 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 48852 22330
rect 1104 22256 48852 22278
rect 12434 22216 12440 22228
rect 12395 22188 12440 22216
rect 12434 22176 12440 22188
rect 12492 22176 12498 22228
rect 14737 22219 14795 22225
rect 14737 22185 14749 22219
rect 14783 22216 14795 22219
rect 14826 22216 14832 22228
rect 14783 22188 14832 22216
rect 14783 22185 14795 22188
rect 14737 22179 14795 22185
rect 14826 22176 14832 22188
rect 14884 22216 14890 22228
rect 15378 22216 15384 22228
rect 14884 22188 15384 22216
rect 14884 22176 14890 22188
rect 15378 22176 15384 22188
rect 15436 22176 15442 22228
rect 18966 22176 18972 22228
rect 19024 22216 19030 22228
rect 19429 22219 19487 22225
rect 19429 22216 19441 22219
rect 19024 22188 19441 22216
rect 19024 22176 19030 22188
rect 19429 22185 19441 22188
rect 19475 22216 19487 22219
rect 19751 22219 19809 22225
rect 19751 22216 19763 22219
rect 19475 22188 19763 22216
rect 19475 22185 19487 22188
rect 19429 22179 19487 22185
rect 19751 22185 19763 22188
rect 19797 22185 19809 22219
rect 19751 22179 19809 22185
rect 20254 22176 20260 22228
rect 20312 22216 20318 22228
rect 23477 22219 23535 22225
rect 23477 22216 23489 22219
rect 20312 22188 23489 22216
rect 20312 22176 20318 22188
rect 23477 22185 23489 22188
rect 23523 22185 23535 22219
rect 23477 22179 23535 22185
rect 23566 22176 23572 22228
rect 23624 22216 23630 22228
rect 23661 22219 23719 22225
rect 23661 22216 23673 22219
rect 23624 22188 23673 22216
rect 23624 22176 23630 22188
rect 23661 22185 23673 22188
rect 23707 22185 23719 22219
rect 28994 22216 29000 22228
rect 28955 22188 29000 22216
rect 23661 22179 23719 22185
rect 28994 22176 29000 22188
rect 29052 22176 29058 22228
rect 29822 22216 29828 22228
rect 29783 22188 29828 22216
rect 29822 22176 29828 22188
rect 29880 22176 29886 22228
rect 30006 22176 30012 22228
rect 30064 22216 30070 22228
rect 30101 22219 30159 22225
rect 30101 22216 30113 22219
rect 30064 22188 30113 22216
rect 30064 22176 30070 22188
rect 30101 22185 30113 22188
rect 30147 22185 30159 22219
rect 31662 22216 31668 22228
rect 31623 22188 31668 22216
rect 30101 22179 30159 22185
rect 31662 22176 31668 22188
rect 31720 22176 31726 22228
rect 34514 22216 34520 22228
rect 34475 22188 34520 22216
rect 34514 22176 34520 22188
rect 34572 22176 34578 22228
rect 34882 22216 34888 22228
rect 34843 22188 34888 22216
rect 34882 22176 34888 22188
rect 34940 22176 34946 22228
rect 35802 22216 35808 22228
rect 35176 22188 35808 22216
rect 12802 22108 12808 22160
rect 12860 22148 12866 22160
rect 13310 22151 13368 22157
rect 13310 22148 13322 22151
rect 12860 22120 13322 22148
rect 12860 22108 12866 22120
rect 13310 22117 13322 22120
rect 13356 22148 13368 22151
rect 14458 22148 14464 22160
rect 13356 22120 14464 22148
rect 13356 22117 13368 22120
rect 13310 22111 13368 22117
rect 14458 22108 14464 22120
rect 14516 22108 14522 22160
rect 15102 22148 15108 22160
rect 15063 22120 15108 22148
rect 15102 22108 15108 22120
rect 15160 22108 15166 22160
rect 15473 22151 15531 22157
rect 15473 22117 15485 22151
rect 15519 22148 15531 22151
rect 15746 22148 15752 22160
rect 15519 22120 15752 22148
rect 15519 22117 15531 22120
rect 15473 22111 15531 22117
rect 15746 22108 15752 22120
rect 15804 22108 15810 22160
rect 15838 22108 15844 22160
rect 15896 22148 15902 22160
rect 16025 22151 16083 22157
rect 16025 22148 16037 22151
rect 15896 22120 16037 22148
rect 15896 22108 15902 22120
rect 16025 22117 16037 22120
rect 16071 22117 16083 22151
rect 17218 22148 17224 22160
rect 17179 22120 17224 22148
rect 16025 22111 16083 22117
rect 17218 22108 17224 22120
rect 17276 22108 17282 22160
rect 17770 22148 17776 22160
rect 17731 22120 17776 22148
rect 17770 22108 17776 22120
rect 17828 22108 17834 22160
rect 18739 22151 18797 22157
rect 18739 22117 18751 22151
rect 18785 22148 18797 22151
rect 19150 22148 19156 22160
rect 18785 22120 19156 22148
rect 18785 22117 18797 22120
rect 18739 22111 18797 22117
rect 19150 22108 19156 22120
rect 19208 22108 19214 22160
rect 21266 22148 21272 22160
rect 21227 22120 21272 22148
rect 21266 22108 21272 22120
rect 21324 22108 21330 22160
rect 26418 22148 26424 22160
rect 23308 22120 26424 22148
rect 10042 22040 10048 22092
rect 10100 22080 10106 22092
rect 11701 22083 11759 22089
rect 11701 22080 11713 22083
rect 10100 22052 11713 22080
rect 10100 22040 10106 22052
rect 11701 22049 11713 22052
rect 11747 22080 11759 22083
rect 11790 22080 11796 22092
rect 11747 22052 11796 22080
rect 11747 22049 11759 22052
rect 11701 22043 11759 22049
rect 11790 22040 11796 22052
rect 11848 22040 11854 22092
rect 11977 22083 12035 22089
rect 11977 22049 11989 22083
rect 12023 22049 12035 22083
rect 12986 22080 12992 22092
rect 12947 22052 12992 22080
rect 11977 22043 12035 22049
rect 11238 21904 11244 21956
rect 11296 21944 11302 21956
rect 11992 21944 12020 22043
rect 12986 22040 12992 22052
rect 13044 22040 13050 22092
rect 18598 22080 18604 22092
rect 18559 22052 18604 22080
rect 18598 22040 18604 22052
rect 18656 22040 18662 22092
rect 19610 22080 19616 22092
rect 19571 22052 19616 22080
rect 19610 22040 19616 22052
rect 19668 22040 19674 22092
rect 22738 22040 22744 22092
rect 22796 22080 22802 22092
rect 23308 22089 23336 22120
rect 26418 22108 26424 22120
rect 26476 22108 26482 22160
rect 28258 22108 28264 22160
rect 28316 22148 28322 22160
rect 28398 22151 28456 22157
rect 28398 22148 28410 22151
rect 28316 22120 28410 22148
rect 28316 22108 28322 22120
rect 28398 22117 28410 22120
rect 28444 22117 28456 22151
rect 33410 22148 33416 22160
rect 28398 22111 28456 22117
rect 30852 22120 32076 22148
rect 33371 22120 33416 22148
rect 23293 22083 23351 22089
rect 23293 22080 23305 22083
rect 22796 22052 23305 22080
rect 22796 22040 22802 22052
rect 23293 22049 23305 22052
rect 23339 22049 23351 22083
rect 24486 22080 24492 22092
rect 24447 22052 24492 22080
rect 23293 22043 23351 22049
rect 24486 22040 24492 22052
rect 24544 22040 24550 22092
rect 24670 22080 24676 22092
rect 24631 22052 24676 22080
rect 24670 22040 24676 22052
rect 24728 22040 24734 22092
rect 26970 22080 26976 22092
rect 26931 22052 26976 22080
rect 26970 22040 26976 22052
rect 27028 22040 27034 22092
rect 30852 22080 30880 22120
rect 27080 22052 30880 22080
rect 27080 22024 27108 22052
rect 30926 22040 30932 22092
rect 30984 22080 30990 22092
rect 31056 22083 31114 22089
rect 31056 22080 31068 22083
rect 30984 22052 31068 22080
rect 30984 22040 30990 22052
rect 31056 22049 31068 22052
rect 31102 22049 31114 22083
rect 32048 22080 32076 22120
rect 33410 22108 33416 22120
rect 33468 22108 33474 22160
rect 35176 22157 35204 22188
rect 35802 22176 35808 22188
rect 35860 22176 35866 22228
rect 38286 22216 38292 22228
rect 38247 22188 38292 22216
rect 38286 22176 38292 22188
rect 38344 22176 38350 22228
rect 38654 22176 38660 22228
rect 38712 22216 38718 22228
rect 38712 22188 41460 22216
rect 38712 22176 38718 22188
rect 35161 22151 35219 22157
rect 35161 22117 35173 22151
rect 35207 22117 35219 22151
rect 35161 22111 35219 22117
rect 35253 22151 35311 22157
rect 35253 22117 35265 22151
rect 35299 22148 35311 22151
rect 35342 22148 35348 22160
rect 35299 22120 35348 22148
rect 35299 22117 35311 22120
rect 35253 22111 35311 22117
rect 35342 22108 35348 22120
rect 35400 22148 35406 22160
rect 35894 22148 35900 22160
rect 35400 22120 35900 22148
rect 35400 22108 35406 22120
rect 35894 22108 35900 22120
rect 35952 22108 35958 22160
rect 40034 22148 40040 22160
rect 39995 22120 40040 22148
rect 40034 22108 40040 22120
rect 40092 22108 40098 22160
rect 41432 22092 41460 22188
rect 43533 22151 43591 22157
rect 43533 22117 43545 22151
rect 43579 22148 43591 22151
rect 43622 22148 43628 22160
rect 43579 22120 43628 22148
rect 43579 22117 43591 22120
rect 43533 22111 43591 22117
rect 43622 22108 43628 22120
rect 43680 22108 43686 22160
rect 32252 22083 32310 22089
rect 32252 22080 32264 22083
rect 32048 22052 32264 22080
rect 31056 22043 31114 22049
rect 32252 22049 32264 22052
rect 32298 22080 32310 22083
rect 32398 22080 32404 22092
rect 32298 22052 32404 22080
rect 32298 22049 32310 22052
rect 32252 22043 32310 22049
rect 32398 22040 32404 22052
rect 32456 22040 32462 22092
rect 36630 22080 36636 22092
rect 36591 22052 36636 22080
rect 36630 22040 36636 22052
rect 36688 22080 36694 22092
rect 36998 22080 37004 22092
rect 36688 22052 37004 22080
rect 36688 22040 36694 22052
rect 36998 22040 37004 22052
rect 37056 22040 37062 22092
rect 37642 22040 37648 22092
rect 37700 22080 37706 22092
rect 37921 22083 37979 22089
rect 37921 22080 37933 22083
rect 37700 22052 37933 22080
rect 37700 22040 37706 22052
rect 37921 22049 37933 22052
rect 37967 22049 37979 22083
rect 41414 22080 41420 22092
rect 41375 22052 41420 22080
rect 37921 22043 37979 22049
rect 41414 22040 41420 22052
rect 41472 22040 41478 22092
rect 41877 22083 41935 22089
rect 41877 22049 41889 22083
rect 41923 22049 41935 22083
rect 41877 22043 41935 22049
rect 12161 22015 12219 22021
rect 12161 21981 12173 22015
rect 12207 22012 12219 22015
rect 12894 22012 12900 22024
rect 12207 21984 12900 22012
rect 12207 21981 12219 21984
rect 12161 21975 12219 21981
rect 12894 21972 12900 21984
rect 12952 21972 12958 22024
rect 14734 21972 14740 22024
rect 14792 22012 14798 22024
rect 15381 22015 15439 22021
rect 15381 22012 15393 22015
rect 14792 21984 15393 22012
rect 14792 21972 14798 21984
rect 15381 21981 15393 21984
rect 15427 22012 15439 22015
rect 16574 22012 16580 22024
rect 15427 21984 16580 22012
rect 15427 21981 15439 21984
rect 15381 21975 15439 21981
rect 16574 21972 16580 21984
rect 16632 21972 16638 22024
rect 17126 22012 17132 22024
rect 17087 21984 17132 22012
rect 17126 21972 17132 21984
rect 17184 21972 17190 22024
rect 19058 21972 19064 22024
rect 19116 22012 19122 22024
rect 21174 22012 21180 22024
rect 19116 21984 21180 22012
rect 19116 21972 19122 21984
rect 21174 21972 21180 21984
rect 21232 21972 21238 22024
rect 21542 22012 21548 22024
rect 21503 21984 21548 22012
rect 21542 21972 21548 21984
rect 21600 21972 21606 22024
rect 24118 21972 24124 22024
rect 24176 22012 24182 22024
rect 27062 22012 27068 22024
rect 24176 21984 27068 22012
rect 24176 21972 24182 21984
rect 27062 21972 27068 21984
rect 27120 21972 27126 22024
rect 27249 22015 27307 22021
rect 27249 21981 27261 22015
rect 27295 22012 27307 22015
rect 27522 22012 27528 22024
rect 27295 21984 27528 22012
rect 27295 21981 27307 21984
rect 27249 21975 27307 21981
rect 27522 21972 27528 21984
rect 27580 22012 27586 22024
rect 27706 22012 27712 22024
rect 27580 21984 27712 22012
rect 27580 21972 27586 21984
rect 27706 21972 27712 21984
rect 27764 21972 27770 22024
rect 28074 22012 28080 22024
rect 27987 21984 28080 22012
rect 28074 21972 28080 21984
rect 28132 22012 28138 22024
rect 28810 22012 28816 22024
rect 28132 21984 28816 22012
rect 28132 21972 28138 21984
rect 28810 21972 28816 21984
rect 28868 21972 28874 22024
rect 31159 22015 31217 22021
rect 31159 21981 31171 22015
rect 31205 22012 31217 22015
rect 31570 22012 31576 22024
rect 31205 21984 31576 22012
rect 31205 21981 31217 21984
rect 31159 21975 31217 21981
rect 31570 21972 31576 21984
rect 31628 21972 31634 22024
rect 33318 22012 33324 22024
rect 33279 21984 33324 22012
rect 33318 21972 33324 21984
rect 33376 21972 33382 22024
rect 33686 22012 33692 22024
rect 33647 21984 33692 22012
rect 33686 21972 33692 21984
rect 33744 21972 33750 22024
rect 35805 22015 35863 22021
rect 35805 21981 35817 22015
rect 35851 22012 35863 22015
rect 36906 22012 36912 22024
rect 35851 21984 36912 22012
rect 35851 21981 35863 21984
rect 35805 21975 35863 21981
rect 36906 21972 36912 21984
rect 36964 21972 36970 22024
rect 39942 22012 39948 22024
rect 39903 21984 39948 22012
rect 39942 21972 39948 21984
rect 40000 21972 40006 22024
rect 40589 22015 40647 22021
rect 40589 21981 40601 22015
rect 40635 22012 40647 22015
rect 41506 22012 41512 22024
rect 40635 21984 41512 22012
rect 40635 21981 40647 21984
rect 40589 21975 40647 21981
rect 41506 21972 41512 21984
rect 41564 21972 41570 22024
rect 12342 21944 12348 21956
rect 11296 21916 12348 21944
rect 11296 21904 11302 21916
rect 12342 21904 12348 21916
rect 12400 21944 12406 21956
rect 12400 21916 19012 21944
rect 12400 21904 12406 21916
rect 18984 21888 19012 21916
rect 21450 21904 21456 21956
rect 21508 21944 21514 21956
rect 23566 21944 23572 21956
rect 21508 21916 23572 21944
rect 21508 21904 21514 21916
rect 23566 21904 23572 21916
rect 23624 21904 23630 21956
rect 27614 21944 27620 21956
rect 24780 21916 27620 21944
rect 13909 21879 13967 21885
rect 13909 21845 13921 21879
rect 13955 21876 13967 21879
rect 15930 21876 15936 21888
rect 13955 21848 15936 21876
rect 13955 21845 13967 21848
rect 13909 21839 13967 21845
rect 15930 21836 15936 21848
rect 15988 21836 15994 21888
rect 18966 21836 18972 21888
rect 19024 21876 19030 21888
rect 19061 21879 19119 21885
rect 19061 21876 19073 21879
rect 19024 21848 19073 21876
rect 19024 21836 19030 21848
rect 19061 21845 19073 21848
rect 19107 21876 19119 21879
rect 19426 21876 19432 21888
rect 19107 21848 19432 21876
rect 19107 21845 19119 21848
rect 19061 21839 19119 21845
rect 19426 21836 19432 21848
rect 19484 21836 19490 21888
rect 23106 21876 23112 21888
rect 23067 21848 23112 21876
rect 23106 21836 23112 21848
rect 23164 21836 23170 21888
rect 24780 21885 24808 21916
rect 27614 21904 27620 21916
rect 27672 21904 27678 21956
rect 29546 21904 29552 21956
rect 29604 21944 29610 21956
rect 34238 21944 34244 21956
rect 29604 21916 34244 21944
rect 29604 21904 29610 21916
rect 34238 21904 34244 21916
rect 34296 21944 34302 21956
rect 34422 21944 34428 21956
rect 34296 21916 34428 21944
rect 34296 21904 34302 21916
rect 34422 21904 34428 21916
rect 34480 21904 34486 21956
rect 41892 21944 41920 22043
rect 42150 22012 42156 22024
rect 42063 21984 42156 22012
rect 42150 21972 42156 21984
rect 42208 22012 42214 22024
rect 42429 22015 42487 22021
rect 42429 22012 42441 22015
rect 42208 21984 42441 22012
rect 42208 21972 42214 21984
rect 42429 21981 42441 21984
rect 42475 21981 42487 22015
rect 43438 22012 43444 22024
rect 43399 21984 43444 22012
rect 42429 21975 42487 21981
rect 43438 21972 43444 21984
rect 43496 21972 43502 22024
rect 43717 22015 43775 22021
rect 43717 22012 43729 22015
rect 43548 21984 43729 22012
rect 42242 21944 42248 21956
rect 37108 21916 42248 21944
rect 37108 21888 37136 21916
rect 42242 21904 42248 21916
rect 42300 21904 42306 21956
rect 43254 21904 43260 21956
rect 43312 21944 43318 21956
rect 43548 21944 43576 21984
rect 43717 21981 43729 21984
rect 43763 21981 43775 22015
rect 43717 21975 43775 21981
rect 43312 21916 43576 21944
rect 43312 21904 43318 21916
rect 23477 21879 23535 21885
rect 23477 21845 23489 21879
rect 23523 21876 23535 21879
rect 24765 21879 24823 21885
rect 24765 21876 24777 21879
rect 23523 21848 24777 21876
rect 23523 21845 23535 21848
rect 23477 21839 23535 21845
rect 24765 21845 24777 21848
rect 24811 21845 24823 21879
rect 24765 21839 24823 21845
rect 32355 21879 32413 21885
rect 32355 21845 32367 21879
rect 32401 21876 32413 21879
rect 32766 21876 32772 21888
rect 32401 21848 32772 21876
rect 32401 21845 32413 21848
rect 32355 21839 32413 21845
rect 32766 21836 32772 21848
rect 32824 21836 32830 21888
rect 33042 21876 33048 21888
rect 33003 21848 33048 21876
rect 33042 21836 33048 21848
rect 33100 21836 33106 21888
rect 36771 21879 36829 21885
rect 36771 21845 36783 21879
rect 36817 21876 36829 21879
rect 36998 21876 37004 21888
rect 36817 21848 37004 21876
rect 36817 21845 36829 21848
rect 36771 21839 36829 21845
rect 36998 21836 37004 21848
rect 37056 21836 37062 21888
rect 37090 21836 37096 21888
rect 37148 21876 37154 21888
rect 38841 21879 38899 21885
rect 37148 21848 37193 21876
rect 37148 21836 37154 21848
rect 38841 21845 38853 21879
rect 38887 21876 38899 21879
rect 39022 21876 39028 21888
rect 38887 21848 39028 21876
rect 38887 21845 38899 21848
rect 38841 21839 38899 21845
rect 39022 21836 39028 21848
rect 39080 21836 39086 21888
rect 1104 21786 48852 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 48852 21786
rect 1104 21712 48852 21734
rect 11238 21672 11244 21684
rect 11199 21644 11244 21672
rect 11238 21632 11244 21644
rect 11296 21632 11302 21684
rect 11885 21675 11943 21681
rect 11885 21641 11897 21675
rect 11931 21672 11943 21675
rect 12710 21672 12716 21684
rect 11931 21644 12716 21672
rect 11931 21641 11943 21644
rect 11885 21635 11943 21641
rect 11900 21604 11928 21635
rect 12710 21632 12716 21644
rect 12768 21632 12774 21684
rect 12802 21632 12808 21684
rect 12860 21672 12866 21684
rect 12860 21644 12905 21672
rect 12860 21632 12866 21644
rect 12986 21632 12992 21684
rect 13044 21672 13050 21684
rect 14093 21675 14151 21681
rect 14093 21672 14105 21675
rect 13044 21644 14105 21672
rect 13044 21632 13050 21644
rect 14093 21641 14105 21644
rect 14139 21641 14151 21675
rect 16574 21672 16580 21684
rect 16535 21644 16580 21672
rect 14093 21635 14151 21641
rect 16574 21632 16580 21644
rect 16632 21632 16638 21684
rect 16899 21675 16957 21681
rect 16899 21641 16911 21675
rect 16945 21672 16957 21675
rect 17126 21672 17132 21684
rect 16945 21644 17132 21672
rect 16945 21641 16957 21644
rect 16899 21635 16957 21641
rect 17126 21632 17132 21644
rect 17184 21632 17190 21684
rect 17218 21632 17224 21684
rect 17276 21672 17282 21684
rect 17586 21672 17592 21684
rect 17276 21644 17592 21672
rect 17276 21632 17282 21644
rect 17586 21632 17592 21644
rect 17644 21632 17650 21684
rect 18598 21672 18604 21684
rect 18559 21644 18604 21672
rect 18598 21632 18604 21644
rect 18656 21632 18662 21684
rect 20441 21675 20499 21681
rect 20441 21641 20453 21675
rect 20487 21672 20499 21675
rect 21266 21672 21272 21684
rect 20487 21644 21272 21672
rect 20487 21641 20499 21644
rect 20441 21635 20499 21641
rect 21266 21632 21272 21644
rect 21324 21672 21330 21684
rect 21821 21675 21879 21681
rect 21821 21672 21833 21675
rect 21324 21644 21833 21672
rect 21324 21632 21330 21644
rect 21821 21641 21833 21644
rect 21867 21641 21879 21675
rect 22738 21672 22744 21684
rect 22699 21644 22744 21672
rect 21821 21635 21879 21641
rect 22738 21632 22744 21644
rect 22796 21632 22802 21684
rect 24486 21672 24492 21684
rect 24447 21644 24492 21672
rect 24486 21632 24492 21644
rect 24544 21632 24550 21684
rect 24670 21632 24676 21684
rect 24728 21672 24734 21684
rect 24857 21675 24915 21681
rect 24857 21672 24869 21675
rect 24728 21644 24869 21672
rect 24728 21632 24734 21644
rect 24857 21641 24869 21644
rect 24903 21641 24915 21675
rect 27154 21672 27160 21684
rect 27115 21644 27160 21672
rect 24857 21635 24915 21641
rect 27154 21632 27160 21644
rect 27212 21672 27218 21684
rect 27755 21675 27813 21681
rect 27755 21672 27767 21675
rect 27212 21644 27767 21672
rect 27212 21632 27218 21644
rect 27755 21641 27767 21644
rect 27801 21641 27813 21675
rect 27755 21635 27813 21641
rect 28258 21632 28264 21684
rect 28316 21672 28322 21684
rect 28629 21675 28687 21681
rect 28629 21672 28641 21675
rect 28316 21644 28641 21672
rect 28316 21632 28322 21644
rect 28629 21641 28641 21644
rect 28675 21672 28687 21675
rect 28813 21675 28871 21681
rect 28813 21672 28825 21675
rect 28675 21644 28825 21672
rect 28675 21641 28687 21644
rect 28629 21635 28687 21641
rect 28813 21641 28825 21644
rect 28859 21641 28871 21675
rect 28813 21635 28871 21641
rect 30837 21675 30895 21681
rect 30837 21641 30849 21675
rect 30883 21672 30895 21675
rect 30926 21672 30932 21684
rect 30883 21644 30932 21672
rect 30883 21641 30895 21644
rect 30837 21635 30895 21641
rect 30926 21632 30932 21644
rect 30984 21632 30990 21684
rect 31202 21632 31208 21684
rect 31260 21672 31266 21684
rect 31389 21675 31447 21681
rect 31389 21672 31401 21675
rect 31260 21644 31401 21672
rect 31260 21632 31266 21644
rect 31389 21641 31401 21644
rect 31435 21641 31447 21675
rect 31389 21635 31447 21641
rect 31849 21675 31907 21681
rect 31849 21641 31861 21675
rect 31895 21672 31907 21675
rect 32490 21672 32496 21684
rect 31895 21644 32496 21672
rect 31895 21641 31907 21644
rect 31849 21635 31907 21641
rect 32490 21632 32496 21644
rect 32548 21672 32554 21684
rect 33318 21672 33324 21684
rect 32548 21644 33324 21672
rect 32548 21632 32554 21644
rect 33318 21632 33324 21644
rect 33376 21632 33382 21684
rect 33410 21632 33416 21684
rect 33468 21672 33474 21684
rect 33965 21675 34023 21681
rect 33965 21672 33977 21675
rect 33468 21644 33977 21672
rect 33468 21632 33474 21644
rect 33965 21641 33977 21644
rect 34011 21672 34023 21675
rect 34054 21672 34060 21684
rect 34011 21644 34060 21672
rect 34011 21641 34023 21644
rect 33965 21635 34023 21641
rect 34054 21632 34060 21644
rect 34112 21632 34118 21684
rect 35894 21672 35900 21684
rect 35855 21644 35900 21672
rect 35894 21632 35900 21644
rect 35952 21632 35958 21684
rect 37642 21632 37648 21684
rect 37700 21672 37706 21684
rect 38289 21675 38347 21681
rect 38289 21672 38301 21675
rect 37700 21644 38301 21672
rect 37700 21632 37706 21644
rect 38289 21641 38301 21644
rect 38335 21641 38347 21675
rect 38289 21635 38347 21641
rect 39942 21632 39948 21684
rect 40000 21672 40006 21684
rect 40221 21675 40279 21681
rect 40221 21672 40233 21675
rect 40000 21644 40233 21672
rect 40000 21632 40006 21644
rect 40221 21641 40233 21644
rect 40267 21672 40279 21675
rect 40635 21675 40693 21681
rect 40635 21672 40647 21675
rect 40267 21644 40647 21672
rect 40267 21641 40279 21644
rect 40221 21635 40279 21641
rect 40635 21641 40647 21644
rect 40681 21641 40693 21675
rect 41414 21672 41420 21684
rect 41375 21644 41420 21672
rect 40635 21635 40693 21641
rect 41414 21632 41420 21644
rect 41472 21632 41478 21684
rect 43438 21632 43444 21684
rect 43496 21672 43502 21684
rect 44913 21675 44971 21681
rect 44913 21672 44925 21675
rect 43496 21644 44925 21672
rect 43496 21632 43502 21644
rect 44913 21641 44925 21644
rect 44959 21641 44971 21675
rect 44913 21635 44971 21641
rect 17310 21604 17316 21616
rect 11399 21576 11928 21604
rect 17271 21576 17316 21604
rect 11399 21477 11427 21576
rect 17310 21564 17316 21576
rect 17368 21564 17374 21616
rect 24213 21607 24271 21613
rect 24213 21573 24225 21607
rect 24259 21604 24271 21607
rect 26142 21604 26148 21616
rect 24259 21576 26148 21604
rect 24259 21573 24271 21576
rect 24213 21567 24271 21573
rect 11471 21539 11529 21545
rect 11471 21505 11483 21539
rect 11517 21536 11529 21539
rect 15289 21539 15347 21545
rect 15289 21536 15301 21539
rect 11517 21508 15301 21536
rect 11517 21505 11529 21508
rect 11471 21499 11529 21505
rect 15289 21505 15301 21508
rect 15335 21536 15347 21539
rect 16209 21539 16267 21545
rect 16209 21536 16221 21539
rect 15335 21508 16221 21536
rect 15335 21505 15347 21508
rect 15289 21499 15347 21505
rect 16209 21505 16221 21508
rect 16255 21505 16267 21539
rect 16209 21499 16267 21505
rect 11384 21471 11442 21477
rect 11384 21437 11396 21471
rect 11430 21437 11442 21471
rect 12894 21468 12900 21480
rect 12855 21440 12900 21468
rect 11384 21431 11442 21437
rect 12894 21428 12900 21440
rect 12952 21428 12958 21480
rect 16828 21471 16886 21477
rect 16828 21437 16840 21471
rect 16874 21468 16886 21471
rect 17328 21468 17356 21564
rect 19426 21496 19432 21548
rect 19484 21536 19490 21548
rect 19978 21536 19984 21548
rect 19484 21508 19984 21536
rect 19484 21496 19490 21508
rect 19978 21496 19984 21508
rect 20036 21496 20042 21548
rect 24118 21536 24124 21548
rect 20732 21508 24124 21536
rect 18782 21468 18788 21480
rect 16874 21440 17356 21468
rect 18743 21440 18788 21468
rect 16874 21437 16886 21440
rect 16828 21431 16886 21437
rect 18782 21428 18788 21440
rect 18840 21428 18846 21480
rect 18966 21428 18972 21480
rect 19024 21468 19030 21480
rect 19245 21471 19303 21477
rect 19245 21468 19257 21471
rect 19024 21440 19257 21468
rect 19024 21428 19030 21440
rect 19245 21437 19257 21440
rect 19291 21468 19303 21471
rect 20530 21468 20536 21480
rect 19291 21440 20536 21468
rect 19291 21437 19303 21440
rect 19245 21431 19303 21437
rect 20530 21428 20536 21440
rect 20588 21428 20594 21480
rect 12802 21360 12808 21412
rect 12860 21400 12866 21412
rect 13218 21403 13276 21409
rect 13218 21400 13230 21403
rect 12860 21372 13230 21400
rect 12860 21360 12866 21372
rect 13218 21369 13230 21372
rect 13264 21369 13276 21403
rect 14737 21403 14795 21409
rect 14737 21400 14749 21403
rect 13218 21363 13276 21369
rect 13832 21372 14749 21400
rect 11790 21292 11796 21344
rect 11848 21332 11854 21344
rect 13832 21341 13860 21372
rect 14737 21369 14749 21372
rect 14783 21400 14795 21403
rect 15105 21403 15163 21409
rect 15105 21400 15117 21403
rect 14783 21372 15117 21400
rect 14783 21369 14795 21372
rect 14737 21363 14795 21369
rect 15105 21369 15117 21372
rect 15151 21400 15163 21403
rect 15381 21403 15439 21409
rect 15381 21400 15393 21403
rect 15151 21372 15393 21400
rect 15151 21369 15163 21372
rect 15105 21363 15163 21369
rect 15381 21369 15393 21372
rect 15427 21400 15439 21403
rect 15746 21400 15752 21412
rect 15427 21372 15752 21400
rect 15427 21369 15439 21372
rect 15381 21363 15439 21369
rect 15746 21360 15752 21372
rect 15804 21360 15810 21412
rect 15933 21403 15991 21409
rect 15933 21369 15945 21403
rect 15979 21400 15991 21403
rect 16022 21400 16028 21412
rect 15979 21372 16028 21400
rect 15979 21369 15991 21372
rect 15933 21363 15991 21369
rect 16022 21360 16028 21372
rect 16080 21360 16086 21412
rect 18230 21360 18236 21412
rect 18288 21400 18294 21412
rect 19610 21400 19616 21412
rect 18288 21372 19616 21400
rect 18288 21360 18294 21372
rect 19610 21360 19616 21372
rect 19668 21400 19674 21412
rect 19705 21403 19763 21409
rect 19705 21400 19717 21403
rect 19668 21372 19717 21400
rect 19668 21360 19674 21372
rect 19705 21369 19717 21372
rect 19751 21400 19763 21403
rect 20732 21400 20760 21508
rect 24118 21496 24124 21508
rect 24176 21496 24182 21548
rect 20901 21471 20959 21477
rect 20901 21437 20913 21471
rect 20947 21468 20959 21471
rect 21358 21468 21364 21480
rect 20947 21440 21364 21468
rect 20947 21437 20959 21440
rect 20901 21431 20959 21437
rect 21358 21428 21364 21440
rect 21416 21468 21422 21480
rect 22097 21471 22155 21477
rect 22097 21468 22109 21471
rect 21416 21440 22109 21468
rect 21416 21428 21422 21440
rect 22097 21437 22109 21440
rect 22143 21437 22155 21471
rect 22097 21431 22155 21437
rect 22370 21428 22376 21480
rect 22428 21468 22434 21480
rect 23728 21471 23786 21477
rect 23728 21468 23740 21471
rect 22428 21440 23740 21468
rect 22428 21428 22434 21440
rect 23728 21437 23740 21440
rect 23774 21468 23786 21471
rect 24228 21468 24256 21567
rect 26142 21564 26148 21576
rect 26200 21564 26206 21616
rect 27522 21564 27528 21616
rect 27580 21604 27586 21616
rect 27890 21604 27896 21616
rect 27580 21576 27896 21604
rect 27580 21564 27586 21576
rect 27890 21564 27896 21576
rect 27948 21564 27954 21616
rect 32079 21607 32137 21613
rect 32079 21573 32091 21607
rect 32125 21604 32137 21607
rect 32125 21576 35020 21604
rect 32125 21573 32137 21576
rect 32079 21567 32137 21573
rect 34992 21548 35020 21576
rect 40494 21564 40500 21616
rect 40552 21604 40558 21616
rect 41230 21604 41236 21616
rect 40552 21576 41236 21604
rect 40552 21564 40558 21576
rect 41230 21564 41236 21576
rect 41288 21604 41294 21616
rect 41969 21607 42027 21613
rect 41969 21604 41981 21607
rect 41288 21576 41981 21604
rect 41288 21564 41294 21576
rect 41969 21573 41981 21576
rect 42015 21573 42027 21607
rect 41969 21567 42027 21573
rect 27706 21496 27712 21548
rect 27764 21536 27770 21548
rect 27985 21539 28043 21545
rect 27985 21536 27997 21539
rect 27764 21508 27997 21536
rect 27764 21496 27770 21508
rect 27985 21505 27997 21508
rect 28031 21505 28043 21539
rect 27985 21499 28043 21505
rect 28353 21539 28411 21545
rect 28353 21505 28365 21539
rect 28399 21536 28411 21539
rect 30650 21536 30656 21548
rect 28399 21508 30656 21536
rect 28399 21505 28411 21508
rect 28353 21499 28411 21505
rect 30650 21496 30656 21508
rect 30708 21496 30714 21548
rect 32398 21536 32404 21548
rect 32359 21508 32404 21536
rect 32398 21496 32404 21508
rect 32456 21496 32462 21548
rect 32766 21496 32772 21548
rect 32824 21536 32830 21548
rect 33045 21539 33103 21545
rect 33045 21536 33057 21539
rect 32824 21508 33057 21536
rect 32824 21496 32830 21508
rect 33045 21505 33057 21508
rect 33091 21505 33103 21539
rect 33686 21536 33692 21548
rect 33647 21508 33692 21536
rect 33045 21499 33103 21505
rect 33686 21496 33692 21508
rect 33744 21496 33750 21548
rect 34974 21536 34980 21548
rect 34887 21508 34980 21536
rect 34974 21496 34980 21508
rect 35032 21496 35038 21548
rect 35250 21536 35256 21548
rect 35211 21508 35256 21536
rect 35250 21496 35256 21508
rect 35308 21496 35314 21548
rect 36909 21539 36967 21545
rect 36909 21505 36921 21539
rect 36955 21536 36967 21539
rect 37182 21536 37188 21548
rect 36955 21508 37188 21536
rect 36955 21505 36967 21508
rect 36909 21499 36967 21505
rect 37182 21496 37188 21508
rect 37240 21496 37246 21548
rect 37274 21496 37280 21548
rect 37332 21536 37338 21548
rect 39945 21539 40003 21545
rect 37332 21508 37377 21536
rect 37332 21496 37338 21508
rect 39945 21505 39957 21539
rect 39991 21536 40003 21539
rect 40034 21536 40040 21548
rect 39991 21508 40040 21536
rect 39991 21505 40003 21508
rect 39945 21499 40003 21505
rect 40034 21496 40040 21508
rect 40092 21496 40098 21548
rect 23774 21440 24256 21468
rect 25409 21471 25467 21477
rect 23774 21437 23786 21440
rect 23728 21431 23786 21437
rect 25409 21437 25421 21471
rect 25455 21468 25467 21471
rect 26142 21468 26148 21480
rect 25455 21440 26148 21468
rect 25455 21437 25467 21440
rect 25409 21431 25467 21437
rect 26142 21428 26148 21440
rect 26200 21428 26206 21480
rect 27614 21468 27620 21480
rect 27575 21440 27620 21468
rect 27614 21428 27620 21440
rect 27672 21428 27678 21480
rect 29089 21471 29147 21477
rect 29089 21437 29101 21471
rect 29135 21468 29147 21471
rect 29546 21468 29552 21480
rect 29135 21440 29552 21468
rect 29135 21437 29147 21440
rect 29089 21431 29147 21437
rect 29546 21428 29552 21440
rect 29604 21428 29610 21480
rect 29730 21468 29736 21480
rect 29691 21440 29736 21468
rect 29730 21428 29736 21440
rect 29788 21428 29794 21480
rect 30996 21471 31054 21477
rect 30996 21437 31008 21471
rect 31042 21468 31054 21471
rect 31202 21468 31208 21480
rect 31042 21440 31208 21468
rect 31042 21437 31054 21440
rect 30996 21431 31054 21437
rect 31202 21428 31208 21440
rect 31260 21428 31266 21480
rect 31478 21428 31484 21480
rect 31536 21468 31542 21480
rect 31976 21471 32034 21477
rect 31976 21468 31988 21471
rect 31536 21440 31988 21468
rect 31536 21428 31542 21440
rect 31976 21437 31988 21440
rect 32022 21468 32034 21471
rect 32858 21468 32864 21480
rect 32022 21440 32864 21468
rect 32022 21437 32034 21440
rect 31976 21431 32034 21437
rect 32858 21428 32864 21440
rect 32916 21428 32922 21480
rect 40310 21428 40316 21480
rect 40368 21468 40374 21480
rect 40532 21471 40590 21477
rect 40532 21468 40544 21471
rect 40368 21440 40544 21468
rect 40368 21428 40374 21440
rect 40532 21437 40544 21440
rect 40578 21468 40590 21471
rect 40957 21471 41015 21477
rect 40957 21468 40969 21471
rect 40578 21440 40969 21468
rect 40578 21437 40590 21440
rect 40532 21431 40590 21437
rect 40957 21437 40969 21440
rect 41003 21437 41015 21471
rect 40957 21431 41015 21437
rect 19751 21372 20760 21400
rect 21222 21403 21280 21409
rect 19751 21369 19763 21372
rect 19705 21363 19763 21369
rect 21222 21369 21234 21403
rect 21268 21369 21280 21403
rect 26234 21400 26240 21412
rect 26195 21372 26240 21400
rect 21222 21363 21280 21369
rect 12161 21335 12219 21341
rect 12161 21332 12173 21335
rect 11848 21304 12173 21332
rect 11848 21292 11854 21304
rect 12161 21301 12173 21304
rect 12207 21301 12219 21335
rect 12161 21295 12219 21301
rect 13817 21335 13875 21341
rect 13817 21301 13829 21335
rect 13863 21301 13875 21335
rect 13817 21295 13875 21301
rect 18138 21292 18144 21344
rect 18196 21332 18202 21344
rect 18506 21332 18512 21344
rect 18196 21304 18512 21332
rect 18196 21292 18202 21304
rect 18506 21292 18512 21304
rect 18564 21292 18570 21344
rect 18966 21332 18972 21344
rect 18927 21304 18972 21332
rect 18966 21292 18972 21304
rect 19024 21292 19030 21344
rect 20714 21332 20720 21344
rect 20675 21304 20720 21332
rect 20714 21292 20720 21304
rect 20772 21332 20778 21344
rect 21237 21332 21265 21363
rect 26234 21360 26240 21372
rect 26292 21360 26298 21412
rect 30006 21400 30012 21412
rect 29967 21372 30012 21400
rect 30006 21360 30012 21372
rect 30064 21360 30070 21412
rect 33137 21403 33195 21409
rect 33137 21369 33149 21403
rect 33183 21400 33195 21403
rect 35069 21403 35127 21409
rect 33183 21372 33217 21400
rect 33796 21372 34744 21400
rect 33183 21369 33195 21372
rect 33137 21363 33195 21369
rect 20772 21304 21265 21332
rect 20772 21292 20778 21304
rect 23566 21292 23572 21344
rect 23624 21332 23630 21344
rect 23799 21335 23857 21341
rect 23799 21332 23811 21335
rect 23624 21304 23811 21332
rect 23624 21292 23630 21304
rect 23799 21301 23811 21304
rect 23845 21301 23857 21335
rect 23799 21295 23857 21301
rect 26605 21335 26663 21341
rect 26605 21301 26617 21335
rect 26651 21332 26663 21335
rect 26970 21332 26976 21344
rect 26651 21304 26976 21332
rect 26651 21301 26663 21304
rect 26605 21295 26663 21301
rect 26970 21292 26976 21304
rect 27028 21292 27034 21344
rect 27522 21332 27528 21344
rect 27483 21304 27528 21332
rect 27522 21292 27528 21304
rect 27580 21292 27586 21344
rect 28813 21335 28871 21341
rect 28813 21301 28825 21335
rect 28859 21332 28871 21335
rect 29822 21332 29828 21344
rect 28859 21304 29828 21332
rect 28859 21301 28871 21304
rect 28813 21295 28871 21301
rect 29822 21292 29828 21304
rect 29880 21292 29886 21344
rect 31067 21335 31125 21341
rect 31067 21301 31079 21335
rect 31113 21332 31125 21335
rect 32122 21332 32128 21344
rect 31113 21304 32128 21332
rect 31113 21301 31125 21304
rect 31067 21295 31125 21301
rect 32122 21292 32128 21304
rect 32180 21292 32186 21344
rect 32950 21292 32956 21344
rect 33008 21332 33014 21344
rect 33152 21332 33180 21363
rect 33796 21332 33824 21372
rect 34716 21341 34744 21372
rect 35069 21369 35081 21403
rect 35115 21369 35127 21403
rect 35069 21363 35127 21369
rect 33008 21304 33824 21332
rect 34701 21335 34759 21341
rect 33008 21292 33014 21304
rect 34701 21301 34713 21335
rect 34747 21332 34759 21335
rect 35084 21332 35112 21363
rect 36906 21360 36912 21412
rect 36964 21400 36970 21412
rect 37001 21403 37059 21409
rect 37001 21400 37013 21403
rect 36964 21372 37013 21400
rect 36964 21360 36970 21372
rect 37001 21369 37013 21372
rect 37047 21369 37059 21403
rect 38930 21400 38936 21412
rect 38891 21372 38936 21400
rect 37001 21363 37059 21369
rect 38930 21360 38936 21372
rect 38988 21360 38994 21412
rect 39022 21360 39028 21412
rect 39080 21400 39086 21412
rect 39574 21400 39580 21412
rect 39080 21372 39125 21400
rect 39535 21372 39580 21400
rect 39080 21360 39086 21372
rect 39574 21360 39580 21372
rect 39632 21360 39638 21412
rect 34747 21304 35112 21332
rect 36357 21335 36415 21341
rect 34747 21301 34759 21304
rect 34701 21295 34759 21301
rect 36357 21301 36369 21335
rect 36403 21332 36415 21335
rect 36446 21332 36452 21344
rect 36403 21304 36452 21332
rect 36403 21301 36415 21304
rect 36357 21295 36415 21301
rect 36446 21292 36452 21304
rect 36504 21292 36510 21344
rect 36630 21332 36636 21344
rect 36591 21304 36636 21332
rect 36630 21292 36636 21304
rect 36688 21292 36694 21344
rect 36814 21292 36820 21344
rect 36872 21332 36878 21344
rect 37921 21335 37979 21341
rect 37921 21332 37933 21335
rect 36872 21304 37933 21332
rect 36872 21292 36878 21304
rect 37921 21301 37933 21304
rect 37967 21332 37979 21335
rect 38286 21332 38292 21344
rect 37967 21304 38292 21332
rect 37967 21301 37979 21304
rect 37921 21295 37979 21301
rect 38286 21292 38292 21304
rect 38344 21292 38350 21344
rect 38749 21335 38807 21341
rect 38749 21301 38761 21335
rect 38795 21332 38807 21335
rect 39040 21332 39068 21360
rect 38795 21304 39068 21332
rect 40972 21332 41000 21431
rect 41984 21400 42012 21567
rect 42150 21536 42156 21548
rect 42111 21508 42156 21536
rect 42150 21496 42156 21508
rect 42208 21496 42214 21548
rect 43714 21496 43720 21548
rect 43772 21536 43778 21548
rect 43993 21539 44051 21545
rect 43993 21536 44005 21539
rect 43772 21508 44005 21536
rect 43772 21496 43778 21508
rect 43993 21505 44005 21508
rect 44039 21505 44051 21539
rect 43993 21499 44051 21505
rect 44174 21496 44180 21548
rect 44232 21536 44238 21548
rect 44269 21539 44327 21545
rect 44269 21536 44281 21539
rect 44232 21508 44281 21536
rect 44232 21496 44238 21508
rect 44269 21505 44281 21508
rect 44315 21505 44327 21539
rect 44269 21499 44327 21505
rect 42474 21403 42532 21409
rect 42474 21400 42486 21403
rect 41984 21372 42486 21400
rect 42474 21369 42486 21372
rect 42520 21369 42532 21403
rect 44085 21403 44143 21409
rect 44085 21400 44097 21403
rect 42474 21363 42532 21369
rect 43732 21372 44097 21400
rect 42978 21332 42984 21344
rect 40972 21304 42984 21332
rect 38795 21301 38807 21304
rect 38749 21295 38807 21301
rect 42978 21292 42984 21304
rect 43036 21292 43042 21344
rect 43073 21335 43131 21341
rect 43073 21301 43085 21335
rect 43119 21332 43131 21335
rect 43441 21335 43499 21341
rect 43441 21332 43453 21335
rect 43119 21304 43453 21332
rect 43119 21301 43131 21304
rect 43073 21295 43131 21301
rect 43441 21301 43453 21304
rect 43487 21332 43499 21335
rect 43622 21332 43628 21344
rect 43487 21304 43628 21332
rect 43487 21301 43499 21304
rect 43441 21295 43499 21301
rect 43622 21292 43628 21304
rect 43680 21332 43686 21344
rect 43732 21341 43760 21372
rect 44085 21369 44097 21372
rect 44131 21369 44143 21403
rect 44085 21363 44143 21369
rect 43717 21335 43775 21341
rect 43717 21332 43729 21335
rect 43680 21304 43729 21332
rect 43680 21292 43686 21304
rect 43717 21301 43729 21304
rect 43763 21301 43775 21335
rect 43717 21295 43775 21301
rect 1104 21242 48852 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 48852 21242
rect 1104 21168 48852 21190
rect 12894 21088 12900 21140
rect 12952 21128 12958 21140
rect 13725 21131 13783 21137
rect 13725 21128 13737 21131
rect 12952 21100 13737 21128
rect 12952 21088 12958 21100
rect 13725 21097 13737 21100
rect 13771 21097 13783 21131
rect 17126 21128 17132 21140
rect 17087 21100 17132 21128
rect 13725 21091 13783 21097
rect 17126 21088 17132 21100
rect 17184 21088 17190 21140
rect 19981 21131 20039 21137
rect 19981 21097 19993 21131
rect 20027 21128 20039 21131
rect 20027 21100 21128 21128
rect 20027 21097 20039 21100
rect 19981 21091 20039 21097
rect 21100 21072 21128 21100
rect 21174 21088 21180 21140
rect 21232 21128 21238 21140
rect 21913 21131 21971 21137
rect 21913 21128 21925 21131
rect 21232 21100 21925 21128
rect 21232 21088 21238 21100
rect 21913 21097 21925 21100
rect 21959 21097 21971 21131
rect 21913 21091 21971 21097
rect 26142 21088 26148 21140
rect 26200 21128 26206 21140
rect 26651 21131 26709 21137
rect 26651 21128 26663 21131
rect 26200 21100 26663 21128
rect 26200 21088 26206 21100
rect 26651 21097 26663 21100
rect 26697 21097 26709 21131
rect 26651 21091 26709 21097
rect 27154 21088 27160 21140
rect 27212 21128 27218 21140
rect 27249 21131 27307 21137
rect 27249 21128 27261 21131
rect 27212 21100 27261 21128
rect 27212 21088 27218 21100
rect 27249 21097 27261 21100
rect 27295 21097 27307 21131
rect 28810 21128 28816 21140
rect 28771 21100 28816 21128
rect 27249 21091 27307 21097
rect 11606 21020 11612 21072
rect 11664 21060 11670 21072
rect 12158 21060 12164 21072
rect 11664 21032 12164 21060
rect 11664 21020 11670 21032
rect 12158 21020 12164 21032
rect 12216 21060 12222 21072
rect 12216 21032 12756 21060
rect 12216 21020 12222 21032
rect 10594 20992 10600 21004
rect 10555 20964 10600 20992
rect 10594 20952 10600 20964
rect 10652 20952 10658 21004
rect 12304 20995 12362 21001
rect 12304 20961 12316 20995
rect 12350 20992 12362 20995
rect 12526 20992 12532 21004
rect 12350 20964 12532 20992
rect 12350 20961 12362 20964
rect 12304 20955 12362 20961
rect 12526 20952 12532 20964
rect 12584 20952 12590 21004
rect 12728 20992 12756 21032
rect 12802 21020 12808 21072
rect 12860 21060 12866 21072
rect 12989 21063 13047 21069
rect 12989 21060 13001 21063
rect 12860 21032 13001 21060
rect 12860 21020 12866 21032
rect 12989 21029 13001 21032
rect 13035 21029 13047 21063
rect 12989 21023 13047 21029
rect 15657 21063 15715 21069
rect 15657 21029 15669 21063
rect 15703 21060 15715 21063
rect 15838 21060 15844 21072
rect 15703 21032 15844 21060
rect 15703 21029 15715 21032
rect 15657 21023 15715 21029
rect 15838 21020 15844 21032
rect 15896 21020 15902 21072
rect 17586 21060 17592 21072
rect 17547 21032 17592 21060
rect 17586 21020 17592 21032
rect 17644 21020 17650 21072
rect 19150 21020 19156 21072
rect 19208 21060 19214 21072
rect 19382 21063 19440 21069
rect 19382 21060 19394 21063
rect 19208 21032 19394 21060
rect 19208 21020 19214 21032
rect 19382 21029 19394 21032
rect 19428 21060 19440 21063
rect 20714 21060 20720 21072
rect 19428 21032 20720 21060
rect 19428 21029 19440 21032
rect 19382 21023 19440 21029
rect 20714 21020 20720 21032
rect 20772 21020 20778 21072
rect 21082 21060 21088 21072
rect 20995 21032 21088 21060
rect 21082 21020 21088 21032
rect 21140 21020 21146 21072
rect 24762 21060 24768 21072
rect 24723 21032 24768 21060
rect 24762 21020 24768 21032
rect 24820 21020 24826 21072
rect 27264 21060 27292 21091
rect 28810 21088 28816 21100
rect 28868 21088 28874 21140
rect 32398 21088 32404 21140
rect 32456 21128 32462 21140
rect 32493 21131 32551 21137
rect 32493 21128 32505 21131
rect 32456 21100 32505 21128
rect 32456 21088 32462 21100
rect 32493 21097 32505 21100
rect 32539 21128 32551 21131
rect 32582 21128 32588 21140
rect 32539 21100 32588 21128
rect 32539 21097 32551 21100
rect 32493 21091 32551 21097
rect 32582 21088 32588 21100
rect 32640 21088 32646 21140
rect 32766 21088 32772 21140
rect 32824 21128 32830 21140
rect 33321 21131 33379 21137
rect 33321 21128 33333 21131
rect 32824 21100 33333 21128
rect 32824 21088 32830 21100
rect 33321 21097 33333 21100
rect 33367 21097 33379 21131
rect 34974 21128 34980 21140
rect 34935 21100 34980 21128
rect 33321 21091 33379 21097
rect 34974 21088 34980 21100
rect 35032 21088 35038 21140
rect 35345 21131 35403 21137
rect 35345 21097 35357 21131
rect 35391 21128 35403 21131
rect 35802 21128 35808 21140
rect 35391 21100 35808 21128
rect 35391 21097 35403 21100
rect 35345 21091 35403 21097
rect 35802 21088 35808 21100
rect 35860 21088 35866 21140
rect 38427 21131 38485 21137
rect 38427 21097 38439 21131
rect 38473 21128 38485 21131
rect 38930 21128 38936 21140
rect 38473 21100 38936 21128
rect 38473 21097 38485 21100
rect 38427 21091 38485 21097
rect 38930 21088 38936 21100
rect 38988 21088 38994 21140
rect 42242 21128 42248 21140
rect 42203 21100 42248 21128
rect 42242 21088 42248 21100
rect 42300 21088 42306 21140
rect 43714 21088 43720 21140
rect 43772 21128 43778 21140
rect 44361 21131 44419 21137
rect 44361 21128 44373 21131
rect 43772 21100 44373 21128
rect 43772 21088 43778 21100
rect 44361 21097 44373 21100
rect 44407 21097 44419 21131
rect 44361 21091 44419 21097
rect 28537 21063 28595 21069
rect 27264 21032 27991 21060
rect 13300 20995 13358 21001
rect 13300 20992 13312 20995
rect 12728 20964 13312 20992
rect 13300 20961 13312 20964
rect 13346 20992 13358 20995
rect 13998 20992 14004 21004
rect 13346 20964 14004 20992
rect 13346 20961 13358 20964
rect 13300 20955 13358 20961
rect 13998 20952 14004 20964
rect 14056 20952 14062 21004
rect 18966 20952 18972 21004
rect 19024 20992 19030 21004
rect 19061 20995 19119 21001
rect 19061 20992 19073 20995
rect 19024 20964 19073 20992
rect 19024 20952 19030 20964
rect 19061 20961 19073 20964
rect 19107 20961 19119 20995
rect 23566 20992 23572 21004
rect 23527 20964 23572 20992
rect 19061 20955 19119 20961
rect 23566 20952 23572 20964
rect 23624 20952 23630 21004
rect 26326 20952 26332 21004
rect 26384 20992 26390 21004
rect 26548 20995 26606 21001
rect 26548 20992 26560 20995
rect 26384 20964 26560 20992
rect 26384 20952 26390 20964
rect 26548 20961 26560 20964
rect 26594 20961 26606 20995
rect 26548 20955 26606 20961
rect 27614 20952 27620 21004
rect 27672 20992 27678 21004
rect 27963 21001 27991 21032
rect 28537 21029 28549 21063
rect 28583 21060 28595 21063
rect 29273 21063 29331 21069
rect 29273 21060 29285 21063
rect 28583 21032 29285 21060
rect 28583 21029 28595 21032
rect 28537 21023 28595 21029
rect 29273 21029 29285 21032
rect 29319 21060 29331 21063
rect 29730 21060 29736 21072
rect 29319 21032 29736 21060
rect 29319 21029 29331 21032
rect 29273 21023 29331 21029
rect 29730 21020 29736 21032
rect 29788 21060 29794 21072
rect 34054 21060 34060 21072
rect 29788 21032 30972 21060
rect 34015 21032 34060 21060
rect 29788 21020 29794 21032
rect 30944 21004 30972 21032
rect 34054 21020 34060 21032
rect 34112 21020 34118 21072
rect 34238 21020 34244 21072
rect 34296 21060 34302 21072
rect 34609 21063 34667 21069
rect 34609 21060 34621 21063
rect 34296 21032 34621 21060
rect 34296 21020 34302 21032
rect 34609 21029 34621 21032
rect 34655 21060 34667 21063
rect 35250 21060 35256 21072
rect 34655 21032 35256 21060
rect 34655 21029 34667 21032
rect 34609 21023 34667 21029
rect 35250 21020 35256 21032
rect 35308 21020 35314 21072
rect 36446 21060 36452 21072
rect 36407 21032 36452 21060
rect 36446 21020 36452 21032
rect 36504 21020 36510 21072
rect 39022 21020 39028 21072
rect 39080 21060 39086 21072
rect 39485 21063 39543 21069
rect 39485 21060 39497 21063
rect 39080 21032 39497 21060
rect 39080 21020 39086 21032
rect 39485 21029 39497 21032
rect 39531 21060 39543 21063
rect 40034 21060 40040 21072
rect 39531 21032 40040 21060
rect 39531 21029 39543 21032
rect 39485 21023 39543 21029
rect 40034 21020 40040 21032
rect 40092 21020 40098 21072
rect 41417 21063 41475 21069
rect 41417 21029 41429 21063
rect 41463 21060 41475 21063
rect 41598 21060 41604 21072
rect 41463 21032 41604 21060
rect 41463 21029 41475 21032
rect 41417 21023 41475 21029
rect 41598 21020 41604 21032
rect 41656 21020 41662 21072
rect 43533 21063 43591 21069
rect 43533 21029 43545 21063
rect 43579 21060 43591 21063
rect 43622 21060 43628 21072
rect 43579 21032 43628 21060
rect 43579 21029 43591 21032
rect 43533 21023 43591 21029
rect 43622 21020 43628 21032
rect 43680 21020 43686 21072
rect 27801 20995 27859 21001
rect 27801 20992 27813 20995
rect 27672 20964 27813 20992
rect 27672 20952 27678 20964
rect 27801 20961 27813 20964
rect 27847 20961 27859 20995
rect 27801 20955 27859 20961
rect 27948 20995 28006 21001
rect 27948 20961 27960 20995
rect 27994 20992 28006 20995
rect 28258 20992 28264 21004
rect 27994 20964 28264 20992
rect 27994 20961 28006 20964
rect 27948 20955 28006 20961
rect 28258 20952 28264 20964
rect 28316 20952 28322 21004
rect 29086 20952 29092 21004
rect 29144 20992 29150 21004
rect 29524 20995 29582 21001
rect 29524 20992 29536 20995
rect 29144 20964 29536 20992
rect 29144 20952 29150 20964
rect 29524 20961 29536 20964
rect 29570 20992 29582 20995
rect 30098 20992 30104 21004
rect 29570 20964 30104 20992
rect 29570 20961 29582 20964
rect 29524 20955 29582 20961
rect 30098 20952 30104 20964
rect 30156 20952 30162 21004
rect 30469 20995 30527 21001
rect 30469 20961 30481 20995
rect 30515 20961 30527 20995
rect 30926 20992 30932 21004
rect 30839 20964 30932 20992
rect 30469 20955 30527 20961
rect 12391 20927 12449 20933
rect 12391 20893 12403 20927
rect 12437 20924 12449 20927
rect 15194 20924 15200 20936
rect 12437 20896 15200 20924
rect 12437 20893 12449 20896
rect 12391 20887 12449 20893
rect 15194 20884 15200 20896
rect 15252 20884 15258 20936
rect 15565 20927 15623 20933
rect 15565 20893 15577 20927
rect 15611 20924 15623 20927
rect 16942 20924 16948 20936
rect 15611 20896 16948 20924
rect 15611 20893 15623 20896
rect 15565 20887 15623 20893
rect 16942 20884 16948 20896
rect 17000 20884 17006 20936
rect 17494 20924 17500 20936
rect 17455 20896 17500 20924
rect 17494 20884 17500 20896
rect 17552 20884 17558 20936
rect 18141 20927 18199 20933
rect 18141 20893 18153 20927
rect 18187 20924 18199 20927
rect 20993 20927 21051 20933
rect 20993 20924 21005 20927
rect 18187 20896 21005 20924
rect 18187 20893 18199 20896
rect 18141 20887 18199 20893
rect 20993 20893 21005 20896
rect 21039 20924 21051 20927
rect 21910 20924 21916 20936
rect 21039 20896 21916 20924
rect 21039 20893 21051 20896
rect 20993 20887 21051 20893
rect 12802 20816 12808 20868
rect 12860 20856 12866 20868
rect 13403 20859 13461 20865
rect 13403 20856 13415 20859
rect 12860 20828 13415 20856
rect 12860 20816 12866 20828
rect 13403 20825 13415 20828
rect 13449 20825 13461 20859
rect 13403 20819 13461 20825
rect 16117 20859 16175 20865
rect 16117 20825 16129 20859
rect 16163 20856 16175 20859
rect 16206 20856 16212 20868
rect 16163 20828 16212 20856
rect 16163 20825 16175 20828
rect 16117 20819 16175 20825
rect 16206 20816 16212 20828
rect 16264 20856 16270 20868
rect 18156 20856 18184 20887
rect 21910 20884 21916 20896
rect 21968 20884 21974 20936
rect 24394 20884 24400 20936
rect 24452 20924 24458 20936
rect 24673 20927 24731 20933
rect 24673 20924 24685 20927
rect 24452 20896 24685 20924
rect 24452 20884 24458 20896
rect 24673 20893 24685 20896
rect 24719 20893 24731 20927
rect 24673 20887 24731 20893
rect 25317 20927 25375 20933
rect 25317 20893 25329 20927
rect 25363 20924 25375 20927
rect 26878 20924 26884 20936
rect 25363 20896 26884 20924
rect 25363 20893 25375 20896
rect 25317 20887 25375 20893
rect 21542 20856 21548 20868
rect 16264 20828 18184 20856
rect 21503 20828 21548 20856
rect 16264 20816 16270 20828
rect 21542 20816 21548 20828
rect 21600 20816 21606 20868
rect 23290 20816 23296 20868
rect 23348 20856 23354 20868
rect 25332 20856 25360 20887
rect 26878 20884 26884 20896
rect 26936 20884 26942 20936
rect 26970 20884 26976 20936
rect 27028 20924 27034 20936
rect 28169 20927 28227 20933
rect 28169 20924 28181 20927
rect 27028 20896 28181 20924
rect 27028 20884 27034 20896
rect 28169 20893 28181 20896
rect 28215 20924 28227 20927
rect 28626 20924 28632 20936
rect 28215 20896 28632 20924
rect 28215 20893 28227 20896
rect 28169 20887 28227 20893
rect 28626 20884 28632 20896
rect 28684 20884 28690 20936
rect 23348 20828 25360 20856
rect 23348 20816 23354 20828
rect 27430 20816 27436 20868
rect 27488 20856 27494 20868
rect 30478 20856 30506 20955
rect 30926 20952 30932 20964
rect 30984 20952 30990 21004
rect 33042 20992 33048 21004
rect 33003 20964 33048 20992
rect 33042 20952 33048 20964
rect 33100 20952 33106 21004
rect 35710 20992 35716 21004
rect 35671 20964 35716 20992
rect 35710 20952 35716 20964
rect 35768 20952 35774 21004
rect 36170 20992 36176 21004
rect 36131 20964 36176 20992
rect 36170 20952 36176 20964
rect 36228 20952 36234 21004
rect 38356 20995 38414 21001
rect 38356 20961 38368 20995
rect 38402 20992 38414 20995
rect 38838 20992 38844 21004
rect 38402 20964 38844 20992
rect 38402 20961 38414 20964
rect 38356 20955 38414 20961
rect 38838 20952 38844 20964
rect 38896 20952 38902 21004
rect 31205 20927 31263 20933
rect 31205 20893 31217 20927
rect 31251 20924 31263 20927
rect 32030 20924 32036 20936
rect 31251 20896 32036 20924
rect 31251 20893 31263 20896
rect 31205 20887 31263 20893
rect 32030 20884 32036 20896
rect 32088 20924 32094 20936
rect 32125 20927 32183 20933
rect 32125 20924 32137 20927
rect 32088 20896 32137 20924
rect 32088 20884 32094 20896
rect 32125 20893 32137 20896
rect 32171 20893 32183 20927
rect 32125 20887 32183 20893
rect 33965 20927 34023 20933
rect 33965 20893 33977 20927
rect 34011 20924 34023 20927
rect 34606 20924 34612 20936
rect 34011 20896 34612 20924
rect 34011 20893 34023 20896
rect 33965 20887 34023 20893
rect 34606 20884 34612 20896
rect 34664 20884 34670 20936
rect 36998 20884 37004 20936
rect 37056 20924 37062 20936
rect 39393 20927 39451 20933
rect 39393 20924 39405 20927
rect 37056 20896 39405 20924
rect 37056 20884 37062 20896
rect 39393 20893 39405 20896
rect 39439 20924 39451 20927
rect 39666 20924 39672 20936
rect 39439 20896 39672 20924
rect 39439 20893 39451 20896
rect 39393 20887 39451 20893
rect 39666 20884 39672 20896
rect 39724 20884 39730 20936
rect 40034 20924 40040 20936
rect 39995 20896 40040 20924
rect 40034 20884 40040 20896
rect 40092 20884 40098 20936
rect 41138 20884 41144 20936
rect 41196 20924 41202 20936
rect 41325 20927 41383 20933
rect 41325 20924 41337 20927
rect 41196 20896 41337 20924
rect 41196 20884 41202 20896
rect 41325 20893 41337 20896
rect 41371 20893 41383 20927
rect 41325 20887 41383 20893
rect 41506 20884 41512 20936
rect 41564 20924 41570 20936
rect 41601 20927 41659 20933
rect 41601 20924 41613 20927
rect 41564 20896 41613 20924
rect 41564 20884 41570 20896
rect 41601 20893 41613 20896
rect 41647 20924 41659 20927
rect 43254 20924 43260 20936
rect 41647 20896 43260 20924
rect 41647 20893 41659 20896
rect 41601 20887 41659 20893
rect 43254 20884 43260 20896
rect 43312 20884 43318 20936
rect 43438 20924 43444 20936
rect 43399 20896 43444 20924
rect 43438 20884 43444 20896
rect 43496 20884 43502 20936
rect 43717 20927 43775 20933
rect 43717 20924 43729 20927
rect 43548 20896 43729 20924
rect 31110 20856 31116 20868
rect 27488 20828 31116 20856
rect 27488 20816 27494 20828
rect 31110 20816 31116 20828
rect 31168 20816 31174 20868
rect 41230 20816 41236 20868
rect 41288 20856 41294 20868
rect 41524 20856 41552 20884
rect 41288 20828 41552 20856
rect 41288 20816 41294 20828
rect 41966 20816 41972 20868
rect 42024 20856 42030 20868
rect 43548 20856 43576 20896
rect 43717 20893 43729 20896
rect 43763 20893 43775 20927
rect 43717 20887 43775 20893
rect 42024 20828 43576 20856
rect 42024 20816 42030 20828
rect 10962 20788 10968 20800
rect 10923 20760 10968 20788
rect 10962 20748 10968 20760
rect 11020 20748 11026 20800
rect 16390 20748 16396 20800
rect 16448 20788 16454 20800
rect 18693 20791 18751 20797
rect 18693 20788 18705 20791
rect 16448 20760 18705 20788
rect 16448 20748 16454 20760
rect 18693 20757 18705 20760
rect 18739 20788 18751 20791
rect 18782 20788 18788 20800
rect 18739 20760 18788 20788
rect 18739 20757 18751 20760
rect 18693 20751 18751 20757
rect 18782 20748 18788 20760
rect 18840 20748 18846 20800
rect 23382 20788 23388 20800
rect 23343 20760 23388 20788
rect 23382 20748 23388 20760
rect 23440 20748 23446 20800
rect 23750 20748 23756 20800
rect 23808 20788 23814 20800
rect 23937 20791 23995 20797
rect 23937 20788 23949 20791
rect 23808 20760 23949 20788
rect 23808 20748 23814 20760
rect 23937 20757 23949 20760
rect 23983 20757 23995 20791
rect 27706 20788 27712 20800
rect 27667 20760 27712 20788
rect 23937 20751 23995 20757
rect 27706 20748 27712 20760
rect 27764 20748 27770 20800
rect 28074 20788 28080 20800
rect 28035 20760 28080 20788
rect 28074 20748 28080 20760
rect 28132 20748 28138 20800
rect 29595 20791 29653 20797
rect 29595 20757 29607 20791
rect 29641 20788 29653 20791
rect 31478 20788 31484 20800
rect 29641 20760 31484 20788
rect 29641 20757 29653 20760
rect 29595 20751 29653 20757
rect 31478 20748 31484 20760
rect 31536 20748 31542 20800
rect 33686 20788 33692 20800
rect 33647 20760 33692 20788
rect 33686 20748 33692 20760
rect 33744 20748 33750 20800
rect 36906 20788 36912 20800
rect 36867 20760 36912 20788
rect 36906 20748 36912 20760
rect 36964 20748 36970 20800
rect 37182 20788 37188 20800
rect 37143 20760 37188 20788
rect 37182 20748 37188 20760
rect 37240 20748 37246 20800
rect 1104 20698 48852 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 48852 20698
rect 1104 20624 48852 20646
rect 10134 20584 10140 20596
rect 10095 20556 10140 20584
rect 10134 20544 10140 20556
rect 10192 20544 10198 20596
rect 12526 20544 12532 20596
rect 12584 20584 12590 20596
rect 12621 20587 12679 20593
rect 12621 20584 12633 20587
rect 12584 20556 12633 20584
rect 12584 20544 12590 20556
rect 12621 20553 12633 20556
rect 12667 20553 12679 20587
rect 13998 20584 14004 20596
rect 13959 20556 14004 20584
rect 12621 20547 12679 20553
rect 13998 20544 14004 20556
rect 14056 20544 14062 20596
rect 14826 20584 14832 20596
rect 14787 20556 14832 20584
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 16942 20584 16948 20596
rect 16903 20556 16948 20584
rect 16942 20544 16948 20556
rect 17000 20544 17006 20596
rect 17497 20587 17555 20593
rect 17497 20553 17509 20587
rect 17543 20584 17555 20587
rect 17586 20584 17592 20596
rect 17543 20556 17592 20584
rect 17543 20553 17555 20556
rect 17497 20547 17555 20553
rect 17586 20544 17592 20556
rect 17644 20584 17650 20596
rect 17773 20587 17831 20593
rect 17773 20584 17785 20587
rect 17644 20556 17785 20584
rect 17644 20544 17650 20556
rect 17773 20553 17785 20556
rect 17819 20553 17831 20587
rect 17773 20547 17831 20553
rect 10152 20448 10180 20544
rect 16206 20516 16212 20528
rect 16167 20488 16212 20516
rect 16206 20476 16212 20488
rect 16264 20476 16270 20528
rect 9727 20420 10180 20448
rect 9727 20389 9755 20420
rect 15838 20408 15844 20460
rect 15896 20448 15902 20460
rect 16577 20451 16635 20457
rect 16577 20448 16589 20451
rect 15896 20420 16589 20448
rect 15896 20408 15902 20420
rect 16577 20417 16589 20420
rect 16623 20417 16635 20451
rect 16577 20411 16635 20417
rect 9712 20383 9770 20389
rect 9712 20349 9724 20383
rect 9758 20349 9770 20383
rect 9712 20343 9770 20349
rect 9815 20383 9873 20389
rect 9815 20349 9827 20383
rect 9861 20380 9873 20383
rect 10597 20383 10655 20389
rect 10597 20380 10609 20383
rect 9861 20352 10609 20380
rect 9861 20349 9873 20352
rect 9815 20343 9873 20349
rect 10597 20349 10609 20352
rect 10643 20380 10655 20383
rect 10781 20383 10839 20389
rect 10781 20380 10793 20383
rect 10643 20352 10793 20380
rect 10643 20349 10655 20352
rect 10597 20343 10655 20349
rect 10781 20349 10793 20352
rect 10827 20349 10839 20383
rect 10781 20343 10839 20349
rect 12253 20383 12311 20389
rect 12253 20349 12265 20383
rect 12299 20380 12311 20383
rect 12618 20380 12624 20392
rect 12299 20352 12624 20380
rect 12299 20349 12311 20352
rect 12253 20343 12311 20349
rect 12618 20340 12624 20352
rect 12676 20380 12682 20392
rect 13081 20383 13139 20389
rect 13081 20380 13093 20383
rect 12676 20352 13093 20380
rect 12676 20340 12682 20352
rect 13081 20349 13093 20352
rect 13127 20349 13139 20383
rect 13081 20343 13139 20349
rect 13170 20340 13176 20392
rect 13228 20380 13234 20392
rect 14620 20383 14678 20389
rect 14620 20380 14632 20383
rect 13228 20352 14632 20380
rect 13228 20340 13234 20352
rect 14620 20349 14632 20352
rect 14666 20380 14678 20383
rect 15013 20383 15071 20389
rect 15013 20380 15025 20383
rect 14666 20352 15025 20380
rect 14666 20349 14678 20352
rect 14620 20343 14678 20349
rect 15013 20349 15025 20352
rect 15059 20349 15071 20383
rect 15013 20343 15071 20349
rect 10686 20312 10692 20324
rect 10647 20284 10692 20312
rect 10686 20272 10692 20284
rect 10744 20272 10750 20324
rect 13722 20312 13728 20324
rect 13683 20284 13728 20312
rect 13722 20272 13728 20284
rect 13780 20272 13786 20324
rect 15657 20315 15715 20321
rect 15657 20281 15669 20315
rect 15703 20281 15715 20315
rect 15657 20275 15715 20281
rect 15378 20244 15384 20256
rect 15339 20216 15384 20244
rect 15378 20204 15384 20216
rect 15436 20244 15442 20256
rect 15672 20244 15700 20275
rect 15746 20272 15752 20324
rect 15804 20312 15810 20324
rect 16298 20312 16304 20324
rect 15804 20284 16304 20312
rect 15804 20272 15810 20284
rect 16298 20272 16304 20284
rect 16356 20272 16362 20324
rect 17788 20312 17816 20547
rect 18966 20544 18972 20596
rect 19024 20584 19030 20596
rect 19429 20587 19487 20593
rect 19429 20584 19441 20587
rect 19024 20556 19441 20584
rect 19024 20544 19030 20556
rect 19429 20553 19441 20556
rect 19475 20553 19487 20587
rect 19429 20547 19487 20553
rect 21082 20544 21088 20596
rect 21140 20584 21146 20596
rect 21545 20587 21603 20593
rect 21545 20584 21557 20587
rect 21140 20556 21557 20584
rect 21140 20544 21146 20556
rect 21545 20553 21557 20556
rect 21591 20553 21603 20587
rect 21910 20584 21916 20596
rect 21871 20556 21916 20584
rect 21545 20547 21603 20553
rect 21910 20544 21916 20556
rect 21968 20544 21974 20596
rect 22235 20587 22293 20593
rect 22235 20553 22247 20587
rect 22281 20584 22293 20587
rect 22370 20584 22376 20596
rect 22281 20556 22376 20584
rect 22281 20553 22293 20556
rect 22235 20547 22293 20553
rect 22370 20544 22376 20556
rect 22428 20544 22434 20596
rect 23382 20584 23388 20596
rect 23343 20556 23388 20584
rect 23382 20544 23388 20556
rect 23440 20544 23446 20596
rect 24762 20584 24768 20596
rect 24723 20556 24768 20584
rect 24762 20544 24768 20556
rect 24820 20584 24826 20596
rect 25498 20584 25504 20596
rect 24820 20556 25504 20584
rect 24820 20544 24826 20556
rect 25498 20544 25504 20556
rect 25556 20584 25562 20596
rect 25685 20587 25743 20593
rect 25685 20584 25697 20587
rect 25556 20556 25697 20584
rect 25556 20544 25562 20556
rect 25685 20553 25697 20556
rect 25731 20553 25743 20587
rect 25685 20547 25743 20553
rect 27782 20587 27840 20593
rect 27782 20553 27794 20587
rect 27828 20584 27840 20587
rect 28258 20584 28264 20596
rect 27828 20556 28264 20584
rect 27828 20553 27840 20556
rect 27782 20547 27840 20553
rect 28258 20544 28264 20556
rect 28316 20544 28322 20596
rect 28626 20584 28632 20596
rect 28587 20556 28632 20584
rect 28626 20544 28632 20556
rect 28684 20544 28690 20596
rect 29086 20584 29092 20596
rect 29047 20556 29092 20584
rect 29086 20544 29092 20556
rect 29144 20544 29150 20596
rect 30926 20544 30932 20596
rect 30984 20584 30990 20596
rect 31481 20587 31539 20593
rect 31481 20584 31493 20587
rect 30984 20556 31493 20584
rect 30984 20544 30990 20556
rect 31481 20553 31493 20556
rect 31527 20553 31539 20587
rect 32030 20584 32036 20596
rect 31991 20556 32036 20584
rect 31481 20547 31539 20553
rect 32030 20544 32036 20556
rect 32088 20544 32094 20596
rect 32490 20584 32496 20596
rect 32451 20556 32496 20584
rect 32490 20544 32496 20556
rect 32548 20544 32554 20596
rect 32674 20544 32680 20596
rect 32732 20584 32738 20596
rect 33045 20587 33103 20593
rect 33045 20584 33057 20587
rect 32732 20556 33057 20584
rect 32732 20544 32738 20556
rect 33045 20553 33057 20556
rect 33091 20553 33103 20587
rect 33045 20547 33103 20553
rect 34054 20544 34060 20596
rect 34112 20584 34118 20596
rect 34241 20587 34299 20593
rect 34241 20584 34253 20587
rect 34112 20556 34253 20584
rect 34112 20544 34118 20556
rect 34241 20553 34253 20556
rect 34287 20553 34299 20587
rect 34606 20584 34612 20596
rect 34567 20556 34612 20584
rect 34241 20547 34299 20553
rect 34606 20544 34612 20556
rect 34664 20584 34670 20596
rect 35023 20587 35081 20593
rect 35023 20584 35035 20587
rect 34664 20556 35035 20584
rect 34664 20544 34670 20556
rect 35023 20553 35035 20556
rect 35069 20553 35081 20587
rect 35434 20584 35440 20596
rect 35395 20556 35440 20584
rect 35023 20547 35081 20553
rect 35434 20544 35440 20556
rect 35492 20544 35498 20596
rect 36170 20544 36176 20596
rect 36228 20584 36234 20596
rect 37369 20587 37427 20593
rect 37369 20584 37381 20587
rect 36228 20556 37381 20584
rect 36228 20544 36234 20556
rect 37369 20553 37381 20556
rect 37415 20553 37427 20587
rect 37369 20547 37427 20553
rect 38838 20544 38844 20596
rect 38896 20584 38902 20596
rect 38933 20587 38991 20593
rect 38933 20584 38945 20587
rect 38896 20556 38945 20584
rect 38896 20544 38902 20556
rect 38933 20553 38945 20556
rect 38979 20553 38991 20587
rect 38933 20547 38991 20553
rect 39022 20544 39028 20596
rect 39080 20584 39086 20596
rect 39301 20587 39359 20593
rect 39301 20584 39313 20587
rect 39080 20556 39313 20584
rect 39080 20544 39086 20556
rect 39301 20553 39313 20556
rect 39347 20553 39359 20587
rect 39666 20584 39672 20596
rect 39627 20556 39672 20584
rect 39301 20547 39359 20553
rect 39666 20544 39672 20556
rect 39724 20544 39730 20596
rect 42705 20587 42763 20593
rect 42705 20553 42717 20587
rect 42751 20584 42763 20587
rect 42935 20587 42993 20593
rect 42935 20584 42947 20587
rect 42751 20556 42947 20584
rect 42751 20553 42763 20556
rect 42705 20547 42763 20553
rect 42935 20553 42947 20556
rect 42981 20584 42993 20587
rect 43438 20584 43444 20596
rect 42981 20556 43444 20584
rect 42981 20553 42993 20556
rect 42935 20547 42993 20553
rect 43438 20544 43444 20556
rect 43496 20544 43502 20596
rect 44266 20584 44272 20596
rect 44227 20556 44272 20584
rect 44266 20544 44272 20556
rect 44324 20544 44330 20596
rect 19150 20516 19156 20528
rect 19111 20488 19156 20516
rect 19150 20476 19156 20488
rect 19208 20476 19214 20528
rect 23017 20519 23075 20525
rect 23017 20485 23029 20519
rect 23063 20516 23075 20519
rect 23566 20516 23572 20528
rect 23063 20488 23572 20516
rect 23063 20485 23075 20488
rect 23017 20479 23075 20485
rect 23566 20476 23572 20488
rect 23624 20476 23630 20528
rect 27430 20476 27436 20528
rect 27488 20516 27494 20528
rect 27893 20519 27951 20525
rect 27893 20516 27905 20519
rect 27488 20488 27905 20516
rect 27488 20476 27494 20488
rect 27893 20485 27905 20488
rect 27939 20516 27951 20519
rect 28074 20516 28080 20528
rect 27939 20488 28080 20516
rect 27939 20485 27951 20488
rect 27893 20479 27951 20485
rect 28074 20476 28080 20488
rect 28132 20476 28138 20528
rect 31110 20516 31116 20528
rect 31071 20488 31116 20516
rect 31110 20476 31116 20488
rect 31168 20476 31174 20528
rect 32766 20476 32772 20528
rect 32824 20516 32830 20528
rect 36630 20516 36636 20528
rect 32824 20488 36636 20516
rect 32824 20476 32830 20488
rect 36630 20476 36636 20488
rect 36688 20476 36694 20528
rect 43898 20516 43904 20528
rect 43272 20488 43904 20516
rect 18141 20451 18199 20457
rect 18141 20417 18153 20451
rect 18187 20448 18199 20451
rect 21269 20451 21327 20457
rect 18187 20420 19932 20448
rect 18187 20417 18199 20420
rect 18141 20411 18199 20417
rect 18233 20315 18291 20321
rect 18233 20312 18245 20315
rect 17788 20284 18245 20312
rect 18233 20281 18245 20284
rect 18279 20281 18291 20315
rect 18233 20275 18291 20281
rect 18785 20315 18843 20321
rect 18785 20281 18797 20315
rect 18831 20312 18843 20315
rect 19058 20312 19064 20324
rect 18831 20284 19064 20312
rect 18831 20281 18843 20284
rect 18785 20275 18843 20281
rect 15436 20216 15700 20244
rect 15436 20204 15442 20216
rect 16022 20204 16028 20256
rect 16080 20244 16086 20256
rect 18800 20244 18828 20275
rect 19058 20272 19064 20284
rect 19116 20272 19122 20324
rect 19904 20253 19932 20420
rect 21269 20417 21281 20451
rect 21315 20448 21327 20451
rect 21358 20448 21364 20460
rect 21315 20420 21364 20448
rect 21315 20417 21327 20420
rect 21269 20411 21327 20417
rect 21358 20408 21364 20420
rect 21416 20408 21422 20460
rect 23198 20408 23204 20460
rect 23256 20448 23262 20460
rect 24029 20451 24087 20457
rect 24029 20448 24041 20451
rect 23256 20420 24041 20448
rect 23256 20408 23262 20420
rect 24029 20417 24041 20420
rect 24075 20417 24087 20451
rect 24029 20411 24087 20417
rect 26510 20408 26516 20460
rect 26568 20448 26574 20460
rect 27985 20451 28043 20457
rect 26568 20420 26832 20448
rect 26568 20408 26574 20420
rect 20533 20383 20591 20389
rect 20533 20349 20545 20383
rect 20579 20349 20591 20383
rect 20533 20343 20591 20349
rect 16080 20216 18828 20244
rect 19889 20247 19947 20253
rect 16080 20204 16086 20216
rect 19889 20213 19901 20247
rect 19935 20244 19947 20247
rect 19978 20244 19984 20256
rect 19935 20216 19984 20244
rect 19935 20213 19947 20216
rect 19889 20207 19947 20213
rect 19978 20204 19984 20216
rect 20036 20204 20042 20256
rect 20346 20244 20352 20256
rect 20307 20216 20352 20244
rect 20346 20204 20352 20216
rect 20404 20244 20410 20256
rect 20548 20244 20576 20343
rect 20622 20340 20628 20392
rect 20680 20380 20686 20392
rect 20993 20383 21051 20389
rect 20993 20380 21005 20383
rect 20680 20352 21005 20380
rect 20680 20340 20686 20352
rect 20993 20349 21005 20352
rect 21039 20349 21051 20383
rect 20993 20343 21051 20349
rect 21542 20340 21548 20392
rect 21600 20380 21606 20392
rect 22132 20383 22190 20389
rect 22132 20380 22144 20383
rect 21600 20352 22144 20380
rect 21600 20340 21606 20352
rect 22132 20349 22144 20352
rect 22178 20380 22190 20383
rect 22557 20383 22615 20389
rect 22557 20380 22569 20383
rect 22178 20352 22569 20380
rect 22178 20349 22190 20352
rect 22132 20343 22190 20349
rect 22557 20349 22569 20352
rect 22603 20349 22615 20383
rect 22557 20343 22615 20349
rect 25317 20383 25375 20389
rect 25317 20349 25329 20383
rect 25363 20380 25375 20383
rect 26053 20383 26111 20389
rect 26053 20380 26065 20383
rect 25363 20352 26065 20380
rect 25363 20349 25375 20352
rect 25317 20343 25375 20349
rect 26053 20349 26065 20352
rect 26099 20380 26111 20383
rect 26694 20380 26700 20392
rect 26099 20352 26700 20380
rect 26099 20349 26111 20352
rect 26053 20343 26111 20349
rect 26694 20340 26700 20352
rect 26752 20340 26758 20392
rect 26804 20389 26832 20420
rect 27985 20417 27997 20451
rect 28031 20417 28043 20451
rect 27985 20411 28043 20417
rect 29917 20451 29975 20457
rect 29917 20417 29929 20451
rect 29963 20448 29975 20451
rect 30006 20448 30012 20460
rect 29963 20420 30012 20448
rect 29963 20417 29975 20420
rect 29917 20411 29975 20417
rect 26789 20383 26847 20389
rect 26789 20349 26801 20383
rect 26835 20380 26847 20383
rect 27617 20383 27675 20389
rect 27617 20380 27629 20383
rect 26835 20352 27629 20380
rect 26835 20349 26847 20352
rect 26789 20343 26847 20349
rect 27617 20349 27629 20352
rect 27663 20349 27675 20383
rect 27617 20343 27675 20349
rect 23750 20312 23756 20324
rect 23711 20284 23756 20312
rect 23750 20272 23756 20284
rect 23808 20272 23814 20324
rect 23845 20315 23903 20321
rect 23845 20281 23857 20315
rect 23891 20281 23903 20315
rect 27706 20312 27712 20324
rect 23845 20275 23903 20281
rect 27080 20284 27712 20312
rect 20404 20216 20576 20244
rect 20404 20204 20410 20216
rect 23382 20204 23388 20256
rect 23440 20244 23446 20256
rect 23860 20244 23888 20275
rect 23440 20216 23888 20244
rect 23440 20204 23446 20216
rect 26142 20204 26148 20256
rect 26200 20244 26206 20256
rect 27080 20253 27108 20284
rect 27706 20272 27712 20284
rect 27764 20312 27770 20324
rect 28000 20312 28028 20411
rect 30006 20408 30012 20420
rect 30064 20408 30070 20460
rect 33321 20451 33379 20457
rect 33321 20417 33333 20451
rect 33367 20448 33379 20451
rect 33686 20448 33692 20460
rect 33367 20420 33692 20448
rect 33367 20417 33379 20420
rect 33321 20411 33379 20417
rect 33686 20408 33692 20420
rect 33744 20408 33750 20460
rect 33778 20408 33784 20460
rect 33836 20448 33842 20460
rect 33836 20420 33881 20448
rect 33836 20408 33842 20420
rect 34698 20408 34704 20460
rect 34756 20448 34762 20460
rect 35989 20451 36047 20457
rect 35989 20448 36001 20451
rect 34756 20420 36001 20448
rect 34756 20408 34762 20420
rect 35989 20417 36001 20420
rect 36035 20417 36047 20451
rect 35989 20411 36047 20417
rect 36173 20451 36231 20457
rect 36173 20417 36185 20451
rect 36219 20448 36231 20451
rect 36446 20448 36452 20460
rect 36219 20420 36452 20448
rect 36219 20417 36231 20420
rect 36173 20411 36231 20417
rect 29822 20340 29828 20392
rect 29880 20380 29886 20392
rect 32284 20383 32342 20389
rect 29880 20352 30328 20380
rect 29880 20340 29886 20352
rect 27764 20284 28028 20312
rect 28353 20315 28411 20321
rect 27764 20272 27770 20284
rect 28353 20281 28365 20315
rect 28399 20312 28411 20315
rect 30098 20312 30104 20324
rect 28399 20284 30104 20312
rect 28399 20281 28411 20284
rect 28353 20275 28411 20281
rect 30098 20272 30104 20284
rect 30156 20272 30162 20324
rect 30300 20321 30328 20352
rect 32284 20349 32296 20383
rect 32330 20380 32342 20383
rect 32674 20380 32680 20392
rect 32330 20352 32680 20380
rect 32330 20349 32342 20352
rect 32284 20343 32342 20349
rect 32674 20340 32680 20352
rect 32732 20340 32738 20392
rect 34952 20383 35010 20389
rect 34952 20349 34964 20383
rect 34998 20380 35010 20383
rect 35434 20380 35440 20392
rect 34998 20352 35440 20380
rect 34998 20349 35010 20352
rect 34952 20343 35010 20349
rect 35434 20340 35440 20352
rect 35492 20340 35498 20392
rect 30279 20315 30337 20321
rect 30279 20281 30291 20315
rect 30325 20312 30337 20315
rect 30325 20284 31064 20312
rect 30325 20281 30337 20284
rect 30279 20275 30337 20281
rect 27065 20247 27123 20253
rect 27065 20244 27077 20247
rect 26200 20216 27077 20244
rect 26200 20204 26206 20216
rect 27065 20213 27077 20216
rect 27111 20213 27123 20247
rect 27430 20244 27436 20256
rect 27391 20216 27436 20244
rect 27065 20207 27123 20213
rect 27430 20204 27436 20216
rect 27488 20204 27494 20256
rect 29825 20247 29883 20253
rect 29825 20213 29837 20247
rect 29871 20244 29883 20247
rect 29914 20244 29920 20256
rect 29871 20216 29920 20244
rect 29871 20213 29883 20216
rect 29825 20207 29883 20213
rect 29914 20204 29920 20216
rect 29972 20204 29978 20256
rect 30650 20204 30656 20256
rect 30708 20244 30714 20256
rect 30837 20247 30895 20253
rect 30837 20244 30849 20247
rect 30708 20216 30849 20244
rect 30708 20204 30714 20216
rect 30837 20213 30849 20216
rect 30883 20213 30895 20247
rect 31036 20244 31064 20284
rect 31110 20272 31116 20324
rect 31168 20312 31174 20324
rect 33318 20312 33324 20324
rect 31168 20284 33324 20312
rect 31168 20272 31174 20284
rect 33318 20272 33324 20284
rect 33376 20272 33382 20324
rect 33413 20315 33471 20321
rect 33413 20281 33425 20315
rect 33459 20281 33471 20315
rect 36004 20312 36032 20411
rect 36446 20408 36452 20420
rect 36504 20408 36510 20460
rect 38013 20451 38071 20457
rect 38013 20417 38025 20451
rect 38059 20448 38071 20451
rect 38102 20448 38108 20460
rect 38059 20420 38108 20448
rect 38059 20417 38071 20420
rect 38013 20411 38071 20417
rect 38102 20408 38108 20420
rect 38160 20408 38166 20460
rect 40034 20408 40040 20460
rect 40092 20448 40098 20460
rect 41601 20451 41659 20457
rect 41601 20448 41613 20451
rect 40092 20420 41613 20448
rect 40092 20408 40098 20420
rect 41601 20417 41613 20420
rect 41647 20448 41659 20451
rect 41966 20448 41972 20460
rect 41647 20420 41972 20448
rect 41647 20417 41659 20420
rect 41601 20411 41659 20417
rect 41966 20408 41972 20420
rect 42024 20408 42030 20460
rect 42886 20389 42892 20392
rect 42864 20383 42892 20389
rect 42864 20380 42876 20383
rect 42799 20352 42876 20380
rect 42864 20349 42876 20352
rect 42944 20380 42950 20392
rect 43272 20389 43300 20488
rect 43898 20476 43904 20488
rect 43956 20476 43962 20528
rect 43257 20383 43315 20389
rect 43257 20380 43269 20383
rect 42944 20352 43269 20380
rect 42864 20343 42892 20349
rect 42886 20340 42892 20343
rect 42944 20340 42950 20352
rect 43257 20349 43269 20352
rect 43303 20349 43315 20383
rect 43806 20380 43812 20392
rect 43770 20352 43812 20380
rect 43257 20343 43315 20349
rect 43806 20340 43812 20352
rect 43864 20389 43870 20392
rect 43864 20383 43918 20389
rect 43864 20349 43872 20383
rect 43906 20380 43918 20383
rect 44266 20380 44272 20392
rect 43906 20352 44272 20380
rect 43906 20349 43918 20352
rect 43864 20343 43918 20349
rect 43864 20340 43870 20343
rect 44266 20340 44272 20352
rect 44324 20340 44330 20392
rect 36494 20315 36552 20321
rect 36494 20312 36506 20315
rect 36004 20284 36506 20312
rect 33413 20275 33471 20281
rect 36494 20281 36506 20284
rect 36540 20312 36552 20315
rect 36814 20312 36820 20324
rect 36540 20284 36820 20312
rect 36540 20281 36552 20284
rect 36494 20275 36552 20281
rect 32398 20244 32404 20256
rect 31036 20216 32404 20244
rect 30837 20207 30895 20213
rect 32398 20204 32404 20216
rect 32456 20244 32462 20256
rect 32677 20247 32735 20253
rect 32677 20244 32689 20247
rect 32456 20216 32689 20244
rect 32456 20204 32462 20216
rect 32677 20213 32689 20216
rect 32723 20213 32735 20247
rect 32677 20207 32735 20213
rect 33134 20204 33140 20256
rect 33192 20244 33198 20256
rect 33428 20244 33456 20275
rect 36814 20272 36820 20284
rect 36872 20272 36878 20324
rect 37737 20315 37795 20321
rect 37737 20312 37749 20315
rect 37108 20284 37749 20312
rect 33192 20216 33456 20244
rect 33192 20204 33198 20216
rect 36262 20204 36268 20256
rect 36320 20244 36326 20256
rect 36906 20244 36912 20256
rect 36320 20216 36912 20244
rect 36320 20204 36326 20216
rect 36906 20204 36912 20216
rect 36964 20244 36970 20256
rect 37108 20253 37136 20284
rect 37737 20281 37749 20284
rect 37783 20281 37795 20315
rect 37737 20275 37795 20281
rect 38105 20315 38163 20321
rect 38105 20281 38117 20315
rect 38151 20281 38163 20315
rect 38105 20275 38163 20281
rect 38657 20315 38715 20321
rect 38657 20281 38669 20315
rect 38703 20312 38715 20315
rect 39206 20312 39212 20324
rect 38703 20284 39212 20312
rect 38703 20281 38715 20284
rect 38657 20275 38715 20281
rect 37093 20247 37151 20253
rect 37093 20244 37105 20247
rect 36964 20216 37105 20244
rect 36964 20204 36970 20216
rect 37093 20213 37105 20216
rect 37139 20213 37151 20247
rect 37752 20244 37780 20275
rect 38120 20244 38148 20275
rect 39206 20272 39212 20284
rect 39264 20272 39270 20324
rect 41322 20312 41328 20324
rect 41283 20284 41328 20312
rect 41322 20272 41328 20284
rect 41380 20272 41386 20324
rect 41417 20315 41475 20321
rect 41417 20281 41429 20315
rect 41463 20312 41475 20315
rect 41598 20312 41604 20324
rect 41463 20284 41604 20312
rect 41463 20281 41475 20284
rect 41417 20275 41475 20281
rect 41598 20272 41604 20284
rect 41656 20272 41662 20324
rect 43438 20272 43444 20324
rect 43496 20312 43502 20324
rect 43947 20315 44005 20321
rect 43947 20312 43959 20315
rect 43496 20284 43959 20312
rect 43496 20272 43502 20284
rect 43947 20281 43959 20284
rect 43993 20281 44005 20315
rect 43947 20275 44005 20281
rect 37752 20216 38148 20244
rect 40773 20247 40831 20253
rect 37093 20207 37151 20213
rect 40773 20213 40785 20247
rect 40819 20244 40831 20247
rect 41046 20244 41052 20256
rect 40819 20216 41052 20244
rect 40819 20213 40831 20216
rect 40773 20207 40831 20213
rect 41046 20204 41052 20216
rect 41104 20204 41110 20256
rect 41138 20204 41144 20256
rect 41196 20244 41202 20256
rect 42245 20247 42303 20253
rect 42245 20244 42257 20247
rect 41196 20216 42257 20244
rect 41196 20204 41202 20216
rect 42245 20213 42257 20216
rect 42291 20213 42303 20247
rect 43622 20244 43628 20256
rect 43583 20216 43628 20244
rect 42245 20207 42303 20213
rect 43622 20204 43628 20216
rect 43680 20204 43686 20256
rect 1104 20154 48852 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 48852 20154
rect 1104 20080 48852 20102
rect 10045 20043 10103 20049
rect 10045 20009 10057 20043
rect 10091 20040 10103 20043
rect 10594 20040 10600 20052
rect 10091 20012 10600 20040
rect 10091 20009 10103 20012
rect 10045 20003 10103 20009
rect 10594 20000 10600 20012
rect 10652 20000 10658 20052
rect 16298 20040 16304 20052
rect 16259 20012 16304 20040
rect 16298 20000 16304 20012
rect 16356 20000 16362 20052
rect 16942 20000 16948 20052
rect 17000 20040 17006 20052
rect 17494 20040 17500 20052
rect 17000 20012 17264 20040
rect 17455 20012 17500 20040
rect 17000 20000 17006 20012
rect 10962 19932 10968 19984
rect 11020 19972 11026 19984
rect 11057 19975 11115 19981
rect 11057 19972 11069 19975
rect 11020 19944 11069 19972
rect 11020 19932 11026 19944
rect 11057 19941 11069 19944
rect 11103 19941 11115 19975
rect 13262 19972 13268 19984
rect 13223 19944 13268 19972
rect 11057 19935 11115 19941
rect 13262 19932 13268 19944
rect 13320 19932 13326 19984
rect 15194 19932 15200 19984
rect 15252 19972 15258 19984
rect 15381 19975 15439 19981
rect 15381 19972 15393 19975
rect 15252 19944 15393 19972
rect 15252 19932 15258 19944
rect 15381 19941 15393 19944
rect 15427 19941 15439 19975
rect 15381 19935 15439 19941
rect 15473 19975 15531 19981
rect 15473 19941 15485 19975
rect 15519 19972 15531 19975
rect 15838 19972 15844 19984
rect 15519 19944 15844 19972
rect 15519 19941 15531 19944
rect 15473 19935 15531 19941
rect 15838 19932 15844 19944
rect 15896 19932 15902 19984
rect 16022 19972 16028 19984
rect 15983 19944 16028 19972
rect 16022 19932 16028 19944
rect 16080 19932 16086 19984
rect 17236 19972 17264 20012
rect 17494 20000 17500 20012
rect 17552 20000 17558 20052
rect 18414 20000 18420 20052
rect 18472 20040 18478 20052
rect 20346 20040 20352 20052
rect 18472 20012 20352 20040
rect 18472 20000 18478 20012
rect 20346 20000 20352 20012
rect 20404 20000 20410 20052
rect 20530 20040 20536 20052
rect 20491 20012 20536 20040
rect 20530 20000 20536 20012
rect 20588 20000 20594 20052
rect 26142 20040 26148 20052
rect 21284 20012 26148 20040
rect 18095 19975 18153 19981
rect 18095 19972 18107 19975
rect 17236 19944 18107 19972
rect 18095 19941 18107 19944
rect 18141 19941 18153 19975
rect 18095 19935 18153 19941
rect 19153 19975 19211 19981
rect 19153 19941 19165 19975
rect 19199 19972 19211 19975
rect 19334 19972 19340 19984
rect 19199 19944 19340 19972
rect 19199 19941 19211 19944
rect 19153 19935 19211 19941
rect 19334 19932 19340 19944
rect 19392 19972 19398 19984
rect 20162 19972 20168 19984
rect 19392 19944 20168 19972
rect 19392 19932 19398 19944
rect 20162 19932 20168 19944
rect 20220 19932 20226 19984
rect 20806 19932 20812 19984
rect 20864 19972 20870 19984
rect 20901 19975 20959 19981
rect 20901 19972 20913 19975
rect 20864 19944 20913 19972
rect 20864 19932 20870 19944
rect 20901 19941 20913 19944
rect 20947 19941 20959 19975
rect 20901 19935 20959 19941
rect 9861 19907 9919 19913
rect 9861 19873 9873 19907
rect 9907 19904 9919 19907
rect 10134 19904 10140 19916
rect 9907 19876 10140 19904
rect 9907 19873 9919 19876
rect 9861 19867 9919 19873
rect 10134 19864 10140 19876
rect 10192 19864 10198 19916
rect 16758 19864 16764 19916
rect 16816 19904 16822 19916
rect 16980 19907 17038 19913
rect 16980 19904 16992 19907
rect 16816 19876 16992 19904
rect 16816 19864 16822 19876
rect 16980 19873 16992 19876
rect 17026 19873 17038 19907
rect 17954 19904 17960 19916
rect 17915 19876 17960 19904
rect 16980 19867 17038 19873
rect 17954 19864 17960 19876
rect 18012 19864 18018 19916
rect 19242 19904 19248 19916
rect 19203 19876 19248 19904
rect 19242 19864 19248 19876
rect 19300 19864 19306 19916
rect 20824 19904 20852 19932
rect 19352 19876 20852 19904
rect 10965 19839 11023 19845
rect 10965 19805 10977 19839
rect 11011 19836 11023 19839
rect 11238 19836 11244 19848
rect 11011 19808 11244 19836
rect 11011 19805 11023 19808
rect 10965 19799 11023 19805
rect 11238 19796 11244 19808
rect 11296 19836 11302 19848
rect 13170 19836 13176 19848
rect 11296 19808 12434 19836
rect 13131 19808 13176 19836
rect 11296 19796 11302 19808
rect 11514 19768 11520 19780
rect 11475 19740 11520 19768
rect 11514 19728 11520 19740
rect 11572 19728 11578 19780
rect 12406 19768 12434 19808
rect 13170 19796 13176 19808
rect 13228 19796 13234 19848
rect 13449 19839 13507 19845
rect 13449 19805 13461 19839
rect 13495 19805 13507 19839
rect 13449 19799 13507 19805
rect 18785 19839 18843 19845
rect 18785 19805 18797 19839
rect 18831 19836 18843 19839
rect 19058 19836 19064 19848
rect 18831 19808 19064 19836
rect 18831 19805 18843 19808
rect 18785 19799 18843 19805
rect 13354 19768 13360 19780
rect 12406 19740 13360 19768
rect 13354 19728 13360 19740
rect 13412 19768 13418 19780
rect 13464 19768 13492 19799
rect 19058 19796 19064 19808
rect 19116 19836 19122 19848
rect 19352 19836 19380 19876
rect 19116 19808 19380 19836
rect 19613 19839 19671 19845
rect 19116 19796 19122 19808
rect 19613 19805 19625 19839
rect 19659 19836 19671 19839
rect 20990 19836 20996 19848
rect 19659 19808 20996 19836
rect 19659 19805 19671 19808
rect 19613 19799 19671 19805
rect 20990 19796 20996 19808
rect 21048 19836 21054 19848
rect 21284 19845 21312 20012
rect 26142 20000 26148 20012
rect 26200 20000 26206 20052
rect 26326 20040 26332 20052
rect 26287 20012 26332 20040
rect 26326 20000 26332 20012
rect 26384 20000 26390 20052
rect 27614 20000 27620 20052
rect 27672 20040 27678 20052
rect 28537 20043 28595 20049
rect 28537 20040 28549 20043
rect 27672 20012 28549 20040
rect 27672 20000 27678 20012
rect 28537 20009 28549 20012
rect 28583 20009 28595 20043
rect 30006 20040 30012 20052
rect 29967 20012 30012 20040
rect 28537 20003 28595 20009
rect 30006 20000 30012 20012
rect 30064 20000 30070 20052
rect 32723 20043 32781 20049
rect 32723 20009 32735 20043
rect 32769 20040 32781 20043
rect 33686 20040 33692 20052
rect 32769 20012 33692 20040
rect 32769 20009 32781 20012
rect 32723 20003 32781 20009
rect 33686 20000 33692 20012
rect 33744 20000 33750 20052
rect 40494 20040 40500 20052
rect 40455 20012 40500 20040
rect 40494 20000 40500 20012
rect 40552 20000 40558 20052
rect 42978 20000 42984 20052
rect 43036 20040 43042 20052
rect 43036 20012 44991 20040
rect 43036 20000 43042 20012
rect 23106 19932 23112 19984
rect 23164 19972 23170 19984
rect 23385 19975 23443 19981
rect 23385 19972 23397 19975
rect 23164 19944 23397 19972
rect 23164 19932 23170 19944
rect 23385 19941 23397 19944
rect 23431 19941 23443 19975
rect 23385 19935 23443 19941
rect 25041 19975 25099 19981
rect 25041 19941 25053 19975
rect 25087 19972 25099 19975
rect 26234 19972 26240 19984
rect 25087 19944 26240 19972
rect 25087 19941 25099 19944
rect 25041 19935 25099 19941
rect 26234 19932 26240 19944
rect 26292 19972 26298 19984
rect 26697 19975 26755 19981
rect 26697 19972 26709 19975
rect 26292 19944 26709 19972
rect 26292 19932 26298 19944
rect 26697 19941 26709 19944
rect 26743 19941 26755 19975
rect 30650 19972 30656 19984
rect 30611 19944 30656 19972
rect 26697 19935 26755 19941
rect 30650 19932 30656 19944
rect 30708 19932 30714 19984
rect 33134 19932 33140 19984
rect 33192 19972 33198 19984
rect 33229 19975 33287 19981
rect 33229 19972 33241 19975
rect 33192 19944 33241 19972
rect 33192 19932 33198 19944
rect 33229 19941 33241 19944
rect 33275 19941 33287 19975
rect 33781 19975 33839 19981
rect 33781 19972 33793 19975
rect 33229 19935 33287 19941
rect 33520 19944 33793 19972
rect 27338 19864 27344 19916
rect 27396 19904 27402 19916
rect 28077 19907 28135 19913
rect 28077 19904 28089 19907
rect 27396 19876 28089 19904
rect 27396 19864 27402 19876
rect 28077 19873 28089 19876
rect 28123 19904 28135 19907
rect 28626 19904 28632 19916
rect 28123 19876 28632 19904
rect 28123 19873 28135 19876
rect 28077 19867 28135 19873
rect 28626 19864 28632 19876
rect 28684 19864 28690 19916
rect 29454 19904 29460 19916
rect 29415 19876 29460 19904
rect 29454 19864 29460 19876
rect 29512 19864 29518 19916
rect 32652 19907 32710 19913
rect 32652 19873 32664 19907
rect 32698 19904 32710 19907
rect 32766 19904 32772 19916
rect 32698 19876 32772 19904
rect 32698 19873 32710 19876
rect 32652 19867 32710 19873
rect 32766 19864 32772 19876
rect 32824 19864 32830 19916
rect 32858 19864 32864 19916
rect 32916 19904 32922 19916
rect 33520 19904 33548 19944
rect 33781 19941 33793 19944
rect 33827 19972 33839 19975
rect 34054 19972 34060 19984
rect 33827 19944 34060 19972
rect 33827 19941 33839 19944
rect 33781 19935 33839 19941
rect 34054 19932 34060 19944
rect 34112 19932 34118 19984
rect 35986 19932 35992 19984
rect 36044 19972 36050 19984
rect 36173 19975 36231 19981
rect 36173 19972 36185 19975
rect 36044 19944 36185 19972
rect 36044 19932 36050 19944
rect 36173 19941 36185 19944
rect 36219 19941 36231 19975
rect 36173 19935 36231 19941
rect 36262 19932 36268 19984
rect 36320 19972 36326 19984
rect 36320 19944 36365 19972
rect 36320 19932 36326 19944
rect 37918 19932 37924 19984
rect 37976 19972 37982 19984
rect 38565 19975 38623 19981
rect 38565 19972 38577 19975
rect 37976 19944 38577 19972
rect 37976 19932 37982 19944
rect 38565 19941 38577 19944
rect 38611 19941 38623 19975
rect 38565 19935 38623 19941
rect 38654 19932 38660 19984
rect 38712 19972 38718 19984
rect 40862 19972 40868 19984
rect 38712 19944 40868 19972
rect 38712 19932 38718 19944
rect 40862 19932 40868 19944
rect 40920 19972 40926 19984
rect 43438 19972 43444 19984
rect 40920 19944 41955 19972
rect 43399 19944 43444 19972
rect 40920 19932 40926 19944
rect 41046 19904 41052 19916
rect 32916 19876 33548 19904
rect 40959 19876 41052 19904
rect 32916 19864 32922 19876
rect 41046 19864 41052 19876
rect 41104 19904 41110 19916
rect 41598 19904 41604 19916
rect 41104 19876 41604 19904
rect 41104 19864 41110 19876
rect 41598 19864 41604 19876
rect 41656 19864 41662 19916
rect 41927 19913 41955 19944
rect 43438 19932 43444 19944
rect 43496 19932 43502 19984
rect 43533 19975 43591 19981
rect 43533 19941 43545 19975
rect 43579 19972 43591 19975
rect 43622 19972 43628 19984
rect 43579 19944 43628 19972
rect 43579 19941 43591 19944
rect 43533 19935 43591 19941
rect 43622 19932 43628 19944
rect 43680 19972 43686 19984
rect 44082 19972 44088 19984
rect 43680 19944 44088 19972
rect 43680 19932 43686 19944
rect 44082 19932 44088 19944
rect 44140 19932 44146 19984
rect 44963 19916 44991 20012
rect 41912 19907 41970 19913
rect 41912 19873 41924 19907
rect 41958 19904 41970 19907
rect 42702 19904 42708 19916
rect 41958 19876 42708 19904
rect 41958 19873 41970 19876
rect 41912 19867 41970 19873
rect 42702 19864 42708 19876
rect 42760 19864 42766 19916
rect 44910 19904 44916 19916
rect 44968 19913 44991 19916
rect 44968 19907 45006 19913
rect 44858 19876 44916 19904
rect 44910 19864 44916 19876
rect 44994 19873 45006 19907
rect 44968 19867 45006 19873
rect 44968 19864 44974 19867
rect 21269 19839 21327 19845
rect 21269 19836 21281 19839
rect 21048 19808 21281 19836
rect 21048 19796 21054 19808
rect 21269 19805 21281 19808
rect 21315 19805 21327 19839
rect 21269 19799 21327 19805
rect 23109 19839 23167 19845
rect 23109 19805 23121 19839
rect 23155 19836 23167 19839
rect 23290 19836 23296 19848
rect 23155 19808 23296 19836
rect 23155 19805 23167 19808
rect 23109 19799 23167 19805
rect 23290 19796 23296 19808
rect 23348 19796 23354 19848
rect 23569 19839 23627 19845
rect 23569 19836 23581 19839
rect 23446 19808 23581 19836
rect 13412 19740 13492 19768
rect 13412 19728 13418 19740
rect 19150 19728 19156 19780
rect 19208 19768 19214 19780
rect 19705 19771 19763 19777
rect 19705 19768 19717 19771
rect 19208 19740 19717 19768
rect 19208 19728 19214 19740
rect 19705 19737 19717 19740
rect 19751 19737 19763 19771
rect 19705 19731 19763 19737
rect 20346 19728 20352 19780
rect 20404 19768 20410 19780
rect 21361 19771 21419 19777
rect 21361 19768 21373 19771
rect 20404 19740 21373 19768
rect 20404 19728 20410 19740
rect 21361 19737 21373 19740
rect 21407 19737 21419 19771
rect 21361 19731 21419 19737
rect 23198 19728 23204 19780
rect 23256 19768 23262 19780
rect 23446 19768 23474 19808
rect 23569 19805 23581 19808
rect 23615 19805 23627 19839
rect 23569 19799 23627 19805
rect 24949 19839 25007 19845
rect 24949 19805 24961 19839
rect 24995 19836 25007 19839
rect 25038 19836 25044 19848
rect 24995 19808 25044 19836
rect 24995 19805 25007 19808
rect 24949 19799 25007 19805
rect 25038 19796 25044 19808
rect 25096 19796 25102 19848
rect 25590 19836 25596 19848
rect 25551 19808 25596 19836
rect 25590 19796 25596 19808
rect 25648 19796 25654 19848
rect 26605 19839 26663 19845
rect 26605 19805 26617 19839
rect 26651 19836 26663 19839
rect 26694 19836 26700 19848
rect 26651 19808 26700 19836
rect 26651 19805 26663 19808
rect 26605 19799 26663 19805
rect 26694 19796 26700 19808
rect 26752 19796 26758 19848
rect 26878 19836 26884 19848
rect 26839 19808 26884 19836
rect 26878 19796 26884 19808
rect 26936 19796 26942 19848
rect 29595 19839 29653 19845
rect 29595 19805 29607 19839
rect 29641 19836 29653 19839
rect 30561 19839 30619 19845
rect 30561 19836 30573 19839
rect 29641 19808 30573 19836
rect 29641 19805 29653 19808
rect 29595 19799 29653 19805
rect 30561 19805 30573 19808
rect 30607 19836 30619 19839
rect 31386 19836 31392 19848
rect 30607 19808 31392 19836
rect 30607 19805 30619 19808
rect 30561 19799 30619 19805
rect 31386 19796 31392 19808
rect 31444 19796 31450 19848
rect 32122 19796 32128 19848
rect 32180 19836 32186 19848
rect 33686 19836 33692 19848
rect 32180 19808 33692 19836
rect 32180 19796 32186 19808
rect 33686 19796 33692 19808
rect 33744 19796 33750 19848
rect 33778 19796 33784 19848
rect 33836 19836 33842 19848
rect 33965 19839 34023 19845
rect 33965 19836 33977 19839
rect 33836 19808 33977 19836
rect 33836 19796 33842 19808
rect 33965 19805 33977 19808
rect 34011 19805 34023 19839
rect 36814 19836 36820 19848
rect 36775 19808 36820 19836
rect 33965 19799 34023 19805
rect 36814 19796 36820 19808
rect 36872 19796 36878 19848
rect 38473 19839 38531 19845
rect 38473 19805 38485 19839
rect 38519 19836 38531 19839
rect 38746 19836 38752 19848
rect 38519 19808 38752 19836
rect 38519 19805 38531 19808
rect 38473 19799 38531 19805
rect 38746 19796 38752 19808
rect 38804 19796 38810 19848
rect 39117 19839 39175 19845
rect 39117 19805 39129 19839
rect 39163 19836 39175 19839
rect 39206 19836 39212 19848
rect 39163 19808 39212 19836
rect 39163 19805 39175 19808
rect 39117 19799 39175 19805
rect 39206 19796 39212 19808
rect 39264 19796 39270 19848
rect 40126 19836 40132 19848
rect 40087 19808 40132 19836
rect 40126 19796 40132 19808
rect 40184 19796 40190 19848
rect 40770 19796 40776 19848
rect 40828 19836 40834 19848
rect 42518 19836 42524 19848
rect 40828 19808 42524 19836
rect 40828 19796 40834 19808
rect 42518 19796 42524 19808
rect 42576 19796 42582 19848
rect 43714 19836 43720 19848
rect 43675 19808 43720 19836
rect 43714 19796 43720 19808
rect 43772 19796 43778 19848
rect 23256 19740 23474 19768
rect 23256 19728 23262 19740
rect 23750 19728 23756 19780
rect 23808 19768 23814 19780
rect 25608 19768 25636 19796
rect 23808 19740 25636 19768
rect 31113 19771 31171 19777
rect 23808 19728 23814 19740
rect 31113 19737 31125 19771
rect 31159 19768 31171 19771
rect 31202 19768 31208 19780
rect 31159 19740 31208 19768
rect 31159 19737 31171 19740
rect 31113 19731 31171 19737
rect 31202 19728 31208 19740
rect 31260 19728 31266 19780
rect 33318 19728 33324 19780
rect 33376 19768 33382 19780
rect 35710 19768 35716 19780
rect 33376 19740 35716 19768
rect 33376 19728 33382 19740
rect 35710 19728 35716 19740
rect 35768 19728 35774 19780
rect 41506 19728 41512 19780
rect 41564 19768 41570 19780
rect 42015 19771 42073 19777
rect 42015 19768 42027 19771
rect 41564 19740 42027 19768
rect 41564 19728 41570 19740
rect 42015 19737 42027 19740
rect 42061 19737 42073 19771
rect 42015 19731 42073 19737
rect 42242 19728 42248 19780
rect 42300 19768 42306 19780
rect 43806 19768 43812 19780
rect 42300 19740 43812 19768
rect 42300 19728 42306 19740
rect 43806 19728 43812 19740
rect 43864 19728 43870 19780
rect 14090 19700 14096 19712
rect 14051 19672 14096 19700
rect 14090 19660 14096 19672
rect 14148 19660 14154 19712
rect 16942 19660 16948 19712
rect 17000 19700 17006 19712
rect 17083 19703 17141 19709
rect 17083 19700 17095 19703
rect 17000 19672 17095 19700
rect 17000 19660 17006 19672
rect 17083 19669 17095 19672
rect 17129 19669 17141 19703
rect 17083 19663 17141 19669
rect 19334 19660 19340 19712
rect 19392 19709 19398 19712
rect 19392 19703 19441 19709
rect 19392 19669 19395 19703
rect 19429 19669 19441 19703
rect 19518 19700 19524 19712
rect 19479 19672 19524 19700
rect 19392 19663 19441 19669
rect 19392 19660 19398 19663
rect 19518 19660 19524 19672
rect 19576 19660 19582 19712
rect 20162 19660 20168 19712
rect 20220 19700 20226 19712
rect 21082 19709 21088 19712
rect 21039 19703 21088 19709
rect 21039 19700 21051 19703
rect 20220 19672 21051 19700
rect 20220 19660 20226 19672
rect 21039 19669 21051 19672
rect 21085 19669 21088 19703
rect 21039 19663 21088 19669
rect 21082 19660 21088 19663
rect 21140 19660 21146 19712
rect 21174 19660 21180 19712
rect 21232 19700 21238 19712
rect 24210 19700 24216 19712
rect 21232 19672 21277 19700
rect 24171 19672 24216 19700
rect 21232 19660 21238 19672
rect 24210 19660 24216 19672
rect 24268 19660 24274 19712
rect 24394 19660 24400 19712
rect 24452 19700 24458 19712
rect 24581 19703 24639 19709
rect 24581 19700 24593 19703
rect 24452 19672 24593 19700
rect 24452 19660 24458 19672
rect 24581 19669 24593 19672
rect 24627 19669 24639 19703
rect 24581 19663 24639 19669
rect 26878 19660 26884 19712
rect 26936 19700 26942 19712
rect 27430 19700 27436 19712
rect 26936 19672 27436 19700
rect 26936 19660 26942 19672
rect 27430 19660 27436 19672
rect 27488 19700 27494 19712
rect 27617 19703 27675 19709
rect 27617 19700 27629 19703
rect 27488 19672 27629 19700
rect 27488 19660 27494 19672
rect 27617 19669 27629 19672
rect 27663 19669 27675 19703
rect 27617 19663 27675 19669
rect 27890 19660 27896 19712
rect 27948 19700 27954 19712
rect 28261 19703 28319 19709
rect 28261 19700 28273 19703
rect 27948 19672 28273 19700
rect 27948 19660 27954 19672
rect 28261 19669 28273 19672
rect 28307 19669 28319 19703
rect 28261 19663 28319 19669
rect 29454 19660 29460 19712
rect 29512 19700 29518 19712
rect 37366 19700 37372 19712
rect 29512 19672 37372 19700
rect 29512 19660 29518 19672
rect 37366 19660 37372 19672
rect 37424 19660 37430 19712
rect 38013 19703 38071 19709
rect 38013 19669 38025 19703
rect 38059 19700 38071 19703
rect 38102 19700 38108 19712
rect 38059 19672 38108 19700
rect 38059 19669 38071 19672
rect 38013 19663 38071 19669
rect 38102 19660 38108 19672
rect 38160 19660 38166 19712
rect 41322 19700 41328 19712
rect 41283 19672 41328 19700
rect 41322 19660 41328 19672
rect 41380 19660 41386 19712
rect 41782 19700 41788 19712
rect 41743 19672 41788 19700
rect 41782 19660 41788 19672
rect 41840 19660 41846 19712
rect 43254 19660 43260 19712
rect 43312 19700 43318 19712
rect 45051 19703 45109 19709
rect 45051 19700 45063 19703
rect 43312 19672 45063 19700
rect 43312 19660 43318 19672
rect 45051 19669 45063 19672
rect 45097 19669 45109 19703
rect 45051 19663 45109 19669
rect 1104 19610 48852 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 48852 19610
rect 1104 19536 48852 19558
rect 9953 19499 10011 19505
rect 9953 19465 9965 19499
rect 9999 19496 10011 19499
rect 10134 19496 10140 19508
rect 9999 19468 10140 19496
rect 9999 19465 10011 19468
rect 9953 19459 10011 19465
rect 10134 19456 10140 19468
rect 10192 19456 10198 19508
rect 10686 19496 10692 19508
rect 10647 19468 10692 19496
rect 10686 19456 10692 19468
rect 10744 19456 10750 19508
rect 12158 19496 12164 19508
rect 12119 19468 12164 19496
rect 12158 19456 12164 19468
rect 12216 19456 12222 19508
rect 12618 19496 12624 19508
rect 12579 19468 12624 19496
rect 12618 19456 12624 19468
rect 12676 19456 12682 19508
rect 15194 19496 15200 19508
rect 15155 19468 15200 19496
rect 15194 19456 15200 19468
rect 15252 19456 15258 19508
rect 15838 19496 15844 19508
rect 15799 19468 15844 19496
rect 15838 19456 15844 19468
rect 15896 19456 15902 19508
rect 16758 19456 16764 19508
rect 16816 19496 16822 19508
rect 17402 19496 17408 19508
rect 16816 19468 17408 19496
rect 16816 19456 16822 19468
rect 17402 19456 17408 19468
rect 17460 19456 17466 19508
rect 17494 19456 17500 19508
rect 17552 19496 17558 19508
rect 18187 19499 18245 19505
rect 18187 19496 18199 19499
rect 17552 19468 18199 19496
rect 17552 19456 17558 19468
rect 18187 19465 18199 19468
rect 18233 19465 18245 19499
rect 18187 19459 18245 19465
rect 18874 19456 18880 19508
rect 18932 19496 18938 19508
rect 19705 19499 19763 19505
rect 19705 19496 19717 19499
rect 18932 19468 19717 19496
rect 18932 19456 18938 19468
rect 19705 19465 19717 19468
rect 19751 19465 19763 19499
rect 19705 19459 19763 19465
rect 19978 19456 19984 19508
rect 20036 19496 20042 19508
rect 20947 19499 21005 19505
rect 20947 19496 20959 19499
rect 20036 19468 20959 19496
rect 20036 19456 20042 19468
rect 20947 19465 20959 19468
rect 20993 19465 21005 19499
rect 20947 19459 21005 19465
rect 21082 19456 21088 19508
rect 21140 19496 21146 19508
rect 22465 19499 22523 19505
rect 22465 19496 22477 19499
rect 21140 19468 22477 19496
rect 21140 19456 21146 19468
rect 22465 19465 22477 19468
rect 22511 19465 22523 19499
rect 23106 19496 23112 19508
rect 23067 19468 23112 19496
rect 22465 19459 22523 19465
rect 23106 19456 23112 19468
rect 23164 19456 23170 19508
rect 24949 19499 25007 19505
rect 24949 19465 24961 19499
rect 24995 19496 25007 19499
rect 26234 19496 26240 19508
rect 24995 19468 26240 19496
rect 24995 19465 25007 19468
rect 24949 19459 25007 19465
rect 26234 19456 26240 19468
rect 26292 19496 26298 19508
rect 26513 19499 26571 19505
rect 26513 19496 26525 19499
rect 26292 19468 26525 19496
rect 26292 19456 26298 19468
rect 26513 19465 26525 19468
rect 26559 19465 26571 19499
rect 28258 19496 28264 19508
rect 28219 19468 28264 19496
rect 26513 19459 26571 19465
rect 28258 19456 28264 19468
rect 28316 19456 28322 19508
rect 28626 19496 28632 19508
rect 28587 19468 28632 19496
rect 28626 19456 28632 19468
rect 28684 19456 28690 19508
rect 29089 19499 29147 19505
rect 29089 19465 29101 19499
rect 29135 19496 29147 19499
rect 29454 19496 29460 19508
rect 29135 19468 29460 19496
rect 29135 19465 29147 19468
rect 29089 19459 29147 19465
rect 29454 19456 29460 19468
rect 29512 19456 29518 19508
rect 31386 19496 31392 19508
rect 31347 19468 31392 19496
rect 31386 19456 31392 19468
rect 31444 19456 31450 19508
rect 32766 19496 32772 19508
rect 32727 19468 32772 19496
rect 32766 19456 32772 19468
rect 32824 19456 32830 19508
rect 33686 19456 33692 19508
rect 33744 19496 33750 19508
rect 34609 19499 34667 19505
rect 34609 19496 34621 19499
rect 33744 19468 34621 19496
rect 33744 19456 33750 19468
rect 34609 19465 34621 19468
rect 34655 19465 34667 19499
rect 34609 19459 34667 19465
rect 35805 19499 35863 19505
rect 35805 19465 35817 19499
rect 35851 19496 35863 19499
rect 35986 19496 35992 19508
rect 35851 19468 35992 19496
rect 35851 19465 35863 19468
rect 35805 19459 35863 19465
rect 35986 19456 35992 19468
rect 36044 19456 36050 19508
rect 36173 19499 36231 19505
rect 36173 19465 36185 19499
rect 36219 19496 36231 19499
rect 36262 19496 36268 19508
rect 36219 19468 36268 19496
rect 36219 19465 36231 19468
rect 36173 19459 36231 19465
rect 36262 19456 36268 19468
rect 36320 19456 36326 19508
rect 37550 19496 37556 19508
rect 36418 19468 37556 19496
rect 14274 19428 14280 19440
rect 14235 19400 14280 19428
rect 14274 19388 14280 19400
rect 14332 19388 14338 19440
rect 19334 19388 19340 19440
rect 19392 19437 19398 19440
rect 19392 19431 19441 19437
rect 19392 19397 19395 19431
rect 19429 19397 19441 19431
rect 19392 19391 19441 19397
rect 20717 19431 20775 19437
rect 20717 19397 20729 19431
rect 20763 19428 20775 19431
rect 20806 19428 20812 19440
rect 20763 19400 20812 19428
rect 20763 19397 20775 19400
rect 20717 19391 20775 19397
rect 19392 19388 19398 19391
rect 20806 19388 20812 19400
rect 20864 19388 20870 19440
rect 30650 19388 30656 19440
rect 30708 19428 30714 19440
rect 31113 19431 31171 19437
rect 31113 19428 31125 19431
rect 30708 19400 31125 19428
rect 30708 19388 30714 19400
rect 31113 19397 31125 19400
rect 31159 19428 31171 19431
rect 32858 19428 32864 19440
rect 31159 19400 32864 19428
rect 31159 19397 31171 19400
rect 31113 19391 31171 19397
rect 32858 19388 32864 19400
rect 32916 19388 32922 19440
rect 33134 19388 33140 19440
rect 33192 19428 33198 19440
rect 33192 19400 34008 19428
rect 33192 19388 33198 19400
rect 10321 19363 10379 19369
rect 10321 19329 10333 19363
rect 10367 19360 10379 19363
rect 10873 19363 10931 19369
rect 10873 19360 10885 19363
rect 10367 19332 10885 19360
rect 10367 19329 10379 19332
rect 10321 19323 10379 19329
rect 10873 19329 10885 19332
rect 10919 19360 10931 19363
rect 11054 19360 11060 19372
rect 10919 19332 11060 19360
rect 10919 19329 10931 19332
rect 10873 19323 10931 19329
rect 11054 19320 11060 19332
rect 11112 19320 11118 19372
rect 11514 19360 11520 19372
rect 11475 19332 11520 19360
rect 11514 19320 11520 19332
rect 11572 19320 11578 19372
rect 15378 19360 15384 19372
rect 15339 19332 15384 19360
rect 15378 19320 15384 19332
rect 15436 19320 15442 19372
rect 19153 19363 19211 19369
rect 19153 19329 19165 19363
rect 19199 19360 19211 19363
rect 19613 19363 19671 19369
rect 19613 19360 19625 19363
rect 19199 19332 19625 19360
rect 19199 19329 19211 19332
rect 19153 19323 19211 19329
rect 19613 19329 19625 19332
rect 19659 19360 19671 19363
rect 19886 19360 19892 19372
rect 19659 19332 19892 19360
rect 19659 19329 19671 19332
rect 19613 19323 19671 19329
rect 19886 19320 19892 19332
rect 19944 19320 19950 19372
rect 21729 19363 21787 19369
rect 21729 19360 21741 19363
rect 20859 19332 21741 19360
rect 12158 19252 12164 19304
rect 12216 19292 12222 19304
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 12216 19264 12449 19292
rect 12216 19252 12222 19264
rect 12437 19261 12449 19264
rect 12483 19261 12495 19295
rect 12437 19255 12495 19261
rect 16301 19295 16359 19301
rect 16301 19261 16313 19295
rect 16347 19292 16359 19295
rect 16942 19292 16948 19304
rect 16347 19264 16948 19292
rect 16347 19261 16359 19264
rect 16301 19255 16359 19261
rect 16942 19252 16948 19264
rect 17000 19252 17006 19304
rect 19518 19301 19524 19304
rect 18084 19295 18142 19301
rect 18084 19292 18096 19295
rect 17788 19264 18096 19292
rect 10965 19227 11023 19233
rect 10965 19193 10977 19227
rect 11011 19193 11023 19227
rect 13725 19227 13783 19233
rect 13725 19224 13737 19227
rect 10965 19187 11023 19193
rect 13648 19196 13737 19224
rect 10686 19116 10692 19168
rect 10744 19156 10750 19168
rect 10980 19156 11008 19187
rect 13648 19168 13676 19196
rect 13725 19193 13737 19196
rect 13771 19193 13783 19227
rect 13725 19187 13783 19193
rect 13814 19184 13820 19236
rect 13872 19224 13878 19236
rect 13872 19196 13917 19224
rect 13872 19184 13878 19196
rect 17034 19184 17040 19236
rect 17092 19224 17098 19236
rect 17129 19227 17187 19233
rect 17129 19224 17141 19227
rect 17092 19196 17141 19224
rect 17092 19184 17098 19196
rect 17129 19193 17141 19196
rect 17175 19193 17187 19227
rect 17129 19187 17187 19193
rect 17788 19168 17816 19264
rect 18084 19261 18096 19264
rect 18130 19261 18142 19295
rect 19475 19295 19524 19301
rect 19475 19292 19487 19295
rect 18084 19255 18142 19261
rect 18800 19264 19487 19292
rect 18800 19168 18828 19264
rect 19475 19261 19487 19264
rect 19521 19261 19524 19295
rect 19475 19255 19524 19261
rect 19518 19252 19524 19255
rect 19576 19252 19582 19304
rect 20070 19252 20076 19304
rect 20128 19292 20134 19304
rect 20859 19301 20887 19332
rect 21729 19329 21741 19332
rect 21775 19329 21787 19363
rect 21729 19323 21787 19329
rect 23753 19363 23811 19369
rect 23753 19329 23765 19363
rect 23799 19360 23811 19363
rect 24210 19360 24216 19372
rect 23799 19332 24216 19360
rect 23799 19329 23811 19332
rect 23753 19323 23811 19329
rect 24210 19320 24216 19332
rect 24268 19320 24274 19372
rect 25590 19320 25596 19372
rect 25648 19360 25654 19372
rect 25685 19363 25743 19369
rect 25685 19360 25697 19363
rect 25648 19332 25697 19360
rect 25648 19320 25654 19332
rect 25685 19329 25697 19332
rect 25731 19329 25743 19363
rect 25685 19323 25743 19329
rect 33042 19320 33048 19372
rect 33100 19360 33106 19372
rect 33594 19360 33600 19372
rect 33100 19332 33600 19360
rect 33100 19320 33106 19332
rect 33594 19320 33600 19332
rect 33652 19320 33658 19372
rect 33980 19360 34008 19400
rect 34054 19388 34060 19440
rect 34112 19428 34118 19440
rect 34241 19431 34299 19437
rect 34241 19428 34253 19431
rect 34112 19400 34253 19428
rect 34112 19388 34118 19400
rect 34241 19397 34253 19400
rect 34287 19397 34299 19431
rect 34241 19391 34299 19397
rect 35161 19431 35219 19437
rect 35161 19397 35173 19431
rect 35207 19428 35219 19431
rect 35437 19431 35495 19437
rect 35437 19428 35449 19431
rect 35207 19400 35449 19428
rect 35207 19397 35219 19400
rect 35161 19391 35219 19397
rect 35437 19397 35449 19400
rect 35483 19428 35495 19431
rect 36418 19428 36446 19468
rect 37550 19456 37556 19468
rect 37608 19496 37614 19508
rect 38654 19496 38660 19508
rect 37608 19468 38660 19496
rect 37608 19456 37614 19468
rect 38654 19456 38660 19468
rect 38712 19456 38718 19508
rect 40221 19499 40279 19505
rect 40221 19465 40233 19499
rect 40267 19496 40279 19499
rect 40494 19496 40500 19508
rect 40267 19468 40500 19496
rect 40267 19465 40279 19468
rect 40221 19459 40279 19465
rect 40494 19456 40500 19468
rect 40552 19456 40558 19508
rect 40819 19499 40877 19505
rect 40819 19465 40831 19499
rect 40865 19496 40877 19499
rect 41138 19496 41144 19508
rect 40865 19468 41144 19496
rect 40865 19465 40877 19468
rect 40819 19459 40877 19465
rect 41138 19456 41144 19468
rect 41196 19456 41202 19508
rect 42702 19496 42708 19508
rect 42663 19468 42708 19496
rect 42702 19456 42708 19468
rect 42760 19456 42766 19508
rect 43165 19499 43223 19505
rect 43165 19465 43177 19499
rect 43211 19496 43223 19499
rect 43438 19496 43444 19508
rect 43211 19468 43444 19496
rect 43211 19465 43223 19468
rect 43165 19459 43223 19465
rect 43438 19456 43444 19468
rect 43496 19456 43502 19508
rect 44082 19496 44088 19508
rect 44043 19468 44088 19496
rect 44082 19456 44088 19468
rect 44140 19456 44146 19508
rect 44910 19496 44916 19508
rect 44871 19468 44916 19496
rect 44910 19456 44916 19468
rect 44968 19456 44974 19508
rect 37274 19428 37280 19440
rect 35483 19400 36446 19428
rect 37235 19400 37280 19428
rect 35483 19397 35495 19400
rect 35437 19391 35495 19397
rect 37274 19388 37280 19400
rect 37332 19388 37338 19440
rect 38562 19388 38568 19440
rect 38620 19428 38626 19440
rect 38749 19431 38807 19437
rect 38749 19428 38761 19431
rect 38620 19400 38761 19428
rect 38620 19388 38626 19400
rect 38749 19397 38761 19400
rect 38795 19397 38807 19431
rect 38749 19391 38807 19397
rect 42337 19431 42395 19437
rect 42337 19397 42349 19431
rect 42383 19428 42395 19431
rect 43714 19428 43720 19440
rect 42383 19400 43720 19428
rect 42383 19397 42395 19400
rect 42337 19391 42395 19397
rect 43714 19388 43720 19400
rect 43772 19388 43778 19440
rect 36906 19360 36912 19372
rect 33980 19332 36912 19360
rect 36906 19320 36912 19332
rect 36964 19360 36970 19372
rect 39482 19360 39488 19372
rect 36964 19332 39488 19360
rect 36964 19320 36970 19332
rect 39482 19320 39488 19332
rect 39540 19360 39546 19372
rect 41141 19363 41199 19369
rect 41141 19360 41153 19363
rect 39540 19332 41153 19360
rect 39540 19320 39546 19332
rect 20844 19295 20902 19301
rect 20844 19292 20856 19295
rect 20128 19264 20856 19292
rect 20128 19252 20134 19264
rect 20844 19261 20856 19264
rect 20890 19261 20902 19295
rect 20844 19255 20902 19261
rect 21634 19252 21640 19304
rect 21692 19292 21698 19304
rect 22002 19292 22008 19304
rect 21692 19264 22008 19292
rect 21692 19252 21698 19264
rect 22002 19252 22008 19264
rect 22060 19252 22066 19304
rect 27157 19295 27215 19301
rect 27157 19261 27169 19295
rect 27203 19292 27215 19295
rect 27890 19292 27896 19304
rect 27203 19264 27896 19292
rect 27203 19261 27215 19264
rect 27157 19255 27215 19261
rect 27890 19252 27896 19264
rect 27948 19252 27954 19304
rect 29822 19292 29828 19304
rect 29783 19264 29828 19292
rect 29822 19252 29828 19264
rect 29880 19252 29886 19304
rect 31754 19252 31760 19304
rect 31812 19292 31818 19304
rect 32252 19295 32310 19301
rect 32252 19292 32264 19295
rect 31812 19264 32264 19292
rect 31812 19252 31818 19264
rect 32252 19261 32264 19264
rect 32298 19292 32310 19295
rect 33134 19292 33140 19304
rect 32298 19264 33140 19292
rect 32298 19261 32310 19264
rect 32252 19255 32310 19261
rect 33134 19252 33140 19264
rect 33192 19252 33198 19304
rect 34952 19295 35010 19301
rect 34952 19261 34964 19295
rect 34998 19292 35010 19295
rect 35161 19295 35219 19301
rect 35161 19292 35173 19295
rect 34998 19264 35173 19292
rect 34998 19261 35010 19264
rect 34952 19255 35010 19261
rect 35161 19261 35173 19264
rect 35207 19261 35219 19295
rect 35161 19255 35219 19261
rect 38562 19252 38568 19304
rect 38620 19292 38626 19304
rect 38841 19295 38899 19301
rect 38841 19292 38853 19295
rect 38620 19264 38853 19292
rect 38620 19252 38626 19264
rect 38841 19261 38853 19264
rect 38887 19261 38899 19295
rect 38841 19255 38899 19261
rect 39301 19295 39359 19301
rect 39301 19261 39313 19295
rect 39347 19261 39359 19295
rect 39301 19255 39359 19261
rect 39577 19295 39635 19301
rect 39577 19261 39589 19295
rect 39623 19292 39635 19295
rect 40126 19292 40132 19304
rect 39623 19264 40132 19292
rect 39623 19261 39635 19264
rect 39577 19255 39635 19261
rect 19245 19227 19303 19233
rect 19245 19193 19257 19227
rect 19291 19193 19303 19227
rect 19536 19224 19564 19252
rect 20257 19227 20315 19233
rect 20257 19224 20269 19227
rect 19536 19196 20269 19224
rect 19245 19187 19303 19193
rect 20257 19193 20269 19196
rect 20303 19224 20315 19227
rect 21174 19224 21180 19236
rect 20303 19196 21180 19224
rect 20303 19193 20315 19196
rect 20257 19187 20315 19193
rect 13078 19156 13084 19168
rect 10744 19128 11008 19156
rect 13039 19128 13084 19156
rect 10744 19116 10750 19128
rect 13078 19116 13084 19128
rect 13136 19156 13142 19168
rect 13262 19156 13268 19168
rect 13136 19128 13268 19156
rect 13136 19116 13142 19128
rect 13262 19116 13268 19128
rect 13320 19156 13326 19168
rect 13449 19159 13507 19165
rect 13449 19156 13461 19159
rect 13320 19128 13461 19156
rect 13320 19116 13326 19128
rect 13449 19125 13461 19128
rect 13495 19125 13507 19159
rect 13449 19119 13507 19125
rect 13630 19116 13636 19168
rect 13688 19116 13694 19168
rect 17770 19156 17776 19168
rect 17731 19128 17776 19156
rect 17770 19116 17776 19128
rect 17828 19116 17834 19168
rect 18782 19156 18788 19168
rect 18743 19128 18788 19156
rect 18782 19116 18788 19128
rect 18840 19116 18846 19168
rect 19058 19116 19064 19168
rect 19116 19156 19122 19168
rect 19260 19156 19288 19187
rect 21174 19184 21180 19196
rect 21232 19224 21238 19236
rect 21269 19227 21327 19233
rect 21269 19224 21281 19227
rect 21232 19196 21281 19224
rect 21232 19184 21238 19196
rect 21269 19193 21281 19196
rect 21315 19224 21327 19227
rect 21315 19196 23520 19224
rect 21315 19193 21327 19196
rect 21269 19187 21327 19193
rect 22186 19156 22192 19168
rect 19116 19128 19288 19156
rect 22147 19128 22192 19156
rect 19116 19116 19122 19128
rect 22186 19116 22192 19128
rect 22244 19116 22250 19168
rect 23382 19156 23388 19168
rect 23343 19128 23388 19156
rect 23382 19116 23388 19128
rect 23440 19116 23446 19168
rect 23492 19156 23520 19196
rect 23566 19184 23572 19236
rect 23624 19224 23630 19236
rect 23845 19227 23903 19233
rect 23845 19224 23857 19227
rect 23624 19196 23857 19224
rect 23624 19184 23630 19196
rect 23845 19193 23857 19196
rect 23891 19193 23903 19227
rect 24394 19224 24400 19236
rect 24355 19196 24400 19224
rect 23845 19187 23903 19193
rect 24394 19184 24400 19196
rect 24452 19184 24458 19236
rect 25406 19224 25412 19236
rect 25367 19196 25412 19224
rect 25406 19184 25412 19196
rect 25464 19184 25470 19236
rect 25498 19184 25504 19236
rect 25556 19224 25562 19236
rect 30147 19227 30205 19233
rect 25556 19196 25601 19224
rect 25556 19184 25562 19196
rect 30147 19193 30159 19227
rect 30193 19193 30205 19227
rect 30147 19187 30205 19193
rect 32355 19227 32413 19233
rect 32355 19193 32367 19227
rect 32401 19224 32413 19227
rect 32858 19224 32864 19236
rect 32401 19196 32864 19224
rect 32401 19193 32413 19196
rect 32355 19187 32413 19193
rect 26878 19156 26884 19168
rect 23492 19128 26884 19156
rect 26878 19116 26884 19128
rect 26936 19116 26942 19168
rect 27430 19116 27436 19168
rect 27488 19156 27494 19168
rect 27525 19159 27583 19165
rect 27525 19156 27537 19159
rect 27488 19128 27537 19156
rect 27488 19116 27494 19128
rect 27525 19125 27537 19128
rect 27571 19125 27583 19159
rect 27525 19119 27583 19125
rect 29733 19159 29791 19165
rect 29733 19125 29745 19159
rect 29779 19156 29791 19159
rect 29914 19156 29920 19168
rect 29779 19128 29920 19156
rect 29779 19125 29791 19128
rect 29733 19119 29791 19125
rect 29914 19116 29920 19128
rect 29972 19156 29978 19168
rect 30162 19156 30190 19187
rect 32858 19184 32864 19196
rect 32916 19224 32922 19236
rect 33321 19227 33379 19233
rect 33321 19224 33333 19227
rect 32916 19196 33333 19224
rect 32916 19184 32922 19196
rect 33321 19193 33333 19196
rect 33367 19193 33379 19227
rect 33321 19187 33379 19193
rect 33413 19227 33471 19233
rect 33413 19193 33425 19227
rect 33459 19224 33471 19227
rect 33686 19224 33692 19236
rect 33459 19196 33692 19224
rect 33459 19193 33471 19196
rect 33413 19187 33471 19193
rect 33686 19184 33692 19196
rect 33744 19184 33750 19236
rect 36722 19224 36728 19236
rect 36683 19196 36728 19224
rect 36722 19184 36728 19196
rect 36780 19184 36786 19236
rect 36817 19227 36875 19233
rect 36817 19193 36829 19227
rect 36863 19193 36875 19227
rect 36817 19187 36875 19193
rect 30558 19156 30564 19168
rect 29972 19128 30564 19156
rect 29972 19116 29978 19128
rect 30558 19116 30564 19128
rect 30616 19116 30622 19168
rect 30745 19159 30803 19165
rect 30745 19125 30757 19159
rect 30791 19156 30803 19159
rect 30834 19156 30840 19168
rect 30791 19128 30840 19156
rect 30791 19125 30803 19128
rect 30745 19119 30803 19125
rect 30834 19116 30840 19128
rect 30892 19116 30898 19168
rect 34698 19116 34704 19168
rect 34756 19156 34762 19168
rect 35023 19159 35081 19165
rect 35023 19156 35035 19159
rect 34756 19128 35035 19156
rect 34756 19116 34762 19128
rect 35023 19125 35035 19128
rect 35069 19125 35081 19159
rect 35023 19119 35081 19125
rect 36541 19159 36599 19165
rect 36541 19125 36553 19159
rect 36587 19156 36599 19159
rect 36832 19156 36860 19187
rect 37090 19184 37096 19236
rect 37148 19224 37154 19236
rect 38289 19227 38347 19233
rect 38289 19224 38301 19227
rect 37148 19196 38301 19224
rect 37148 19184 37154 19196
rect 38289 19193 38301 19196
rect 38335 19224 38347 19227
rect 38470 19224 38476 19236
rect 38335 19196 38476 19224
rect 38335 19193 38347 19196
rect 38289 19187 38347 19193
rect 38470 19184 38476 19196
rect 38528 19224 38534 19236
rect 39316 19224 39344 19255
rect 40126 19252 40132 19264
rect 40184 19252 40190 19304
rect 40731 19301 40759 19332
rect 41141 19329 41153 19332
rect 41187 19329 41199 19363
rect 41782 19360 41788 19372
rect 41743 19332 41788 19360
rect 41141 19323 41199 19329
rect 41782 19320 41788 19332
rect 41840 19360 41846 19372
rect 41840 19334 42656 19360
rect 41840 19332 42748 19334
rect 41840 19320 41846 19332
rect 42628 19306 42748 19332
rect 40716 19295 40774 19301
rect 40716 19261 40728 19295
rect 40762 19261 40774 19295
rect 40716 19255 40774 19261
rect 38528 19196 39344 19224
rect 41877 19227 41935 19233
rect 38528 19184 38534 19196
rect 41877 19193 41889 19227
rect 41923 19193 41935 19227
rect 42720 19224 42748 19306
rect 43308 19295 43366 19301
rect 43308 19261 43320 19295
rect 43354 19292 43366 19295
rect 43354 19264 43530 19292
rect 43354 19261 43366 19264
rect 43308 19255 43366 19261
rect 43395 19227 43453 19233
rect 43395 19224 43407 19227
rect 42720 19196 43407 19224
rect 41877 19187 41935 19193
rect 43395 19193 43407 19196
rect 43441 19193 43453 19227
rect 43395 19187 43453 19193
rect 37918 19156 37924 19168
rect 36587 19128 37924 19156
rect 36587 19125 36599 19128
rect 36541 19119 36599 19125
rect 37918 19116 37924 19128
rect 37976 19116 37982 19168
rect 41598 19156 41604 19168
rect 41559 19128 41604 19156
rect 41598 19116 41604 19128
rect 41656 19156 41662 19168
rect 41892 19156 41920 19187
rect 41656 19128 41920 19156
rect 41656 19116 41662 19128
rect 42518 19116 42524 19168
rect 42576 19156 42582 19168
rect 43502 19156 43530 19264
rect 43717 19159 43775 19165
rect 43717 19156 43729 19159
rect 42576 19128 43729 19156
rect 42576 19116 42582 19128
rect 43717 19125 43729 19128
rect 43763 19125 43775 19159
rect 43717 19119 43775 19125
rect 1104 19066 48852 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 48852 19066
rect 1104 18992 48852 19014
rect 10962 18952 10968 18964
rect 10923 18924 10968 18952
rect 10962 18912 10968 18924
rect 11020 18912 11026 18964
rect 11238 18952 11244 18964
rect 11199 18924 11244 18952
rect 11238 18912 11244 18924
rect 11296 18912 11302 18964
rect 13170 18952 13176 18964
rect 13131 18924 13176 18952
rect 13170 18912 13176 18924
rect 13228 18912 13234 18964
rect 13814 18952 13820 18964
rect 13556 18924 13820 18952
rect 12713 18887 12771 18893
rect 12713 18853 12725 18887
rect 12759 18884 12771 18887
rect 13078 18884 13084 18896
rect 12759 18856 13084 18884
rect 12759 18853 12771 18856
rect 12713 18847 12771 18853
rect 13078 18844 13084 18856
rect 13136 18884 13142 18896
rect 13556 18884 13584 18924
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 18966 18912 18972 18964
rect 19024 18952 19030 18964
rect 19153 18955 19211 18961
rect 19153 18952 19165 18955
rect 19024 18924 19165 18952
rect 19024 18912 19030 18924
rect 19153 18921 19165 18924
rect 19199 18952 19211 18955
rect 19334 18952 19340 18964
rect 19199 18924 19340 18952
rect 19199 18921 19211 18924
rect 19153 18915 19211 18921
rect 19334 18912 19340 18924
rect 19392 18912 19398 18964
rect 20714 18952 20720 18964
rect 20675 18924 20720 18952
rect 20714 18912 20720 18924
rect 20772 18912 20778 18964
rect 20898 18912 20904 18964
rect 20956 18952 20962 18964
rect 21085 18955 21143 18961
rect 21085 18952 21097 18955
rect 20956 18924 21097 18952
rect 20956 18912 20962 18924
rect 21085 18921 21097 18924
rect 21131 18921 21143 18955
rect 22002 18952 22008 18964
rect 21963 18924 22008 18952
rect 21085 18915 21143 18921
rect 22002 18912 22008 18924
rect 22060 18912 22066 18964
rect 23658 18952 23664 18964
rect 23619 18924 23664 18952
rect 23658 18912 23664 18924
rect 23716 18912 23722 18964
rect 25406 18912 25412 18964
rect 25464 18952 25470 18964
rect 25685 18955 25743 18961
rect 25685 18952 25697 18955
rect 25464 18924 25697 18952
rect 25464 18912 25470 18924
rect 25685 18921 25697 18924
rect 25731 18921 25743 18955
rect 32858 18952 32864 18964
rect 32819 18924 32864 18952
rect 25685 18915 25743 18921
rect 32858 18912 32864 18924
rect 32916 18912 32922 18964
rect 33778 18912 33784 18964
rect 33836 18952 33842 18964
rect 33836 18924 35848 18952
rect 33836 18912 33842 18924
rect 13722 18884 13728 18896
rect 13136 18856 13584 18884
rect 13683 18856 13728 18884
rect 13136 18844 13142 18856
rect 13722 18844 13728 18856
rect 13780 18844 13786 18896
rect 14274 18884 14280 18896
rect 14235 18856 14280 18884
rect 14274 18844 14280 18856
rect 14332 18844 14338 18896
rect 18598 18844 18604 18896
rect 18656 18884 18662 18896
rect 18785 18887 18843 18893
rect 18785 18884 18797 18887
rect 18656 18856 18797 18884
rect 18656 18844 18662 18856
rect 18785 18853 18797 18856
rect 18831 18884 18843 18887
rect 19242 18884 19248 18896
rect 18831 18856 19248 18884
rect 18831 18853 18843 18856
rect 18785 18847 18843 18853
rect 19242 18844 19248 18856
rect 19300 18844 19306 18896
rect 22020 18884 22048 18912
rect 21422 18856 22048 18884
rect 23109 18887 23167 18893
rect 21422 18828 21450 18856
rect 23109 18853 23121 18887
rect 23155 18884 23167 18887
rect 23382 18884 23388 18896
rect 23155 18856 23388 18884
rect 23155 18853 23167 18856
rect 23109 18847 23167 18853
rect 23382 18844 23388 18856
rect 23440 18884 23446 18896
rect 23566 18884 23572 18896
rect 23440 18856 23572 18884
rect 23440 18844 23446 18856
rect 23566 18844 23572 18856
rect 23624 18844 23630 18896
rect 29641 18887 29699 18893
rect 29641 18853 29653 18887
rect 29687 18884 29699 18887
rect 29822 18884 29828 18896
rect 29687 18856 29828 18884
rect 29687 18853 29699 18856
rect 29641 18847 29699 18853
rect 29822 18844 29828 18856
rect 29880 18884 29886 18896
rect 29917 18887 29975 18893
rect 29917 18884 29929 18887
rect 29880 18856 29929 18884
rect 29880 18844 29886 18856
rect 29917 18853 29929 18856
rect 29963 18853 29975 18887
rect 29917 18847 29975 18853
rect 30653 18887 30711 18893
rect 30653 18853 30665 18887
rect 30699 18884 30711 18887
rect 30834 18884 30840 18896
rect 30699 18856 30840 18884
rect 30699 18853 30711 18856
rect 30653 18847 30711 18853
rect 30834 18844 30840 18856
rect 30892 18844 30898 18896
rect 31202 18884 31208 18896
rect 31163 18856 31208 18884
rect 31202 18844 31208 18856
rect 31260 18844 31266 18896
rect 33321 18887 33379 18893
rect 33321 18853 33333 18887
rect 33367 18884 33379 18887
rect 33686 18884 33692 18896
rect 33367 18856 33692 18884
rect 33367 18853 33379 18856
rect 33321 18847 33379 18853
rect 33686 18844 33692 18856
rect 33744 18844 33750 18896
rect 34238 18884 34244 18896
rect 34199 18856 34244 18884
rect 34238 18844 34244 18856
rect 34296 18844 34302 18896
rect 34606 18844 34612 18896
rect 34664 18884 34670 18896
rect 35161 18887 35219 18893
rect 35161 18884 35173 18887
rect 34664 18856 35173 18884
rect 34664 18844 34670 18856
rect 35161 18853 35173 18856
rect 35207 18853 35219 18887
rect 35161 18847 35219 18853
rect 35250 18844 35256 18896
rect 35308 18884 35314 18896
rect 35820 18893 35848 18924
rect 38746 18912 38752 18964
rect 38804 18952 38810 18964
rect 39117 18955 39175 18961
rect 39117 18952 39129 18955
rect 38804 18924 39129 18952
rect 38804 18912 38810 18924
rect 39117 18921 39129 18924
rect 39163 18921 39175 18955
rect 40126 18952 40132 18964
rect 40087 18924 40132 18952
rect 39117 18915 39175 18921
rect 40126 18912 40132 18924
rect 40184 18912 40190 18964
rect 40543 18955 40601 18961
rect 40543 18921 40555 18955
rect 40589 18952 40601 18955
rect 41322 18952 41328 18964
rect 40589 18924 41328 18952
rect 40589 18921 40601 18924
rect 40543 18915 40601 18921
rect 41322 18912 41328 18924
rect 41380 18912 41386 18964
rect 35805 18887 35863 18893
rect 35308 18856 35353 18884
rect 35308 18844 35314 18856
rect 35805 18853 35817 18887
rect 35851 18853 35863 18887
rect 35805 18847 35863 18853
rect 37642 18844 37648 18896
rect 37700 18884 37706 18896
rect 38289 18887 38347 18893
rect 38289 18884 38301 18887
rect 37700 18856 38301 18884
rect 37700 18844 37706 18856
rect 38289 18853 38301 18856
rect 38335 18853 38347 18887
rect 41506 18884 41512 18896
rect 41467 18856 41512 18884
rect 38289 18847 38347 18853
rect 41506 18844 41512 18856
rect 41564 18844 41570 18896
rect 41598 18844 41604 18896
rect 41656 18884 41662 18896
rect 41656 18856 41701 18884
rect 41656 18844 41662 18856
rect 10480 18819 10538 18825
rect 10480 18785 10492 18819
rect 10526 18816 10538 18819
rect 10870 18816 10876 18828
rect 10526 18788 10876 18816
rect 10526 18785 10538 18788
rect 10480 18779 10538 18785
rect 10870 18776 10876 18788
rect 10928 18816 10934 18828
rect 11514 18816 11520 18828
rect 10928 18788 11520 18816
rect 10928 18776 10934 18788
rect 11514 18776 11520 18788
rect 11572 18776 11578 18828
rect 12066 18776 12072 18828
rect 12124 18816 12130 18828
rect 12621 18819 12679 18825
rect 12621 18816 12633 18819
rect 12124 18788 12633 18816
rect 12124 18776 12130 18788
rect 12621 18785 12633 18788
rect 12667 18816 12679 18819
rect 12802 18816 12808 18828
rect 12667 18788 12808 18816
rect 12667 18785 12679 18788
rect 12621 18779 12679 18785
rect 12802 18776 12808 18788
rect 12860 18776 12866 18828
rect 15632 18819 15690 18825
rect 15632 18785 15644 18819
rect 15678 18816 15690 18819
rect 15838 18816 15844 18828
rect 15678 18788 15844 18816
rect 15678 18785 15690 18788
rect 15632 18779 15690 18785
rect 15838 18776 15844 18788
rect 15896 18776 15902 18828
rect 17218 18816 17224 18828
rect 17179 18788 17224 18816
rect 17218 18776 17224 18788
rect 17276 18776 17282 18828
rect 17402 18776 17408 18828
rect 17460 18816 17466 18828
rect 18141 18819 18199 18825
rect 18141 18816 18153 18819
rect 17460 18788 18153 18816
rect 17460 18776 17466 18788
rect 18141 18785 18153 18788
rect 18187 18785 18199 18819
rect 21358 18816 21364 18828
rect 21317 18788 21364 18816
rect 18141 18779 18199 18785
rect 21358 18776 21364 18788
rect 21416 18825 21450 18828
rect 21416 18819 21465 18825
rect 21416 18785 21419 18819
rect 21453 18785 21465 18819
rect 21416 18779 21465 18785
rect 21499 18819 21557 18825
rect 21499 18785 21511 18819
rect 21545 18816 21557 18819
rect 22465 18819 22523 18825
rect 22465 18816 22477 18819
rect 21545 18788 22477 18816
rect 21545 18785 21557 18788
rect 21499 18779 21557 18785
rect 22465 18785 22477 18788
rect 22511 18816 22523 18819
rect 23014 18816 23020 18828
rect 22511 18788 23020 18816
rect 22511 18785 22523 18788
rect 22465 18779 22523 18785
rect 21416 18776 21422 18779
rect 23014 18776 23020 18788
rect 23072 18776 23078 18828
rect 24578 18816 24584 18828
rect 23446 18788 24584 18816
rect 13630 18748 13636 18760
rect 13591 18720 13636 18748
rect 13630 18708 13636 18720
rect 13688 18708 13694 18760
rect 16574 18748 16580 18760
rect 16535 18720 16580 18748
rect 16574 18708 16580 18720
rect 16632 18708 16638 18760
rect 19392 18751 19450 18757
rect 19392 18717 19404 18751
rect 19438 18748 19450 18751
rect 19518 18748 19524 18760
rect 19438 18720 19524 18748
rect 19438 18717 19450 18720
rect 19392 18711 19450 18717
rect 19518 18708 19524 18720
rect 19576 18708 19582 18760
rect 19613 18751 19671 18757
rect 19613 18717 19625 18751
rect 19659 18748 19671 18751
rect 19886 18748 19892 18760
rect 19659 18720 19892 18748
rect 19659 18717 19671 18720
rect 19613 18711 19671 18717
rect 19886 18708 19892 18720
rect 19944 18708 19950 18760
rect 19981 18751 20039 18757
rect 19981 18717 19993 18751
rect 20027 18748 20039 18751
rect 20714 18748 20720 18760
rect 20027 18720 20720 18748
rect 20027 18717 20039 18720
rect 19981 18711 20039 18717
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 22186 18708 22192 18760
rect 22244 18748 22250 18760
rect 23446 18748 23474 18788
rect 24578 18776 24584 18788
rect 24636 18776 24642 18828
rect 25409 18819 25467 18825
rect 25409 18785 25421 18819
rect 25455 18816 25467 18819
rect 25498 18816 25504 18828
rect 25455 18788 25504 18816
rect 25455 18785 25467 18788
rect 25409 18779 25467 18785
rect 25498 18776 25504 18788
rect 25556 18776 25562 18828
rect 27062 18816 27068 18828
rect 27023 18788 27068 18816
rect 27062 18776 27068 18788
rect 27120 18776 27126 18828
rect 29178 18816 29184 18828
rect 29139 18788 29184 18816
rect 29178 18776 29184 18788
rect 29236 18776 29242 18828
rect 29457 18819 29515 18825
rect 29457 18785 29469 18819
rect 29503 18816 29515 18819
rect 29730 18816 29736 18828
rect 29503 18788 29736 18816
rect 29503 18785 29515 18788
rect 29457 18779 29515 18785
rect 29730 18776 29736 18788
rect 29788 18776 29794 18828
rect 32033 18819 32091 18825
rect 32033 18785 32045 18819
rect 32079 18816 32091 18819
rect 32122 18816 32128 18828
rect 32079 18788 32128 18816
rect 32079 18785 32091 18788
rect 32033 18779 32091 18785
rect 32122 18776 32128 18788
rect 32180 18776 32186 18828
rect 36684 18819 36742 18825
rect 36684 18785 36696 18819
rect 36730 18816 36742 18819
rect 36906 18816 36912 18828
rect 36730 18788 36912 18816
rect 36730 18785 36742 18788
rect 36684 18779 36742 18785
rect 36906 18776 36912 18788
rect 36964 18776 36970 18828
rect 40218 18776 40224 18828
rect 40276 18816 40282 18828
rect 40440 18819 40498 18825
rect 40440 18816 40452 18819
rect 40276 18788 40452 18816
rect 40276 18776 40282 18788
rect 40440 18785 40452 18788
rect 40486 18785 40498 18819
rect 40440 18779 40498 18785
rect 43416 18819 43474 18825
rect 43416 18785 43428 18819
rect 43462 18816 43474 18819
rect 43990 18816 43996 18828
rect 43462 18788 43996 18816
rect 43462 18785 43474 18788
rect 43416 18779 43474 18785
rect 43990 18776 43996 18788
rect 44048 18776 44054 18828
rect 22244 18720 23474 18748
rect 24673 18751 24731 18757
rect 22244 18708 22250 18720
rect 24673 18717 24685 18751
rect 24719 18748 24731 18751
rect 24854 18748 24860 18760
rect 24719 18720 24860 18748
rect 24719 18717 24731 18720
rect 24673 18711 24731 18717
rect 24854 18708 24860 18720
rect 24912 18708 24918 18760
rect 27709 18751 27767 18757
rect 27709 18717 27721 18751
rect 27755 18748 27767 18751
rect 28534 18748 28540 18760
rect 27755 18720 28540 18748
rect 27755 18717 27767 18720
rect 27709 18711 27767 18717
rect 28534 18708 28540 18720
rect 28592 18708 28598 18760
rect 30377 18751 30435 18757
rect 30377 18717 30389 18751
rect 30423 18748 30435 18751
rect 30561 18751 30619 18757
rect 30561 18748 30573 18751
rect 30423 18720 30573 18748
rect 30423 18717 30435 18720
rect 30377 18711 30435 18717
rect 30561 18717 30573 18720
rect 30607 18748 30619 18751
rect 32263 18751 32321 18757
rect 32263 18748 32275 18751
rect 30607 18720 32275 18748
rect 30607 18717 30619 18720
rect 30561 18711 30619 18717
rect 32263 18717 32275 18720
rect 32309 18717 32321 18751
rect 33594 18748 33600 18760
rect 33507 18720 33600 18748
rect 32263 18711 32321 18717
rect 33594 18708 33600 18720
rect 33652 18748 33658 18760
rect 34698 18748 34704 18760
rect 33652 18720 34704 18748
rect 33652 18708 33658 18720
rect 34698 18708 34704 18720
rect 34756 18708 34762 18760
rect 36771 18751 36829 18757
rect 36771 18717 36783 18751
rect 36817 18748 36829 18751
rect 38197 18751 38255 18757
rect 38197 18748 38209 18751
rect 36817 18720 38209 18748
rect 36817 18717 36829 18720
rect 36771 18711 36829 18717
rect 38197 18717 38209 18720
rect 38243 18748 38255 18751
rect 38838 18748 38844 18760
rect 38243 18720 38844 18748
rect 38243 18717 38255 18720
rect 38197 18711 38255 18717
rect 38838 18708 38844 18720
rect 38896 18708 38902 18760
rect 40586 18708 40592 18760
rect 40644 18748 40650 18760
rect 41785 18751 41843 18757
rect 41785 18748 41797 18751
rect 40644 18720 41797 18748
rect 40644 18708 40650 18720
rect 41785 18717 41797 18720
rect 41831 18748 41843 18751
rect 44174 18748 44180 18760
rect 41831 18720 44180 18748
rect 41831 18717 41843 18720
rect 41785 18711 41843 18717
rect 44174 18708 44180 18720
rect 44232 18708 44238 18760
rect 8386 18640 8392 18692
rect 8444 18680 8450 18692
rect 9398 18680 9404 18692
rect 8444 18652 9404 18680
rect 8444 18640 8450 18652
rect 9398 18640 9404 18652
rect 9456 18640 9462 18692
rect 11054 18640 11060 18692
rect 11112 18680 11118 18692
rect 14274 18680 14280 18692
rect 11112 18652 14280 18680
rect 11112 18640 11118 18652
rect 14274 18640 14280 18652
rect 14332 18640 14338 18692
rect 16758 18640 16764 18692
rect 16816 18680 16822 18692
rect 17954 18680 17960 18692
rect 16816 18652 17960 18680
rect 16816 18640 16822 18652
rect 17954 18640 17960 18652
rect 18012 18640 18018 18692
rect 33106 18652 34100 18680
rect 8754 18572 8760 18624
rect 8812 18612 8818 18624
rect 10551 18615 10609 18621
rect 10551 18612 10563 18615
rect 8812 18584 10563 18612
rect 8812 18572 8818 18584
rect 10551 18581 10563 18584
rect 10597 18581 10609 18615
rect 10551 18575 10609 18581
rect 15703 18615 15761 18621
rect 15703 18581 15715 18615
rect 15749 18612 15761 18615
rect 16482 18612 16488 18624
rect 15749 18584 16488 18612
rect 15749 18581 15761 18584
rect 15703 18575 15761 18581
rect 16482 18572 16488 18584
rect 16540 18572 16546 18624
rect 18322 18612 18328 18624
rect 18283 18584 18328 18612
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 19518 18612 19524 18624
rect 19479 18584 19524 18612
rect 19518 18572 19524 18584
rect 19576 18572 19582 18624
rect 25038 18612 25044 18624
rect 24999 18584 25044 18612
rect 25038 18572 25044 18584
rect 25096 18572 25102 18624
rect 26694 18612 26700 18624
rect 26655 18584 26700 18612
rect 26694 18572 26700 18584
rect 26752 18572 26758 18624
rect 31478 18572 31484 18624
rect 31536 18612 31542 18624
rect 33106 18612 33134 18652
rect 31536 18584 33134 18612
rect 34072 18612 34100 18652
rect 36078 18640 36084 18692
rect 36136 18680 36142 18692
rect 38562 18680 38568 18692
rect 36136 18652 38568 18680
rect 36136 18640 36142 18652
rect 38562 18640 38568 18652
rect 38620 18640 38626 18692
rect 38749 18683 38807 18689
rect 38749 18649 38761 18683
rect 38795 18680 38807 18683
rect 39206 18680 39212 18692
rect 38795 18652 39212 18680
rect 38795 18649 38807 18652
rect 38749 18643 38807 18649
rect 39206 18640 39212 18652
rect 39264 18640 39270 18692
rect 36722 18612 36728 18624
rect 34072 18584 36728 18612
rect 31536 18572 31542 18584
rect 36722 18572 36728 18584
rect 36780 18612 36786 18624
rect 37093 18615 37151 18621
rect 37093 18612 37105 18615
rect 36780 18584 37105 18612
rect 36780 18572 36786 18584
rect 37093 18581 37105 18584
rect 37139 18581 37151 18615
rect 43070 18612 43076 18624
rect 42983 18584 43076 18612
rect 37093 18575 37151 18581
rect 43070 18572 43076 18584
rect 43128 18612 43134 18624
rect 43487 18615 43545 18621
rect 43487 18612 43499 18615
rect 43128 18584 43499 18612
rect 43128 18572 43134 18584
rect 43487 18581 43499 18584
rect 43533 18581 43545 18615
rect 43487 18575 43545 18581
rect 1104 18522 48852 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 48852 18522
rect 1104 18448 48852 18470
rect 10870 18408 10876 18420
rect 10831 18380 10876 18408
rect 10870 18368 10876 18380
rect 10928 18368 10934 18420
rect 12066 18408 12072 18420
rect 12027 18380 12072 18408
rect 12066 18368 12072 18380
rect 12124 18368 12130 18420
rect 13630 18368 13636 18420
rect 13688 18408 13694 18420
rect 13688 18380 14412 18408
rect 13688 18368 13694 18380
rect 12805 18343 12863 18349
rect 12805 18309 12817 18343
rect 12851 18340 12863 18343
rect 13078 18340 13084 18352
rect 12851 18312 13084 18340
rect 12851 18309 12863 18312
rect 12805 18303 12863 18309
rect 13078 18300 13084 18312
rect 13136 18340 13142 18352
rect 13722 18340 13728 18352
rect 13136 18312 13728 18340
rect 13136 18300 13142 18312
rect 13722 18300 13728 18312
rect 13780 18300 13786 18352
rect 13354 18272 13360 18284
rect 13315 18244 13360 18272
rect 13354 18232 13360 18244
rect 13412 18232 13418 18284
rect 9677 18207 9735 18213
rect 9677 18173 9689 18207
rect 9723 18204 9735 18207
rect 10042 18204 10048 18216
rect 9723 18176 10048 18204
rect 9723 18173 9735 18176
rect 9677 18167 9735 18173
rect 10042 18164 10048 18176
rect 10100 18164 10106 18216
rect 10318 18204 10324 18216
rect 10279 18176 10324 18204
rect 10318 18164 10324 18176
rect 10376 18164 10382 18216
rect 11368 18207 11426 18213
rect 11368 18204 11380 18207
rect 11164 18176 11380 18204
rect 10502 18136 10508 18148
rect 10463 18108 10508 18136
rect 10502 18096 10508 18108
rect 10560 18096 10566 18148
rect 9214 18068 9220 18080
rect 9175 18040 9220 18068
rect 9214 18028 9220 18040
rect 9272 18028 9278 18080
rect 10870 18028 10876 18080
rect 10928 18068 10934 18080
rect 11164 18077 11192 18176
rect 11368 18173 11380 18176
rect 11414 18173 11426 18207
rect 11368 18167 11426 18173
rect 12986 18136 12992 18148
rect 12947 18108 12992 18136
rect 12986 18096 12992 18108
rect 13044 18096 13050 18148
rect 13078 18096 13084 18148
rect 13136 18136 13142 18148
rect 14384 18145 14412 18380
rect 17218 18368 17224 18420
rect 17276 18408 17282 18420
rect 17497 18411 17555 18417
rect 17497 18408 17509 18411
rect 17276 18380 17509 18408
rect 17276 18368 17282 18380
rect 17497 18377 17509 18380
rect 17543 18408 17555 18411
rect 18322 18408 18328 18420
rect 17543 18380 18328 18408
rect 17543 18377 17555 18380
rect 17497 18371 17555 18377
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 18598 18408 18604 18420
rect 18559 18380 18604 18408
rect 18598 18368 18604 18380
rect 18656 18368 18662 18420
rect 18966 18408 18972 18420
rect 18927 18380 18972 18408
rect 18966 18368 18972 18380
rect 19024 18368 19030 18420
rect 19337 18411 19395 18417
rect 19337 18377 19349 18411
rect 19383 18408 19395 18411
rect 19886 18408 19892 18420
rect 19383 18380 19892 18408
rect 19383 18377 19395 18380
rect 19337 18371 19395 18377
rect 19886 18368 19892 18380
rect 19944 18368 19950 18420
rect 21358 18408 21364 18420
rect 21319 18380 21364 18408
rect 21358 18368 21364 18380
rect 21416 18368 21422 18420
rect 23014 18408 23020 18420
rect 22975 18380 23020 18408
rect 23014 18368 23020 18380
rect 23072 18368 23078 18420
rect 23477 18411 23535 18417
rect 23477 18377 23489 18411
rect 23523 18408 23535 18411
rect 23842 18408 23848 18420
rect 23523 18380 23848 18408
rect 23523 18377 23535 18380
rect 23477 18371 23535 18377
rect 23842 18368 23848 18380
rect 23900 18368 23906 18420
rect 24578 18368 24584 18420
rect 24636 18408 24642 18420
rect 24673 18411 24731 18417
rect 24673 18408 24685 18411
rect 24636 18380 24685 18408
rect 24636 18368 24642 18380
rect 24673 18377 24685 18380
rect 24719 18377 24731 18411
rect 27062 18408 27068 18420
rect 27023 18380 27068 18408
rect 24673 18371 24731 18377
rect 27062 18368 27068 18380
rect 27120 18368 27126 18420
rect 28997 18411 29055 18417
rect 28997 18377 29009 18411
rect 29043 18408 29055 18411
rect 29178 18408 29184 18420
rect 29043 18380 29184 18408
rect 29043 18377 29055 18380
rect 28997 18371 29055 18377
rect 29178 18368 29184 18380
rect 29236 18368 29242 18420
rect 29730 18408 29736 18420
rect 29691 18380 29736 18408
rect 29730 18368 29736 18380
rect 29788 18368 29794 18420
rect 33045 18411 33103 18417
rect 33045 18377 33057 18411
rect 33091 18408 33103 18411
rect 33594 18408 33600 18420
rect 33091 18380 33600 18408
rect 33091 18377 33103 18380
rect 33045 18371 33103 18377
rect 33594 18368 33600 18380
rect 33652 18368 33658 18420
rect 33686 18368 33692 18420
rect 33744 18408 33750 18420
rect 34057 18411 34115 18417
rect 34057 18408 34069 18411
rect 33744 18380 34069 18408
rect 33744 18368 33750 18380
rect 34057 18377 34069 18380
rect 34103 18408 34115 18411
rect 35250 18408 35256 18420
rect 34103 18380 35256 18408
rect 34103 18377 34115 18380
rect 34057 18371 34115 18377
rect 35250 18368 35256 18380
rect 35308 18408 35314 18420
rect 35713 18411 35771 18417
rect 35713 18408 35725 18411
rect 35308 18380 35725 18408
rect 35308 18368 35314 18380
rect 35713 18377 35725 18380
rect 35759 18377 35771 18411
rect 35713 18371 35771 18377
rect 36449 18411 36507 18417
rect 36449 18377 36461 18411
rect 36495 18408 36507 18411
rect 36906 18408 36912 18420
rect 36495 18380 36912 18408
rect 36495 18377 36507 18380
rect 36449 18371 36507 18377
rect 36906 18368 36912 18380
rect 36964 18368 36970 18420
rect 37642 18408 37648 18420
rect 37603 18380 37648 18408
rect 37642 18368 37648 18380
rect 37700 18368 37706 18420
rect 39574 18368 39580 18420
rect 39632 18408 39638 18420
rect 39853 18411 39911 18417
rect 39853 18408 39865 18411
rect 39632 18380 39865 18408
rect 39632 18368 39638 18380
rect 39853 18377 39865 18380
rect 39899 18408 39911 18411
rect 40586 18408 40592 18420
rect 39899 18380 40592 18408
rect 39899 18377 39911 18380
rect 39853 18371 39911 18377
rect 40586 18368 40592 18380
rect 40644 18368 40650 18420
rect 41506 18368 41512 18420
rect 41564 18408 41570 18420
rect 41877 18411 41935 18417
rect 41877 18408 41889 18411
rect 41564 18380 41889 18408
rect 41564 18368 41570 18380
rect 41877 18377 41889 18380
rect 41923 18377 41935 18411
rect 43990 18408 43996 18420
rect 41877 18371 41935 18377
rect 42766 18380 43996 18408
rect 17402 18300 17408 18352
rect 17460 18340 17466 18352
rect 17773 18343 17831 18349
rect 17773 18340 17785 18343
rect 17460 18312 17785 18340
rect 17460 18300 17466 18312
rect 17773 18309 17785 18312
rect 17819 18309 17831 18343
rect 17773 18303 17831 18309
rect 23658 18300 23664 18352
rect 23716 18340 23722 18352
rect 25501 18343 25559 18349
rect 23716 18312 23796 18340
rect 23716 18300 23722 18312
rect 16482 18272 16488 18284
rect 16443 18244 16488 18272
rect 16482 18232 16488 18244
rect 16540 18232 16546 18284
rect 20438 18272 20444 18284
rect 20399 18244 20444 18272
rect 20438 18232 20444 18244
rect 20496 18232 20502 18284
rect 23768 18281 23796 18312
rect 25501 18309 25513 18343
rect 25547 18340 25559 18343
rect 25547 18312 26372 18340
rect 25547 18309 25559 18312
rect 25501 18303 25559 18309
rect 23753 18275 23811 18281
rect 23753 18241 23765 18275
rect 23799 18241 23811 18275
rect 24210 18272 24216 18284
rect 24171 18244 24216 18272
rect 23753 18235 23811 18241
rect 24210 18232 24216 18244
rect 24268 18232 24274 18284
rect 25406 18232 25412 18284
rect 25464 18272 25470 18284
rect 25866 18272 25872 18284
rect 25464 18244 25872 18272
rect 25464 18232 25470 18244
rect 25866 18232 25872 18244
rect 25924 18272 25930 18284
rect 25961 18275 26019 18281
rect 25961 18272 25973 18275
rect 25924 18244 25973 18272
rect 25924 18232 25930 18244
rect 25961 18241 25973 18244
rect 26007 18241 26019 18275
rect 25961 18235 26019 18241
rect 14458 18164 14464 18216
rect 14516 18204 14522 18216
rect 14620 18207 14678 18213
rect 14620 18204 14632 18207
rect 14516 18176 14632 18204
rect 14516 18164 14522 18176
rect 14620 18173 14632 18176
rect 14666 18204 14678 18207
rect 15102 18204 15108 18216
rect 14666 18176 15108 18204
rect 14666 18173 14678 18176
rect 14620 18167 14678 18173
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 17954 18204 17960 18216
rect 17915 18176 17960 18204
rect 17954 18164 17960 18176
rect 18012 18164 18018 18216
rect 18230 18164 18236 18216
rect 18288 18204 18294 18216
rect 18782 18204 18788 18216
rect 18288 18176 18788 18204
rect 18288 18164 18294 18176
rect 18782 18164 18788 18176
rect 18840 18204 18846 18216
rect 19518 18204 19524 18216
rect 18840 18176 19524 18204
rect 18840 18164 18846 18176
rect 19518 18164 19524 18176
rect 19576 18204 19582 18216
rect 19613 18207 19671 18213
rect 19613 18204 19625 18207
rect 19576 18176 19625 18204
rect 19576 18164 19582 18176
rect 19613 18173 19625 18176
rect 19659 18173 19671 18207
rect 19978 18204 19984 18216
rect 19939 18176 19984 18204
rect 19613 18167 19671 18173
rect 19978 18164 19984 18176
rect 20036 18164 20042 18216
rect 20254 18164 20260 18216
rect 20312 18204 20318 18216
rect 20349 18207 20407 18213
rect 20349 18204 20361 18207
rect 20312 18176 20361 18204
rect 20312 18164 20318 18176
rect 20349 18173 20361 18176
rect 20395 18173 20407 18207
rect 20349 18167 20407 18173
rect 14369 18139 14427 18145
rect 13136 18108 13181 18136
rect 13136 18096 13142 18108
rect 14369 18105 14381 18139
rect 14415 18136 14427 18139
rect 16022 18136 16028 18148
rect 14415 18108 16028 18136
rect 14415 18105 14427 18108
rect 14369 18099 14427 18105
rect 16022 18096 16028 18108
rect 16080 18096 16086 18148
rect 16301 18139 16359 18145
rect 16301 18105 16313 18139
rect 16347 18136 16359 18139
rect 16574 18136 16580 18148
rect 16347 18108 16580 18136
rect 16347 18105 16359 18108
rect 16301 18099 16359 18105
rect 16574 18096 16580 18108
rect 16632 18096 16638 18148
rect 17126 18136 17132 18148
rect 17087 18108 17132 18136
rect 17126 18096 17132 18108
rect 17184 18096 17190 18148
rect 22097 18139 22155 18145
rect 22097 18105 22109 18139
rect 22143 18105 22155 18139
rect 22097 18099 22155 18105
rect 11149 18071 11207 18077
rect 11149 18068 11161 18071
rect 10928 18040 11161 18068
rect 10928 18028 10934 18040
rect 11149 18037 11161 18040
rect 11195 18037 11207 18071
rect 11149 18031 11207 18037
rect 11471 18071 11529 18077
rect 11471 18037 11483 18071
rect 11517 18068 11529 18071
rect 11882 18068 11888 18080
rect 11517 18040 11888 18068
rect 11517 18037 11529 18040
rect 11471 18031 11529 18037
rect 11882 18028 11888 18040
rect 11940 18028 11946 18080
rect 13722 18028 13728 18080
rect 13780 18068 13786 18080
rect 13909 18071 13967 18077
rect 13909 18068 13921 18071
rect 13780 18040 13921 18068
rect 13780 18028 13786 18040
rect 13909 18037 13921 18040
rect 13955 18037 13967 18071
rect 13909 18031 13967 18037
rect 14691 18071 14749 18077
rect 14691 18037 14703 18071
rect 14737 18068 14749 18071
rect 14918 18068 14924 18080
rect 14737 18040 14924 18068
rect 14737 18037 14749 18040
rect 14691 18031 14749 18037
rect 14918 18028 14924 18040
rect 14976 18028 14982 18080
rect 15657 18071 15715 18077
rect 15657 18037 15669 18071
rect 15703 18068 15715 18071
rect 15838 18068 15844 18080
rect 15703 18040 15844 18068
rect 15703 18037 15715 18040
rect 15657 18031 15715 18037
rect 15838 18028 15844 18040
rect 15896 18028 15902 18080
rect 17862 18028 17868 18080
rect 17920 18068 17926 18080
rect 18187 18071 18245 18077
rect 18187 18068 18199 18071
rect 17920 18040 18199 18068
rect 17920 18028 17926 18040
rect 18187 18037 18199 18040
rect 18233 18037 18245 18071
rect 21910 18068 21916 18080
rect 21871 18040 21916 18068
rect 18187 18031 18245 18037
rect 21910 18028 21916 18040
rect 21968 18028 21974 18080
rect 22002 18028 22008 18080
rect 22060 18068 22066 18080
rect 22112 18068 22140 18099
rect 22186 18096 22192 18148
rect 22244 18136 22250 18148
rect 22741 18139 22799 18145
rect 22244 18108 22289 18136
rect 22244 18096 22250 18108
rect 22741 18105 22753 18139
rect 22787 18136 22799 18139
rect 22787 18108 23796 18136
rect 22787 18105 22799 18108
rect 22741 18099 22799 18105
rect 22060 18040 22140 18068
rect 23768 18068 23796 18108
rect 23842 18096 23848 18148
rect 23900 18136 23906 18148
rect 24946 18136 24952 18148
rect 23900 18108 24952 18136
rect 23900 18096 23906 18108
rect 24946 18096 24952 18108
rect 25004 18096 25010 18148
rect 25133 18139 25191 18145
rect 25133 18105 25145 18139
rect 25179 18136 25191 18139
rect 25685 18139 25743 18145
rect 25685 18136 25697 18139
rect 25179 18108 25697 18136
rect 25179 18105 25191 18108
rect 25133 18099 25191 18105
rect 25685 18105 25697 18108
rect 25731 18105 25743 18139
rect 25685 18099 25743 18105
rect 25777 18139 25835 18145
rect 25777 18105 25789 18139
rect 25823 18136 25835 18139
rect 26344 18136 26372 18312
rect 36814 18300 36820 18352
rect 36872 18340 36878 18352
rect 40218 18340 40224 18352
rect 36872 18312 38516 18340
rect 40179 18312 40224 18340
rect 36872 18300 36878 18312
rect 27985 18275 28043 18281
rect 27985 18272 27997 18275
rect 26988 18244 27997 18272
rect 26786 18136 26792 18148
rect 25823 18108 26792 18136
rect 25823 18105 25835 18108
rect 25777 18099 25835 18105
rect 24210 18068 24216 18080
rect 23768 18040 24216 18068
rect 22060 18028 22066 18040
rect 24210 18028 24216 18040
rect 24268 18028 24274 18080
rect 25700 18068 25728 18099
rect 26786 18096 26792 18108
rect 26844 18096 26850 18148
rect 26988 18068 27016 18244
rect 27985 18241 27997 18244
rect 28031 18272 28043 18275
rect 28718 18272 28724 18284
rect 28031 18244 28724 18272
rect 28031 18241 28043 18244
rect 27985 18235 28043 18241
rect 28718 18232 28724 18244
rect 28776 18232 28782 18284
rect 33502 18232 33508 18284
rect 33560 18272 33566 18284
rect 36633 18275 36691 18281
rect 33560 18244 34979 18272
rect 33560 18232 33566 18244
rect 28810 18164 28816 18216
rect 28868 18204 28874 18216
rect 29308 18207 29366 18213
rect 29308 18204 29320 18207
rect 28868 18176 29320 18204
rect 28868 18164 28874 18176
rect 29308 18173 29320 18176
rect 29354 18204 29366 18207
rect 30101 18207 30159 18213
rect 30101 18204 30113 18207
rect 29354 18176 30113 18204
rect 29354 18173 29366 18176
rect 29308 18167 29366 18173
rect 30101 18173 30113 18176
rect 30147 18173 30159 18207
rect 30650 18204 30656 18216
rect 30611 18176 30656 18204
rect 30101 18167 30159 18173
rect 30650 18164 30656 18176
rect 30708 18164 30714 18216
rect 33172 18207 33230 18213
rect 33172 18173 33184 18207
rect 33218 18173 33230 18207
rect 33172 18167 33230 18173
rect 33275 18207 33333 18213
rect 33275 18173 33287 18207
rect 33321 18204 33333 18207
rect 34698 18204 34704 18216
rect 33321 18176 34704 18204
rect 33321 18173 33333 18176
rect 33275 18167 33333 18173
rect 27706 18136 27712 18148
rect 27667 18108 27712 18136
rect 27706 18096 27712 18108
rect 27764 18096 27770 18148
rect 27801 18139 27859 18145
rect 27801 18105 27813 18139
rect 27847 18105 27859 18139
rect 30974 18139 31032 18145
rect 30974 18136 30986 18139
rect 27801 18099 27859 18105
rect 30576 18108 30986 18136
rect 27430 18068 27436 18080
rect 25700 18040 27016 18068
rect 27391 18040 27436 18068
rect 27430 18028 27436 18040
rect 27488 18068 27494 18080
rect 27816 18068 27844 18099
rect 30576 18080 30604 18108
rect 30974 18105 30986 18108
rect 31020 18105 31032 18139
rect 32214 18136 32220 18148
rect 32175 18108 32220 18136
rect 30974 18099 31032 18105
rect 32214 18096 32220 18108
rect 32272 18096 32278 18148
rect 33187 18136 33215 18167
rect 34698 18164 34704 18176
rect 34756 18164 34762 18216
rect 34951 18213 34979 18244
rect 36633 18241 36645 18275
rect 36679 18272 36691 18275
rect 37366 18272 37372 18284
rect 36679 18244 37372 18272
rect 36679 18241 36691 18244
rect 36633 18235 36691 18241
rect 37366 18232 37372 18244
rect 37424 18232 37430 18284
rect 38488 18281 38516 18312
rect 40218 18300 40224 18312
rect 40276 18300 40282 18352
rect 40604 18281 40632 18368
rect 41598 18340 41604 18352
rect 41559 18312 41604 18340
rect 41598 18300 41604 18312
rect 41656 18300 41662 18352
rect 41690 18300 41696 18352
rect 41748 18340 41754 18352
rect 42766 18340 42794 18380
rect 43990 18368 43996 18380
rect 44048 18368 44054 18420
rect 41748 18312 42794 18340
rect 41748 18300 41754 18312
rect 38473 18275 38531 18281
rect 38473 18241 38485 18275
rect 38519 18241 38531 18275
rect 38473 18235 38531 18241
rect 40589 18275 40647 18281
rect 40589 18241 40601 18275
rect 40635 18241 40647 18275
rect 43070 18272 43076 18284
rect 43031 18244 43076 18272
rect 40589 18235 40647 18241
rect 43070 18232 43076 18244
rect 43128 18232 43134 18284
rect 43717 18275 43775 18281
rect 43717 18241 43729 18275
rect 43763 18272 43775 18275
rect 44174 18272 44180 18284
rect 43763 18244 44180 18272
rect 43763 18241 43775 18244
rect 43717 18235 43775 18241
rect 44174 18232 44180 18244
rect 44232 18232 44238 18284
rect 34936 18207 34994 18213
rect 34936 18173 34948 18207
rect 34982 18204 34994 18207
rect 35342 18204 35348 18216
rect 34982 18176 35348 18204
rect 34982 18173 34994 18176
rect 34936 18167 34994 18173
rect 35342 18164 35348 18176
rect 35400 18164 35406 18216
rect 33187 18108 33272 18136
rect 33244 18080 33272 18108
rect 33502 18096 33508 18148
rect 33560 18136 33566 18148
rect 35023 18139 35081 18145
rect 35023 18136 35035 18139
rect 33560 18108 35035 18136
rect 33560 18096 33566 18108
rect 35023 18105 35035 18108
rect 35069 18105 35081 18139
rect 35023 18099 35081 18105
rect 36725 18139 36783 18145
rect 36725 18105 36737 18139
rect 36771 18136 36783 18139
rect 37090 18136 37096 18148
rect 36771 18108 37096 18136
rect 36771 18105 36783 18108
rect 36725 18099 36783 18105
rect 37090 18096 37096 18108
rect 37148 18096 37154 18148
rect 37274 18136 37280 18148
rect 37235 18108 37280 18136
rect 37274 18096 37280 18108
rect 37332 18096 37338 18148
rect 38194 18136 38200 18148
rect 38155 18108 38200 18136
rect 38194 18096 38200 18108
rect 38252 18096 38258 18148
rect 38289 18139 38347 18145
rect 38289 18105 38301 18139
rect 38335 18105 38347 18139
rect 38289 18099 38347 18105
rect 27488 18040 27844 18068
rect 27488 18028 27494 18040
rect 28994 18028 29000 18080
rect 29052 18068 29058 18080
rect 29411 18071 29469 18077
rect 29411 18068 29423 18071
rect 29052 18040 29423 18068
rect 29052 18028 29058 18040
rect 29411 18037 29423 18040
rect 29457 18037 29469 18071
rect 30558 18068 30564 18080
rect 30519 18040 30564 18068
rect 29411 18031 29469 18037
rect 30558 18028 30564 18040
rect 30616 18028 30622 18080
rect 31110 18028 31116 18080
rect 31168 18068 31174 18080
rect 31573 18071 31631 18077
rect 31573 18068 31585 18071
rect 31168 18040 31585 18068
rect 31168 18028 31174 18040
rect 31573 18037 31585 18040
rect 31619 18037 31631 18071
rect 33226 18068 33232 18080
rect 33139 18040 33232 18068
rect 31573 18031 31631 18037
rect 33226 18028 33232 18040
rect 33284 18068 33290 18080
rect 33689 18071 33747 18077
rect 33689 18068 33701 18071
rect 33284 18040 33701 18068
rect 33284 18028 33290 18040
rect 33689 18037 33701 18040
rect 33735 18068 33747 18071
rect 33962 18068 33968 18080
rect 33735 18040 33968 18068
rect 33735 18037 33747 18040
rect 33689 18031 33747 18037
rect 33962 18028 33968 18040
rect 34020 18028 34026 18080
rect 34606 18068 34612 18080
rect 34567 18040 34612 18068
rect 34606 18028 34612 18040
rect 34664 18028 34670 18080
rect 37918 18068 37924 18080
rect 37879 18040 37924 18068
rect 37918 18028 37924 18040
rect 37976 18068 37982 18080
rect 38304 18068 38332 18099
rect 40678 18096 40684 18148
rect 40736 18136 40742 18148
rect 41230 18136 41236 18148
rect 40736 18108 40781 18136
rect 41191 18108 41236 18136
rect 40736 18096 40742 18108
rect 41230 18096 41236 18108
rect 41288 18096 41294 18148
rect 42889 18139 42947 18145
rect 42889 18105 42901 18139
rect 42935 18136 42947 18139
rect 43165 18139 43223 18145
rect 43165 18136 43177 18139
rect 42935 18108 43177 18136
rect 42935 18105 42947 18108
rect 42889 18099 42947 18105
rect 43165 18105 43177 18108
rect 43211 18136 43223 18139
rect 43530 18136 43536 18148
rect 43211 18108 43536 18136
rect 43211 18105 43223 18108
rect 43165 18099 43223 18105
rect 43530 18096 43536 18108
rect 43588 18096 43594 18148
rect 37976 18040 38332 18068
rect 37976 18028 37982 18040
rect 38562 18028 38568 18080
rect 38620 18068 38626 18080
rect 39117 18071 39175 18077
rect 39117 18068 39129 18071
rect 38620 18040 39129 18068
rect 38620 18028 38626 18040
rect 39117 18037 39129 18040
rect 39163 18037 39175 18071
rect 39117 18031 39175 18037
rect 1104 17978 48852 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 48852 17978
rect 1104 17904 48852 17926
rect 9858 17864 9864 17876
rect 9819 17836 9864 17864
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 10318 17864 10324 17876
rect 9968 17836 10324 17864
rect 9214 17756 9220 17808
rect 9272 17796 9278 17808
rect 9968 17796 9996 17836
rect 10318 17824 10324 17836
rect 10376 17824 10382 17876
rect 10502 17824 10508 17876
rect 10560 17864 10566 17876
rect 10781 17867 10839 17873
rect 10781 17864 10793 17867
rect 10560 17836 10793 17864
rect 10560 17824 10566 17836
rect 10781 17833 10793 17836
rect 10827 17833 10839 17867
rect 12986 17864 12992 17876
rect 12947 17836 12992 17864
rect 10781 17827 10839 17833
rect 12986 17824 12992 17836
rect 13044 17824 13050 17876
rect 16482 17864 16488 17876
rect 16443 17836 16488 17864
rect 16482 17824 16488 17836
rect 16540 17824 16546 17876
rect 18969 17867 19027 17873
rect 18969 17833 18981 17867
rect 19015 17864 19027 17867
rect 19242 17864 19248 17876
rect 19015 17836 19248 17864
rect 19015 17833 19027 17836
rect 18969 17827 19027 17833
rect 19242 17824 19248 17836
rect 19300 17824 19306 17876
rect 19978 17864 19984 17876
rect 19939 17836 19984 17864
rect 19978 17824 19984 17836
rect 20036 17824 20042 17876
rect 21266 17864 21272 17876
rect 21227 17836 21272 17864
rect 21266 17824 21272 17836
rect 21324 17824 21330 17876
rect 23446 17836 24900 17864
rect 11698 17796 11704 17808
rect 9272 17768 9996 17796
rect 11659 17768 11704 17796
rect 9272 17756 9278 17768
rect 11698 17756 11704 17768
rect 11756 17756 11762 17808
rect 11882 17756 11888 17808
rect 11940 17796 11946 17808
rect 13170 17796 13176 17808
rect 11940 17768 13176 17796
rect 11940 17756 11946 17768
rect 13170 17756 13176 17768
rect 13228 17756 13234 17808
rect 13265 17799 13323 17805
rect 13265 17765 13277 17799
rect 13311 17796 13323 17799
rect 13446 17796 13452 17808
rect 13311 17768 13452 17796
rect 13311 17765 13323 17768
rect 13265 17759 13323 17765
rect 13446 17756 13452 17768
rect 13504 17756 13510 17808
rect 15473 17799 15531 17805
rect 15473 17765 15485 17799
rect 15519 17796 15531 17799
rect 15562 17796 15568 17808
rect 15519 17768 15568 17796
rect 15519 17765 15531 17768
rect 15473 17759 15531 17765
rect 15562 17756 15568 17768
rect 15620 17756 15626 17808
rect 17034 17796 17040 17808
rect 16995 17768 17040 17796
rect 17034 17756 17040 17768
rect 17092 17756 17098 17808
rect 23290 17796 23296 17808
rect 23251 17768 23296 17796
rect 23290 17756 23296 17768
rect 23348 17796 23354 17808
rect 23446 17796 23474 17836
rect 24872 17808 24900 17836
rect 27062 17824 27068 17876
rect 27120 17873 27126 17876
rect 27120 17867 27169 17873
rect 27120 17833 27123 17867
rect 27157 17833 27169 17867
rect 27120 17827 27169 17833
rect 27120 17824 27126 17827
rect 30834 17824 30840 17876
rect 30892 17864 30898 17876
rect 31113 17867 31171 17873
rect 31113 17864 31125 17867
rect 30892 17836 31125 17864
rect 30892 17824 30898 17836
rect 31113 17833 31125 17836
rect 31159 17864 31171 17867
rect 33686 17864 33692 17876
rect 31159 17836 33692 17864
rect 31159 17833 31171 17836
rect 31113 17827 31171 17833
rect 33686 17824 33692 17836
rect 33744 17824 33750 17876
rect 36679 17867 36737 17873
rect 36679 17833 36691 17867
rect 36725 17864 36737 17867
rect 37182 17864 37188 17876
rect 36725 17836 37188 17864
rect 36725 17833 36737 17836
rect 36679 17827 36737 17833
rect 37182 17824 37188 17836
rect 37240 17824 37246 17876
rect 37366 17864 37372 17876
rect 37327 17836 37372 17864
rect 37366 17824 37372 17836
rect 37424 17824 37430 17876
rect 38102 17824 38108 17876
rect 38160 17864 38166 17876
rect 38562 17864 38568 17876
rect 38160 17836 38568 17864
rect 38160 17824 38166 17836
rect 38562 17824 38568 17836
rect 38620 17824 38626 17876
rect 38838 17864 38844 17876
rect 38799 17836 38844 17864
rect 38838 17824 38844 17836
rect 38896 17824 38902 17876
rect 45051 17867 45109 17873
rect 45051 17864 45063 17867
rect 43456 17836 45063 17864
rect 23348 17768 23474 17796
rect 23845 17799 23903 17805
rect 23348 17756 23354 17768
rect 23845 17765 23857 17799
rect 23891 17796 23903 17799
rect 24394 17796 24400 17808
rect 23891 17768 24400 17796
rect 23891 17765 23903 17768
rect 23845 17759 23903 17765
rect 24394 17756 24400 17768
rect 24452 17756 24458 17808
rect 24854 17796 24860 17808
rect 24815 17768 24860 17796
rect 24854 17756 24860 17768
rect 24912 17756 24918 17808
rect 28169 17799 28227 17805
rect 28169 17765 28181 17799
rect 28215 17796 28227 17799
rect 28534 17796 28540 17808
rect 28215 17768 28540 17796
rect 28215 17765 28227 17768
rect 28169 17759 28227 17765
rect 28534 17756 28540 17768
rect 28592 17756 28598 17808
rect 28718 17796 28724 17808
rect 28679 17768 28724 17796
rect 28718 17756 28724 17768
rect 28776 17756 28782 17808
rect 29730 17756 29736 17808
rect 29788 17796 29794 17808
rect 29788 17768 30512 17796
rect 29788 17756 29794 17768
rect 30484 17740 30512 17768
rect 30650 17756 30656 17808
rect 30708 17796 30714 17808
rect 30745 17799 30803 17805
rect 30745 17796 30757 17799
rect 30708 17768 30757 17796
rect 30708 17756 30714 17768
rect 30745 17765 30757 17768
rect 30791 17796 30803 17799
rect 31389 17799 31447 17805
rect 31389 17796 31401 17799
rect 30791 17768 31401 17796
rect 30791 17765 30803 17768
rect 30745 17759 30803 17765
rect 31389 17765 31401 17768
rect 31435 17765 31447 17799
rect 31389 17759 31447 17765
rect 33321 17799 33379 17805
rect 33321 17765 33333 17799
rect 33367 17796 33379 17799
rect 33502 17796 33508 17808
rect 33367 17768 33508 17796
rect 33367 17765 33379 17768
rect 33321 17759 33379 17765
rect 33502 17756 33508 17768
rect 33560 17756 33566 17808
rect 33594 17756 33600 17808
rect 33652 17796 33658 17808
rect 34330 17796 34336 17808
rect 33652 17768 34336 17796
rect 33652 17756 33658 17768
rect 34330 17756 34336 17768
rect 34388 17796 34394 17808
rect 35161 17799 35219 17805
rect 35161 17796 35173 17799
rect 34388 17768 35173 17796
rect 34388 17756 34394 17768
rect 35161 17765 35173 17768
rect 35207 17765 35219 17799
rect 35161 17759 35219 17765
rect 36354 17756 36360 17808
rect 36412 17796 36418 17808
rect 37090 17796 37096 17808
rect 36412 17768 36722 17796
rect 37003 17768 37096 17796
rect 36412 17756 36418 17768
rect 10045 17731 10103 17737
rect 10045 17697 10057 17731
rect 10091 17728 10103 17731
rect 10318 17728 10324 17740
rect 10091 17700 10180 17728
rect 10279 17700 10324 17728
rect 10091 17697 10103 17700
rect 10045 17691 10103 17697
rect 9674 17484 9680 17536
rect 9732 17524 9738 17536
rect 10152 17524 10180 17700
rect 10318 17688 10324 17700
rect 10376 17688 10382 17740
rect 17954 17688 17960 17740
rect 18012 17728 18018 17740
rect 18141 17731 18199 17737
rect 18141 17728 18153 17731
rect 18012 17700 18153 17728
rect 18012 17688 18018 17700
rect 18141 17697 18153 17700
rect 18187 17728 18199 17731
rect 19521 17731 19579 17737
rect 19521 17728 19533 17731
rect 18187 17700 19533 17728
rect 18187 17697 18199 17700
rect 18141 17691 18199 17697
rect 19521 17697 19533 17700
rect 19567 17697 19579 17731
rect 19521 17691 19579 17697
rect 27040 17731 27098 17737
rect 27040 17697 27052 17731
rect 27086 17728 27098 17731
rect 27338 17728 27344 17740
rect 27086 17700 27344 17728
rect 27086 17697 27098 17700
rect 27040 17691 27098 17697
rect 27338 17688 27344 17700
rect 27396 17688 27402 17740
rect 30282 17728 30288 17740
rect 30243 17700 30288 17728
rect 30282 17688 30288 17700
rect 30340 17688 30346 17740
rect 30466 17728 30472 17740
rect 30379 17700 30472 17728
rect 30466 17688 30472 17700
rect 30524 17688 30530 17740
rect 36538 17728 36544 17740
rect 36499 17700 36544 17728
rect 36538 17688 36544 17700
rect 36596 17688 36602 17740
rect 36694 17728 36722 17768
rect 37090 17756 37096 17768
rect 37148 17796 37154 17808
rect 37642 17796 37648 17808
rect 37148 17768 37648 17796
rect 37148 17756 37154 17768
rect 37642 17756 37648 17768
rect 37700 17756 37706 17808
rect 39482 17756 39488 17808
rect 39540 17796 39546 17808
rect 41506 17805 41512 17808
rect 39714 17799 39772 17805
rect 39714 17796 39726 17799
rect 39540 17768 39726 17796
rect 39540 17756 39546 17768
rect 39714 17765 39726 17768
rect 39760 17796 39772 17799
rect 41462 17799 41512 17805
rect 41462 17796 41474 17799
rect 39760 17768 41474 17796
rect 39760 17765 39772 17768
rect 39714 17759 39772 17765
rect 41462 17765 41474 17768
rect 41508 17765 41512 17799
rect 41462 17759 41512 17765
rect 41506 17756 41512 17759
rect 41564 17756 41570 17808
rect 43456 17805 43484 17836
rect 45051 17833 45063 17836
rect 45097 17833 45109 17867
rect 45051 17827 45109 17833
rect 43165 17799 43223 17805
rect 43165 17765 43177 17799
rect 43211 17796 43223 17799
rect 43441 17799 43499 17805
rect 43441 17796 43453 17799
rect 43211 17768 43453 17796
rect 43211 17765 43223 17768
rect 43165 17759 43223 17765
rect 43441 17765 43453 17768
rect 43487 17765 43499 17799
rect 43441 17759 43499 17765
rect 43530 17756 43536 17808
rect 43588 17796 43594 17808
rect 43588 17768 43633 17796
rect 43588 17756 43594 17768
rect 37826 17728 37832 17740
rect 36694 17700 37832 17728
rect 37826 17688 37832 17700
rect 37884 17688 37890 17740
rect 38381 17731 38439 17737
rect 38381 17697 38393 17731
rect 38427 17728 38439 17731
rect 38470 17728 38476 17740
rect 38427 17700 38476 17728
rect 38427 17697 38439 17700
rect 38381 17691 38439 17697
rect 38470 17688 38476 17700
rect 38528 17688 38534 17740
rect 40678 17728 40684 17740
rect 40591 17700 40684 17728
rect 40678 17688 40684 17700
rect 40736 17728 40742 17740
rect 42061 17731 42119 17737
rect 42061 17728 42073 17731
rect 40736 17700 42073 17728
rect 40736 17688 40742 17700
rect 42061 17697 42073 17700
rect 42107 17697 42119 17731
rect 42061 17691 42119 17697
rect 44980 17731 45038 17737
rect 44980 17697 44992 17731
rect 45026 17728 45038 17731
rect 45186 17728 45192 17740
rect 45026 17700 45192 17728
rect 45026 17697 45038 17700
rect 44980 17691 45038 17697
rect 45186 17688 45192 17700
rect 45244 17688 45250 17740
rect 11330 17620 11336 17672
rect 11388 17660 11394 17672
rect 11609 17663 11667 17669
rect 11609 17660 11621 17663
rect 11388 17632 11621 17660
rect 11388 17620 11394 17632
rect 11609 17629 11621 17632
rect 11655 17629 11667 17663
rect 13449 17663 13507 17669
rect 13449 17660 13461 17663
rect 11609 17623 11667 17629
rect 13366 17632 13461 17660
rect 12161 17595 12219 17601
rect 12161 17561 12173 17595
rect 12207 17592 12219 17595
rect 12526 17592 12532 17604
rect 12207 17564 12532 17592
rect 12207 17561 12219 17564
rect 12161 17555 12219 17561
rect 12526 17552 12532 17564
rect 12584 17592 12590 17604
rect 12621 17595 12679 17601
rect 12621 17592 12633 17595
rect 12584 17564 12633 17592
rect 12584 17552 12590 17564
rect 12621 17561 12633 17564
rect 12667 17592 12679 17595
rect 13366 17592 13394 17632
rect 13449 17629 13461 17632
rect 13495 17629 13507 17663
rect 13449 17623 13507 17629
rect 15102 17620 15108 17672
rect 15160 17660 15166 17672
rect 15381 17663 15439 17669
rect 15381 17660 15393 17663
rect 15160 17632 15393 17660
rect 15160 17620 15166 17632
rect 15381 17629 15393 17632
rect 15427 17629 15439 17663
rect 16022 17660 16028 17672
rect 15983 17632 16028 17660
rect 15381 17623 15439 17629
rect 12667 17564 13394 17592
rect 15396 17592 15424 17623
rect 16022 17620 16028 17632
rect 16080 17620 16086 17672
rect 16945 17663 17003 17669
rect 16945 17629 16957 17663
rect 16991 17660 17003 17663
rect 17402 17660 17408 17672
rect 16991 17632 17408 17660
rect 16991 17629 17003 17632
rect 16945 17623 17003 17629
rect 17402 17620 17408 17632
rect 17460 17660 17466 17672
rect 17862 17660 17868 17672
rect 17460 17632 17868 17660
rect 17460 17620 17466 17632
rect 17862 17620 17868 17632
rect 17920 17620 17926 17672
rect 18598 17660 18604 17672
rect 18559 17632 18604 17660
rect 18598 17620 18604 17632
rect 18656 17620 18662 17672
rect 20622 17620 20628 17672
rect 20680 17660 20686 17672
rect 20901 17663 20959 17669
rect 20901 17660 20913 17663
rect 20680 17632 20913 17660
rect 20680 17620 20686 17632
rect 20901 17629 20913 17632
rect 20947 17629 20959 17663
rect 23198 17660 23204 17672
rect 23159 17632 23204 17660
rect 20901 17623 20959 17629
rect 23198 17620 23204 17632
rect 23256 17620 23262 17672
rect 24762 17660 24768 17672
rect 24723 17632 24768 17660
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 25038 17660 25044 17672
rect 24999 17632 25044 17660
rect 25038 17620 25044 17632
rect 25096 17620 25102 17672
rect 28077 17663 28135 17669
rect 28077 17629 28089 17663
rect 28123 17660 28135 17663
rect 28994 17660 29000 17672
rect 28123 17632 29000 17660
rect 28123 17629 28135 17632
rect 28077 17623 28135 17629
rect 28994 17620 29000 17632
rect 29052 17620 29058 17672
rect 31202 17620 31208 17672
rect 31260 17660 31266 17672
rect 32125 17663 32183 17669
rect 32125 17660 32137 17663
rect 31260 17632 32137 17660
rect 31260 17620 31266 17632
rect 32125 17629 32137 17632
rect 32171 17629 32183 17663
rect 33778 17660 33784 17672
rect 33739 17632 33784 17660
rect 32125 17623 32183 17629
rect 33778 17620 33784 17632
rect 33836 17620 33842 17672
rect 34698 17620 34704 17672
rect 34756 17660 34762 17672
rect 35069 17663 35127 17669
rect 35069 17660 35081 17663
rect 34756 17632 35081 17660
rect 34756 17620 34762 17632
rect 35069 17629 35081 17632
rect 35115 17660 35127 17663
rect 35434 17660 35440 17672
rect 35115 17632 35440 17660
rect 35115 17629 35127 17632
rect 35069 17623 35127 17629
rect 35434 17620 35440 17632
rect 35492 17620 35498 17672
rect 38565 17663 38623 17669
rect 38565 17629 38577 17663
rect 38611 17660 38623 17663
rect 39393 17663 39451 17669
rect 39393 17660 39405 17663
rect 38611 17632 39405 17660
rect 38611 17629 38623 17632
rect 38565 17623 38623 17629
rect 39393 17629 39405 17632
rect 39439 17660 39451 17663
rect 39850 17660 39856 17672
rect 39439 17632 39856 17660
rect 39439 17629 39451 17632
rect 39393 17623 39451 17629
rect 39850 17620 39856 17632
rect 39908 17620 39914 17672
rect 41046 17620 41052 17672
rect 41104 17660 41110 17672
rect 41141 17663 41199 17669
rect 41141 17660 41153 17663
rect 41104 17632 41153 17660
rect 41104 17620 41110 17632
rect 41141 17629 41153 17632
rect 41187 17629 41199 17663
rect 43717 17663 43775 17669
rect 43717 17660 43729 17663
rect 41141 17623 41199 17629
rect 43548 17632 43729 17660
rect 17126 17592 17132 17604
rect 15396 17564 17132 17592
rect 12667 17561 12679 17564
rect 12621 17555 12679 17561
rect 17126 17552 17132 17564
rect 17184 17592 17190 17604
rect 17497 17595 17555 17601
rect 17497 17592 17509 17595
rect 17184 17564 17509 17592
rect 17184 17552 17190 17564
rect 17497 17561 17509 17564
rect 17543 17561 17555 17595
rect 17497 17555 17555 17561
rect 17604 17564 18552 17592
rect 14550 17524 14556 17536
rect 9732 17496 14556 17524
rect 9732 17484 9738 17496
rect 14550 17484 14556 17496
rect 14608 17524 14614 17536
rect 17604 17524 17632 17564
rect 14608 17496 17632 17524
rect 14608 17484 14614 17496
rect 18138 17484 18144 17536
rect 18196 17524 18202 17536
rect 18417 17527 18475 17533
rect 18417 17524 18429 17527
rect 18196 17496 18429 17524
rect 18196 17484 18202 17496
rect 18417 17493 18429 17496
rect 18463 17493 18475 17527
rect 18524 17524 18552 17564
rect 20070 17552 20076 17604
rect 20128 17592 20134 17604
rect 21821 17595 21879 17601
rect 21821 17592 21833 17595
rect 20128 17564 21833 17592
rect 20128 17552 20134 17564
rect 21821 17561 21833 17564
rect 21867 17561 21879 17595
rect 21821 17555 21879 17561
rect 34238 17552 34244 17604
rect 34296 17592 34302 17604
rect 35621 17595 35679 17601
rect 35621 17592 35633 17595
rect 34296 17564 35633 17592
rect 34296 17552 34302 17564
rect 35621 17561 35633 17564
rect 35667 17561 35679 17595
rect 35621 17555 35679 17561
rect 40586 17552 40592 17604
rect 40644 17592 40650 17604
rect 41966 17592 41972 17604
rect 40644 17564 41972 17592
rect 40644 17552 40650 17564
rect 41966 17552 41972 17564
rect 42024 17592 42030 17604
rect 43548 17592 43576 17632
rect 43717 17629 43729 17632
rect 43763 17629 43775 17663
rect 43717 17623 43775 17629
rect 42024 17564 43576 17592
rect 42024 17552 42030 17564
rect 20254 17524 20260 17536
rect 18524 17496 20260 17524
rect 18417 17487 18475 17493
rect 20254 17484 20260 17496
rect 20312 17484 20318 17536
rect 22002 17484 22008 17536
rect 22060 17524 22066 17536
rect 22097 17527 22155 17533
rect 22097 17524 22109 17527
rect 22060 17496 22109 17524
rect 22060 17484 22066 17496
rect 22097 17493 22109 17496
rect 22143 17493 22155 17527
rect 22097 17487 22155 17493
rect 25590 17484 25596 17536
rect 25648 17524 25654 17536
rect 25685 17527 25743 17533
rect 25685 17524 25697 17527
rect 25648 17496 25697 17524
rect 25648 17484 25654 17496
rect 25685 17493 25697 17496
rect 25731 17493 25743 17527
rect 27706 17524 27712 17536
rect 27619 17496 27712 17524
rect 25685 17487 25743 17493
rect 27706 17484 27712 17496
rect 27764 17524 27770 17536
rect 29086 17524 29092 17536
rect 27764 17496 29092 17524
rect 27764 17484 27770 17496
rect 29086 17484 29092 17496
rect 29144 17484 29150 17536
rect 40310 17524 40316 17536
rect 40271 17496 40316 17524
rect 40310 17484 40316 17496
rect 40368 17484 40374 17536
rect 1104 17434 48852 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 48852 17434
rect 1104 17360 48852 17382
rect 9674 17320 9680 17332
rect 9635 17292 9680 17320
rect 9674 17280 9680 17292
rect 9732 17280 9738 17332
rect 13170 17280 13176 17332
rect 13228 17320 13234 17332
rect 13817 17323 13875 17329
rect 13817 17320 13829 17323
rect 13228 17292 13829 17320
rect 13228 17280 13234 17292
rect 13817 17289 13829 17292
rect 13863 17289 13875 17323
rect 13817 17283 13875 17289
rect 14918 17280 14924 17332
rect 14976 17320 14982 17332
rect 15749 17323 15807 17329
rect 15749 17320 15761 17323
rect 14976 17292 15761 17320
rect 14976 17280 14982 17292
rect 15749 17289 15761 17292
rect 15795 17289 15807 17323
rect 17402 17320 17408 17332
rect 17363 17292 17408 17320
rect 15749 17283 15807 17289
rect 13446 17252 13452 17264
rect 13407 17224 13452 17252
rect 13446 17212 13452 17224
rect 13504 17212 13510 17264
rect 10137 17187 10195 17193
rect 10137 17153 10149 17187
rect 10183 17184 10195 17187
rect 10502 17184 10508 17196
rect 10183 17156 10508 17184
rect 10183 17153 10195 17156
rect 10137 17147 10195 17153
rect 10502 17144 10508 17156
rect 10560 17144 10566 17196
rect 12526 17184 12532 17196
rect 12487 17156 12532 17184
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 12986 17184 12992 17196
rect 12947 17156 12992 17184
rect 12986 17144 12992 17156
rect 13044 17144 13050 17196
rect 14274 17116 14280 17128
rect 14187 17088 14280 17116
rect 14274 17076 14280 17088
rect 14332 17116 14338 17128
rect 14461 17119 14519 17125
rect 14461 17116 14473 17119
rect 14332 17088 14473 17116
rect 14332 17076 14338 17088
rect 14461 17085 14473 17088
rect 14507 17085 14519 17119
rect 15764 17116 15792 17283
rect 17402 17280 17408 17292
rect 17460 17280 17466 17332
rect 19242 17320 19248 17332
rect 19203 17292 19248 17320
rect 19242 17280 19248 17292
rect 19300 17280 19306 17332
rect 21361 17323 21419 17329
rect 21361 17289 21373 17323
rect 21407 17320 21419 17323
rect 21450 17320 21456 17332
rect 21407 17292 21456 17320
rect 21407 17289 21419 17292
rect 21361 17283 21419 17289
rect 21450 17280 21456 17292
rect 21508 17280 21514 17332
rect 23109 17323 23167 17329
rect 23109 17289 23121 17323
rect 23155 17320 23167 17323
rect 23290 17320 23296 17332
rect 23155 17292 23296 17320
rect 23155 17289 23167 17292
rect 23109 17283 23167 17289
rect 23290 17280 23296 17292
rect 23348 17280 23354 17332
rect 24765 17323 24823 17329
rect 24765 17289 24777 17323
rect 24811 17320 24823 17323
rect 24854 17320 24860 17332
rect 24811 17292 24860 17320
rect 24811 17289 24823 17292
rect 24765 17283 24823 17289
rect 24854 17280 24860 17292
rect 24912 17320 24918 17332
rect 25317 17323 25375 17329
rect 25317 17320 25329 17323
rect 24912 17292 25329 17320
rect 24912 17280 24918 17292
rect 25317 17289 25329 17292
rect 25363 17320 25375 17323
rect 25682 17320 25688 17332
rect 25363 17292 25688 17320
rect 25363 17289 25375 17292
rect 25317 17283 25375 17289
rect 25682 17280 25688 17292
rect 25740 17280 25746 17332
rect 28994 17320 29000 17332
rect 28955 17292 29000 17320
rect 28994 17280 29000 17292
rect 29052 17280 29058 17332
rect 29086 17280 29092 17332
rect 29144 17320 29150 17332
rect 29411 17323 29469 17329
rect 29411 17320 29423 17323
rect 29144 17292 29423 17320
rect 29144 17280 29150 17292
rect 29411 17289 29423 17292
rect 29457 17289 29469 17323
rect 30466 17320 30472 17332
rect 30427 17292 30472 17320
rect 29411 17283 29469 17289
rect 30466 17280 30472 17292
rect 30524 17280 30530 17332
rect 33134 17280 33140 17332
rect 33192 17320 33198 17332
rect 33870 17320 33876 17332
rect 33192 17292 33876 17320
rect 33192 17280 33198 17292
rect 33870 17280 33876 17292
rect 33928 17280 33934 17332
rect 34330 17320 34336 17332
rect 34291 17292 34336 17320
rect 34330 17280 34336 17292
rect 34388 17280 34394 17332
rect 35986 17280 35992 17332
rect 36044 17320 36050 17332
rect 39482 17320 39488 17332
rect 36044 17292 39488 17320
rect 36044 17280 36050 17292
rect 39482 17280 39488 17292
rect 39540 17280 39546 17332
rect 39850 17320 39856 17332
rect 39811 17292 39856 17320
rect 39850 17280 39856 17292
rect 39908 17280 39914 17332
rect 40310 17320 40316 17332
rect 40271 17292 40316 17320
rect 40310 17280 40316 17292
rect 40368 17280 40374 17332
rect 41506 17320 41512 17332
rect 41467 17292 41512 17320
rect 41506 17280 41512 17292
rect 41564 17320 41570 17332
rect 42245 17323 42303 17329
rect 42245 17320 42257 17323
rect 41564 17292 42257 17320
rect 41564 17280 41570 17292
rect 42245 17289 42257 17292
rect 42291 17320 42303 17323
rect 43254 17320 43260 17332
rect 42291 17292 43260 17320
rect 42291 17289 42303 17292
rect 42245 17283 42303 17289
rect 15838 17212 15844 17264
rect 15896 17252 15902 17264
rect 18969 17255 19027 17261
rect 18969 17252 18981 17255
rect 15896 17224 18981 17252
rect 15896 17212 15902 17224
rect 18969 17221 18981 17224
rect 19015 17221 19027 17255
rect 18969 17215 19027 17221
rect 20806 17212 20812 17264
rect 20864 17252 20870 17264
rect 22511 17255 22569 17261
rect 22511 17252 22523 17255
rect 20864 17224 22523 17252
rect 20864 17212 20870 17224
rect 22511 17221 22523 17224
rect 22557 17221 22569 17255
rect 22511 17215 22569 17221
rect 31110 17212 31116 17264
rect 31168 17252 31174 17264
rect 32677 17255 32735 17261
rect 32677 17252 32689 17255
rect 31168 17224 32689 17252
rect 31168 17212 31174 17224
rect 32677 17221 32689 17224
rect 32723 17252 32735 17255
rect 33594 17252 33600 17264
rect 32723 17224 33600 17252
rect 32723 17221 32735 17224
rect 32677 17215 32735 17221
rect 33594 17212 33600 17224
rect 33652 17212 33658 17264
rect 36538 17252 36544 17264
rect 36499 17224 36544 17252
rect 36538 17212 36544 17224
rect 36596 17212 36602 17264
rect 36814 17212 36820 17264
rect 36872 17252 36878 17264
rect 37277 17255 37335 17261
rect 37277 17252 37289 17255
rect 36872 17224 37289 17252
rect 36872 17212 36878 17224
rect 37277 17221 37289 17224
rect 37323 17221 37335 17255
rect 37826 17252 37832 17264
rect 37787 17224 37832 17252
rect 37277 17215 37335 17221
rect 37826 17212 37832 17224
rect 37884 17212 37890 17264
rect 38378 17252 38384 17264
rect 38339 17224 38384 17252
rect 38378 17212 38384 17224
rect 38436 17212 38442 17264
rect 41141 17255 41199 17261
rect 41141 17221 41153 17255
rect 41187 17252 41199 17255
rect 41230 17252 41236 17264
rect 41187 17224 41236 17252
rect 41187 17221 41199 17224
rect 41141 17215 41199 17221
rect 41230 17212 41236 17224
rect 41288 17212 41294 17264
rect 20438 17184 20444 17196
rect 20399 17156 20444 17184
rect 20438 17144 20444 17156
rect 20496 17144 20502 17196
rect 22281 17187 22339 17193
rect 22281 17153 22293 17187
rect 22327 17184 22339 17187
rect 23106 17184 23112 17196
rect 22327 17156 23112 17184
rect 22327 17153 22339 17156
rect 22281 17147 22339 17153
rect 16025 17119 16083 17125
rect 16025 17116 16037 17119
rect 15764 17088 16037 17116
rect 14461 17079 14519 17085
rect 16025 17085 16037 17088
rect 16071 17085 16083 17119
rect 16025 17079 16083 17085
rect 18049 17119 18107 17125
rect 18049 17085 18061 17119
rect 18095 17116 18107 17119
rect 18138 17116 18144 17128
rect 18095 17088 18144 17116
rect 18095 17085 18107 17088
rect 18049 17079 18107 17085
rect 18138 17076 18144 17088
rect 18196 17076 18202 17128
rect 22455 17125 22483 17156
rect 23106 17144 23112 17156
rect 23164 17144 23170 17196
rect 24397 17187 24455 17193
rect 24397 17153 24409 17187
rect 24443 17184 24455 17187
rect 25038 17184 25044 17196
rect 24443 17156 25044 17184
rect 24443 17153 24455 17156
rect 24397 17147 24455 17153
rect 25038 17144 25044 17156
rect 25096 17144 25102 17196
rect 25866 17184 25872 17196
rect 25827 17156 25872 17184
rect 25866 17144 25872 17156
rect 25924 17144 25930 17196
rect 27065 17187 27123 17193
rect 27065 17153 27077 17187
rect 27111 17184 27123 17187
rect 27338 17184 27344 17196
rect 27111 17156 27344 17184
rect 27111 17153 27123 17156
rect 27065 17147 27123 17153
rect 27338 17144 27344 17156
rect 27396 17144 27402 17196
rect 31021 17187 31079 17193
rect 31021 17153 31033 17187
rect 31067 17184 31079 17187
rect 31202 17184 31208 17196
rect 31067 17156 31208 17184
rect 31067 17153 31079 17156
rect 31021 17147 31079 17153
rect 31202 17144 31208 17156
rect 31260 17144 31266 17196
rect 31294 17144 31300 17196
rect 31352 17184 31358 17196
rect 31481 17187 31539 17193
rect 31481 17184 31493 17187
rect 31352 17156 31493 17184
rect 31352 17144 31358 17156
rect 31481 17153 31493 17156
rect 31527 17153 31539 17187
rect 31481 17147 31539 17153
rect 33042 17144 33048 17196
rect 33100 17184 33106 17196
rect 33689 17187 33747 17193
rect 33689 17184 33701 17187
rect 33100 17156 33701 17184
rect 33100 17144 33106 17156
rect 33689 17153 33701 17156
rect 33735 17184 33747 17187
rect 33962 17184 33968 17196
rect 33735 17156 33968 17184
rect 33735 17153 33747 17156
rect 33689 17147 33747 17153
rect 33962 17144 33968 17156
rect 34020 17144 34026 17196
rect 36725 17187 36783 17193
rect 36725 17153 36737 17187
rect 36771 17184 36783 17187
rect 37090 17184 37096 17196
rect 36771 17156 37096 17184
rect 36771 17153 36783 17156
rect 36725 17147 36783 17153
rect 37090 17144 37096 17156
rect 37148 17144 37154 17196
rect 22440 17119 22498 17125
rect 22440 17116 22452 17119
rect 22418 17088 22452 17116
rect 22440 17085 22452 17088
rect 22486 17085 22498 17119
rect 22440 17079 22498 17085
rect 27525 17119 27583 17125
rect 27525 17085 27537 17119
rect 27571 17085 27583 17119
rect 27525 17079 27583 17085
rect 10045 17051 10103 17057
rect 10045 17017 10057 17051
rect 10091 17048 10103 17051
rect 10318 17048 10324 17060
rect 10091 17020 10324 17048
rect 10091 17017 10103 17020
rect 10045 17011 10103 17017
rect 10318 17008 10324 17020
rect 10376 17048 10382 17060
rect 10458 17051 10516 17057
rect 10458 17048 10470 17051
rect 10376 17020 10470 17048
rect 10376 17008 10382 17020
rect 10458 17017 10470 17020
rect 10504 17017 10516 17051
rect 10458 17011 10516 17017
rect 12253 17051 12311 17057
rect 12253 17017 12265 17051
rect 12299 17048 12311 17051
rect 12618 17048 12624 17060
rect 12299 17020 12624 17048
rect 12299 17017 12311 17020
rect 12253 17011 12311 17017
rect 12618 17008 12624 17020
rect 12676 17008 12682 17060
rect 15105 17051 15163 17057
rect 15105 17017 15117 17051
rect 15151 17048 15163 17051
rect 15470 17048 15476 17060
rect 15151 17020 15476 17048
rect 15151 17017 15163 17020
rect 15105 17011 15163 17017
rect 15470 17008 15476 17020
rect 15528 17008 15534 17060
rect 15933 17051 15991 17057
rect 15933 17017 15945 17051
rect 15979 17017 15991 17051
rect 15933 17011 15991 17017
rect 9214 16980 9220 16992
rect 9175 16952 9220 16980
rect 9214 16940 9220 16952
rect 9272 16940 9278 16992
rect 11054 16980 11060 16992
rect 11015 16952 11060 16980
rect 11054 16940 11060 16952
rect 11112 16940 11118 16992
rect 11609 16983 11667 16989
rect 11609 16949 11621 16983
rect 11655 16980 11667 16983
rect 11698 16980 11704 16992
rect 11655 16952 11704 16980
rect 11655 16949 11667 16952
rect 11609 16943 11667 16949
rect 11698 16940 11704 16952
rect 11756 16980 11762 16992
rect 11882 16980 11888 16992
rect 11756 16952 11888 16980
rect 11756 16940 11762 16952
rect 11882 16940 11888 16952
rect 11940 16940 11946 16992
rect 15381 16983 15439 16989
rect 15381 16949 15393 16983
rect 15427 16980 15439 16983
rect 15562 16980 15568 16992
rect 15427 16952 15568 16980
rect 15427 16949 15439 16952
rect 15381 16943 15439 16949
rect 15562 16940 15568 16952
rect 15620 16980 15626 16992
rect 15948 16980 15976 17011
rect 19242 17008 19248 17060
rect 19300 17048 19306 17060
rect 20257 17051 20315 17057
rect 20257 17048 20269 17051
rect 19300 17020 20269 17048
rect 19300 17008 19306 17020
rect 20257 17017 20269 17020
rect 20303 17048 20315 17051
rect 20762 17051 20820 17057
rect 20762 17048 20774 17051
rect 20303 17020 20774 17048
rect 20303 17017 20315 17020
rect 20257 17011 20315 17017
rect 20762 17017 20774 17020
rect 20808 17048 20820 17051
rect 21266 17048 21272 17060
rect 20808 17020 21272 17048
rect 20808 17017 20820 17020
rect 20762 17011 20820 17017
rect 21266 17008 21272 17020
rect 21324 17048 21330 17060
rect 21637 17051 21695 17057
rect 21637 17048 21649 17051
rect 21324 17020 21649 17048
rect 21324 17008 21330 17020
rect 21637 17017 21649 17020
rect 21683 17017 21695 17051
rect 23750 17048 23756 17060
rect 23711 17020 23756 17048
rect 21637 17011 21695 17017
rect 23750 17008 23756 17020
rect 23808 17008 23814 17060
rect 23845 17051 23903 17057
rect 23845 17017 23857 17051
rect 23891 17017 23903 17051
rect 25590 17048 25596 17060
rect 25551 17020 25596 17048
rect 23845 17011 23903 17017
rect 17034 16980 17040 16992
rect 15620 16952 15976 16980
rect 16995 16952 17040 16980
rect 15620 16940 15626 16952
rect 17034 16940 17040 16952
rect 17092 16940 17098 16992
rect 17865 16983 17923 16989
rect 17865 16949 17877 16983
rect 17911 16980 17923 16983
rect 18322 16980 18328 16992
rect 17911 16952 18328 16980
rect 17911 16949 17923 16952
rect 17865 16943 17923 16949
rect 18322 16940 18328 16952
rect 18380 16980 18386 16992
rect 18417 16983 18475 16989
rect 18417 16980 18429 16983
rect 18380 16952 18429 16980
rect 18380 16940 18386 16952
rect 18417 16949 18429 16952
rect 18463 16980 18475 16983
rect 19260 16980 19288 17008
rect 18463 16952 19288 16980
rect 23477 16983 23535 16989
rect 18463 16949 18475 16952
rect 18417 16943 18475 16949
rect 23477 16949 23489 16983
rect 23523 16980 23535 16983
rect 23566 16980 23572 16992
rect 23523 16952 23572 16980
rect 23523 16949 23535 16952
rect 23477 16943 23535 16949
rect 23566 16940 23572 16952
rect 23624 16980 23630 16992
rect 23860 16980 23888 17011
rect 25590 17008 25596 17020
rect 25648 17008 25654 17060
rect 25682 17008 25688 17060
rect 25740 17048 25746 17060
rect 25740 17020 25785 17048
rect 25740 17008 25746 17020
rect 26786 16980 26792 16992
rect 23624 16952 26792 16980
rect 23624 16940 23630 16952
rect 26786 16940 26792 16952
rect 26844 16940 26850 16992
rect 27154 16940 27160 16992
rect 27212 16980 27218 16992
rect 27341 16983 27399 16989
rect 27341 16980 27353 16983
rect 27212 16952 27353 16980
rect 27212 16940 27218 16952
rect 27341 16949 27353 16952
rect 27387 16980 27399 16983
rect 27540 16980 27568 17079
rect 27614 17076 27620 17128
rect 27672 17116 27678 17128
rect 27985 17119 28043 17125
rect 27985 17116 27997 17119
rect 27672 17088 27997 17116
rect 27672 17076 27678 17088
rect 27985 17085 27997 17088
rect 28031 17085 28043 17119
rect 27985 17079 28043 17085
rect 29178 17076 29184 17128
rect 29236 17116 29242 17128
rect 29308 17119 29366 17125
rect 29308 17116 29320 17119
rect 29236 17088 29320 17116
rect 29236 17076 29242 17088
rect 29308 17085 29320 17088
rect 29354 17085 29366 17119
rect 29308 17079 29366 17085
rect 33134 17076 33140 17128
rect 33192 17076 33198 17128
rect 34422 17076 34428 17128
rect 34480 17116 34486 17128
rect 34701 17119 34759 17125
rect 34701 17116 34713 17119
rect 34480 17088 34713 17116
rect 34480 17076 34486 17088
rect 34701 17085 34713 17088
rect 34747 17116 34759 17119
rect 35069 17119 35127 17125
rect 35069 17116 35081 17119
rect 34747 17088 35081 17116
rect 34747 17085 34759 17088
rect 34701 17079 34759 17085
rect 35069 17085 35081 17088
rect 35115 17085 35127 17119
rect 35069 17079 35127 17085
rect 35250 17076 35256 17128
rect 35308 17116 35314 17128
rect 35529 17119 35587 17125
rect 35529 17116 35541 17119
rect 35308 17088 35541 17116
rect 35308 17076 35314 17088
rect 35529 17085 35541 17088
rect 35575 17085 35587 17119
rect 35529 17079 35587 17085
rect 37550 17076 37556 17128
rect 37608 17116 37614 17128
rect 38396 17116 38424 17212
rect 39209 17187 39267 17193
rect 39209 17153 39221 17187
rect 39255 17184 39267 17187
rect 41046 17184 41052 17196
rect 39255 17156 41052 17184
rect 39255 17153 39267 17156
rect 39209 17147 39267 17153
rect 41046 17144 41052 17156
rect 41104 17184 41110 17196
rect 41877 17187 41935 17193
rect 41877 17184 41889 17187
rect 41104 17156 41889 17184
rect 41104 17144 41110 17156
rect 41877 17153 41889 17156
rect 41923 17153 41935 17187
rect 41877 17147 41935 17153
rect 38473 17119 38531 17125
rect 38473 17116 38485 17119
rect 37608 17088 38485 17116
rect 37608 17076 37614 17088
rect 38473 17085 38485 17088
rect 38519 17085 38531 17119
rect 38473 17079 38531 17085
rect 38562 17076 38568 17128
rect 38620 17116 38626 17128
rect 38933 17119 38991 17125
rect 38933 17116 38945 17119
rect 38620 17088 38945 17116
rect 38620 17076 38626 17088
rect 38933 17085 38945 17088
rect 38979 17085 38991 17119
rect 42426 17116 42432 17128
rect 42387 17088 42432 17116
rect 38933 17079 38991 17085
rect 42426 17076 42432 17088
rect 42484 17076 42490 17128
rect 30101 17051 30159 17057
rect 30101 17017 30113 17051
rect 30147 17048 30159 17051
rect 30282 17048 30288 17060
rect 30147 17020 30288 17048
rect 30147 17017 30159 17020
rect 30101 17011 30159 17017
rect 30282 17008 30288 17020
rect 30340 17048 30346 17060
rect 30340 17020 31064 17048
rect 30340 17008 30346 17020
rect 27798 16980 27804 16992
rect 27387 16952 27568 16980
rect 27759 16952 27804 16980
rect 27387 16949 27399 16952
rect 27341 16943 27399 16949
rect 27798 16940 27804 16952
rect 27856 16940 27862 16992
rect 28626 16980 28632 16992
rect 28587 16952 28632 16980
rect 28626 16940 28632 16952
rect 28684 16940 28690 16992
rect 31036 16980 31064 17020
rect 31202 17008 31208 17060
rect 31260 17048 31266 17060
rect 31297 17051 31355 17057
rect 31297 17048 31309 17051
rect 31260 17020 31309 17048
rect 31260 17008 31266 17020
rect 31297 17017 31309 17020
rect 31343 17017 31355 17051
rect 33152 17048 33180 17076
rect 33318 17048 33324 17060
rect 31297 17011 31355 17017
rect 31404 17020 33180 17048
rect 33279 17020 33324 17048
rect 31404 16980 31432 17020
rect 33318 17008 33324 17020
rect 33376 17008 33382 17060
rect 33413 17051 33471 17057
rect 33413 17017 33425 17051
rect 33459 17048 33471 17051
rect 33594 17048 33600 17060
rect 33459 17020 33600 17048
rect 33459 17017 33471 17020
rect 33413 17011 33471 17017
rect 31036 16952 31432 16980
rect 33137 16983 33195 16989
rect 33137 16949 33149 16983
rect 33183 16980 33195 16983
rect 33428 16980 33456 17011
rect 33594 17008 33600 17020
rect 33652 17008 33658 17060
rect 35802 17048 35808 17060
rect 35763 17020 35808 17048
rect 35802 17008 35808 17020
rect 35860 17008 35866 17060
rect 36173 17051 36231 17057
rect 36173 17017 36185 17051
rect 36219 17048 36231 17051
rect 36817 17051 36875 17057
rect 36817 17048 36829 17051
rect 36219 17020 36829 17048
rect 36219 17017 36231 17020
rect 36173 17011 36231 17017
rect 36817 17017 36829 17020
rect 36863 17048 36875 17051
rect 36998 17048 37004 17060
rect 36863 17020 37004 17048
rect 36863 17017 36875 17020
rect 36817 17011 36875 17017
rect 36998 17008 37004 17020
rect 37056 17008 37062 17060
rect 40586 17048 40592 17060
rect 40547 17020 40592 17048
rect 40586 17008 40592 17020
rect 40644 17008 40650 17060
rect 42766 17057 42794 17292
rect 43254 17280 43260 17292
rect 43312 17280 43318 17332
rect 43349 17323 43407 17329
rect 43349 17289 43361 17323
rect 43395 17320 43407 17323
rect 43530 17320 43536 17332
rect 43395 17292 43536 17320
rect 43395 17289 43407 17292
rect 43349 17283 43407 17289
rect 43530 17280 43536 17292
rect 43588 17320 43594 17332
rect 43625 17323 43683 17329
rect 43625 17320 43637 17323
rect 43588 17292 43637 17320
rect 43588 17280 43594 17292
rect 43625 17289 43637 17292
rect 43671 17320 43683 17323
rect 44358 17320 44364 17332
rect 43671 17292 44364 17320
rect 43671 17289 43683 17292
rect 43625 17283 43683 17289
rect 44358 17280 44364 17292
rect 44416 17280 44422 17332
rect 45186 17320 45192 17332
rect 45147 17292 45192 17320
rect 45186 17280 45192 17292
rect 45244 17280 45250 17332
rect 43714 17144 43720 17196
rect 43772 17184 43778 17196
rect 44545 17187 44603 17193
rect 44545 17184 44557 17187
rect 43772 17156 44557 17184
rect 43772 17144 43778 17156
rect 44545 17153 44557 17156
rect 44591 17153 44603 17187
rect 44545 17147 44603 17153
rect 40681 17051 40739 17057
rect 40681 17017 40693 17051
rect 40727 17017 40739 17051
rect 40681 17011 40739 17017
rect 42751 17051 42809 17057
rect 42751 17017 42763 17051
rect 42797 17017 42809 17051
rect 42751 17011 42809 17017
rect 44269 17051 44327 17057
rect 44269 17017 44281 17051
rect 44315 17017 44327 17051
rect 44269 17011 44327 17017
rect 33183 16952 33456 16980
rect 33183 16949 33195 16952
rect 33137 16943 33195 16949
rect 40310 16940 40316 16992
rect 40368 16980 40374 16992
rect 40696 16980 40724 17011
rect 40368 16952 40724 16980
rect 40368 16940 40374 16952
rect 43806 16940 43812 16992
rect 43864 16980 43870 16992
rect 43993 16983 44051 16989
rect 43993 16980 44005 16983
rect 43864 16952 44005 16980
rect 43864 16940 43870 16952
rect 43993 16949 44005 16952
rect 44039 16980 44051 16983
rect 44284 16980 44312 17011
rect 44358 17008 44364 17060
rect 44416 17048 44422 17060
rect 44416 17020 44461 17048
rect 44416 17008 44422 17020
rect 44039 16952 44312 16980
rect 44039 16949 44051 16952
rect 43993 16943 44051 16949
rect 1104 16890 48852 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 48852 16890
rect 1104 16816 48852 16838
rect 10318 16776 10324 16788
rect 10279 16748 10324 16776
rect 10318 16736 10324 16748
rect 10376 16736 10382 16788
rect 10870 16776 10876 16788
rect 10831 16748 10876 16776
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 14274 16736 14280 16788
rect 14332 16776 14338 16788
rect 14369 16779 14427 16785
rect 14369 16776 14381 16779
rect 14332 16748 14381 16776
rect 14332 16736 14338 16748
rect 14369 16745 14381 16748
rect 14415 16745 14427 16779
rect 15102 16776 15108 16788
rect 15063 16748 15108 16776
rect 14369 16739 14427 16745
rect 15102 16736 15108 16748
rect 15160 16736 15166 16788
rect 18598 16776 18604 16788
rect 18559 16748 18604 16776
rect 18598 16736 18604 16748
rect 18656 16776 18662 16788
rect 18877 16779 18935 16785
rect 18877 16776 18889 16779
rect 18656 16748 18889 16776
rect 18656 16736 18662 16748
rect 18877 16745 18889 16748
rect 18923 16745 18935 16779
rect 20438 16776 20444 16788
rect 20399 16748 20444 16776
rect 18877 16739 18935 16745
rect 20438 16736 20444 16748
rect 20496 16736 20502 16788
rect 23198 16776 23204 16788
rect 23032 16748 23204 16776
rect 12710 16708 12716 16720
rect 12671 16680 12716 16708
rect 12710 16668 12716 16680
rect 12768 16668 12774 16720
rect 15470 16708 15476 16720
rect 15431 16680 15476 16708
rect 15470 16668 15476 16680
rect 15528 16668 15534 16720
rect 16022 16708 16028 16720
rect 15983 16680 16028 16708
rect 16022 16668 16028 16680
rect 16080 16668 16086 16720
rect 16574 16668 16580 16720
rect 16632 16708 16638 16720
rect 17037 16711 17095 16717
rect 17037 16708 17049 16711
rect 16632 16680 17049 16708
rect 16632 16668 16638 16680
rect 17037 16677 17049 16680
rect 17083 16708 17095 16711
rect 17402 16708 17408 16720
rect 17083 16680 17408 16708
rect 17083 16677 17095 16680
rect 17037 16671 17095 16677
rect 17402 16668 17408 16680
rect 17460 16668 17466 16720
rect 22465 16711 22523 16717
rect 22465 16677 22477 16711
rect 22511 16708 22523 16711
rect 22830 16708 22836 16720
rect 22511 16680 22836 16708
rect 22511 16677 22523 16680
rect 22465 16671 22523 16677
rect 22830 16668 22836 16680
rect 22888 16668 22894 16720
rect 23032 16717 23060 16748
rect 23198 16736 23204 16748
rect 23256 16776 23262 16788
rect 23293 16779 23351 16785
rect 23293 16776 23305 16779
rect 23256 16748 23305 16776
rect 23256 16736 23262 16748
rect 23293 16745 23305 16748
rect 23339 16745 23351 16779
rect 23750 16776 23756 16788
rect 23711 16748 23756 16776
rect 23293 16739 23351 16745
rect 23750 16736 23756 16748
rect 23808 16736 23814 16788
rect 24762 16776 24768 16788
rect 24723 16748 24768 16776
rect 24762 16736 24768 16748
rect 24820 16736 24826 16788
rect 28810 16776 28816 16788
rect 28771 16748 28816 16776
rect 28810 16736 28816 16748
rect 28868 16736 28874 16788
rect 31202 16776 31208 16788
rect 31163 16748 31208 16776
rect 31202 16736 31208 16748
rect 31260 16736 31266 16788
rect 32631 16779 32689 16785
rect 32631 16745 32643 16779
rect 32677 16776 32689 16779
rect 33318 16776 33324 16788
rect 32677 16748 33324 16776
rect 32677 16745 32689 16748
rect 32631 16739 32689 16745
rect 33318 16736 33324 16748
rect 33376 16736 33382 16788
rect 34146 16776 34152 16788
rect 33612 16748 34152 16776
rect 23017 16711 23075 16717
rect 23017 16677 23029 16711
rect 23063 16677 23075 16711
rect 25038 16708 25044 16720
rect 24999 16680 25044 16708
rect 23017 16671 23075 16677
rect 25038 16668 25044 16680
rect 25096 16668 25102 16720
rect 28255 16711 28313 16717
rect 28255 16677 28267 16711
rect 28301 16708 28313 16711
rect 28534 16708 28540 16720
rect 28301 16680 28540 16708
rect 28301 16677 28313 16680
rect 28255 16671 28313 16677
rect 28534 16668 28540 16680
rect 28592 16668 28598 16720
rect 33410 16668 33416 16720
rect 33468 16708 33474 16720
rect 33612 16717 33640 16748
rect 34146 16736 34152 16748
rect 34204 16736 34210 16788
rect 34514 16736 34520 16788
rect 34572 16776 34578 16788
rect 35069 16779 35127 16785
rect 35069 16776 35081 16779
rect 34572 16748 35081 16776
rect 34572 16736 34578 16748
rect 35069 16745 35081 16748
rect 35115 16776 35127 16779
rect 35250 16776 35256 16788
rect 35115 16748 35256 16776
rect 35115 16745 35127 16748
rect 35069 16739 35127 16745
rect 35250 16736 35256 16748
rect 35308 16736 35314 16788
rect 35434 16776 35440 16788
rect 35395 16748 35440 16776
rect 35434 16736 35440 16748
rect 35492 16736 35498 16788
rect 36817 16779 36875 16785
rect 36817 16745 36829 16779
rect 36863 16776 36875 16779
rect 36998 16776 37004 16788
rect 36863 16748 37004 16776
rect 36863 16745 36875 16748
rect 36817 16739 36875 16745
rect 36998 16736 37004 16748
rect 37056 16736 37062 16788
rect 37366 16736 37372 16788
rect 37424 16776 37430 16788
rect 37875 16779 37933 16785
rect 37875 16776 37887 16779
rect 37424 16748 37887 16776
rect 37424 16736 37430 16748
rect 37875 16745 37887 16748
rect 37921 16745 37933 16779
rect 37875 16739 37933 16745
rect 38197 16779 38255 16785
rect 38197 16745 38209 16779
rect 38243 16776 38255 16779
rect 38562 16776 38568 16788
rect 38243 16748 38568 16776
rect 38243 16745 38255 16748
rect 38197 16739 38255 16745
rect 38562 16736 38568 16748
rect 38620 16736 38626 16788
rect 40586 16736 40592 16788
rect 40644 16776 40650 16788
rect 40865 16779 40923 16785
rect 40865 16776 40877 16779
rect 40644 16748 40877 16776
rect 40644 16736 40650 16748
rect 40865 16745 40877 16748
rect 40911 16745 40923 16779
rect 42426 16776 42432 16788
rect 42387 16748 42432 16776
rect 40865 16739 40923 16745
rect 42426 16736 42432 16748
rect 42484 16736 42490 16788
rect 33597 16711 33655 16717
rect 33597 16708 33609 16711
rect 33468 16680 33609 16708
rect 33468 16668 33474 16680
rect 33597 16677 33609 16680
rect 33643 16677 33655 16711
rect 33597 16671 33655 16677
rect 33689 16711 33747 16717
rect 33689 16677 33701 16711
rect 33735 16708 33747 16711
rect 34238 16708 34244 16720
rect 33735 16680 34244 16708
rect 33735 16677 33747 16680
rect 33689 16671 33747 16677
rect 34238 16668 34244 16680
rect 34296 16668 34302 16720
rect 35986 16668 35992 16720
rect 36044 16708 36050 16720
rect 36218 16711 36276 16717
rect 36218 16708 36230 16711
rect 36044 16680 36230 16708
rect 36044 16668 36050 16680
rect 36218 16677 36230 16680
rect 36264 16677 36276 16711
rect 37016 16708 37044 16736
rect 38286 16708 38292 16720
rect 37016 16680 38292 16708
rect 36218 16671 36276 16677
rect 38286 16668 38292 16680
rect 38344 16668 38350 16720
rect 38580 16708 38608 16736
rect 41230 16708 41236 16720
rect 38580 16680 39896 16708
rect 41191 16680 41236 16708
rect 39868 16652 39896 16680
rect 41230 16668 41236 16680
rect 41288 16668 41294 16720
rect 43530 16717 43536 16720
rect 43165 16711 43223 16717
rect 43165 16677 43177 16711
rect 43211 16708 43223 16711
rect 43510 16711 43536 16717
rect 43510 16708 43522 16711
rect 43211 16680 43522 16708
rect 43211 16677 43223 16680
rect 43165 16671 43223 16677
rect 43510 16677 43522 16680
rect 43510 16671 43536 16677
rect 43530 16668 43536 16671
rect 43588 16668 43594 16720
rect 9306 16600 9312 16652
rect 9364 16640 9370 16652
rect 9858 16640 9864 16652
rect 9364 16612 9864 16640
rect 9364 16600 9370 16612
rect 9858 16600 9864 16612
rect 9916 16640 9922 16652
rect 9953 16643 10011 16649
rect 9953 16640 9965 16643
rect 9916 16612 9965 16640
rect 9916 16600 9922 16612
rect 9953 16609 9965 16612
rect 9999 16609 10011 16643
rect 9953 16603 10011 16609
rect 14185 16643 14243 16649
rect 14185 16609 14197 16643
rect 14231 16640 14243 16643
rect 14458 16640 14464 16652
rect 14231 16612 14464 16640
rect 14231 16609 14243 16612
rect 14185 16603 14243 16609
rect 14458 16600 14464 16612
rect 14516 16600 14522 16652
rect 18969 16643 19027 16649
rect 18969 16609 18981 16643
rect 19015 16609 19027 16643
rect 18969 16603 19027 16609
rect 12250 16532 12256 16584
rect 12308 16572 12314 16584
rect 12621 16575 12679 16581
rect 12621 16572 12633 16575
rect 12308 16544 12633 16572
rect 12308 16532 12314 16544
rect 12621 16541 12633 16544
rect 12667 16541 12679 16575
rect 12986 16572 12992 16584
rect 12947 16544 12992 16572
rect 12621 16535 12679 16541
rect 12986 16532 12992 16544
rect 13044 16532 13050 16584
rect 14918 16532 14924 16584
rect 14976 16572 14982 16584
rect 15381 16575 15439 16581
rect 15381 16572 15393 16575
rect 14976 16544 15393 16572
rect 14976 16532 14982 16544
rect 15381 16541 15393 16544
rect 15427 16572 15439 16575
rect 16942 16572 16948 16584
rect 15427 16544 16252 16572
rect 16903 16544 16948 16572
rect 15427 16541 15439 16544
rect 15381 16535 15439 16541
rect 10042 16464 10048 16516
rect 10100 16504 10106 16516
rect 14642 16504 14648 16516
rect 10100 16476 14648 16504
rect 10100 16464 10106 16476
rect 14642 16464 14648 16476
rect 14700 16464 14706 16516
rect 16224 16504 16252 16544
rect 16942 16532 16948 16544
rect 17000 16532 17006 16584
rect 17126 16532 17132 16584
rect 17184 16572 17190 16584
rect 17221 16575 17279 16581
rect 17221 16572 17233 16575
rect 17184 16544 17233 16572
rect 17184 16532 17190 16544
rect 17221 16541 17233 16544
rect 17267 16541 17279 16575
rect 18984 16572 19012 16603
rect 19058 16600 19064 16652
rect 19116 16640 19122 16652
rect 19245 16643 19303 16649
rect 19245 16640 19257 16643
rect 19116 16612 19257 16640
rect 19116 16600 19122 16612
rect 19245 16609 19257 16612
rect 19291 16609 19303 16643
rect 19245 16603 19303 16609
rect 21269 16643 21327 16649
rect 21269 16609 21281 16643
rect 21315 16640 21327 16643
rect 21358 16640 21364 16652
rect 21315 16612 21364 16640
rect 21315 16609 21327 16612
rect 21269 16603 21327 16609
rect 21358 16600 21364 16612
rect 21416 16600 21422 16652
rect 23382 16600 23388 16652
rect 23440 16640 23446 16652
rect 23880 16643 23938 16649
rect 23880 16640 23892 16643
rect 23440 16612 23892 16640
rect 23440 16600 23446 16612
rect 23880 16609 23892 16612
rect 23926 16609 23938 16643
rect 23880 16603 23938 16609
rect 26418 16600 26424 16652
rect 26476 16640 26482 16652
rect 26548 16643 26606 16649
rect 26548 16640 26560 16643
rect 26476 16612 26560 16640
rect 26476 16600 26482 16612
rect 26548 16609 26560 16612
rect 26594 16609 26606 16643
rect 26548 16603 26606 16609
rect 27798 16600 27804 16652
rect 27856 16640 27862 16652
rect 27893 16643 27951 16649
rect 27893 16640 27905 16643
rect 27856 16612 27905 16640
rect 27856 16600 27862 16612
rect 27893 16609 27905 16612
rect 27939 16609 27951 16643
rect 29638 16640 29644 16652
rect 29599 16612 29644 16640
rect 27893 16603 27951 16609
rect 29638 16600 29644 16612
rect 29696 16600 29702 16652
rect 29730 16600 29736 16652
rect 29788 16640 29794 16652
rect 30101 16643 30159 16649
rect 30101 16640 30113 16643
rect 29788 16612 30113 16640
rect 29788 16600 29794 16612
rect 30101 16609 30113 16612
rect 30147 16640 30159 16643
rect 30466 16640 30472 16652
rect 30147 16612 30472 16640
rect 30147 16609 30159 16612
rect 30101 16603 30159 16609
rect 30466 16600 30472 16612
rect 30524 16600 30530 16652
rect 32560 16643 32618 16649
rect 32560 16609 32572 16643
rect 32606 16640 32618 16643
rect 32950 16640 32956 16652
rect 32606 16612 32956 16640
rect 32606 16609 32618 16612
rect 32560 16603 32618 16609
rect 32950 16600 32956 16612
rect 33008 16600 33014 16652
rect 37642 16600 37648 16652
rect 37700 16640 37706 16652
rect 37772 16643 37830 16649
rect 37772 16640 37784 16643
rect 37700 16612 37784 16640
rect 37700 16600 37706 16612
rect 37772 16609 37784 16612
rect 37818 16609 37830 16643
rect 39390 16640 39396 16652
rect 39351 16612 39396 16640
rect 37772 16603 37830 16609
rect 39390 16600 39396 16612
rect 39448 16600 39454 16652
rect 39850 16640 39856 16652
rect 39763 16612 39856 16640
rect 39850 16600 39856 16612
rect 39908 16600 39914 16652
rect 22373 16575 22431 16581
rect 18984 16544 19288 16572
rect 17221 16535 17279 16541
rect 17144 16504 17172 16532
rect 19260 16516 19288 16544
rect 22373 16541 22385 16575
rect 22419 16541 22431 16575
rect 22373 16535 22431 16541
rect 24949 16575 25007 16581
rect 24949 16541 24961 16575
rect 24995 16541 25007 16575
rect 25590 16572 25596 16584
rect 25551 16544 25596 16572
rect 24949 16535 25007 16541
rect 16224 16476 17172 16504
rect 17236 16476 18736 16504
rect 11330 16396 11336 16448
rect 11388 16436 11394 16448
rect 11517 16439 11575 16445
rect 11517 16436 11529 16439
rect 11388 16408 11529 16436
rect 11388 16396 11394 16408
rect 11517 16405 11529 16408
rect 11563 16405 11575 16439
rect 14660 16436 14688 16464
rect 17236 16436 17264 16476
rect 14660 16408 17264 16436
rect 18141 16439 18199 16445
rect 11517 16399 11575 16405
rect 18141 16405 18153 16439
rect 18187 16436 18199 16439
rect 18598 16436 18604 16448
rect 18187 16408 18604 16436
rect 18187 16405 18199 16408
rect 18141 16399 18199 16405
rect 18598 16396 18604 16408
rect 18656 16396 18662 16448
rect 18708 16436 18736 16476
rect 19242 16464 19248 16516
rect 19300 16464 19306 16516
rect 21407 16507 21465 16513
rect 21407 16473 21419 16507
rect 21453 16504 21465 16507
rect 22278 16504 22284 16516
rect 21453 16476 22284 16504
rect 21453 16473 21465 16476
rect 21407 16467 21465 16473
rect 22278 16464 22284 16476
rect 22336 16504 22342 16516
rect 22388 16504 22416 16535
rect 23983 16507 24041 16513
rect 23983 16504 23995 16507
rect 22336 16476 22416 16504
rect 22526 16476 23995 16504
rect 22336 16464 22342 16476
rect 19889 16439 19947 16445
rect 19889 16436 19901 16439
rect 18708 16408 19901 16436
rect 19889 16405 19901 16408
rect 19935 16436 19947 16439
rect 20254 16436 20260 16448
rect 19935 16408 20260 16436
rect 19935 16405 19947 16408
rect 19889 16399 19947 16405
rect 20254 16396 20260 16408
rect 20312 16396 20318 16448
rect 20622 16396 20628 16448
rect 20680 16436 20686 16448
rect 21085 16439 21143 16445
rect 21085 16436 21097 16439
rect 20680 16408 21097 16436
rect 20680 16396 20686 16408
rect 21085 16405 21097 16408
rect 21131 16405 21143 16439
rect 22094 16436 22100 16448
rect 22007 16408 22100 16436
rect 21085 16399 21143 16405
rect 22094 16396 22100 16408
rect 22152 16436 22158 16448
rect 22526 16436 22554 16476
rect 23983 16473 23995 16476
rect 24029 16473 24041 16507
rect 24964 16504 24992 16535
rect 25590 16532 25596 16544
rect 25648 16532 25654 16584
rect 30190 16572 30196 16584
rect 30151 16544 30196 16572
rect 30190 16532 30196 16544
rect 30248 16532 30254 16584
rect 33870 16572 33876 16584
rect 33831 16544 33876 16572
rect 33870 16532 33876 16544
rect 33928 16532 33934 16584
rect 35894 16572 35900 16584
rect 35855 16544 35900 16572
rect 35894 16532 35900 16544
rect 35952 16532 35958 16584
rect 40129 16575 40187 16581
rect 40129 16541 40141 16575
rect 40175 16572 40187 16575
rect 40494 16572 40500 16584
rect 40175 16544 40500 16572
rect 40175 16541 40187 16544
rect 40129 16535 40187 16541
rect 40494 16532 40500 16544
rect 40552 16532 40558 16584
rect 41138 16572 41144 16584
rect 41099 16544 41144 16572
rect 41138 16532 41144 16544
rect 41196 16532 41202 16584
rect 41322 16532 41328 16584
rect 41380 16572 41386 16584
rect 41417 16575 41475 16581
rect 41417 16572 41429 16575
rect 41380 16544 41429 16572
rect 41380 16532 41386 16544
rect 41417 16541 41429 16544
rect 41463 16541 41475 16575
rect 43438 16572 43444 16584
rect 43399 16544 43444 16572
rect 41417 16535 41475 16541
rect 43438 16532 43444 16544
rect 43496 16532 43502 16584
rect 43717 16575 43775 16581
rect 43717 16572 43729 16575
rect 43548 16544 43729 16572
rect 25406 16504 25412 16516
rect 24964 16476 25412 16504
rect 23983 16467 24041 16473
rect 25406 16464 25412 16476
rect 25464 16504 25470 16516
rect 26651 16507 26709 16513
rect 26651 16504 26663 16507
rect 25464 16476 26663 16504
rect 25464 16464 25470 16476
rect 26651 16473 26663 16476
rect 26697 16473 26709 16507
rect 26651 16467 26709 16473
rect 34054 16464 34060 16516
rect 34112 16504 34118 16516
rect 41046 16504 41052 16516
rect 34112 16476 41052 16504
rect 34112 16464 34118 16476
rect 41046 16464 41052 16476
rect 41104 16464 41110 16516
rect 41156 16504 41184 16532
rect 43548 16504 43576 16544
rect 43717 16541 43729 16544
rect 43763 16541 43775 16575
rect 43717 16535 43775 16541
rect 41156 16476 43576 16504
rect 22152 16408 22554 16436
rect 22152 16396 22158 16408
rect 23290 16396 23296 16448
rect 23348 16436 23354 16448
rect 23750 16436 23756 16448
rect 23348 16408 23756 16436
rect 23348 16396 23354 16408
rect 23750 16396 23756 16408
rect 23808 16396 23814 16448
rect 24302 16436 24308 16448
rect 24263 16408 24308 16436
rect 24302 16396 24308 16408
rect 24360 16396 24366 16448
rect 27522 16436 27528 16448
rect 27483 16408 27528 16436
rect 27522 16396 27528 16408
rect 27580 16396 27586 16448
rect 29178 16396 29184 16448
rect 29236 16436 29242 16448
rect 29273 16439 29331 16445
rect 29273 16436 29285 16439
rect 29236 16408 29285 16436
rect 29236 16396 29242 16408
rect 29273 16405 29285 16408
rect 29319 16405 29331 16439
rect 37090 16436 37096 16448
rect 37051 16408 37096 16436
rect 29273 16399 29331 16405
rect 37090 16396 37096 16408
rect 37148 16396 37154 16448
rect 39022 16436 39028 16448
rect 38983 16408 39028 16436
rect 39022 16396 39028 16408
rect 39080 16396 39086 16448
rect 1104 16346 48852 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 48852 16346
rect 1104 16272 48852 16294
rect 9306 16232 9312 16244
rect 9267 16204 9312 16232
rect 9306 16192 9312 16204
rect 9364 16192 9370 16244
rect 9677 16235 9735 16241
rect 9677 16201 9689 16235
rect 9723 16232 9735 16235
rect 11054 16232 11060 16244
rect 9723 16204 11060 16232
rect 9723 16201 9735 16204
rect 9677 16195 9735 16201
rect 9851 16037 9879 16204
rect 11054 16192 11060 16204
rect 11112 16192 11118 16244
rect 11698 16232 11704 16244
rect 11440 16204 11704 16232
rect 9907 16167 9965 16173
rect 9907 16133 9919 16167
rect 9953 16164 9965 16167
rect 11330 16164 11336 16176
rect 9953 16136 11336 16164
rect 9953 16133 9965 16136
rect 9907 16127 9965 16133
rect 11330 16124 11336 16136
rect 11388 16124 11394 16176
rect 11440 16173 11468 16204
rect 11698 16192 11704 16204
rect 11756 16232 11762 16244
rect 12250 16232 12256 16244
rect 11756 16204 12256 16232
rect 11756 16192 11762 16204
rect 12250 16192 12256 16204
rect 12308 16192 12314 16244
rect 12710 16232 12716 16244
rect 12671 16204 12716 16232
rect 12710 16192 12716 16204
rect 12768 16232 12774 16244
rect 12989 16235 13047 16241
rect 12989 16232 13001 16235
rect 12768 16204 13001 16232
rect 12768 16192 12774 16204
rect 12989 16201 13001 16204
rect 13035 16232 13047 16235
rect 13354 16232 13360 16244
rect 13035 16204 13360 16232
rect 13035 16201 13047 16204
rect 12989 16195 13047 16201
rect 13354 16192 13360 16204
rect 13412 16192 13418 16244
rect 14277 16235 14335 16241
rect 14277 16201 14289 16235
rect 14323 16232 14335 16235
rect 14458 16232 14464 16244
rect 14323 16204 14464 16232
rect 14323 16201 14335 16204
rect 14277 16195 14335 16201
rect 14458 16192 14464 16204
rect 14516 16192 14522 16244
rect 14918 16232 14924 16244
rect 14879 16204 14924 16232
rect 14918 16192 14924 16204
rect 14976 16192 14982 16244
rect 15470 16232 15476 16244
rect 15028 16204 15476 16232
rect 11425 16167 11483 16173
rect 11425 16133 11437 16167
rect 11471 16133 11483 16167
rect 11425 16127 11483 16133
rect 13262 16056 13268 16108
rect 13320 16096 13326 16108
rect 13541 16099 13599 16105
rect 13541 16096 13553 16099
rect 13320 16068 13553 16096
rect 13320 16056 13326 16068
rect 13541 16065 13553 16068
rect 13587 16065 13599 16099
rect 13541 16059 13599 16065
rect 9836 16031 9894 16037
rect 9836 15997 9848 16031
rect 9882 15997 9894 16031
rect 9836 15991 9894 15997
rect 10870 15960 10876 15972
rect 10831 15932 10876 15960
rect 10870 15920 10876 15932
rect 10928 15920 10934 15972
rect 10965 15963 11023 15969
rect 10965 15929 10977 15963
rect 11011 15960 11023 15963
rect 11882 15960 11888 15972
rect 11011 15932 11888 15960
rect 11011 15929 11023 15932
rect 10965 15923 11023 15929
rect 10318 15892 10324 15904
rect 10279 15864 10324 15892
rect 10318 15852 10324 15864
rect 10376 15852 10382 15904
rect 10689 15895 10747 15901
rect 10689 15861 10701 15895
rect 10735 15892 10747 15895
rect 10980 15892 11008 15923
rect 11882 15920 11888 15932
rect 11940 15920 11946 15972
rect 13262 15960 13268 15972
rect 13223 15932 13268 15960
rect 13262 15920 13268 15932
rect 13320 15920 13326 15972
rect 13354 15920 13360 15972
rect 13412 15960 13418 15972
rect 14550 15960 14556 15972
rect 13412 15932 14556 15960
rect 13412 15920 13418 15932
rect 14550 15920 14556 15932
rect 14608 15960 14614 15972
rect 15028 15960 15056 16204
rect 15470 16192 15476 16204
rect 15528 16232 15534 16244
rect 15841 16235 15899 16241
rect 15841 16232 15853 16235
rect 15528 16204 15853 16232
rect 15528 16192 15534 16204
rect 15841 16201 15853 16204
rect 15887 16201 15899 16235
rect 17402 16232 17408 16244
rect 17363 16204 17408 16232
rect 15841 16195 15899 16201
rect 17402 16192 17408 16204
rect 17460 16192 17466 16244
rect 19797 16235 19855 16241
rect 19797 16201 19809 16235
rect 19843 16232 19855 16235
rect 19978 16232 19984 16244
rect 19843 16204 19984 16232
rect 19843 16201 19855 16204
rect 19797 16195 19855 16201
rect 19978 16192 19984 16204
rect 20036 16192 20042 16244
rect 24121 16235 24179 16241
rect 24121 16201 24133 16235
rect 24167 16232 24179 16235
rect 24394 16232 24400 16244
rect 24167 16204 24400 16232
rect 24167 16201 24179 16204
rect 24121 16195 24179 16201
rect 24394 16192 24400 16204
rect 24452 16232 24458 16244
rect 24854 16232 24860 16244
rect 24452 16204 24860 16232
rect 24452 16192 24458 16204
rect 24854 16192 24860 16204
rect 24912 16192 24918 16244
rect 25038 16192 25044 16244
rect 25096 16232 25102 16244
rect 25317 16235 25375 16241
rect 25317 16232 25329 16235
rect 25096 16204 25329 16232
rect 25096 16192 25102 16204
rect 25317 16201 25329 16204
rect 25363 16232 25375 16235
rect 27430 16232 27436 16244
rect 25363 16204 27436 16232
rect 25363 16201 25375 16204
rect 25317 16195 25375 16201
rect 27430 16192 27436 16204
rect 27488 16192 27494 16244
rect 29638 16232 29644 16244
rect 29599 16204 29644 16232
rect 29638 16192 29644 16204
rect 29696 16192 29702 16244
rect 33321 16235 33379 16241
rect 33321 16201 33333 16235
rect 33367 16232 33379 16235
rect 33410 16232 33416 16244
rect 33367 16204 33416 16232
rect 33367 16201 33379 16204
rect 33321 16195 33379 16201
rect 33410 16192 33416 16204
rect 33468 16192 33474 16244
rect 33551 16235 33609 16241
rect 33551 16201 33563 16235
rect 33597 16232 33609 16235
rect 34606 16232 34612 16244
rect 33597 16204 34612 16232
rect 33597 16201 33609 16204
rect 33551 16195 33609 16201
rect 34606 16192 34612 16204
rect 34664 16192 34670 16244
rect 35207 16235 35265 16241
rect 35207 16201 35219 16235
rect 35253 16232 35265 16235
rect 37090 16232 37096 16244
rect 35253 16204 37096 16232
rect 35253 16201 35265 16204
rect 35207 16195 35265 16201
rect 37090 16192 37096 16204
rect 37148 16192 37154 16244
rect 37642 16192 37648 16244
rect 37700 16232 37706 16244
rect 37737 16235 37795 16241
rect 37737 16232 37749 16235
rect 37700 16204 37749 16232
rect 37700 16192 37706 16204
rect 37737 16201 37749 16204
rect 37783 16201 37795 16235
rect 37737 16195 37795 16201
rect 39482 16192 39488 16244
rect 39540 16232 39546 16244
rect 40221 16235 40279 16241
rect 40221 16232 40233 16235
rect 39540 16204 40233 16232
rect 39540 16192 39546 16204
rect 40221 16201 40233 16204
rect 40267 16201 40279 16235
rect 40221 16195 40279 16201
rect 15289 16167 15347 16173
rect 15289 16133 15301 16167
rect 15335 16164 15347 16167
rect 18782 16164 18788 16176
rect 15335 16136 18788 16164
rect 15335 16133 15347 16136
rect 15289 16127 15347 16133
rect 15442 16037 15470 16136
rect 18782 16124 18788 16136
rect 18840 16124 18846 16176
rect 22922 16124 22928 16176
rect 22980 16164 22986 16176
rect 25056 16164 25084 16192
rect 22980 16136 25084 16164
rect 22980 16124 22986 16136
rect 32766 16124 32772 16176
rect 32824 16164 32830 16176
rect 35529 16167 35587 16173
rect 35529 16164 35541 16167
rect 32824 16136 35541 16164
rect 32824 16124 32830 16136
rect 35529 16133 35541 16136
rect 35575 16164 35587 16167
rect 35986 16164 35992 16176
rect 35575 16136 35992 16164
rect 35575 16133 35587 16136
rect 35529 16127 35587 16133
rect 15519 16099 15577 16105
rect 15519 16065 15531 16099
rect 15565 16096 15577 16099
rect 16942 16096 16948 16108
rect 15565 16068 16948 16096
rect 15565 16065 15577 16068
rect 15519 16059 15577 16065
rect 16942 16056 16948 16068
rect 17000 16056 17006 16108
rect 17126 16096 17132 16108
rect 17087 16068 17132 16096
rect 17126 16056 17132 16068
rect 17184 16056 17190 16108
rect 20622 16096 20628 16108
rect 20583 16068 20628 16096
rect 20622 16056 20628 16068
rect 20680 16056 20686 16108
rect 22094 16096 22100 16108
rect 22055 16068 22100 16096
rect 22094 16056 22100 16068
rect 22152 16056 22158 16108
rect 22741 16099 22799 16105
rect 22741 16065 22753 16099
rect 22787 16096 22799 16099
rect 23198 16096 23204 16108
rect 22787 16068 23204 16096
rect 22787 16065 22799 16068
rect 22741 16059 22799 16065
rect 23198 16056 23204 16068
rect 23256 16056 23262 16108
rect 25590 16056 25596 16108
rect 25648 16096 25654 16108
rect 26145 16099 26203 16105
rect 26145 16096 26157 16099
rect 25648 16068 26157 16096
rect 25648 16056 25654 16068
rect 26145 16065 26157 16068
rect 26191 16065 26203 16099
rect 26145 16059 26203 16065
rect 30101 16099 30159 16105
rect 30101 16065 30113 16099
rect 30147 16096 30159 16099
rect 30190 16096 30196 16108
rect 30147 16068 30196 16096
rect 30147 16065 30159 16068
rect 30101 16059 30159 16065
rect 30190 16056 30196 16068
rect 30248 16056 30254 16108
rect 31294 16056 31300 16108
rect 31352 16096 31358 16108
rect 31938 16096 31944 16108
rect 31352 16068 31944 16096
rect 31352 16056 31358 16068
rect 31938 16056 31944 16068
rect 31996 16056 32002 16108
rect 32585 16099 32643 16105
rect 32585 16065 32597 16099
rect 32631 16096 32643 16099
rect 33870 16096 33876 16108
rect 32631 16068 33876 16096
rect 32631 16065 32643 16068
rect 32585 16059 32643 16065
rect 33870 16056 33876 16068
rect 33928 16096 33934 16108
rect 34514 16096 34520 16108
rect 33928 16068 34520 16096
rect 33928 16056 33934 16068
rect 34514 16056 34520 16068
rect 34572 16056 34578 16108
rect 15427 16031 15485 16037
rect 15427 15997 15439 16031
rect 15473 15997 15485 16031
rect 15427 15991 15485 15997
rect 17865 16031 17923 16037
rect 17865 15997 17877 16031
rect 17911 16028 17923 16031
rect 18046 16028 18052 16040
rect 17911 16000 18052 16028
rect 17911 15997 17923 16000
rect 17865 15991 17923 15997
rect 18046 15988 18052 16000
rect 18104 15988 18110 16040
rect 18598 16028 18604 16040
rect 18511 16000 18604 16028
rect 18598 15988 18604 16000
rect 18656 16028 18662 16040
rect 19058 16028 19064 16040
rect 18656 16000 19064 16028
rect 18656 15988 18662 16000
rect 19058 15988 19064 16000
rect 19116 15988 19122 16040
rect 19978 16028 19984 16040
rect 19939 16000 19984 16028
rect 19978 15988 19984 16000
rect 20036 15988 20042 16040
rect 20254 15988 20260 16040
rect 20312 16028 20318 16040
rect 20349 16031 20407 16037
rect 20349 16028 20361 16031
rect 20312 16000 20361 16028
rect 20312 15988 20318 16000
rect 20349 15997 20361 16000
rect 20395 15997 20407 16031
rect 27617 16031 27675 16037
rect 27617 16028 27629 16031
rect 20349 15991 20407 15997
rect 27448 16000 27629 16028
rect 16482 15960 16488 15972
rect 14608 15932 15056 15960
rect 16443 15932 16488 15960
rect 14608 15920 14614 15932
rect 16482 15920 16488 15932
rect 16540 15920 16546 15972
rect 16577 15963 16635 15969
rect 16577 15929 16589 15963
rect 16623 15929 16635 15963
rect 21910 15960 21916 15972
rect 21823 15932 21916 15960
rect 16577 15923 16635 15929
rect 10735 15864 11008 15892
rect 16301 15895 16359 15901
rect 10735 15861 10747 15864
rect 10689 15855 10747 15861
rect 16301 15861 16313 15895
rect 16347 15892 16359 15895
rect 16592 15892 16620 15923
rect 21910 15920 21916 15932
rect 21968 15960 21974 15972
rect 22189 15963 22247 15969
rect 22189 15960 22201 15963
rect 21968 15932 22201 15960
rect 21968 15920 21974 15932
rect 22189 15929 22201 15932
rect 22235 15960 22247 15963
rect 22738 15960 22744 15972
rect 22235 15932 22744 15960
rect 22235 15929 22247 15932
rect 22189 15923 22247 15929
rect 22738 15920 22744 15932
rect 22796 15920 22802 15972
rect 24302 15960 24308 15972
rect 24263 15932 24308 15960
rect 24302 15920 24308 15932
rect 24360 15920 24366 15972
rect 24394 15920 24400 15972
rect 24452 15960 24458 15972
rect 24946 15960 24952 15972
rect 24452 15932 24497 15960
rect 24907 15932 24952 15960
rect 24452 15920 24458 15932
rect 24946 15920 24952 15932
rect 25004 15920 25010 15972
rect 25866 15960 25872 15972
rect 25827 15932 25872 15960
rect 25866 15920 25872 15932
rect 25924 15920 25930 15972
rect 25961 15963 26019 15969
rect 25961 15929 25973 15963
rect 26007 15960 26019 15963
rect 26326 15960 26332 15972
rect 26007 15932 26332 15960
rect 26007 15929 26019 15932
rect 25961 15923 26019 15929
rect 17034 15892 17040 15904
rect 16347 15864 17040 15892
rect 16347 15861 16359 15864
rect 16301 15855 16359 15861
rect 17034 15852 17040 15864
rect 17092 15852 17098 15904
rect 18138 15892 18144 15904
rect 18099 15864 18144 15892
rect 18138 15852 18144 15864
rect 18196 15852 18202 15904
rect 18966 15852 18972 15904
rect 19024 15892 19030 15904
rect 19153 15895 19211 15901
rect 19153 15892 19165 15895
rect 19024 15864 19165 15892
rect 19024 15852 19030 15864
rect 19153 15861 19165 15864
rect 19199 15892 19211 15895
rect 19242 15892 19248 15904
rect 19199 15864 19248 15892
rect 19199 15861 19211 15864
rect 19153 15855 19211 15861
rect 19242 15852 19248 15864
rect 19300 15852 19306 15904
rect 21358 15892 21364 15904
rect 21319 15864 21364 15892
rect 21358 15852 21364 15864
rect 21416 15852 21422 15904
rect 22922 15852 22928 15904
rect 22980 15892 22986 15904
rect 23017 15895 23075 15901
rect 23017 15892 23029 15895
rect 22980 15864 23029 15892
rect 22980 15852 22986 15864
rect 23017 15861 23029 15864
rect 23063 15861 23075 15895
rect 23382 15892 23388 15904
rect 23343 15864 23388 15892
rect 23017 15855 23075 15861
rect 23382 15852 23388 15864
rect 23440 15852 23446 15904
rect 25685 15895 25743 15901
rect 25685 15861 25697 15895
rect 25731 15892 25743 15895
rect 25976 15892 26004 15923
rect 26326 15920 26332 15932
rect 26384 15920 26390 15972
rect 25731 15864 26004 15892
rect 25731 15861 25743 15864
rect 25685 15855 25743 15861
rect 26418 15852 26424 15904
rect 26476 15892 26482 15904
rect 26789 15895 26847 15901
rect 26789 15892 26801 15895
rect 26476 15864 26801 15892
rect 26476 15852 26482 15864
rect 26789 15861 26801 15864
rect 26835 15861 26847 15895
rect 26789 15855 26847 15861
rect 27154 15852 27160 15904
rect 27212 15892 27218 15904
rect 27448 15901 27476 16000
rect 27617 15997 27629 16000
rect 27663 15997 27675 16031
rect 28074 16028 28080 16040
rect 28035 16000 28080 16028
rect 27617 15991 27675 15997
rect 28074 15988 28080 16000
rect 28132 15988 28138 16040
rect 33480 16031 33538 16037
rect 33480 15997 33492 16031
rect 33526 16028 33538 16031
rect 33965 16031 34023 16037
rect 33965 16028 33977 16031
rect 33526 16000 33977 16028
rect 33526 15997 33538 16000
rect 33480 15991 33538 15997
rect 33965 15997 33977 16000
rect 34011 16028 34023 16031
rect 34698 16028 34704 16040
rect 34011 16000 34704 16028
rect 34011 15997 34023 16000
rect 33965 15991 34023 15997
rect 34698 15988 34704 16000
rect 34756 16028 34762 16040
rect 35104 16031 35162 16037
rect 35104 16028 35116 16031
rect 34756 16000 35116 16028
rect 34756 15988 34762 16000
rect 35104 15997 35116 16000
rect 35150 15997 35162 16031
rect 35104 15991 35162 15997
rect 35728 15972 35756 16136
rect 35986 16124 35992 16136
rect 36044 16124 36050 16176
rect 39850 16164 39856 16176
rect 39811 16136 39856 16164
rect 39850 16124 39856 16136
rect 39908 16124 39914 16176
rect 35894 16056 35900 16108
rect 35952 16096 35958 16108
rect 37277 16099 37335 16105
rect 37277 16096 37289 16099
rect 35952 16068 37289 16096
rect 35952 16056 35958 16068
rect 37277 16065 37289 16068
rect 37323 16065 37335 16099
rect 37277 16059 37335 16065
rect 38197 16099 38255 16105
rect 38197 16065 38209 16099
rect 38243 16096 38255 16099
rect 39022 16096 39028 16108
rect 38243 16068 39028 16096
rect 38243 16065 38255 16068
rect 38197 16059 38255 16065
rect 39022 16056 39028 16068
rect 39080 16056 39086 16108
rect 35802 15988 35808 16040
rect 35860 16028 35866 16040
rect 36081 16031 36139 16037
rect 36081 16028 36093 16031
rect 35860 16000 36093 16028
rect 35860 15988 35866 16000
rect 36081 15997 36093 16000
rect 36127 15997 36139 16031
rect 36081 15991 36139 15997
rect 28258 15920 28264 15972
rect 28316 15960 28322 15972
rect 28353 15963 28411 15969
rect 28353 15960 28365 15963
rect 28316 15932 28365 15960
rect 28316 15920 28322 15932
rect 28353 15929 28365 15932
rect 28399 15929 28411 15963
rect 30422 15963 30480 15969
rect 30422 15960 30434 15963
rect 28353 15923 28411 15929
rect 29932 15932 30434 15960
rect 27433 15895 27491 15901
rect 27433 15892 27445 15895
rect 27212 15864 27445 15892
rect 27212 15852 27218 15864
rect 27433 15861 27445 15864
rect 27479 15861 27491 15895
rect 27433 15855 27491 15861
rect 28534 15852 28540 15904
rect 28592 15892 28598 15904
rect 29932 15901 29960 15932
rect 30422 15929 30434 15932
rect 30468 15960 30480 15963
rect 30558 15960 30564 15972
rect 30468 15932 30564 15960
rect 30468 15929 30480 15932
rect 30422 15923 30480 15929
rect 30558 15920 30564 15932
rect 30616 15960 30622 15972
rect 31754 15960 31760 15972
rect 30616 15932 31760 15960
rect 30616 15920 30622 15932
rect 31754 15920 31760 15932
rect 31812 15920 31818 15972
rect 32033 15963 32091 15969
rect 32033 15929 32045 15963
rect 32079 15929 32091 15963
rect 35710 15960 35716 15972
rect 35623 15932 35716 15960
rect 32033 15923 32091 15929
rect 28629 15895 28687 15901
rect 28629 15892 28641 15895
rect 28592 15864 28641 15892
rect 28592 15852 28598 15864
rect 28629 15861 28641 15864
rect 28675 15892 28687 15895
rect 29917 15895 29975 15901
rect 29917 15892 29929 15895
rect 28675 15864 29929 15892
rect 28675 15861 28687 15864
rect 28629 15855 28687 15861
rect 29917 15861 29929 15864
rect 29963 15861 29975 15895
rect 29917 15855 29975 15861
rect 31021 15895 31079 15901
rect 31021 15861 31033 15895
rect 31067 15892 31079 15895
rect 31665 15895 31723 15901
rect 31665 15892 31677 15895
rect 31067 15864 31677 15892
rect 31067 15861 31079 15864
rect 31021 15855 31079 15861
rect 31665 15861 31677 15864
rect 31711 15892 31723 15895
rect 32048 15892 32076 15923
rect 35710 15920 35716 15932
rect 35768 15960 35774 15972
rect 36402 15963 36460 15969
rect 36402 15960 36414 15963
rect 35768 15932 36414 15960
rect 35768 15920 35774 15932
rect 36402 15929 36414 15932
rect 36448 15929 36460 15963
rect 38286 15960 38292 15972
rect 38247 15932 38292 15960
rect 36402 15923 36460 15929
rect 38286 15920 38292 15932
rect 38344 15920 38350 15972
rect 38838 15960 38844 15972
rect 38799 15932 38844 15960
rect 38838 15920 38844 15932
rect 38896 15920 38902 15972
rect 40236 15960 40264 16195
rect 41230 16192 41236 16244
rect 41288 16232 41294 16244
rect 41417 16235 41475 16241
rect 41417 16232 41429 16235
rect 41288 16204 41429 16232
rect 41288 16192 41294 16204
rect 41417 16201 41429 16204
rect 41463 16232 41475 16235
rect 41693 16235 41751 16241
rect 41693 16232 41705 16235
rect 41463 16204 41705 16232
rect 41463 16201 41475 16204
rect 41417 16195 41475 16201
rect 41693 16201 41705 16204
rect 41739 16201 41751 16235
rect 41693 16195 41751 16201
rect 43441 16235 43499 16241
rect 43441 16201 43453 16235
rect 43487 16232 43499 16235
rect 43530 16232 43536 16244
rect 43487 16204 43536 16232
rect 43487 16201 43499 16204
rect 43441 16195 43499 16201
rect 43530 16192 43536 16204
rect 43588 16192 43594 16244
rect 41046 16124 41052 16176
rect 41104 16164 41110 16176
rect 42061 16167 42119 16173
rect 42061 16164 42073 16167
rect 41104 16136 42073 16164
rect 41104 16124 41110 16136
rect 42061 16133 42073 16136
rect 42107 16133 42119 16167
rect 42061 16127 42119 16133
rect 40494 16096 40500 16108
rect 40455 16068 40500 16096
rect 40494 16056 40500 16068
rect 40552 16056 40558 16108
rect 42076 16028 42104 16127
rect 43806 16096 43812 16108
rect 43767 16068 43812 16096
rect 43806 16056 43812 16068
rect 43864 16056 43870 16108
rect 42245 16031 42303 16037
rect 42245 16028 42257 16031
rect 42076 16000 42257 16028
rect 42245 15997 42257 16000
rect 42291 15997 42303 16031
rect 42702 16028 42708 16040
rect 42663 16000 42708 16028
rect 42245 15991 42303 15997
rect 42702 15988 42708 16000
rect 42760 15988 42766 16040
rect 40818 15963 40876 15969
rect 40818 15960 40830 15963
rect 40236 15932 40830 15960
rect 40818 15929 40830 15932
rect 40864 15960 40876 15963
rect 41046 15960 41052 15972
rect 40864 15932 41052 15960
rect 40864 15929 40876 15932
rect 40818 15923 40876 15929
rect 41046 15920 41052 15932
rect 41104 15920 41110 15972
rect 43438 15920 43444 15972
rect 43496 15960 43502 15972
rect 44269 15963 44327 15969
rect 44269 15960 44281 15963
rect 43496 15932 44281 15960
rect 43496 15920 43502 15932
rect 44269 15929 44281 15932
rect 44315 15929 44327 15963
rect 44269 15923 44327 15929
rect 32950 15892 32956 15904
rect 31711 15864 32076 15892
rect 32911 15864 32956 15892
rect 31711 15861 31723 15864
rect 31665 15855 31723 15861
rect 32950 15852 32956 15864
rect 33008 15852 33014 15904
rect 34238 15892 34244 15904
rect 34199 15864 34244 15892
rect 34238 15852 34244 15864
rect 34296 15852 34302 15904
rect 36998 15892 37004 15904
rect 36959 15864 37004 15892
rect 36998 15852 37004 15864
rect 37056 15852 37062 15904
rect 38378 15852 38384 15904
rect 38436 15892 38442 15904
rect 39390 15892 39396 15904
rect 38436 15864 39396 15892
rect 38436 15852 38442 15864
rect 39390 15852 39396 15864
rect 39448 15852 39454 15904
rect 42337 15895 42395 15901
rect 42337 15861 42349 15895
rect 42383 15892 42395 15895
rect 42426 15892 42432 15904
rect 42383 15864 42432 15892
rect 42383 15861 42395 15864
rect 42337 15855 42395 15861
rect 42426 15852 42432 15864
rect 42484 15852 42490 15904
rect 1104 15802 48852 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 48852 15802
rect 1104 15728 48852 15750
rect 13262 15648 13268 15700
rect 13320 15688 13326 15700
rect 13541 15691 13599 15697
rect 13541 15688 13553 15691
rect 13320 15660 13553 15688
rect 13320 15648 13326 15660
rect 13541 15657 13553 15660
rect 13587 15657 13599 15691
rect 13541 15651 13599 15657
rect 16942 15648 16948 15700
rect 17000 15688 17006 15700
rect 17313 15691 17371 15697
rect 17313 15688 17325 15691
rect 17000 15660 17325 15688
rect 17000 15648 17006 15660
rect 17313 15657 17325 15660
rect 17359 15657 17371 15691
rect 18782 15688 18788 15700
rect 18743 15660 18788 15688
rect 17313 15651 17371 15657
rect 18782 15648 18788 15660
rect 18840 15648 18846 15700
rect 21266 15688 21272 15700
rect 21227 15660 21272 15688
rect 21266 15648 21272 15660
rect 21324 15648 21330 15700
rect 21358 15648 21364 15700
rect 21416 15688 21422 15700
rect 21821 15691 21879 15697
rect 21821 15688 21833 15691
rect 21416 15660 21833 15688
rect 21416 15648 21422 15660
rect 21821 15657 21833 15660
rect 21867 15657 21879 15691
rect 22278 15688 22284 15700
rect 22239 15660 22284 15688
rect 21821 15651 21879 15657
rect 22278 15648 22284 15660
rect 22336 15648 22342 15700
rect 25406 15688 25412 15700
rect 25367 15660 25412 15688
rect 25406 15648 25412 15660
rect 25464 15648 25470 15700
rect 27798 15648 27804 15700
rect 27856 15688 27862 15700
rect 27985 15691 28043 15697
rect 27985 15688 27997 15691
rect 27856 15660 27997 15688
rect 27856 15648 27862 15660
rect 27985 15657 27997 15660
rect 28031 15657 28043 15691
rect 27985 15651 28043 15657
rect 28534 15648 28540 15700
rect 28592 15688 28598 15700
rect 28629 15691 28687 15697
rect 28629 15688 28641 15691
rect 28592 15660 28641 15688
rect 28592 15648 28598 15660
rect 28629 15657 28641 15660
rect 28675 15657 28687 15691
rect 29178 15688 29184 15700
rect 29139 15660 29184 15688
rect 28629 15651 28687 15657
rect 29178 15648 29184 15660
rect 29236 15648 29242 15700
rect 29730 15688 29736 15700
rect 29691 15660 29736 15688
rect 29730 15648 29736 15660
rect 29788 15648 29794 15700
rect 30190 15688 30196 15700
rect 30151 15660 30196 15688
rect 30190 15648 30196 15660
rect 30248 15648 30254 15700
rect 31938 15688 31944 15700
rect 31899 15660 31944 15688
rect 31938 15648 31944 15660
rect 31996 15648 32002 15700
rect 33321 15691 33379 15697
rect 33321 15657 33333 15691
rect 33367 15688 33379 15691
rect 34238 15688 34244 15700
rect 33367 15660 34244 15688
rect 33367 15657 33379 15660
rect 33321 15651 33379 15657
rect 34238 15648 34244 15660
rect 34296 15648 34302 15700
rect 35894 15648 35900 15700
rect 35952 15688 35958 15700
rect 35989 15691 36047 15697
rect 35989 15688 36001 15691
rect 35952 15660 36001 15688
rect 35952 15648 35958 15660
rect 35989 15657 36001 15660
rect 36035 15657 36047 15691
rect 35989 15651 36047 15657
rect 38197 15691 38255 15697
rect 38197 15657 38209 15691
rect 38243 15688 38255 15691
rect 38286 15688 38292 15700
rect 38243 15660 38292 15688
rect 38243 15657 38255 15660
rect 38197 15651 38255 15657
rect 38286 15648 38292 15660
rect 38344 15648 38350 15700
rect 40405 15691 40463 15697
rect 40405 15657 40417 15691
rect 40451 15688 40463 15691
rect 41138 15688 41144 15700
rect 40451 15660 41144 15688
rect 40451 15657 40463 15660
rect 40405 15651 40463 15657
rect 41138 15648 41144 15660
rect 41196 15648 41202 15700
rect 43438 15648 43444 15700
rect 43496 15697 43502 15700
rect 43496 15691 43545 15697
rect 43496 15657 43499 15691
rect 43533 15657 43545 15691
rect 43496 15651 43545 15657
rect 43496 15648 43502 15651
rect 11146 15620 11152 15632
rect 11107 15592 11152 15620
rect 11146 15580 11152 15592
rect 11204 15580 11210 15632
rect 11698 15620 11704 15632
rect 11659 15592 11704 15620
rect 11698 15580 11704 15592
rect 11756 15580 11762 15632
rect 12618 15580 12624 15632
rect 12676 15620 12682 15632
rect 12713 15623 12771 15629
rect 12713 15620 12725 15623
rect 12676 15592 12725 15620
rect 12676 15580 12682 15592
rect 12713 15589 12725 15592
rect 12759 15620 12771 15623
rect 15473 15623 15531 15629
rect 15473 15620 15485 15623
rect 12759 15592 15485 15620
rect 12759 15589 12771 15592
rect 12713 15583 12771 15589
rect 15473 15589 15485 15592
rect 15519 15620 15531 15623
rect 15562 15620 15568 15632
rect 15519 15592 15568 15620
rect 15519 15589 15531 15592
rect 15473 15583 15531 15589
rect 15562 15580 15568 15592
rect 15620 15580 15626 15632
rect 18227 15623 18285 15629
rect 18227 15589 18239 15623
rect 18273 15620 18285 15623
rect 18322 15620 18328 15632
rect 18273 15592 18328 15620
rect 18273 15589 18285 15592
rect 18227 15583 18285 15589
rect 18322 15580 18328 15592
rect 18380 15580 18386 15632
rect 21284 15620 21312 15648
rect 24442 15623 24500 15629
rect 24442 15620 24454 15623
rect 21284 15592 24454 15620
rect 24442 15589 24454 15592
rect 24488 15620 24500 15623
rect 24670 15620 24676 15632
rect 24488 15592 24676 15620
rect 24488 15589 24500 15592
rect 24442 15583 24500 15589
rect 24670 15580 24676 15592
rect 24728 15580 24734 15632
rect 26697 15623 26755 15629
rect 26697 15589 26709 15623
rect 26743 15620 26755 15623
rect 26786 15620 26792 15632
rect 26743 15592 26792 15620
rect 26743 15589 26755 15592
rect 26697 15583 26755 15589
rect 26786 15580 26792 15592
rect 26844 15580 26850 15632
rect 29748 15620 29776 15648
rect 29748 15592 30972 15620
rect 9950 15552 9956 15564
rect 9911 15524 9956 15552
rect 9950 15512 9956 15524
rect 10008 15512 10014 15564
rect 16920 15555 16978 15561
rect 16920 15521 16932 15555
rect 16966 15552 16978 15555
rect 17218 15552 17224 15564
rect 16966 15524 17224 15552
rect 16966 15521 16978 15524
rect 16920 15515 16978 15521
rect 17218 15512 17224 15524
rect 17276 15512 17282 15564
rect 19680 15555 19738 15561
rect 19680 15521 19692 15555
rect 19726 15552 19738 15555
rect 19794 15552 19800 15564
rect 19726 15524 19800 15552
rect 19726 15521 19738 15524
rect 19680 15515 19738 15521
rect 19794 15512 19800 15524
rect 19852 15512 19858 15564
rect 22554 15512 22560 15564
rect 22612 15552 22618 15564
rect 22684 15555 22742 15561
rect 22684 15552 22696 15555
rect 22612 15524 22696 15552
rect 22612 15512 22618 15524
rect 22684 15521 22696 15524
rect 22730 15521 22742 15555
rect 22684 15515 22742 15521
rect 25041 15555 25099 15561
rect 25041 15521 25053 15555
rect 25087 15552 25099 15555
rect 26418 15552 26424 15564
rect 25087 15524 26424 15552
rect 25087 15521 25099 15524
rect 25041 15515 25099 15521
rect 26418 15512 26424 15524
rect 26476 15512 26482 15564
rect 30944 15561 30972 15592
rect 31754 15580 31760 15632
rect 31812 15620 31818 15632
rect 32766 15629 32772 15632
rect 32722 15623 32772 15629
rect 32722 15620 32734 15623
rect 31812 15592 32734 15620
rect 31812 15580 31818 15592
rect 32722 15589 32734 15592
rect 32768 15589 32772 15623
rect 32722 15583 32772 15589
rect 32766 15580 32772 15583
rect 32824 15580 32830 15632
rect 33962 15620 33968 15632
rect 33923 15592 33968 15620
rect 33962 15580 33968 15592
rect 34020 15580 34026 15632
rect 34330 15620 34336 15632
rect 34291 15592 34336 15620
rect 34330 15580 34336 15592
rect 34388 15580 34394 15632
rect 35802 15580 35808 15632
rect 35860 15620 35866 15632
rect 36725 15623 36783 15629
rect 36725 15620 36737 15623
rect 35860 15592 36737 15620
rect 35860 15580 35866 15592
rect 36725 15589 36737 15592
rect 36771 15589 36783 15623
rect 36725 15583 36783 15589
rect 36998 15580 37004 15632
rect 37056 15620 37062 15632
rect 37918 15620 37924 15632
rect 37056 15592 37924 15620
rect 37056 15580 37062 15592
rect 37918 15580 37924 15592
rect 37976 15620 37982 15632
rect 38473 15623 38531 15629
rect 38473 15620 38485 15623
rect 37976 15592 38485 15620
rect 37976 15580 37982 15592
rect 38473 15589 38485 15592
rect 38519 15620 38531 15623
rect 39114 15620 39120 15632
rect 38519 15592 39120 15620
rect 38519 15589 38531 15592
rect 38473 15583 38531 15589
rect 39114 15580 39120 15592
rect 39172 15580 39178 15632
rect 30745 15555 30803 15561
rect 30745 15521 30757 15555
rect 30791 15521 30803 15555
rect 30745 15515 30803 15521
rect 30929 15555 30987 15561
rect 30929 15521 30941 15555
rect 30975 15552 30987 15555
rect 31110 15552 31116 15564
rect 30975 15524 31116 15552
rect 30975 15521 30987 15524
rect 30929 15515 30987 15521
rect 10091 15487 10149 15493
rect 10091 15453 10103 15487
rect 10137 15484 10149 15487
rect 11057 15487 11115 15493
rect 11057 15484 11069 15487
rect 10137 15456 11069 15484
rect 10137 15453 10149 15456
rect 10091 15447 10149 15453
rect 11057 15453 11069 15456
rect 11103 15484 11115 15487
rect 11514 15484 11520 15496
rect 11103 15456 11520 15484
rect 11103 15453 11115 15456
rect 11057 15447 11115 15453
rect 11514 15444 11520 15456
rect 11572 15444 11578 15496
rect 12158 15444 12164 15496
rect 12216 15484 12222 15496
rect 12621 15487 12679 15493
rect 12621 15484 12633 15487
rect 12216 15456 12633 15484
rect 12216 15444 12222 15456
rect 12621 15453 12633 15456
rect 12667 15453 12679 15487
rect 12621 15447 12679 15453
rect 15381 15487 15439 15493
rect 15381 15453 15393 15487
rect 15427 15484 15439 15487
rect 16022 15484 16028 15496
rect 15427 15456 16028 15484
rect 15427 15453 15439 15456
rect 15381 15447 15439 15453
rect 16022 15444 16028 15456
rect 16080 15444 16086 15496
rect 17494 15444 17500 15496
rect 17552 15484 17558 15496
rect 17865 15487 17923 15493
rect 17865 15484 17877 15487
rect 17552 15456 17877 15484
rect 17552 15444 17558 15456
rect 17865 15453 17877 15456
rect 17911 15453 17923 15487
rect 20898 15484 20904 15496
rect 20859 15456 20904 15484
rect 17865 15447 17923 15453
rect 20898 15444 20904 15456
rect 20956 15444 20962 15496
rect 24121 15487 24179 15493
rect 24121 15453 24133 15487
rect 24167 15484 24179 15487
rect 24210 15484 24216 15496
rect 24167 15456 24216 15484
rect 24167 15453 24179 15456
rect 24121 15447 24179 15453
rect 24210 15444 24216 15456
rect 24268 15444 24274 15496
rect 26602 15484 26608 15496
rect 26563 15456 26608 15484
rect 26602 15444 26608 15456
rect 26660 15444 26666 15496
rect 26878 15444 26884 15496
rect 26936 15484 26942 15496
rect 27617 15487 27675 15493
rect 27617 15484 27629 15487
rect 26936 15456 27629 15484
rect 26936 15444 26942 15456
rect 27617 15453 27629 15456
rect 27663 15484 27675 15487
rect 28074 15484 28080 15496
rect 27663 15456 28080 15484
rect 27663 15453 27675 15456
rect 27617 15447 27675 15453
rect 28074 15444 28080 15456
rect 28132 15444 28138 15496
rect 28258 15484 28264 15496
rect 28219 15456 28264 15484
rect 28258 15444 28264 15456
rect 28316 15444 28322 15496
rect 13170 15416 13176 15428
rect 13131 15388 13176 15416
rect 13170 15376 13176 15388
rect 13228 15376 13234 15428
rect 15930 15416 15936 15428
rect 15891 15388 15936 15416
rect 15930 15376 15936 15388
rect 15988 15376 15994 15428
rect 16482 15416 16488 15428
rect 16395 15388 16488 15416
rect 16482 15376 16488 15388
rect 16540 15416 16546 15428
rect 19751 15419 19809 15425
rect 19751 15416 19763 15419
rect 16540 15388 19763 15416
rect 16540 15376 16546 15388
rect 19751 15385 19763 15388
rect 19797 15385 19809 15419
rect 19751 15379 19809 15385
rect 24946 15376 24952 15428
rect 25004 15416 25010 15428
rect 26694 15416 26700 15428
rect 25004 15388 26700 15416
rect 25004 15376 25010 15388
rect 26694 15376 26700 15388
rect 26752 15416 26758 15428
rect 27157 15419 27215 15425
rect 27157 15416 27169 15419
rect 26752 15388 27169 15416
rect 26752 15376 26758 15388
rect 27157 15385 27169 15388
rect 27203 15385 27215 15419
rect 27157 15379 27215 15385
rect 30282 15376 30288 15428
rect 30340 15416 30346 15428
rect 30760 15416 30788 15515
rect 31110 15512 31116 15524
rect 31168 15512 31174 15564
rect 31205 15487 31263 15493
rect 31205 15453 31217 15487
rect 31251 15484 31263 15487
rect 32401 15487 32459 15493
rect 32401 15484 32413 15487
rect 31251 15456 32413 15484
rect 31251 15453 31263 15456
rect 31205 15447 31263 15453
rect 32401 15453 32413 15456
rect 32447 15484 32459 15487
rect 33870 15484 33876 15496
rect 32447 15456 33876 15484
rect 32447 15453 32459 15456
rect 32401 15447 32459 15453
rect 33870 15444 33876 15456
rect 33928 15444 33934 15496
rect 33980 15484 34008 15580
rect 35989 15555 36047 15561
rect 35989 15521 36001 15555
rect 36035 15552 36047 15555
rect 36078 15552 36084 15564
rect 36035 15524 36084 15552
rect 36035 15521 36047 15524
rect 35989 15515 36047 15521
rect 36078 15512 36084 15524
rect 36136 15512 36142 15564
rect 36173 15555 36231 15561
rect 36173 15521 36185 15555
rect 36219 15521 36231 15555
rect 40494 15552 40500 15564
rect 40455 15524 40500 15552
rect 36173 15515 36231 15521
rect 34241 15487 34299 15493
rect 34241 15484 34253 15487
rect 33980 15456 34253 15484
rect 34241 15453 34253 15456
rect 34287 15453 34299 15487
rect 34514 15484 34520 15496
rect 34475 15456 34520 15484
rect 34241 15447 34299 15453
rect 34514 15444 34520 15456
rect 34572 15444 34578 15496
rect 35250 15444 35256 15496
rect 35308 15484 35314 15496
rect 36188 15484 36216 15515
rect 40494 15512 40500 15524
rect 40552 15512 40558 15564
rect 40957 15555 41015 15561
rect 40957 15521 40969 15555
rect 41003 15552 41015 15555
rect 42245 15555 42303 15561
rect 42245 15552 42257 15555
rect 41003 15524 42257 15552
rect 41003 15521 41015 15524
rect 40957 15515 41015 15521
rect 42245 15521 42257 15524
rect 42291 15552 42303 15555
rect 42702 15552 42708 15564
rect 42291 15524 42708 15552
rect 42291 15521 42303 15524
rect 42245 15515 42303 15521
rect 36262 15484 36268 15496
rect 35308 15456 36268 15484
rect 35308 15444 35314 15456
rect 36262 15444 36268 15456
rect 36320 15444 36326 15496
rect 38381 15487 38439 15493
rect 38381 15453 38393 15487
rect 38427 15484 38439 15487
rect 38470 15484 38476 15496
rect 38427 15456 38476 15484
rect 38427 15453 38439 15456
rect 38381 15447 38439 15453
rect 38470 15444 38476 15456
rect 38528 15444 38534 15496
rect 38838 15484 38844 15496
rect 38799 15456 38844 15484
rect 38838 15444 38844 15456
rect 38896 15444 38902 15496
rect 39850 15444 39856 15496
rect 39908 15484 39914 15496
rect 40972 15484 41000 15515
rect 42702 15512 42708 15524
rect 42760 15512 42766 15564
rect 43257 15555 43315 15561
rect 43257 15521 43269 15555
rect 43303 15552 43315 15555
rect 43346 15552 43352 15564
rect 43303 15524 43352 15552
rect 43303 15521 43315 15524
rect 43257 15515 43315 15521
rect 43346 15512 43352 15524
rect 43404 15512 43410 15564
rect 41138 15484 41144 15496
rect 39908 15456 41000 15484
rect 41099 15456 41144 15484
rect 39908 15444 39914 15456
rect 41138 15444 41144 15456
rect 41196 15444 41202 15496
rect 35342 15416 35348 15428
rect 30340 15388 35348 15416
rect 30340 15376 30346 15388
rect 35342 15376 35348 15388
rect 35400 15416 35406 15428
rect 37550 15416 37556 15428
rect 35400 15388 37556 15416
rect 35400 15376 35406 15388
rect 37550 15376 37556 15388
rect 37608 15376 37614 15428
rect 10870 15348 10876 15360
rect 10831 15320 10876 15348
rect 10870 15308 10876 15320
rect 10928 15308 10934 15360
rect 15654 15308 15660 15360
rect 15712 15348 15718 15360
rect 16991 15351 17049 15357
rect 16991 15348 17003 15351
rect 15712 15320 17003 15348
rect 15712 15308 15718 15320
rect 16991 15317 17003 15320
rect 17037 15317 17049 15351
rect 19058 15348 19064 15360
rect 19019 15320 19064 15348
rect 16991 15311 17049 15317
rect 19058 15308 19064 15320
rect 19116 15308 19122 15360
rect 22646 15308 22652 15360
rect 22704 15348 22710 15360
rect 22787 15351 22845 15357
rect 22787 15348 22799 15351
rect 22704 15320 22799 15348
rect 22704 15308 22710 15320
rect 22787 15317 22799 15320
rect 22833 15317 22845 15351
rect 25866 15348 25872 15360
rect 25779 15320 25872 15348
rect 22787 15311 22845 15317
rect 25866 15308 25872 15320
rect 25924 15348 25930 15360
rect 27338 15348 27344 15360
rect 25924 15320 27344 15348
rect 25924 15308 25930 15320
rect 27338 15308 27344 15320
rect 27396 15308 27402 15360
rect 37182 15348 37188 15360
rect 37143 15320 37188 15348
rect 37182 15308 37188 15320
rect 37240 15308 37246 15360
rect 41874 15348 41880 15360
rect 41835 15320 41880 15348
rect 41874 15308 41880 15320
rect 41932 15308 41938 15360
rect 1104 15258 48852 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 48852 15258
rect 1104 15184 48852 15206
rect 9493 15147 9551 15153
rect 9493 15113 9505 15147
rect 9539 15144 9551 15147
rect 9950 15144 9956 15156
rect 9539 15116 9956 15144
rect 9539 15113 9551 15116
rect 9493 15107 9551 15113
rect 9950 15104 9956 15116
rect 10008 15144 10014 15156
rect 10873 15147 10931 15153
rect 10873 15144 10885 15147
rect 10008 15116 10885 15144
rect 10008 15104 10014 15116
rect 10873 15113 10885 15116
rect 10919 15113 10931 15147
rect 11514 15144 11520 15156
rect 11475 15116 11520 15144
rect 10873 15107 10931 15113
rect 11514 15104 11520 15116
rect 11572 15104 11578 15156
rect 12618 15144 12624 15156
rect 12579 15116 12624 15144
rect 12618 15104 12624 15116
rect 12676 15104 12682 15156
rect 14550 15144 14556 15156
rect 14511 15116 14556 15144
rect 14550 15104 14556 15116
rect 14608 15104 14614 15156
rect 15562 15104 15568 15156
rect 15620 15144 15626 15156
rect 15657 15147 15715 15153
rect 15657 15144 15669 15147
rect 15620 15116 15669 15144
rect 15620 15104 15626 15116
rect 15657 15113 15669 15116
rect 15703 15113 15715 15147
rect 16022 15144 16028 15156
rect 15983 15116 16028 15144
rect 15657 15107 15715 15113
rect 16022 15104 16028 15116
rect 16080 15104 16086 15156
rect 17865 15147 17923 15153
rect 17865 15113 17877 15147
rect 17911 15144 17923 15147
rect 18322 15144 18328 15156
rect 17911 15116 18328 15144
rect 17911 15113 17923 15116
rect 17865 15107 17923 15113
rect 18322 15104 18328 15116
rect 18380 15104 18386 15156
rect 19337 15147 19395 15153
rect 19337 15113 19349 15147
rect 19383 15144 19395 15147
rect 19705 15147 19763 15153
rect 19705 15144 19717 15147
rect 19383 15116 19717 15144
rect 19383 15113 19395 15116
rect 19337 15107 19395 15113
rect 19705 15113 19717 15116
rect 19751 15144 19763 15147
rect 19794 15144 19800 15156
rect 19751 15116 19800 15144
rect 19751 15113 19763 15116
rect 19705 15107 19763 15113
rect 19794 15104 19800 15116
rect 19852 15104 19858 15156
rect 21913 15147 21971 15153
rect 21913 15113 21925 15147
rect 21959 15144 21971 15147
rect 23382 15144 23388 15156
rect 21959 15116 23388 15144
rect 21959 15113 21971 15116
rect 21913 15107 21971 15113
rect 23382 15104 23388 15116
rect 23440 15104 23446 15156
rect 24670 15144 24676 15156
rect 24631 15116 24676 15144
rect 24670 15104 24676 15116
rect 24728 15144 24734 15156
rect 25409 15147 25467 15153
rect 25409 15144 25421 15147
rect 24728 15116 25421 15144
rect 24728 15104 24734 15116
rect 25409 15113 25421 15116
rect 25455 15113 25467 15147
rect 25409 15107 25467 15113
rect 14090 14968 14096 15020
rect 14148 15008 14154 15020
rect 15013 15011 15071 15017
rect 15013 15008 15025 15011
rect 14148 14980 15025 15008
rect 14148 14968 14154 14980
rect 15013 14977 15025 14980
rect 15059 15008 15071 15011
rect 15930 15008 15936 15020
rect 15059 14980 15936 15008
rect 15059 14977 15071 14980
rect 15013 14971 15071 14977
rect 15930 14968 15936 14980
rect 15988 14968 15994 15020
rect 18417 15011 18475 15017
rect 18417 14977 18429 15011
rect 18463 15008 18475 15011
rect 18690 15008 18696 15020
rect 18463 14980 18696 15008
rect 18463 14977 18475 14980
rect 18417 14971 18475 14977
rect 18690 14968 18696 14980
rect 18748 14968 18754 15020
rect 20898 14968 20904 15020
rect 20956 15008 20962 15020
rect 22189 15011 22247 15017
rect 22189 15008 22201 15011
rect 20956 14980 22201 15008
rect 20956 14968 20962 14980
rect 22189 14977 22201 14980
rect 22235 14977 22247 15011
rect 24210 15008 24216 15020
rect 24171 14980 24216 15008
rect 22189 14971 22247 14977
rect 24210 14968 24216 14980
rect 24268 14968 24274 15020
rect 25424 15008 25452 15107
rect 26602 15104 26608 15156
rect 26660 15144 26666 15156
rect 27157 15147 27215 15153
rect 27157 15144 27169 15147
rect 26660 15116 27169 15144
rect 26660 15104 26666 15116
rect 27157 15113 27169 15116
rect 27203 15144 27215 15147
rect 27246 15144 27252 15156
rect 27203 15116 27252 15144
rect 27203 15113 27215 15116
rect 27157 15107 27215 15113
rect 27246 15104 27252 15116
rect 27304 15104 27310 15156
rect 27338 15104 27344 15156
rect 27396 15144 27402 15156
rect 27479 15147 27537 15153
rect 27479 15144 27491 15147
rect 27396 15116 27491 15144
rect 27396 15104 27402 15116
rect 27479 15113 27491 15116
rect 27525 15113 27537 15147
rect 27479 15107 27537 15113
rect 28258 15104 28264 15156
rect 28316 15144 28322 15156
rect 28629 15147 28687 15153
rect 28629 15144 28641 15147
rect 28316 15116 28641 15144
rect 28316 15104 28322 15116
rect 28629 15113 28641 15116
rect 28675 15113 28687 15147
rect 28629 15107 28687 15113
rect 29730 15104 29736 15156
rect 29788 15144 29794 15156
rect 29825 15147 29883 15153
rect 29825 15144 29837 15147
rect 29788 15116 29837 15144
rect 29788 15104 29794 15116
rect 29825 15113 29837 15116
rect 29871 15113 29883 15147
rect 30282 15144 30288 15156
rect 30243 15116 30288 15144
rect 29825 15107 29883 15113
rect 30282 15104 30288 15116
rect 30340 15104 30346 15156
rect 31754 15144 31760 15156
rect 31715 15116 31760 15144
rect 31754 15104 31760 15116
rect 31812 15144 31818 15156
rect 32033 15147 32091 15153
rect 32033 15144 32045 15147
rect 31812 15116 32045 15144
rect 31812 15104 31818 15116
rect 32033 15113 32045 15116
rect 32079 15144 32091 15147
rect 32125 15147 32183 15153
rect 32125 15144 32137 15147
rect 32079 15116 32137 15144
rect 32079 15113 32091 15116
rect 32033 15107 32091 15113
rect 32125 15113 32137 15116
rect 32171 15113 32183 15147
rect 33870 15144 33876 15156
rect 33831 15116 33876 15144
rect 32125 15107 32183 15113
rect 33870 15104 33876 15116
rect 33928 15104 33934 15156
rect 34054 15104 34060 15156
rect 34112 15144 34118 15156
rect 34517 15147 34575 15153
rect 34517 15144 34529 15147
rect 34112 15116 34529 15144
rect 34112 15104 34118 15116
rect 34517 15113 34529 15116
rect 34563 15144 34575 15147
rect 34609 15147 34667 15153
rect 34609 15144 34621 15147
rect 34563 15116 34621 15144
rect 34563 15113 34575 15116
rect 34517 15107 34575 15113
rect 34609 15113 34621 15116
rect 34655 15113 34667 15147
rect 34609 15107 34667 15113
rect 35989 15147 36047 15153
rect 35989 15113 36001 15147
rect 36035 15144 36047 15147
rect 36078 15144 36084 15156
rect 36035 15116 36084 15144
rect 36035 15113 36047 15116
rect 35989 15107 36047 15113
rect 36078 15104 36084 15116
rect 36136 15104 36142 15156
rect 36262 15144 36268 15156
rect 36223 15116 36268 15144
rect 36262 15104 36268 15116
rect 36320 15104 36326 15156
rect 37182 15104 37188 15156
rect 37240 15144 37246 15156
rect 38427 15147 38485 15153
rect 38427 15144 38439 15147
rect 37240 15116 38439 15144
rect 37240 15104 37246 15116
rect 38427 15113 38439 15116
rect 38473 15113 38485 15147
rect 38427 15107 38485 15113
rect 39022 15104 39028 15156
rect 39080 15144 39086 15156
rect 39439 15147 39497 15153
rect 39439 15144 39451 15147
rect 39080 15116 39451 15144
rect 39080 15104 39086 15116
rect 39439 15113 39451 15116
rect 39485 15113 39497 15147
rect 39439 15107 39497 15113
rect 39850 15104 39856 15156
rect 39908 15144 39914 15156
rect 40221 15147 40279 15153
rect 40221 15144 40233 15147
rect 39908 15116 40233 15144
rect 39908 15104 39914 15116
rect 40221 15113 40233 15116
rect 40267 15113 40279 15147
rect 40221 15107 40279 15113
rect 40494 15104 40500 15156
rect 40552 15144 40558 15156
rect 41417 15147 41475 15153
rect 41417 15144 41429 15147
rect 40552 15116 41429 15144
rect 40552 15104 40558 15116
rect 41417 15113 41429 15116
rect 41463 15113 41475 15147
rect 43346 15144 43352 15156
rect 43307 15116 43352 15144
rect 41417 15107 41475 15113
rect 43346 15104 43352 15116
rect 43404 15104 43410 15156
rect 26786 15076 26792 15088
rect 26747 15048 26792 15076
rect 26786 15036 26792 15048
rect 26844 15036 26850 15088
rect 28261 15011 28319 15017
rect 28261 15008 28273 15011
rect 25424 14980 28273 15008
rect 9125 14943 9183 14949
rect 9125 14909 9137 14943
rect 9171 14940 9183 14943
rect 9858 14940 9864 14952
rect 9171 14912 9864 14940
rect 9171 14909 9183 14912
rect 9125 14903 9183 14909
rect 9858 14900 9864 14912
rect 9916 14940 9922 14952
rect 9953 14943 10011 14949
rect 9953 14940 9965 14943
rect 9916 14912 9965 14940
rect 9916 14900 9922 14912
rect 9953 14909 9965 14912
rect 9999 14909 10011 14943
rect 9953 14903 10011 14909
rect 13424 14943 13482 14949
rect 13424 14909 13436 14943
rect 13470 14940 13482 14943
rect 13470 14912 13814 14940
rect 13470 14909 13482 14912
rect 13424 14903 13482 14909
rect 12158 14832 12164 14884
rect 12216 14872 12222 14884
rect 12989 14875 13047 14881
rect 12989 14872 13001 14875
rect 12216 14844 13001 14872
rect 12216 14832 12222 14844
rect 12989 14841 13001 14844
rect 13035 14841 13047 14875
rect 12989 14835 13047 14841
rect 9861 14807 9919 14813
rect 9861 14773 9873 14807
rect 9907 14804 9919 14807
rect 10318 14804 10324 14816
rect 9907 14776 10324 14804
rect 9907 14773 9919 14776
rect 9861 14767 9919 14773
rect 10318 14764 10324 14776
rect 10376 14764 10382 14816
rect 11146 14764 11152 14816
rect 11204 14804 11210 14816
rect 11241 14807 11299 14813
rect 11241 14804 11253 14807
rect 11204 14776 11253 14804
rect 11204 14764 11210 14776
rect 11241 14773 11253 14776
rect 11287 14804 11299 14807
rect 11974 14804 11980 14816
rect 11287 14776 11980 14804
rect 11287 14773 11299 14776
rect 11241 14767 11299 14773
rect 11974 14764 11980 14776
rect 12032 14764 12038 14816
rect 13354 14764 13360 14816
rect 13412 14804 13418 14816
rect 13495 14807 13553 14813
rect 13495 14804 13507 14807
rect 13412 14776 13507 14804
rect 13412 14764 13418 14776
rect 13495 14773 13507 14776
rect 13541 14773 13553 14807
rect 13786 14804 13814 14912
rect 15838 14900 15844 14952
rect 15896 14940 15902 14952
rect 16244 14943 16302 14949
rect 16244 14940 16256 14943
rect 15896 14912 16256 14940
rect 15896 14900 15902 14912
rect 16244 14909 16256 14912
rect 16290 14940 16302 14943
rect 16669 14943 16727 14949
rect 16669 14940 16681 14943
rect 16290 14912 16681 14940
rect 16290 14909 16302 14912
rect 16244 14903 16302 14909
rect 16669 14909 16681 14912
rect 16715 14909 16727 14943
rect 16669 14903 16727 14909
rect 20165 14943 20223 14949
rect 20165 14909 20177 14943
rect 20211 14940 20223 14943
rect 20990 14940 20996 14952
rect 20211 14912 20996 14940
rect 20211 14909 20223 14912
rect 20165 14903 20223 14909
rect 20990 14900 20996 14912
rect 21048 14900 21054 14952
rect 21082 14900 21088 14952
rect 21140 14940 21146 14952
rect 23382 14940 23388 14952
rect 21140 14912 23388 14940
rect 21140 14900 21146 14912
rect 23382 14900 23388 14912
rect 23440 14940 23446 14952
rect 23661 14943 23719 14949
rect 23661 14940 23673 14943
rect 23440 14912 23673 14940
rect 23440 14900 23446 14912
rect 23661 14909 23673 14912
rect 23707 14909 23719 14943
rect 23661 14903 23719 14909
rect 23750 14900 23756 14952
rect 23808 14940 23814 14952
rect 24121 14943 24179 14949
rect 24121 14940 24133 14943
rect 23808 14912 24133 14940
rect 23808 14900 23814 14912
rect 24121 14909 24133 14912
rect 24167 14909 24179 14943
rect 25130 14940 25136 14952
rect 25043 14912 25136 14940
rect 24121 14903 24179 14909
rect 25130 14900 25136 14912
rect 25188 14940 25194 14952
rect 25593 14943 25651 14949
rect 25593 14940 25605 14943
rect 25188 14912 25605 14940
rect 25188 14900 25194 14912
rect 25593 14909 25605 14912
rect 25639 14909 25651 14943
rect 25593 14903 25651 14909
rect 14734 14872 14740 14884
rect 14695 14844 14740 14872
rect 14734 14832 14740 14844
rect 14792 14832 14798 14884
rect 14829 14875 14887 14881
rect 14829 14841 14841 14875
rect 14875 14841 14887 14875
rect 14829 14835 14887 14841
rect 13909 14807 13967 14813
rect 13909 14804 13921 14807
rect 13786 14776 13921 14804
rect 13495 14767 13553 14773
rect 13909 14773 13921 14776
rect 13955 14804 13967 14807
rect 14090 14804 14096 14816
rect 13955 14776 14096 14804
rect 13955 14773 13967 14776
rect 13909 14767 13967 14773
rect 14090 14764 14096 14776
rect 14148 14764 14154 14816
rect 14550 14764 14556 14816
rect 14608 14804 14614 14816
rect 14844 14804 14872 14835
rect 18322 14832 18328 14884
rect 18380 14872 18386 14884
rect 18738 14875 18796 14881
rect 18738 14872 18750 14875
rect 18380 14844 18750 14872
rect 18380 14832 18386 14844
rect 18738 14841 18750 14844
rect 18784 14872 18796 14875
rect 20441 14875 20499 14881
rect 20441 14872 20453 14875
rect 18784 14844 20453 14872
rect 18784 14841 18796 14844
rect 18738 14835 18796 14841
rect 20441 14841 20453 14844
rect 20487 14872 20499 14875
rect 20809 14875 20867 14881
rect 20809 14872 20821 14875
rect 20487 14844 20821 14872
rect 20487 14841 20499 14844
rect 20441 14835 20499 14841
rect 20809 14841 20821 14844
rect 20855 14872 20867 14875
rect 21266 14872 21272 14884
rect 20855 14844 21272 14872
rect 20855 14841 20867 14844
rect 20809 14835 20867 14841
rect 21266 14832 21272 14844
rect 21324 14881 21330 14884
rect 25929 14881 25957 14980
rect 28261 14977 28273 14980
rect 28307 15008 28319 15011
rect 28534 15008 28540 15020
rect 28307 14980 28540 15008
rect 28307 14977 28319 14980
rect 28261 14971 28319 14977
rect 28534 14968 28540 14980
rect 28592 14968 28598 15020
rect 36354 15008 36360 15020
rect 31036 14980 36360 15008
rect 26513 14943 26571 14949
rect 26513 14909 26525 14943
rect 26559 14940 26571 14943
rect 27376 14943 27434 14949
rect 27376 14940 27388 14943
rect 26559 14912 27388 14940
rect 26559 14909 26571 14912
rect 26513 14903 26571 14909
rect 27376 14909 27388 14912
rect 27422 14940 27434 14943
rect 27801 14943 27859 14949
rect 27801 14940 27813 14943
rect 27422 14912 27813 14940
rect 27422 14909 27434 14912
rect 27376 14903 27434 14909
rect 27801 14909 27813 14912
rect 27847 14909 27859 14943
rect 27801 14903 27859 14909
rect 29089 14943 29147 14949
rect 29089 14909 29101 14943
rect 29135 14940 29147 14943
rect 29178 14940 29184 14952
rect 29135 14912 29184 14940
rect 29135 14909 29147 14912
rect 29089 14903 29147 14909
rect 29178 14900 29184 14912
rect 29236 14940 29242 14952
rect 31036 14949 31064 14980
rect 36354 14968 36360 14980
rect 36412 14968 36418 15020
rect 36817 15011 36875 15017
rect 36817 14977 36829 15011
rect 36863 15008 36875 15011
rect 37200 15008 37228 15104
rect 39114 15076 39120 15088
rect 39075 15048 39120 15076
rect 39114 15036 39120 15048
rect 39172 15036 39178 15088
rect 39577 15079 39635 15085
rect 39577 15045 39589 15079
rect 39623 15076 39635 15079
rect 39761 15079 39819 15085
rect 39761 15076 39773 15079
rect 39623 15048 39773 15076
rect 39623 15045 39635 15048
rect 39577 15039 39635 15045
rect 39761 15045 39773 15048
rect 39807 15076 39819 15079
rect 40770 15076 40776 15088
rect 39807 15048 40776 15076
rect 39807 15045 39819 15048
rect 39761 15039 39819 15045
rect 40770 15036 40776 15048
rect 40828 15036 40834 15088
rect 40954 15076 40960 15088
rect 40915 15048 40960 15076
rect 40954 15036 40960 15048
rect 41012 15036 41018 15088
rect 41322 15036 41328 15088
rect 41380 15076 41386 15088
rect 42429 15079 42487 15085
rect 42429 15076 42441 15079
rect 41380 15048 42441 15076
rect 41380 15036 41386 15048
rect 42429 15045 42441 15048
rect 42475 15045 42487 15079
rect 42889 15079 42947 15085
rect 42889 15076 42901 15079
rect 42429 15039 42487 15045
rect 42766 15048 42901 15076
rect 36863 14980 37228 15008
rect 38197 15011 38255 15017
rect 36863 14977 36875 14980
rect 36817 14971 36875 14977
rect 38197 14977 38209 15011
rect 38243 15008 38255 15011
rect 38470 15008 38476 15020
rect 38243 14980 38476 15008
rect 38243 14977 38255 14980
rect 38197 14971 38255 14977
rect 38470 14968 38476 14980
rect 38528 15008 38534 15020
rect 40635 15011 40693 15017
rect 40635 15008 40647 15011
rect 38528 14980 40647 15008
rect 38528 14968 38534 14980
rect 40635 14977 40647 14980
rect 40681 14977 40693 15011
rect 40635 14971 40693 14977
rect 29308 14943 29366 14949
rect 29308 14940 29320 14943
rect 29236 14912 29320 14940
rect 29236 14900 29242 14912
rect 29308 14909 29320 14912
rect 29354 14909 29366 14943
rect 29308 14903 29366 14909
rect 30653 14943 30711 14949
rect 30653 14909 30665 14943
rect 30699 14940 30711 14943
rect 31021 14943 31079 14949
rect 31021 14940 31033 14943
rect 30699 14912 31033 14940
rect 30699 14909 30711 14912
rect 30653 14903 30711 14909
rect 31021 14909 31033 14912
rect 31067 14909 31079 14943
rect 31021 14903 31079 14909
rect 31110 14900 31116 14952
rect 31168 14940 31174 14952
rect 31205 14943 31263 14949
rect 31205 14940 31217 14943
rect 31168 14912 31217 14940
rect 31168 14900 31174 14912
rect 31205 14909 31217 14912
rect 31251 14909 31263 14943
rect 31205 14903 31263 14909
rect 31481 14943 31539 14949
rect 31481 14909 31493 14943
rect 31527 14940 31539 14943
rect 32309 14943 32367 14949
rect 32309 14940 32321 14943
rect 31527 14912 32321 14940
rect 31527 14909 31539 14912
rect 31481 14903 31539 14909
rect 32309 14909 32321 14912
rect 32355 14940 32367 14943
rect 33505 14943 33563 14949
rect 33505 14940 33517 14943
rect 32355 14912 33517 14940
rect 32355 14909 32367 14912
rect 32309 14903 32367 14909
rect 33505 14909 33517 14912
rect 33551 14909 33563 14943
rect 33505 14903 33563 14909
rect 34517 14943 34575 14949
rect 34517 14909 34529 14943
rect 34563 14940 34575 14943
rect 34885 14943 34943 14949
rect 34885 14940 34897 14943
rect 34563 14912 34897 14940
rect 34563 14909 34575 14912
rect 34517 14903 34575 14909
rect 34885 14909 34897 14912
rect 34931 14909 34943 14943
rect 34885 14903 34943 14909
rect 35250 14900 35256 14952
rect 35308 14940 35314 14952
rect 35345 14943 35403 14949
rect 35345 14940 35357 14943
rect 35308 14912 35357 14940
rect 35308 14900 35314 14912
rect 35345 14909 35357 14912
rect 35391 14909 35403 14943
rect 38324 14943 38382 14949
rect 38324 14940 38336 14943
rect 35345 14903 35403 14909
rect 38028 14912 38336 14940
rect 21324 14875 21372 14881
rect 21324 14841 21326 14875
rect 21360 14841 21372 14875
rect 21324 14835 21372 14841
rect 25914 14875 25972 14881
rect 25914 14841 25926 14875
rect 25960 14841 25972 14875
rect 25914 14835 25972 14841
rect 32033 14875 32091 14881
rect 32033 14841 32045 14875
rect 32079 14872 32091 14875
rect 32490 14872 32496 14884
rect 32079 14844 32496 14872
rect 32079 14841 32091 14844
rect 32033 14835 32091 14841
rect 21324 14832 21330 14835
rect 32490 14832 32496 14844
rect 32548 14872 32554 14884
rect 32630 14875 32688 14881
rect 32630 14872 32642 14875
rect 32548 14844 32642 14872
rect 32548 14832 32554 14844
rect 32630 14841 32642 14844
rect 32676 14841 32688 14875
rect 32630 14835 32688 14841
rect 33134 14832 33140 14884
rect 33192 14872 33198 14884
rect 35618 14872 35624 14884
rect 33192 14844 35388 14872
rect 35579 14844 35624 14872
rect 33192 14832 33198 14844
rect 14608 14776 14872 14804
rect 14608 14764 14614 14776
rect 16206 14764 16212 14816
rect 16264 14804 16270 14816
rect 16347 14807 16405 14813
rect 16347 14804 16359 14807
rect 16264 14776 16359 14804
rect 16264 14764 16270 14776
rect 16347 14773 16359 14776
rect 16393 14773 16405 14807
rect 16347 14767 16405 14773
rect 17129 14807 17187 14813
rect 17129 14773 17141 14807
rect 17175 14804 17187 14807
rect 17218 14804 17224 14816
rect 17175 14776 17224 14804
rect 17175 14773 17187 14776
rect 17129 14767 17187 14773
rect 17218 14764 17224 14776
rect 17276 14764 17282 14816
rect 17494 14804 17500 14816
rect 17455 14776 17500 14804
rect 17494 14764 17500 14776
rect 17552 14764 17558 14816
rect 22554 14764 22560 14816
rect 22612 14804 22618 14816
rect 22649 14807 22707 14813
rect 22649 14804 22661 14807
rect 22612 14776 22661 14804
rect 22612 14764 22618 14776
rect 22649 14773 22661 14776
rect 22695 14773 22707 14807
rect 22649 14767 22707 14773
rect 28350 14764 28356 14816
rect 28408 14804 28414 14816
rect 29411 14807 29469 14813
rect 29411 14804 29423 14807
rect 28408 14776 29423 14804
rect 28408 14764 28414 14776
rect 29411 14773 29423 14776
rect 29457 14773 29469 14807
rect 33226 14804 33232 14816
rect 33187 14776 33232 14804
rect 29411 14767 29469 14773
rect 33226 14764 33232 14776
rect 33284 14764 33290 14816
rect 34238 14804 34244 14816
rect 34199 14776 34244 14804
rect 34238 14764 34244 14776
rect 34296 14764 34302 14816
rect 35360 14804 35388 14844
rect 35618 14832 35624 14844
rect 35676 14832 35682 14884
rect 36906 14872 36912 14884
rect 36867 14844 36912 14872
rect 36906 14832 36912 14844
rect 36964 14832 36970 14884
rect 37274 14832 37280 14884
rect 37332 14872 37338 14884
rect 37461 14875 37519 14881
rect 37461 14872 37473 14875
rect 37332 14844 37473 14872
rect 37332 14832 37338 14844
rect 37461 14841 37473 14844
rect 37507 14872 37519 14875
rect 37918 14872 37924 14884
rect 37507 14844 37924 14872
rect 37507 14841 37519 14844
rect 37461 14835 37519 14841
rect 37918 14832 37924 14844
rect 37976 14832 37982 14884
rect 38028 14804 38056 14912
rect 38324 14909 38336 14912
rect 38370 14940 38382 14943
rect 38749 14943 38807 14949
rect 38749 14940 38761 14943
rect 38370 14912 38761 14940
rect 38370 14909 38382 14912
rect 38324 14903 38382 14909
rect 38749 14909 38761 14912
rect 38795 14909 38807 14943
rect 38749 14903 38807 14909
rect 39368 14943 39426 14949
rect 39368 14909 39380 14943
rect 39414 14940 39426 14943
rect 39577 14943 39635 14949
rect 39577 14940 39589 14943
rect 39414 14912 39589 14940
rect 39414 14909 39426 14912
rect 39368 14903 39426 14909
rect 39577 14909 39589 14912
rect 39623 14909 39635 14943
rect 39577 14903 39635 14909
rect 40548 14943 40606 14949
rect 40548 14909 40560 14943
rect 40594 14940 40606 14943
rect 40972 14940 41000 15036
rect 41877 15011 41935 15017
rect 41877 14977 41889 15011
rect 41923 15008 41935 15011
rect 42766 15008 42794 15048
rect 42889 15045 42901 15048
rect 42935 15076 42947 15079
rect 43714 15076 43720 15088
rect 42935 15048 43720 15076
rect 42935 15045 42947 15048
rect 42889 15039 42947 15045
rect 43714 15036 43720 15048
rect 43772 15036 43778 15088
rect 41923 14980 42794 15008
rect 41923 14977 41935 14980
rect 41877 14971 41935 14977
rect 41230 14940 41236 14952
rect 40594 14912 41236 14940
rect 40594 14909 40606 14912
rect 40548 14903 40606 14909
rect 38764 14872 38792 14903
rect 41230 14900 41236 14912
rect 41288 14900 41294 14952
rect 41690 14872 41696 14884
rect 38764 14844 41696 14872
rect 41690 14832 41696 14844
rect 41748 14832 41754 14884
rect 41874 14832 41880 14884
rect 41932 14872 41938 14884
rect 41969 14875 42027 14881
rect 41969 14872 41981 14875
rect 41932 14844 41981 14872
rect 41932 14832 41938 14844
rect 41969 14841 41981 14844
rect 42015 14841 42027 14875
rect 41969 14835 42027 14841
rect 35360 14776 38056 14804
rect 1104 14714 48852 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 48852 14714
rect 1104 14640 48852 14662
rect 10318 14560 10324 14612
rect 10376 14600 10382 14612
rect 10413 14603 10471 14609
rect 10413 14600 10425 14603
rect 10376 14572 10425 14600
rect 10376 14560 10382 14572
rect 10413 14569 10425 14572
rect 10459 14569 10471 14603
rect 10413 14563 10471 14569
rect 13354 14560 13360 14612
rect 13412 14600 13418 14612
rect 13412 14572 13492 14600
rect 13412 14560 13418 14572
rect 11974 14532 11980 14544
rect 11935 14504 11980 14532
rect 11974 14492 11980 14504
rect 12032 14492 12038 14544
rect 13464 14541 13492 14572
rect 17494 14560 17500 14612
rect 17552 14600 17558 14612
rect 18417 14603 18475 14609
rect 18417 14600 18429 14603
rect 17552 14572 18429 14600
rect 17552 14560 17558 14572
rect 18417 14569 18429 14572
rect 18463 14569 18475 14603
rect 20990 14600 20996 14612
rect 20951 14572 20996 14600
rect 18417 14563 18475 14569
rect 20990 14560 20996 14572
rect 21048 14560 21054 14612
rect 23750 14600 23756 14612
rect 23711 14572 23756 14600
rect 23750 14560 23756 14572
rect 23808 14560 23814 14612
rect 24210 14600 24216 14612
rect 24171 14572 24216 14600
rect 24210 14560 24216 14572
rect 24268 14560 24274 14612
rect 25130 14600 25136 14612
rect 25091 14572 25136 14600
rect 25130 14560 25136 14572
rect 25188 14560 25194 14612
rect 27522 14560 27528 14612
rect 27580 14600 27586 14612
rect 30377 14603 30435 14609
rect 27580 14572 28488 14600
rect 27580 14560 27586 14572
rect 13449 14535 13507 14541
rect 13449 14501 13461 14535
rect 13495 14501 13507 14535
rect 13449 14495 13507 14501
rect 13538 14492 13544 14544
rect 13596 14532 13602 14544
rect 15654 14532 15660 14544
rect 13596 14504 13641 14532
rect 15615 14504 15660 14532
rect 13596 14492 13602 14504
rect 15654 14492 15660 14504
rect 15712 14492 15718 14544
rect 15746 14492 15752 14544
rect 15804 14532 15810 14544
rect 16574 14532 16580 14544
rect 15804 14504 16580 14532
rect 15804 14492 15810 14504
rect 16574 14492 16580 14504
rect 16632 14492 16638 14544
rect 22649 14535 22707 14541
rect 22649 14501 22661 14535
rect 22695 14532 22707 14535
rect 22738 14532 22744 14544
rect 22695 14504 22744 14532
rect 22695 14501 22707 14504
rect 22649 14495 22707 14501
rect 22738 14492 22744 14504
rect 22796 14492 22802 14544
rect 23201 14535 23259 14541
rect 23201 14501 23213 14535
rect 23247 14532 23259 14535
rect 23290 14532 23296 14544
rect 23247 14504 23296 14532
rect 23247 14501 23259 14504
rect 23201 14495 23259 14501
rect 23290 14492 23296 14504
rect 23348 14492 23354 14544
rect 26418 14492 26424 14544
rect 26476 14532 26482 14544
rect 26697 14535 26755 14541
rect 26697 14532 26709 14535
rect 26476 14504 26709 14532
rect 26476 14492 26482 14504
rect 26697 14501 26709 14504
rect 26743 14501 26755 14535
rect 27246 14532 27252 14544
rect 27207 14504 27252 14532
rect 26697 14495 26755 14501
rect 27246 14492 27252 14504
rect 27304 14492 27310 14544
rect 28350 14532 28356 14544
rect 28311 14504 28356 14532
rect 28350 14492 28356 14504
rect 28408 14492 28414 14544
rect 28460 14541 28488 14572
rect 30377 14569 30389 14603
rect 30423 14600 30435 14603
rect 31110 14600 31116 14612
rect 30423 14572 31116 14600
rect 30423 14569 30435 14572
rect 30377 14563 30435 14569
rect 28445 14535 28503 14541
rect 28445 14501 28457 14535
rect 28491 14501 28503 14535
rect 28445 14495 28503 14501
rect 17380 14467 17438 14473
rect 17380 14433 17392 14467
rect 17426 14464 17438 14467
rect 17862 14464 17868 14476
rect 17426 14436 17868 14464
rect 17426 14433 17438 14436
rect 17380 14427 17438 14433
rect 17862 14424 17868 14436
rect 17920 14424 17926 14476
rect 18230 14424 18236 14476
rect 18288 14464 18294 14476
rect 18325 14467 18383 14473
rect 18325 14464 18337 14467
rect 18288 14436 18337 14464
rect 18288 14424 18294 14436
rect 18325 14433 18337 14436
rect 18371 14433 18383 14467
rect 18325 14427 18383 14433
rect 18785 14467 18843 14473
rect 18785 14433 18797 14467
rect 18831 14464 18843 14467
rect 19058 14464 19064 14476
rect 18831 14436 19064 14464
rect 18831 14433 18843 14436
rect 18785 14427 18843 14433
rect 10045 14399 10103 14405
rect 10045 14396 10057 14399
rect 9876 14368 10057 14396
rect 9674 14220 9680 14272
rect 9732 14260 9738 14272
rect 9876 14269 9904 14368
rect 10045 14365 10057 14368
rect 10091 14365 10103 14399
rect 10045 14359 10103 14365
rect 11146 14356 11152 14408
rect 11204 14396 11210 14408
rect 11885 14399 11943 14405
rect 11885 14396 11897 14399
rect 11204 14368 11897 14396
rect 11204 14356 11210 14368
rect 11885 14365 11897 14368
rect 11931 14365 11943 14399
rect 12158 14396 12164 14408
rect 12119 14368 12164 14396
rect 11885 14359 11943 14365
rect 12158 14356 12164 14368
rect 12216 14356 12222 14408
rect 13262 14356 13268 14408
rect 13320 14396 13326 14408
rect 13538 14396 13544 14408
rect 13320 14368 13544 14396
rect 13320 14356 13326 14368
rect 13538 14356 13544 14368
rect 13596 14396 13602 14408
rect 13725 14399 13783 14405
rect 13725 14396 13737 14399
rect 13596 14368 13737 14396
rect 13596 14356 13602 14368
rect 13725 14365 13737 14368
rect 13771 14365 13783 14399
rect 15930 14396 15936 14408
rect 15891 14368 15936 14396
rect 13725 14359 13783 14365
rect 15930 14356 15936 14368
rect 15988 14356 15994 14408
rect 17586 14356 17592 14408
rect 17644 14396 17650 14408
rect 18800 14396 18828 14427
rect 19058 14424 19064 14436
rect 19116 14424 19122 14476
rect 19978 14424 19984 14476
rect 20036 14464 20042 14476
rect 20901 14467 20959 14473
rect 20901 14464 20913 14467
rect 20036 14436 20913 14464
rect 20036 14424 20042 14436
rect 20901 14433 20913 14436
rect 20947 14464 20959 14467
rect 21082 14464 21088 14476
rect 20947 14436 21088 14464
rect 20947 14433 20959 14436
rect 20901 14427 20959 14433
rect 21082 14424 21088 14436
rect 21140 14424 21146 14476
rect 21453 14467 21511 14473
rect 21453 14433 21465 14467
rect 21499 14464 21511 14467
rect 21726 14464 21732 14476
rect 21499 14436 21732 14464
rect 21499 14433 21511 14436
rect 21453 14427 21511 14433
rect 21726 14424 21732 14436
rect 21784 14424 21790 14476
rect 23382 14424 23388 14476
rect 23440 14464 23446 14476
rect 24857 14467 24915 14473
rect 24857 14464 24869 14467
rect 23440 14436 24869 14464
rect 23440 14424 23446 14436
rect 24857 14433 24869 14436
rect 24903 14464 24915 14467
rect 24946 14464 24952 14476
rect 24903 14436 24952 14464
rect 24903 14433 24915 14436
rect 24857 14427 24915 14433
rect 24946 14424 24952 14436
rect 25004 14424 25010 14476
rect 25314 14464 25320 14476
rect 25275 14436 25320 14464
rect 25314 14424 25320 14436
rect 25372 14424 25378 14476
rect 30742 14464 30748 14476
rect 30703 14436 30748 14464
rect 30742 14424 30748 14436
rect 30800 14424 30806 14476
rect 30944 14473 30972 14572
rect 31110 14560 31116 14572
rect 31168 14560 31174 14612
rect 32490 14600 32496 14612
rect 32451 14572 32496 14600
rect 32490 14560 32496 14572
rect 32548 14560 32554 14612
rect 33045 14603 33103 14609
rect 33045 14569 33057 14603
rect 33091 14600 33103 14603
rect 34238 14600 34244 14612
rect 33091 14572 34244 14600
rect 33091 14569 33103 14572
rect 33045 14563 33103 14569
rect 34238 14560 34244 14572
rect 34296 14560 34302 14612
rect 34977 14603 35035 14609
rect 34977 14569 34989 14603
rect 35023 14600 35035 14603
rect 35250 14600 35256 14612
rect 35023 14572 35256 14600
rect 35023 14569 35035 14572
rect 34977 14563 35035 14569
rect 35250 14560 35256 14572
rect 35308 14600 35314 14612
rect 35526 14600 35532 14612
rect 35308 14572 35532 14600
rect 35308 14560 35314 14572
rect 35526 14560 35532 14572
rect 35584 14560 35590 14612
rect 41874 14560 41880 14612
rect 41932 14600 41938 14612
rect 42061 14603 42119 14609
rect 42061 14600 42073 14603
rect 41932 14572 42073 14600
rect 41932 14560 41938 14572
rect 42061 14569 42073 14572
rect 42107 14569 42119 14603
rect 42061 14563 42119 14569
rect 33226 14492 33232 14544
rect 33284 14532 33290 14544
rect 34057 14535 34115 14541
rect 34057 14532 34069 14535
rect 33284 14504 34069 14532
rect 33284 14492 33290 14504
rect 34057 14501 34069 14504
rect 34103 14532 34115 14535
rect 34146 14532 34152 14544
rect 34103 14504 34152 14532
rect 34103 14501 34115 14504
rect 34057 14495 34115 14501
rect 34146 14492 34152 14504
rect 34204 14492 34210 14544
rect 36265 14535 36323 14541
rect 36265 14501 36277 14535
rect 36311 14532 36323 14535
rect 36906 14532 36912 14544
rect 36311 14504 36912 14532
rect 36311 14501 36323 14504
rect 36265 14495 36323 14501
rect 36906 14492 36912 14504
rect 36964 14532 36970 14544
rect 37185 14535 37243 14541
rect 37185 14532 37197 14535
rect 36964 14504 37197 14532
rect 36964 14492 36970 14504
rect 37185 14501 37197 14504
rect 37231 14532 37243 14535
rect 38470 14532 38476 14544
rect 37231 14504 38476 14532
rect 37231 14501 37243 14504
rect 37185 14495 37243 14501
rect 38470 14492 38476 14504
rect 38528 14532 38534 14544
rect 38565 14535 38623 14541
rect 38565 14532 38577 14535
rect 38528 14504 38577 14532
rect 38528 14492 38534 14504
rect 38565 14501 38577 14504
rect 38611 14501 38623 14535
rect 38565 14495 38623 14501
rect 41046 14492 41052 14544
rect 41104 14532 41110 14544
rect 41462 14535 41520 14541
rect 41462 14532 41474 14535
rect 41104 14504 41474 14532
rect 41104 14492 41110 14504
rect 41462 14501 41474 14504
rect 41508 14501 41520 14535
rect 41462 14495 41520 14501
rect 30929 14467 30987 14473
rect 30929 14433 30941 14467
rect 30975 14433 30987 14467
rect 30929 14427 30987 14433
rect 36814 14424 36820 14476
rect 36872 14464 36878 14476
rect 41138 14464 41144 14476
rect 36872 14436 36917 14464
rect 41099 14436 41144 14464
rect 36872 14424 36878 14436
rect 41138 14424 41144 14436
rect 41196 14424 41202 14476
rect 17644 14368 18828 14396
rect 17644 14356 17650 14368
rect 22278 14356 22284 14408
rect 22336 14396 22342 14408
rect 22557 14399 22615 14405
rect 22557 14396 22569 14399
rect 22336 14368 22569 14396
rect 22336 14356 22342 14368
rect 22557 14365 22569 14368
rect 22603 14365 22615 14399
rect 22557 14359 22615 14365
rect 22738 14356 22744 14408
rect 22796 14396 22802 14408
rect 23198 14396 23204 14408
rect 22796 14368 23204 14396
rect 22796 14356 22802 14368
rect 23198 14356 23204 14368
rect 23256 14356 23262 14408
rect 26602 14396 26608 14408
rect 26563 14368 26608 14396
rect 26602 14356 26608 14368
rect 26660 14356 26666 14408
rect 28997 14399 29055 14405
rect 28997 14365 29009 14399
rect 29043 14396 29055 14399
rect 29638 14396 29644 14408
rect 29043 14368 29644 14396
rect 29043 14365 29055 14368
rect 28997 14359 29055 14365
rect 14734 14328 14740 14340
rect 14647 14300 14740 14328
rect 14734 14288 14740 14300
rect 14792 14328 14798 14340
rect 15948 14328 15976 14356
rect 14792 14300 15976 14328
rect 14792 14288 14798 14300
rect 24302 14288 24308 14340
rect 24360 14328 24366 14340
rect 29012 14328 29040 14359
rect 29638 14356 29644 14368
rect 29696 14356 29702 14408
rect 31205 14399 31263 14405
rect 31205 14365 31217 14399
rect 31251 14396 31263 14399
rect 31662 14396 31668 14408
rect 31251 14368 31668 14396
rect 31251 14365 31263 14368
rect 31205 14359 31263 14365
rect 31662 14356 31668 14368
rect 31720 14396 31726 14408
rect 32125 14399 32183 14405
rect 32125 14396 32137 14399
rect 31720 14368 32137 14396
rect 31720 14356 31726 14368
rect 32125 14365 32137 14368
rect 32171 14365 32183 14399
rect 32125 14359 32183 14365
rect 33594 14356 33600 14408
rect 33652 14396 33658 14408
rect 33778 14396 33784 14408
rect 33652 14368 33784 14396
rect 33652 14356 33658 14368
rect 33778 14356 33784 14368
rect 33836 14396 33842 14408
rect 33965 14399 34023 14405
rect 33965 14396 33977 14399
rect 33836 14368 33977 14396
rect 33836 14356 33842 14368
rect 33965 14365 33977 14368
rect 34011 14365 34023 14399
rect 36170 14396 36176 14408
rect 36131 14368 36176 14396
rect 33965 14359 34023 14365
rect 36170 14356 36176 14368
rect 36228 14356 36234 14408
rect 38470 14396 38476 14408
rect 38431 14368 38476 14396
rect 38470 14356 38476 14368
rect 38528 14356 38534 14408
rect 39117 14399 39175 14405
rect 39117 14365 39129 14399
rect 39163 14396 39175 14399
rect 39206 14396 39212 14408
rect 39163 14368 39212 14396
rect 39163 14365 39175 14368
rect 39117 14359 39175 14365
rect 39206 14356 39212 14368
rect 39264 14356 39270 14408
rect 34514 14328 34520 14340
rect 24360 14300 29040 14328
rect 34475 14300 34520 14328
rect 24360 14288 24366 14300
rect 34514 14288 34520 14300
rect 34572 14288 34578 14340
rect 9861 14263 9919 14269
rect 9861 14260 9873 14263
rect 9732 14232 9873 14260
rect 9732 14220 9738 14232
rect 9861 14229 9873 14232
rect 9907 14229 9919 14263
rect 10962 14260 10968 14272
rect 10923 14232 10968 14260
rect 9861 14223 9919 14229
rect 10962 14220 10968 14232
rect 11020 14220 11026 14272
rect 13262 14260 13268 14272
rect 13223 14232 13268 14260
rect 13262 14220 13268 14232
rect 13320 14220 13326 14272
rect 16390 14220 16396 14272
rect 16448 14260 16454 14272
rect 16577 14263 16635 14269
rect 16577 14260 16589 14263
rect 16448 14232 16589 14260
rect 16448 14220 16454 14232
rect 16577 14229 16589 14232
rect 16623 14229 16635 14263
rect 16577 14223 16635 14229
rect 16850 14220 16856 14272
rect 16908 14260 16914 14272
rect 17451 14263 17509 14269
rect 17451 14260 17463 14263
rect 16908 14232 17463 14260
rect 16908 14220 16914 14232
rect 17451 14229 17463 14232
rect 17497 14229 17509 14263
rect 17451 14223 17509 14229
rect 18233 14263 18291 14269
rect 18233 14229 18245 14263
rect 18279 14260 18291 14263
rect 18690 14260 18696 14272
rect 18279 14232 18696 14260
rect 18279 14229 18291 14232
rect 18233 14223 18291 14229
rect 18690 14220 18696 14232
rect 18748 14220 18754 14272
rect 29362 14260 29368 14272
rect 29323 14232 29368 14260
rect 29362 14220 29368 14232
rect 29420 14220 29426 14272
rect 1104 14170 48852 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 48852 14170
rect 1104 14096 48852 14118
rect 10870 14016 10876 14068
rect 10928 14056 10934 14068
rect 11471 14059 11529 14065
rect 11471 14056 11483 14059
rect 10928 14028 11483 14056
rect 10928 14016 10934 14028
rect 11471 14025 11483 14028
rect 11517 14025 11529 14059
rect 11471 14019 11529 14025
rect 12713 14059 12771 14065
rect 12713 14025 12725 14059
rect 12759 14056 12771 14059
rect 13354 14056 13360 14068
rect 12759 14028 13360 14056
rect 12759 14025 12771 14028
rect 12713 14019 12771 14025
rect 13354 14016 13360 14028
rect 13412 14016 13418 14068
rect 13446 14016 13452 14068
rect 13504 14056 13510 14068
rect 14277 14059 14335 14065
rect 14277 14056 14289 14059
rect 13504 14028 14289 14056
rect 13504 14016 13510 14028
rect 14277 14025 14289 14028
rect 14323 14056 14335 14059
rect 15746 14056 15752 14068
rect 14323 14028 15752 14056
rect 14323 14025 14335 14028
rect 14277 14019 14335 14025
rect 15746 14016 15752 14028
rect 15804 14056 15810 14068
rect 16117 14059 16175 14065
rect 16117 14056 16129 14059
rect 15804 14028 16129 14056
rect 15804 14016 15810 14028
rect 16117 14025 16129 14028
rect 16163 14025 16175 14059
rect 16117 14019 16175 14025
rect 19978 14016 19984 14068
rect 20036 14056 20042 14068
rect 20165 14059 20223 14065
rect 20165 14056 20177 14059
rect 20036 14028 20177 14056
rect 20036 14016 20042 14028
rect 20165 14025 20177 14028
rect 20211 14025 20223 14059
rect 20165 14019 20223 14025
rect 11885 13991 11943 13997
rect 11885 13957 11897 13991
rect 11931 13988 11943 13991
rect 11974 13988 11980 14000
rect 11931 13960 11980 13988
rect 11931 13957 11943 13960
rect 11885 13951 11943 13957
rect 11974 13948 11980 13960
rect 12032 13988 12038 14000
rect 13464 13988 13492 14016
rect 12032 13960 13492 13988
rect 15381 13991 15439 13997
rect 12032 13948 12038 13960
rect 15381 13957 15393 13991
rect 15427 13988 15439 13991
rect 15930 13988 15936 14000
rect 15427 13960 15936 13988
rect 15427 13957 15439 13960
rect 15381 13951 15439 13957
rect 15930 13948 15936 13960
rect 15988 13948 15994 14000
rect 16022 13948 16028 14000
rect 16080 13988 16086 14000
rect 16080 13960 16712 13988
rect 16080 13948 16086 13960
rect 9214 13880 9220 13932
rect 9272 13920 9278 13932
rect 9309 13923 9367 13929
rect 9309 13920 9321 13923
rect 9272 13892 9321 13920
rect 9272 13880 9278 13892
rect 9309 13889 9321 13892
rect 9355 13920 9367 13923
rect 12161 13923 12219 13929
rect 12161 13920 12173 13923
rect 9355 13892 10272 13920
rect 9355 13889 9367 13892
rect 9309 13883 9367 13889
rect 10244 13864 10272 13892
rect 11383 13892 12173 13920
rect 10045 13855 10103 13861
rect 10045 13852 10057 13855
rect 9600 13824 10057 13852
rect 9600 13725 9628 13824
rect 10045 13821 10057 13824
rect 10091 13852 10103 13855
rect 10091 13824 10180 13852
rect 10091 13821 10103 13824
rect 10045 13815 10103 13821
rect 10152 13796 10180 13824
rect 10226 13812 10232 13864
rect 10284 13852 10290 13864
rect 10284 13824 10329 13852
rect 10284 13812 10290 13824
rect 10962 13812 10968 13864
rect 11020 13852 11026 13864
rect 11383 13861 11411 13892
rect 12161 13889 12173 13892
rect 12207 13889 12219 13923
rect 12161 13883 12219 13889
rect 13081 13923 13139 13929
rect 13081 13889 13093 13923
rect 13127 13920 13139 13923
rect 13354 13920 13360 13932
rect 13127 13892 13360 13920
rect 13127 13889 13139 13892
rect 13081 13883 13139 13889
rect 11368 13855 11426 13861
rect 11368 13852 11380 13855
rect 11020 13824 11380 13852
rect 11020 13812 11026 13824
rect 11368 13821 11380 13824
rect 11414 13821 11426 13855
rect 11368 13815 11426 13821
rect 11974 13812 11980 13864
rect 12032 13852 12038 13864
rect 13096 13852 13124 13883
rect 13354 13880 13360 13892
rect 13412 13880 13418 13932
rect 13538 13920 13544 13932
rect 13499 13892 13544 13920
rect 13538 13880 13544 13892
rect 13596 13880 13602 13932
rect 14826 13920 14832 13932
rect 14739 13892 14832 13920
rect 14826 13880 14832 13892
rect 14884 13920 14890 13932
rect 16206 13920 16212 13932
rect 14884 13892 16212 13920
rect 14884 13880 14890 13892
rect 16206 13880 16212 13892
rect 16264 13880 16270 13932
rect 16684 13929 16712 13960
rect 18874 13948 18880 14000
rect 18932 13988 18938 14000
rect 19426 13988 19432 14000
rect 18932 13960 19432 13988
rect 18932 13948 18938 13960
rect 19426 13948 19432 13960
rect 19484 13948 19490 14000
rect 16669 13923 16727 13929
rect 16669 13889 16681 13923
rect 16715 13920 16727 13923
rect 17126 13920 17132 13932
rect 16715 13892 17132 13920
rect 16715 13889 16727 13892
rect 16669 13883 16727 13889
rect 17126 13880 17132 13892
rect 17184 13880 17190 13932
rect 12032 13824 13124 13852
rect 18877 13855 18935 13861
rect 12032 13812 12038 13824
rect 18877 13821 18889 13855
rect 18923 13821 18935 13855
rect 18877 13815 18935 13821
rect 19061 13855 19119 13861
rect 19061 13821 19073 13855
rect 19107 13852 19119 13855
rect 20180 13852 20208 14019
rect 20254 14016 20260 14068
rect 20312 14056 20318 14068
rect 24946 14056 24952 14068
rect 20312 14028 23474 14056
rect 24907 14028 24952 14056
rect 20312 14016 20318 14028
rect 21082 13948 21088 14000
rect 21140 13988 21146 14000
rect 21361 13991 21419 13997
rect 21361 13988 21373 13991
rect 21140 13960 21373 13988
rect 21140 13948 21146 13960
rect 21361 13957 21373 13960
rect 21407 13957 21419 13991
rect 23446 13988 23474 14028
rect 24946 14016 24952 14028
rect 25004 14016 25010 14068
rect 25639 14059 25697 14065
rect 25639 14025 25651 14059
rect 25685 14056 25697 14059
rect 26602 14056 26608 14068
rect 25685 14028 26608 14056
rect 25685 14025 25697 14028
rect 25639 14019 25697 14025
rect 26602 14016 26608 14028
rect 26660 14056 26666 14068
rect 27525 14059 27583 14065
rect 27525 14056 27537 14059
rect 26660 14028 27537 14056
rect 26660 14016 26666 14028
rect 27525 14025 27537 14028
rect 27571 14025 27583 14059
rect 27525 14019 27583 14025
rect 27985 14059 28043 14065
rect 27985 14025 27997 14059
rect 28031 14056 28043 14059
rect 28350 14056 28356 14068
rect 28031 14028 28356 14056
rect 28031 14025 28043 14028
rect 27985 14019 28043 14025
rect 28350 14016 28356 14028
rect 28408 14016 28414 14068
rect 30929 14059 30987 14065
rect 30929 14025 30941 14059
rect 30975 14056 30987 14059
rect 31110 14056 31116 14068
rect 30975 14028 31116 14056
rect 30975 14025 30987 14028
rect 30929 14019 30987 14025
rect 31110 14016 31116 14028
rect 31168 14016 31174 14068
rect 31662 14056 31668 14068
rect 31623 14028 31668 14056
rect 31662 14016 31668 14028
rect 31720 14016 31726 14068
rect 32401 14059 32459 14065
rect 32401 14025 32413 14059
rect 32447 14056 32459 14059
rect 32490 14056 32496 14068
rect 32447 14028 32496 14056
rect 32447 14025 32459 14028
rect 32401 14019 32459 14025
rect 32490 14016 32496 14028
rect 32548 14016 32554 14068
rect 33594 14056 33600 14068
rect 33555 14028 33600 14056
rect 33594 14016 33600 14028
rect 33652 14016 33658 14068
rect 34146 14056 34152 14068
rect 34107 14028 34152 14056
rect 34146 14016 34152 14028
rect 34204 14016 34210 14068
rect 34514 14056 34520 14068
rect 34475 14028 34520 14056
rect 34514 14016 34520 14028
rect 34572 14016 34578 14068
rect 35529 14059 35587 14065
rect 35529 14025 35541 14059
rect 35575 14056 35587 14059
rect 35710 14056 35716 14068
rect 35575 14028 35716 14056
rect 35575 14025 35587 14028
rect 35529 14019 35587 14025
rect 35710 14016 35716 14028
rect 35768 14056 35774 14068
rect 35986 14056 35992 14068
rect 35768 14028 35992 14056
rect 35768 14016 35774 14028
rect 35986 14016 35992 14028
rect 36044 14016 36050 14068
rect 36170 14016 36176 14068
rect 36228 14056 36234 14068
rect 36906 14056 36912 14068
rect 36228 14028 36912 14056
rect 36228 14016 36234 14028
rect 36906 14016 36912 14028
rect 36964 14056 36970 14068
rect 37185 14059 37243 14065
rect 37185 14056 37197 14059
rect 36964 14028 37197 14056
rect 36964 14016 36970 14028
rect 37185 14025 37197 14028
rect 37231 14025 37243 14059
rect 37185 14019 37243 14025
rect 41138 14016 41144 14068
rect 41196 14056 41202 14068
rect 41509 14059 41567 14065
rect 41509 14056 41521 14059
rect 41196 14028 41521 14056
rect 41196 14016 41202 14028
rect 41509 14025 41521 14028
rect 41555 14025 41567 14059
rect 41509 14019 41567 14025
rect 25314 13988 25320 14000
rect 23446 13960 25320 13988
rect 21361 13951 21419 13957
rect 25314 13948 25320 13960
rect 25372 13948 25378 14000
rect 26418 13988 26424 14000
rect 26331 13960 26424 13988
rect 26418 13948 26424 13960
rect 26476 13988 26482 14000
rect 30561 13991 30619 13997
rect 26476 13960 28396 13988
rect 26476 13948 26482 13960
rect 20898 13920 20904 13932
rect 20859 13892 20904 13920
rect 20898 13880 20904 13892
rect 20956 13880 20962 13932
rect 24673 13923 24731 13929
rect 24673 13889 24685 13923
rect 24719 13920 24731 13923
rect 24762 13920 24768 13932
rect 24719 13892 24768 13920
rect 24719 13889 24731 13892
rect 24673 13883 24731 13889
rect 24762 13880 24768 13892
rect 24820 13880 24826 13932
rect 26053 13923 26111 13929
rect 26053 13889 26065 13923
rect 26099 13920 26111 13923
rect 26694 13920 26700 13932
rect 26099 13892 26700 13920
rect 26099 13889 26111 13892
rect 26053 13883 26111 13889
rect 26694 13880 26700 13892
rect 26752 13880 26758 13932
rect 27246 13920 27252 13932
rect 27207 13892 27252 13920
rect 27246 13880 27252 13892
rect 27304 13880 27310 13932
rect 20349 13855 20407 13861
rect 20349 13852 20361 13855
rect 19107 13824 19141 13852
rect 20180 13824 20361 13852
rect 19107 13821 19119 13824
rect 19061 13815 19119 13821
rect 20349 13821 20361 13824
rect 20395 13821 20407 13855
rect 20349 13815 20407 13821
rect 10134 13744 10140 13796
rect 10192 13744 10198 13796
rect 10318 13744 10324 13796
rect 10376 13784 10382 13796
rect 10873 13787 10931 13793
rect 10873 13784 10885 13787
rect 10376 13756 10885 13784
rect 10376 13744 10382 13756
rect 10873 13753 10885 13756
rect 10919 13784 10931 13787
rect 13262 13784 13268 13796
rect 10919 13756 11928 13784
rect 13223 13756 13268 13784
rect 10919 13753 10931 13756
rect 10873 13747 10931 13753
rect 9585 13719 9643 13725
rect 9585 13685 9597 13719
rect 9631 13685 9643 13719
rect 9858 13716 9864 13728
rect 9819 13688 9864 13716
rect 9585 13679 9643 13685
rect 9858 13676 9864 13688
rect 9916 13676 9922 13728
rect 11146 13716 11152 13728
rect 11107 13688 11152 13716
rect 11146 13676 11152 13688
rect 11204 13676 11210 13728
rect 11900 13716 11928 13756
rect 13262 13744 13268 13756
rect 13320 13744 13326 13796
rect 13354 13744 13360 13796
rect 13412 13784 13418 13796
rect 14553 13787 14611 13793
rect 14553 13784 14565 13787
rect 13412 13756 14565 13784
rect 13412 13744 13418 13756
rect 14553 13753 14565 13756
rect 14599 13784 14611 13787
rect 14921 13787 14979 13793
rect 14921 13784 14933 13787
rect 14599 13756 14933 13784
rect 14599 13753 14611 13756
rect 14553 13747 14611 13753
rect 14921 13753 14933 13756
rect 14967 13784 14979 13787
rect 16206 13784 16212 13796
rect 14967 13756 16212 13784
rect 14967 13753 14979 13756
rect 14921 13747 14979 13753
rect 16206 13744 16212 13756
rect 16264 13744 16270 13796
rect 16390 13784 16396 13796
rect 16351 13756 16396 13784
rect 16390 13744 16396 13756
rect 16448 13744 16454 13796
rect 16485 13787 16543 13793
rect 16485 13753 16497 13787
rect 16531 13784 16543 13787
rect 16574 13784 16580 13796
rect 16531 13756 16580 13784
rect 16531 13753 16543 13756
rect 16485 13747 16543 13753
rect 16574 13744 16580 13756
rect 16632 13744 16638 13796
rect 13630 13716 13636 13728
rect 11900 13688 13636 13716
rect 13630 13676 13636 13688
rect 13688 13676 13694 13728
rect 17402 13716 17408 13728
rect 17363 13688 17408 13716
rect 17402 13676 17408 13688
rect 17460 13716 17466 13728
rect 17586 13716 17592 13728
rect 17460 13688 17592 13716
rect 17460 13676 17466 13688
rect 17586 13676 17592 13688
rect 17644 13716 17650 13728
rect 17773 13719 17831 13725
rect 17773 13716 17785 13719
rect 17644 13688 17785 13716
rect 17644 13676 17650 13688
rect 17773 13685 17785 13688
rect 17819 13685 17831 13719
rect 17773 13679 17831 13685
rect 18230 13676 18236 13728
rect 18288 13716 18294 13728
rect 18325 13719 18383 13725
rect 18325 13716 18337 13719
rect 18288 13688 18337 13716
rect 18288 13676 18294 13688
rect 18325 13685 18337 13688
rect 18371 13685 18383 13719
rect 18690 13716 18696 13728
rect 18651 13688 18696 13716
rect 18325 13679 18383 13685
rect 18690 13676 18696 13688
rect 18748 13676 18754 13728
rect 18892 13716 18920 13815
rect 18966 13744 18972 13796
rect 19024 13784 19030 13796
rect 19076 13784 19104 13815
rect 20530 13812 20536 13864
rect 20588 13852 20594 13864
rect 20809 13855 20867 13861
rect 20809 13852 20821 13855
rect 20588 13824 20821 13852
rect 20588 13812 20594 13824
rect 20809 13821 20821 13824
rect 20855 13821 20867 13855
rect 20809 13815 20867 13821
rect 22624 13855 22682 13861
rect 22624 13821 22636 13855
rect 22670 13852 22682 13855
rect 22738 13852 22744 13864
rect 22670 13824 22744 13852
rect 22670 13821 22682 13824
rect 22624 13815 22682 13821
rect 22738 13812 22744 13824
rect 22796 13812 22802 13864
rect 25406 13812 25412 13864
rect 25464 13852 25470 13864
rect 25536 13855 25594 13861
rect 25536 13852 25548 13855
rect 25464 13824 25548 13852
rect 25464 13812 25470 13824
rect 25536 13821 25548 13824
rect 25582 13821 25594 13855
rect 25536 13815 25594 13821
rect 26418 13812 26424 13864
rect 26476 13812 26482 13864
rect 28144 13855 28202 13861
rect 28144 13821 28156 13855
rect 28190 13852 28202 13855
rect 28258 13852 28264 13864
rect 28190 13824 28264 13852
rect 28190 13821 28202 13824
rect 28144 13815 28202 13821
rect 28258 13812 28264 13824
rect 28316 13812 28322 13864
rect 28368 13852 28396 13960
rect 30561 13957 30573 13991
rect 30607 13988 30619 13991
rect 30742 13988 30748 14000
rect 30607 13960 30748 13988
rect 30607 13957 30619 13960
rect 30561 13951 30619 13957
rect 30742 13948 30748 13960
rect 30800 13988 30806 14000
rect 38286 13988 38292 14000
rect 30800 13960 38292 13988
rect 30800 13948 30806 13960
rect 38286 13948 38292 13960
rect 38344 13948 38350 14000
rect 40313 13991 40371 13997
rect 40313 13957 40325 13991
rect 40359 13988 40371 13991
rect 41322 13988 41328 14000
rect 40359 13960 41328 13988
rect 40359 13957 40371 13960
rect 40313 13951 40371 13957
rect 29638 13920 29644 13932
rect 29599 13892 29644 13920
rect 29638 13880 29644 13892
rect 29696 13880 29702 13932
rect 32677 13923 32735 13929
rect 32677 13920 32689 13923
rect 31899 13892 32689 13920
rect 28626 13852 28632 13864
rect 28368 13824 28632 13852
rect 28626 13812 28632 13824
rect 28684 13852 28690 13864
rect 29086 13852 29092 13864
rect 28684 13824 29092 13852
rect 28684 13812 28690 13824
rect 29086 13812 29092 13824
rect 29144 13812 29150 13864
rect 31202 13812 31208 13864
rect 31260 13852 31266 13864
rect 31899 13861 31927 13892
rect 32677 13889 32689 13892
rect 32723 13889 32735 13923
rect 35618 13920 35624 13932
rect 35579 13892 35624 13920
rect 32677 13883 32735 13889
rect 35618 13880 35624 13892
rect 35676 13880 35682 13932
rect 38838 13920 38844 13932
rect 38799 13892 38844 13920
rect 38838 13880 38844 13892
rect 38896 13880 38902 13932
rect 31884 13855 31942 13861
rect 31884 13852 31896 13855
rect 31260 13824 31896 13852
rect 31260 13812 31266 13824
rect 31884 13821 31896 13824
rect 31930 13821 31942 13855
rect 31884 13815 31942 13821
rect 33756 13855 33814 13861
rect 33756 13821 33768 13855
rect 33802 13852 33814 13855
rect 34514 13852 34520 13864
rect 33802 13824 34520 13852
rect 33802 13821 33814 13824
rect 33756 13815 33814 13821
rect 34514 13812 34520 13824
rect 34572 13812 34578 13864
rect 40579 13861 40607 13960
rect 41322 13948 41328 13960
rect 41380 13948 41386 14000
rect 41046 13880 41052 13932
rect 41104 13920 41110 13932
rect 41141 13923 41199 13929
rect 41141 13920 41153 13923
rect 41104 13892 41153 13920
rect 41104 13880 41110 13892
rect 41141 13889 41153 13892
rect 41187 13920 41199 13923
rect 41598 13920 41604 13932
rect 41187 13892 41604 13920
rect 41187 13889 41199 13892
rect 41141 13883 41199 13889
rect 41598 13880 41604 13892
rect 41656 13880 41662 13932
rect 40564 13855 40622 13861
rect 40564 13821 40576 13855
rect 40610 13821 40622 13855
rect 40564 13815 40622 13821
rect 19024 13756 19104 13784
rect 23477 13787 23535 13793
rect 19024 13744 19030 13756
rect 23477 13753 23489 13787
rect 23523 13784 23535 13787
rect 24026 13784 24032 13796
rect 23523 13756 24032 13784
rect 23523 13753 23535 13756
rect 23477 13747 23535 13753
rect 24026 13744 24032 13756
rect 24084 13744 24090 13796
rect 24118 13744 24124 13796
rect 24176 13784 24182 13796
rect 26436 13784 26464 13812
rect 24176 13756 26464 13784
rect 26605 13787 26663 13793
rect 24176 13744 24182 13756
rect 26605 13753 26617 13787
rect 26651 13753 26663 13787
rect 26605 13747 26663 13753
rect 19242 13716 19248 13728
rect 18892 13688 19248 13716
rect 19242 13676 19248 13688
rect 19300 13716 19306 13728
rect 20254 13716 20260 13728
rect 19300 13688 20260 13716
rect 19300 13676 19306 13688
rect 20254 13676 20260 13688
rect 20312 13676 20318 13728
rect 21726 13716 21732 13728
rect 21687 13688 21732 13716
rect 21726 13676 21732 13688
rect 21784 13676 21790 13728
rect 22278 13676 22284 13728
rect 22336 13716 22342 13728
rect 22373 13719 22431 13725
rect 22373 13716 22385 13719
rect 22336 13688 22385 13716
rect 22336 13676 22342 13688
rect 22373 13685 22385 13688
rect 22419 13685 22431 13719
rect 22373 13679 22431 13685
rect 22695 13719 22753 13725
rect 22695 13685 22707 13719
rect 22741 13716 22753 13719
rect 23014 13716 23020 13728
rect 22741 13688 23020 13716
rect 22741 13685 22753 13688
rect 22695 13679 22753 13685
rect 23014 13676 23020 13688
rect 23072 13676 23078 13728
rect 23109 13719 23167 13725
rect 23109 13685 23121 13719
rect 23155 13716 23167 13719
rect 23198 13716 23204 13728
rect 23155 13688 23204 13716
rect 23155 13685 23167 13688
rect 23109 13679 23167 13685
rect 23198 13676 23204 13688
rect 23256 13716 23262 13728
rect 24136 13716 24164 13744
rect 23256 13688 24164 13716
rect 23256 13676 23262 13688
rect 26326 13676 26332 13728
rect 26384 13716 26390 13728
rect 26620 13716 26648 13747
rect 26694 13744 26700 13796
rect 26752 13784 26758 13796
rect 27522 13784 27528 13796
rect 26752 13756 27528 13784
rect 26752 13744 26758 13756
rect 27522 13744 27528 13756
rect 27580 13784 27586 13796
rect 28537 13787 28595 13793
rect 28537 13784 28549 13787
rect 27580 13756 28549 13784
rect 27580 13744 27586 13756
rect 28537 13753 28549 13756
rect 28583 13753 28595 13787
rect 29362 13784 29368 13796
rect 29323 13756 29368 13784
rect 28537 13747 28595 13753
rect 29362 13744 29368 13756
rect 29420 13744 29426 13796
rect 29457 13787 29515 13793
rect 29457 13753 29469 13787
rect 29503 13753 29515 13787
rect 29457 13747 29515 13753
rect 37369 13787 37427 13793
rect 37369 13753 37381 13787
rect 37415 13784 37427 13787
rect 38197 13787 38255 13793
rect 38197 13784 38209 13787
rect 37415 13756 38209 13784
rect 37415 13753 37427 13756
rect 37369 13747 37427 13753
rect 38197 13753 38209 13756
rect 38243 13784 38255 13787
rect 38473 13787 38531 13793
rect 38473 13784 38485 13787
rect 38243 13756 38485 13784
rect 38243 13753 38255 13756
rect 38197 13747 38255 13753
rect 38473 13753 38485 13756
rect 38519 13753 38531 13787
rect 38473 13747 38531 13753
rect 38565 13787 38623 13793
rect 38565 13753 38577 13787
rect 38611 13753 38623 13787
rect 38565 13747 38623 13753
rect 28215 13719 28273 13725
rect 28215 13716 28227 13719
rect 26384 13688 28227 13716
rect 26384 13676 26390 13688
rect 28215 13685 28227 13688
rect 28261 13685 28273 13719
rect 28215 13679 28273 13685
rect 29086 13676 29092 13728
rect 29144 13716 29150 13728
rect 29472 13716 29500 13747
rect 29144 13688 29500 13716
rect 31987 13719 32045 13725
rect 29144 13676 29150 13688
rect 31987 13685 31999 13719
rect 32033 13716 32045 13719
rect 32674 13716 32680 13728
rect 32033 13688 32680 13716
rect 32033 13685 32045 13688
rect 31987 13679 32045 13685
rect 32674 13676 32680 13688
rect 32732 13676 32738 13728
rect 33594 13676 33600 13728
rect 33652 13716 33658 13728
rect 33827 13719 33885 13725
rect 33827 13716 33839 13719
rect 33652 13688 33839 13716
rect 33652 13676 33658 13688
rect 33827 13685 33839 13688
rect 33873 13685 33885 13719
rect 35986 13716 35992 13728
rect 35947 13688 35992 13716
rect 33827 13679 33885 13685
rect 35986 13676 35992 13688
rect 36044 13676 36050 13728
rect 36541 13719 36599 13725
rect 36541 13685 36553 13719
rect 36587 13716 36599 13719
rect 36909 13719 36967 13725
rect 36909 13716 36921 13719
rect 36587 13688 36921 13716
rect 36587 13685 36599 13688
rect 36541 13679 36599 13685
rect 36909 13685 36921 13688
rect 36955 13716 36967 13719
rect 37921 13719 37979 13725
rect 37921 13716 37933 13719
rect 36955 13688 37933 13716
rect 36955 13685 36967 13688
rect 36909 13679 36967 13685
rect 37921 13685 37933 13688
rect 37967 13716 37979 13719
rect 38378 13716 38384 13728
rect 37967 13688 38384 13716
rect 37967 13685 37979 13688
rect 37921 13679 37979 13685
rect 38378 13676 38384 13688
rect 38436 13716 38442 13728
rect 38580 13716 38608 13747
rect 38436 13688 38608 13716
rect 38436 13676 38442 13688
rect 38654 13676 38660 13728
rect 38712 13716 38718 13728
rect 39393 13719 39451 13725
rect 39393 13716 39405 13719
rect 38712 13688 39405 13716
rect 38712 13676 38718 13688
rect 39393 13685 39405 13688
rect 39439 13685 39451 13719
rect 39393 13679 39451 13685
rect 39574 13676 39580 13728
rect 39632 13716 39638 13728
rect 40635 13719 40693 13725
rect 40635 13716 40647 13719
rect 39632 13688 40647 13716
rect 39632 13676 39638 13688
rect 40635 13685 40647 13688
rect 40681 13685 40693 13719
rect 40635 13679 40693 13685
rect 1104 13626 48852 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 48852 13626
rect 1104 13552 48852 13574
rect 9674 13472 9680 13524
rect 9732 13512 9738 13524
rect 9861 13515 9919 13521
rect 9861 13512 9873 13515
rect 9732 13484 9873 13512
rect 9732 13472 9738 13484
rect 9861 13481 9873 13484
rect 9907 13481 9919 13515
rect 9861 13475 9919 13481
rect 13262 13472 13268 13524
rect 13320 13512 13326 13524
rect 14090 13512 14096 13524
rect 13320 13484 13814 13512
rect 14051 13484 14096 13512
rect 13320 13472 13326 13484
rect 11514 13404 11520 13456
rect 11572 13444 11578 13456
rect 11609 13447 11667 13453
rect 11609 13444 11621 13447
rect 11572 13416 11621 13444
rect 11572 13404 11578 13416
rect 11609 13413 11621 13416
rect 11655 13444 11667 13447
rect 11974 13444 11980 13456
rect 11655 13416 11980 13444
rect 11655 13413 11667 13416
rect 11609 13407 11667 13413
rect 11974 13404 11980 13416
rect 12032 13404 12038 13456
rect 12158 13444 12164 13456
rect 12119 13416 12164 13444
rect 12158 13404 12164 13416
rect 12216 13404 12222 13456
rect 13535 13447 13593 13453
rect 13535 13413 13547 13447
rect 13581 13444 13593 13447
rect 13630 13444 13636 13456
rect 13581 13416 13636 13444
rect 13581 13413 13593 13416
rect 13535 13407 13593 13413
rect 13630 13404 13636 13416
rect 13688 13404 13694 13456
rect 13786 13444 13814 13484
rect 14090 13472 14096 13484
rect 14148 13472 14154 13524
rect 14826 13512 14832 13524
rect 14787 13484 14832 13512
rect 14826 13472 14832 13484
rect 14884 13472 14890 13524
rect 15654 13472 15660 13524
rect 15712 13512 15718 13524
rect 15749 13515 15807 13521
rect 15749 13512 15761 13515
rect 15712 13484 15761 13512
rect 15712 13472 15718 13484
rect 15749 13481 15761 13484
rect 15795 13481 15807 13515
rect 15749 13475 15807 13481
rect 18693 13515 18751 13521
rect 18693 13481 18705 13515
rect 18739 13512 18751 13515
rect 19153 13515 19211 13521
rect 19153 13512 19165 13515
rect 18739 13484 19165 13512
rect 18739 13481 18751 13484
rect 18693 13475 18751 13481
rect 19153 13481 19165 13484
rect 19199 13512 19211 13515
rect 19242 13512 19248 13524
rect 19199 13484 19248 13512
rect 19199 13481 19211 13484
rect 19153 13475 19211 13481
rect 19242 13472 19248 13484
rect 19300 13472 19306 13524
rect 20990 13512 20996 13524
rect 20951 13484 20996 13512
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 22646 13472 22652 13524
rect 22704 13512 22710 13524
rect 24029 13515 24087 13521
rect 22704 13484 22784 13512
rect 22704 13472 22710 13484
rect 15427 13447 15485 13453
rect 15427 13444 15439 13447
rect 13786 13416 15439 13444
rect 15427 13413 15439 13416
rect 15473 13413 15485 13447
rect 15427 13407 15485 13413
rect 16206 13404 16212 13456
rect 16264 13444 16270 13456
rect 16945 13447 17003 13453
rect 16945 13444 16957 13447
rect 16264 13416 16957 13444
rect 16264 13404 16270 13416
rect 16945 13413 16957 13416
rect 16991 13444 17003 13447
rect 17034 13444 17040 13456
rect 16991 13416 17040 13444
rect 16991 13413 17003 13416
rect 16945 13407 17003 13413
rect 17034 13404 17040 13416
rect 17092 13404 17098 13456
rect 22756 13453 22784 13484
rect 22848 13484 23704 13512
rect 22848 13456 22876 13484
rect 22741 13447 22799 13453
rect 22741 13413 22753 13447
rect 22787 13413 22799 13447
rect 22741 13407 22799 13413
rect 22830 13404 22836 13456
rect 22888 13444 22894 13456
rect 22888 13416 22933 13444
rect 22888 13404 22894 13416
rect 23014 13404 23020 13456
rect 23072 13444 23078 13456
rect 23676 13444 23704 13484
rect 24029 13481 24041 13515
rect 24075 13512 24087 13515
rect 24118 13512 24124 13524
rect 24075 13484 24124 13512
rect 24075 13481 24087 13484
rect 24029 13475 24087 13481
rect 24118 13472 24124 13484
rect 24176 13472 24182 13524
rect 26326 13512 26332 13524
rect 26287 13484 26332 13512
rect 26326 13472 26332 13484
rect 26384 13472 26390 13524
rect 27433 13515 27491 13521
rect 27433 13481 27445 13515
rect 27479 13512 27491 13515
rect 28169 13515 28227 13521
rect 28169 13512 28181 13515
rect 27479 13484 28181 13512
rect 27479 13481 27491 13484
rect 27433 13475 27491 13481
rect 28169 13481 28181 13484
rect 28215 13512 28227 13515
rect 28258 13512 28264 13524
rect 28215 13484 28264 13512
rect 28215 13481 28227 13484
rect 28169 13475 28227 13481
rect 28258 13472 28264 13484
rect 28316 13472 28322 13524
rect 28626 13512 28632 13524
rect 28587 13484 28632 13512
rect 28626 13472 28632 13484
rect 28684 13472 28690 13524
rect 29362 13472 29368 13524
rect 29420 13512 29426 13524
rect 30147 13515 30205 13521
rect 30147 13512 30159 13515
rect 29420 13484 30159 13512
rect 29420 13472 29426 13484
rect 30147 13481 30159 13484
rect 30193 13481 30205 13515
rect 35618 13512 35624 13524
rect 35579 13484 35624 13512
rect 30147 13475 30205 13481
rect 35618 13472 35624 13484
rect 35676 13472 35682 13524
rect 38378 13472 38384 13524
rect 38436 13512 38442 13524
rect 38749 13515 38807 13521
rect 38749 13512 38761 13515
rect 38436 13484 38761 13512
rect 38436 13472 38442 13484
rect 38749 13481 38761 13484
rect 38795 13481 38807 13515
rect 38749 13475 38807 13481
rect 24397 13447 24455 13453
rect 24397 13444 24409 13447
rect 23072 13416 23474 13444
rect 23676 13416 24409 13444
rect 23072 13404 23078 13416
rect 10042 13376 10048 13388
rect 10003 13348 10048 13376
rect 10042 13336 10048 13348
rect 10100 13336 10106 13388
rect 10226 13376 10232 13388
rect 10187 13348 10232 13376
rect 10226 13336 10232 13348
rect 10284 13336 10290 13388
rect 15194 13376 15200 13388
rect 15155 13348 15200 13376
rect 15194 13336 15200 13348
rect 15252 13336 15258 13388
rect 18690 13336 18696 13388
rect 18748 13376 18754 13388
rect 18877 13379 18935 13385
rect 18877 13376 18889 13379
rect 18748 13348 18889 13376
rect 18748 13336 18754 13348
rect 18877 13345 18889 13348
rect 18923 13345 18935 13379
rect 18877 13339 18935 13345
rect 19061 13379 19119 13385
rect 19061 13345 19073 13379
rect 19107 13376 19119 13379
rect 19242 13376 19248 13388
rect 19107 13348 19248 13376
rect 19107 13345 19119 13348
rect 19061 13339 19119 13345
rect 19242 13336 19248 13348
rect 19300 13336 19306 13388
rect 20438 13336 20444 13388
rect 20496 13376 20502 13388
rect 20901 13379 20959 13385
rect 20901 13376 20913 13379
rect 20496 13348 20913 13376
rect 20496 13336 20502 13348
rect 20901 13345 20913 13348
rect 20947 13376 20959 13379
rect 21082 13376 21088 13388
rect 20947 13348 21088 13376
rect 20947 13345 20959 13348
rect 20901 13339 20959 13345
rect 21082 13336 21088 13348
rect 21140 13336 21146 13388
rect 21174 13336 21180 13388
rect 21232 13376 21238 13388
rect 21361 13379 21419 13385
rect 21361 13376 21373 13379
rect 21232 13348 21373 13376
rect 21232 13336 21238 13348
rect 21361 13345 21373 13348
rect 21407 13345 21419 13379
rect 21361 13339 21419 13345
rect 11330 13268 11336 13320
rect 11388 13308 11394 13320
rect 11517 13311 11575 13317
rect 11517 13308 11529 13311
rect 11388 13280 11529 13308
rect 11388 13268 11394 13280
rect 11517 13277 11529 13280
rect 11563 13277 11575 13311
rect 11517 13271 11575 13277
rect 13173 13311 13231 13317
rect 13173 13277 13185 13311
rect 13219 13308 13231 13311
rect 13906 13308 13912 13320
rect 13219 13280 13912 13308
rect 13219 13277 13231 13280
rect 13173 13271 13231 13277
rect 13906 13268 13912 13280
rect 13964 13268 13970 13320
rect 16114 13268 16120 13320
rect 16172 13308 16178 13320
rect 16850 13308 16856 13320
rect 16172 13280 16856 13308
rect 16172 13268 16178 13280
rect 16850 13268 16856 13280
rect 16908 13268 16914 13320
rect 17126 13308 17132 13320
rect 17087 13280 17132 13308
rect 17126 13268 17132 13280
rect 17184 13268 17190 13320
rect 23106 13308 23112 13320
rect 23067 13280 23112 13308
rect 23106 13268 23112 13280
rect 23164 13268 23170 13320
rect 23446 13308 23474 13416
rect 24397 13413 24409 13416
rect 24443 13413 24455 13447
rect 24397 13407 24455 13413
rect 26875 13447 26933 13453
rect 26875 13413 26887 13447
rect 26921 13444 26933 13447
rect 26970 13444 26976 13456
rect 26921 13416 26976 13444
rect 26921 13413 26933 13416
rect 26875 13407 26933 13413
rect 26970 13404 26976 13416
rect 27028 13404 27034 13456
rect 35345 13447 35403 13453
rect 35345 13413 35357 13447
rect 35391 13444 35403 13447
rect 35526 13444 35532 13456
rect 35391 13416 35532 13444
rect 35391 13413 35403 13416
rect 35345 13407 35403 13413
rect 35526 13404 35532 13416
rect 35584 13404 35590 13456
rect 35986 13404 35992 13456
rect 36044 13444 36050 13456
rect 36167 13447 36225 13453
rect 36167 13444 36179 13447
rect 36044 13416 36179 13444
rect 36044 13404 36050 13416
rect 36167 13413 36179 13416
rect 36213 13413 36225 13447
rect 36167 13407 36225 13413
rect 37642 13404 37648 13456
rect 37700 13444 37706 13456
rect 37921 13447 37979 13453
rect 37921 13444 37933 13447
rect 37700 13416 37933 13444
rect 37700 13404 37706 13416
rect 37921 13413 37933 13416
rect 37967 13413 37979 13447
rect 39482 13444 39488 13456
rect 39443 13416 39488 13444
rect 37921 13407 37979 13413
rect 39482 13404 39488 13416
rect 39540 13404 39546 13456
rect 29181 13379 29239 13385
rect 29181 13345 29193 13379
rect 29227 13376 29239 13379
rect 30044 13379 30102 13385
rect 30044 13376 30056 13379
rect 29227 13348 30056 13376
rect 29227 13345 29239 13348
rect 29181 13339 29239 13345
rect 30044 13345 30056 13348
rect 30090 13376 30102 13379
rect 30466 13376 30472 13388
rect 30090 13348 30472 13376
rect 30090 13345 30102 13348
rect 30044 13339 30102 13345
rect 30466 13336 30472 13348
rect 30524 13336 30530 13388
rect 32192 13379 32250 13385
rect 32192 13345 32204 13379
rect 32238 13376 32250 13379
rect 33134 13376 33140 13388
rect 32238 13348 33140 13376
rect 32238 13345 32250 13348
rect 32192 13339 32250 13345
rect 33134 13336 33140 13348
rect 33192 13376 33198 13388
rect 33192 13348 33285 13376
rect 33192 13336 33198 13348
rect 34698 13336 34704 13388
rect 34756 13376 34762 13388
rect 34828 13379 34886 13385
rect 34828 13376 34840 13379
rect 34756 13348 34840 13376
rect 34756 13336 34762 13348
rect 34828 13345 34840 13348
rect 34874 13345 34886 13379
rect 34828 13339 34886 13345
rect 24305 13311 24363 13317
rect 24305 13308 24317 13311
rect 23446 13280 24317 13308
rect 24305 13277 24317 13280
rect 24351 13308 24363 13311
rect 24578 13308 24584 13320
rect 24351 13280 24584 13308
rect 24351 13277 24363 13280
rect 24305 13271 24363 13277
rect 24578 13268 24584 13280
rect 24636 13268 24642 13320
rect 24762 13308 24768 13320
rect 24723 13280 24768 13308
rect 24762 13268 24768 13280
rect 24820 13268 24826 13320
rect 26510 13308 26516 13320
rect 26471 13280 26516 13308
rect 26510 13268 26516 13280
rect 26568 13268 26574 13320
rect 28258 13308 28264 13320
rect 28219 13280 28264 13308
rect 28258 13268 28264 13280
rect 28316 13268 28322 13320
rect 35802 13308 35808 13320
rect 35763 13280 35808 13308
rect 35802 13268 35808 13280
rect 35860 13268 35866 13320
rect 37829 13311 37887 13317
rect 37829 13277 37841 13311
rect 37875 13308 37887 13311
rect 37918 13308 37924 13320
rect 37875 13280 37924 13308
rect 37875 13277 37887 13280
rect 37829 13271 37887 13277
rect 37918 13268 37924 13280
rect 37976 13268 37982 13320
rect 39206 13268 39212 13320
rect 39264 13308 39270 13320
rect 39393 13311 39451 13317
rect 39393 13308 39405 13311
rect 39264 13280 39405 13308
rect 39264 13268 39270 13280
rect 39393 13277 39405 13280
rect 39439 13308 39451 13311
rect 40218 13308 40224 13320
rect 39439 13280 40224 13308
rect 39439 13277 39451 13280
rect 39393 13271 39451 13277
rect 40218 13268 40224 13280
rect 40276 13268 40282 13320
rect 34931 13243 34989 13249
rect 34931 13209 34943 13243
rect 34977 13240 34989 13243
rect 38102 13240 38108 13252
rect 34977 13212 38108 13240
rect 34977 13209 34989 13212
rect 34931 13203 34989 13209
rect 38102 13200 38108 13212
rect 38160 13200 38166 13252
rect 38378 13240 38384 13252
rect 38339 13212 38384 13240
rect 38378 13200 38384 13212
rect 38436 13240 38442 13252
rect 39945 13243 40003 13249
rect 39945 13240 39957 13243
rect 38436 13212 39957 13240
rect 38436 13200 38442 13212
rect 39945 13209 39957 13212
rect 39991 13209 40003 13243
rect 39945 13203 40003 13209
rect 10134 13132 10140 13184
rect 10192 13172 10198 13184
rect 10781 13175 10839 13181
rect 10781 13172 10793 13175
rect 10192 13144 10793 13172
rect 10192 13132 10198 13144
rect 10781 13141 10793 13144
rect 10827 13141 10839 13175
rect 16574 13172 16580 13184
rect 16535 13144 16580 13172
rect 10781 13135 10839 13141
rect 16574 13132 16580 13144
rect 16632 13132 16638 13184
rect 17862 13172 17868 13184
rect 17823 13144 17868 13172
rect 17862 13132 17868 13144
rect 17920 13132 17926 13184
rect 20441 13175 20499 13181
rect 20441 13141 20453 13175
rect 20487 13172 20499 13175
rect 20530 13172 20536 13184
rect 20487 13144 20536 13172
rect 20487 13141 20499 13144
rect 20441 13135 20499 13141
rect 20530 13132 20536 13144
rect 20588 13132 20594 13184
rect 22557 13175 22615 13181
rect 22557 13141 22569 13175
rect 22603 13172 22615 13175
rect 22738 13172 22744 13184
rect 22603 13144 22744 13172
rect 22603 13141 22615 13144
rect 22557 13135 22615 13141
rect 22738 13132 22744 13144
rect 22796 13172 22802 13184
rect 22922 13172 22928 13184
rect 22796 13144 22928 13172
rect 22796 13132 22802 13144
rect 22922 13132 22928 13144
rect 22980 13132 22986 13184
rect 25590 13172 25596 13184
rect 25551 13144 25596 13172
rect 25590 13132 25596 13144
rect 25648 13132 25654 13184
rect 27798 13172 27804 13184
rect 27759 13144 27804 13172
rect 27798 13132 27804 13144
rect 27856 13132 27862 13184
rect 29454 13172 29460 13184
rect 29415 13144 29460 13172
rect 29454 13132 29460 13144
rect 29512 13132 29518 13184
rect 31018 13172 31024 13184
rect 30979 13144 31024 13172
rect 31018 13132 31024 13144
rect 31076 13132 31082 13184
rect 32263 13175 32321 13181
rect 32263 13141 32275 13175
rect 32309 13172 32321 13175
rect 32582 13172 32588 13184
rect 32309 13144 32588 13172
rect 32309 13141 32321 13144
rect 32263 13135 32321 13141
rect 32582 13132 32588 13144
rect 32640 13132 32646 13184
rect 33318 13172 33324 13184
rect 33279 13144 33324 13172
rect 33318 13132 33324 13144
rect 33376 13132 33382 13184
rect 36725 13175 36783 13181
rect 36725 13141 36737 13175
rect 36771 13172 36783 13175
rect 37642 13172 37648 13184
rect 36771 13144 37648 13172
rect 36771 13141 36783 13144
rect 36725 13135 36783 13141
rect 37642 13132 37648 13144
rect 37700 13132 37706 13184
rect 37826 13132 37832 13184
rect 37884 13172 37890 13184
rect 40402 13172 40408 13184
rect 37884 13144 40408 13172
rect 37884 13132 37890 13144
rect 40402 13132 40408 13144
rect 40460 13132 40466 13184
rect 1104 13082 48852 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 48852 13082
rect 1104 13008 48852 13030
rect 9263 12971 9321 12977
rect 9263 12937 9275 12971
rect 9309 12968 9321 12971
rect 11330 12968 11336 12980
rect 9309 12940 11336 12968
rect 9309 12937 9321 12940
rect 9263 12931 9321 12937
rect 11330 12928 11336 12940
rect 11388 12928 11394 12980
rect 11514 12968 11520 12980
rect 11475 12940 11520 12968
rect 11514 12928 11520 12940
rect 11572 12928 11578 12980
rect 13081 12971 13139 12977
rect 13081 12937 13093 12971
rect 13127 12968 13139 12971
rect 13630 12968 13636 12980
rect 13127 12940 13636 12968
rect 13127 12937 13139 12940
rect 13081 12931 13139 12937
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 16114 12968 16120 12980
rect 16075 12940 16120 12968
rect 16114 12928 16120 12940
rect 16172 12928 16178 12980
rect 16206 12928 16212 12980
rect 16264 12968 16270 12980
rect 16393 12971 16451 12977
rect 16393 12968 16405 12971
rect 16264 12940 16405 12968
rect 16264 12928 16270 12940
rect 16393 12937 16405 12940
rect 16439 12937 16451 12971
rect 16393 12931 16451 12937
rect 17862 12928 17868 12980
rect 17920 12968 17926 12980
rect 19337 12971 19395 12977
rect 19337 12968 19349 12971
rect 17920 12940 19349 12968
rect 17920 12928 17926 12940
rect 19337 12937 19349 12940
rect 19383 12937 19395 12971
rect 19337 12931 19395 12937
rect 22646 12928 22652 12980
rect 22704 12968 22710 12980
rect 23017 12971 23075 12977
rect 23017 12968 23029 12971
rect 22704 12940 23029 12968
rect 22704 12928 22710 12940
rect 23017 12937 23029 12940
rect 23063 12937 23075 12971
rect 23017 12931 23075 12937
rect 23799 12971 23857 12977
rect 23799 12937 23811 12971
rect 23845 12968 23857 12971
rect 24026 12968 24032 12980
rect 23845 12940 24032 12968
rect 23845 12937 23857 12940
rect 23799 12931 23857 12937
rect 24026 12928 24032 12940
rect 24084 12928 24090 12980
rect 24578 12968 24584 12980
rect 24539 12940 24584 12968
rect 24578 12928 24584 12940
rect 24636 12928 24642 12980
rect 25590 12928 25596 12980
rect 25648 12968 25654 12980
rect 26513 12971 26571 12977
rect 26513 12968 26525 12971
rect 25648 12940 26525 12968
rect 25648 12928 25654 12940
rect 26513 12937 26525 12940
rect 26559 12937 26571 12971
rect 26513 12931 26571 12937
rect 29178 12928 29184 12980
rect 29236 12968 29242 12980
rect 30193 12971 30251 12977
rect 30193 12968 30205 12971
rect 29236 12940 30205 12968
rect 29236 12928 29242 12940
rect 30193 12937 30205 12940
rect 30239 12937 30251 12971
rect 30466 12968 30472 12980
rect 30427 12940 30472 12968
rect 30193 12931 30251 12937
rect 30466 12928 30472 12940
rect 30524 12928 30530 12980
rect 32582 12968 32588 12980
rect 32543 12940 32588 12968
rect 32582 12928 32588 12940
rect 32640 12928 32646 12980
rect 36771 12971 36829 12977
rect 36771 12937 36783 12971
rect 36817 12968 36829 12971
rect 36906 12968 36912 12980
rect 36817 12940 36912 12968
rect 36817 12937 36829 12940
rect 36771 12931 36829 12937
rect 36906 12928 36912 12940
rect 36964 12928 36970 12980
rect 37642 12968 37648 12980
rect 37603 12940 37648 12968
rect 37642 12928 37648 12940
rect 37700 12928 37706 12980
rect 38194 12928 38200 12980
rect 38252 12968 38258 12980
rect 38289 12971 38347 12977
rect 38289 12968 38301 12971
rect 38252 12940 38301 12968
rect 38252 12928 38258 12940
rect 38289 12937 38301 12940
rect 38335 12937 38347 12971
rect 38289 12931 38347 12937
rect 39482 12928 39488 12980
rect 39540 12968 39546 12980
rect 39853 12971 39911 12977
rect 39853 12968 39865 12971
rect 39540 12940 39865 12968
rect 39540 12928 39546 12940
rect 39853 12937 39865 12940
rect 39899 12968 39911 12971
rect 39942 12968 39948 12980
rect 39899 12940 39948 12968
rect 39899 12937 39911 12940
rect 39853 12931 39911 12937
rect 39942 12928 39948 12940
rect 40000 12928 40006 12980
rect 40218 12968 40224 12980
rect 40179 12940 40224 12968
rect 40218 12928 40224 12940
rect 40276 12928 40282 12980
rect 8251 12903 8309 12909
rect 8251 12869 8263 12903
rect 8297 12900 8309 12903
rect 11146 12900 11152 12912
rect 8297 12872 11152 12900
rect 8297 12869 8309 12872
rect 8251 12863 8309 12869
rect 11146 12860 11152 12872
rect 11204 12860 11210 12912
rect 11348 12900 11376 12928
rect 12161 12903 12219 12909
rect 12161 12900 12173 12903
rect 11348 12872 12173 12900
rect 12161 12869 12173 12872
rect 12207 12869 12219 12903
rect 14090 12900 14096 12912
rect 12161 12863 12219 12869
rect 13786 12872 14096 12900
rect 9861 12835 9919 12841
rect 9861 12801 9873 12835
rect 9907 12832 9919 12835
rect 10042 12832 10048 12844
rect 9907 12804 10048 12832
rect 9907 12801 9919 12804
rect 9861 12795 9919 12801
rect 10042 12792 10048 12804
rect 10100 12832 10106 12844
rect 13786 12832 13814 12872
rect 14090 12860 14096 12872
rect 14148 12860 14154 12912
rect 18322 12900 18328 12912
rect 18283 12872 18328 12900
rect 18322 12860 18328 12872
rect 18380 12860 18386 12912
rect 22741 12903 22799 12909
rect 22741 12869 22753 12903
rect 22787 12900 22799 12903
rect 22830 12900 22836 12912
rect 22787 12872 22836 12900
rect 22787 12869 22799 12872
rect 22741 12863 22799 12869
rect 22830 12860 22836 12872
rect 22888 12900 22894 12912
rect 24213 12903 24271 12909
rect 24213 12900 24225 12903
rect 22888 12872 24225 12900
rect 22888 12860 22894 12872
rect 24213 12869 24225 12872
rect 24259 12869 24271 12903
rect 24213 12863 24271 12869
rect 25501 12903 25559 12909
rect 25501 12869 25513 12903
rect 25547 12900 25559 12903
rect 26881 12903 26939 12909
rect 26881 12900 26893 12903
rect 25547 12872 26893 12900
rect 25547 12869 25559 12872
rect 25501 12863 25559 12869
rect 13906 12832 13912 12844
rect 10100 12804 13814 12832
rect 13867 12804 13912 12832
rect 10100 12792 10106 12804
rect 13906 12792 13912 12804
rect 13964 12792 13970 12844
rect 17129 12835 17187 12841
rect 17129 12801 17141 12835
rect 17175 12832 17187 12835
rect 18230 12832 18236 12844
rect 17175 12804 18236 12832
rect 17175 12801 17187 12804
rect 17129 12795 17187 12801
rect 18230 12792 18236 12804
rect 18288 12792 18294 12844
rect 20073 12835 20131 12841
rect 20073 12801 20085 12835
rect 20119 12832 20131 12835
rect 20901 12835 20959 12841
rect 20901 12832 20913 12835
rect 20119 12804 20913 12832
rect 20119 12801 20131 12804
rect 20073 12795 20131 12801
rect 20901 12801 20913 12804
rect 20947 12832 20959 12835
rect 20990 12832 20996 12844
rect 20947 12804 20996 12832
rect 20947 12801 20959 12804
rect 20901 12795 20959 12801
rect 20990 12792 20996 12804
rect 21048 12792 21054 12844
rect 8180 12767 8238 12773
rect 8180 12733 8192 12767
rect 8226 12764 8238 12767
rect 9030 12764 9036 12776
rect 8226 12736 8708 12764
rect 8991 12736 9036 12764
rect 8226 12733 8238 12736
rect 8180 12727 8238 12733
rect 8680 12640 8708 12736
rect 9030 12724 9036 12736
rect 9088 12764 9094 12776
rect 9160 12767 9218 12773
rect 9160 12764 9172 12767
rect 9088 12736 9172 12764
rect 9088 12724 9094 12736
rect 9160 12733 9172 12736
rect 9206 12733 9218 12767
rect 9160 12727 9218 12733
rect 9674 12724 9680 12776
rect 9732 12764 9738 12776
rect 10134 12764 10140 12776
rect 9732 12736 10140 12764
rect 9732 12724 9738 12736
rect 10134 12724 10140 12736
rect 10192 12724 10198 12776
rect 10226 12724 10232 12776
rect 10284 12764 10290 12776
rect 10597 12767 10655 12773
rect 10597 12764 10609 12767
rect 10284 12736 10609 12764
rect 10284 12724 10290 12736
rect 10597 12733 10609 12736
rect 10643 12764 10655 12767
rect 11793 12767 11851 12773
rect 11793 12764 11805 12767
rect 10643 12736 11805 12764
rect 10643 12733 10655 12736
rect 10597 12727 10655 12733
rect 11793 12733 11805 12736
rect 11839 12733 11851 12767
rect 11793 12727 11851 12733
rect 12713 12767 12771 12773
rect 12713 12733 12725 12767
rect 12759 12764 12771 12767
rect 12894 12764 12900 12776
rect 12759 12736 12900 12764
rect 12759 12733 12771 12736
rect 12713 12727 12771 12733
rect 11808 12696 11836 12727
rect 12894 12724 12900 12736
rect 12952 12764 12958 12776
rect 13173 12767 13231 12773
rect 13173 12764 13185 12767
rect 12952 12736 13185 12764
rect 12952 12724 12958 12736
rect 13173 12733 13185 12736
rect 13219 12733 13231 12767
rect 13173 12727 13231 12733
rect 13633 12767 13691 12773
rect 13633 12733 13645 12767
rect 13679 12764 13691 12767
rect 14182 12764 14188 12776
rect 13679 12736 14188 12764
rect 13679 12733 13691 12736
rect 13633 12727 13691 12733
rect 12802 12696 12808 12708
rect 11808 12668 12808 12696
rect 12802 12656 12808 12668
rect 12860 12696 12866 12708
rect 13648 12696 13676 12727
rect 14182 12724 14188 12736
rect 14240 12724 14246 12776
rect 14829 12767 14887 12773
rect 14829 12733 14841 12767
rect 14875 12764 14887 12767
rect 14921 12767 14979 12773
rect 14921 12764 14933 12767
rect 14875 12736 14933 12764
rect 14875 12733 14887 12736
rect 14829 12727 14887 12733
rect 14921 12733 14933 12736
rect 14967 12733 14979 12767
rect 15378 12764 15384 12776
rect 15339 12736 15384 12764
rect 14921 12727 14979 12733
rect 12860 12668 13676 12696
rect 14936 12696 14964 12727
rect 15378 12724 15384 12736
rect 15436 12724 15442 12776
rect 16761 12767 16819 12773
rect 16761 12733 16773 12767
rect 16807 12764 16819 12767
rect 17865 12767 17923 12773
rect 16807 12736 17540 12764
rect 16807 12733 16819 12736
rect 16761 12727 16819 12733
rect 15746 12696 15752 12708
rect 14936 12668 15752 12696
rect 12860 12656 12866 12668
rect 15746 12656 15752 12668
rect 15804 12656 15810 12708
rect 16574 12696 16580 12708
rect 16535 12668 16580 12696
rect 16574 12656 16580 12668
rect 16632 12656 16638 12708
rect 17512 12696 17540 12736
rect 17865 12733 17877 12767
rect 17911 12764 17923 12767
rect 18417 12767 18475 12773
rect 18417 12764 18429 12767
rect 17911 12736 18429 12764
rect 17911 12733 17923 12736
rect 17865 12727 17923 12733
rect 18417 12733 18429 12736
rect 18463 12764 18475 12767
rect 18506 12764 18512 12776
rect 18463 12736 18512 12764
rect 18463 12733 18475 12736
rect 18417 12727 18475 12733
rect 18506 12724 18512 12736
rect 18564 12724 18570 12776
rect 23477 12767 23535 12773
rect 23477 12733 23489 12767
rect 23523 12764 23535 12767
rect 23696 12767 23754 12773
rect 23696 12764 23708 12767
rect 23523 12736 23708 12764
rect 23523 12733 23535 12736
rect 23477 12727 23535 12733
rect 23696 12733 23708 12736
rect 23742 12764 23754 12767
rect 23934 12764 23940 12776
rect 23742 12736 23940 12764
rect 23742 12733 23754 12736
rect 23696 12727 23754 12733
rect 23934 12724 23940 12736
rect 23992 12724 23998 12776
rect 25130 12764 25136 12776
rect 25043 12736 25136 12764
rect 25130 12724 25136 12736
rect 25188 12764 25194 12776
rect 25593 12767 25651 12773
rect 25593 12764 25605 12767
rect 25188 12736 25605 12764
rect 25188 12724 25194 12736
rect 25593 12733 25605 12736
rect 25639 12733 25651 12767
rect 25593 12727 25651 12733
rect 21266 12705 21272 12708
rect 18738 12699 18796 12705
rect 17512 12668 18368 12696
rect 17512 12640 17540 12668
rect 8662 12628 8668 12640
rect 8623 12600 8668 12628
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 10226 12628 10232 12640
rect 10187 12600 10232 12628
rect 10226 12588 10232 12600
rect 10284 12588 10290 12640
rect 15010 12628 15016 12640
rect 14971 12600 15016 12628
rect 15010 12588 15016 12600
rect 15068 12588 15074 12640
rect 17494 12628 17500 12640
rect 17455 12600 17500 12628
rect 17494 12588 17500 12600
rect 17552 12588 17558 12640
rect 18340 12628 18368 12668
rect 18738 12665 18750 12699
rect 18784 12696 18796 12699
rect 20717 12699 20775 12705
rect 20717 12696 20729 12699
rect 18784 12668 20729 12696
rect 18784 12665 18796 12668
rect 18738 12659 18796 12665
rect 20717 12665 20729 12668
rect 20763 12696 20775 12699
rect 21222 12699 21272 12705
rect 21222 12696 21234 12699
rect 20763 12668 21234 12696
rect 20763 12665 20775 12668
rect 20717 12659 20775 12665
rect 21222 12665 21234 12668
rect 21268 12665 21272 12699
rect 21222 12659 21272 12665
rect 21266 12656 21272 12659
rect 21324 12656 21330 12708
rect 25929 12705 25957 12872
rect 26881 12869 26893 12872
rect 26927 12900 26939 12903
rect 26970 12900 26976 12912
rect 26927 12872 26976 12900
rect 26927 12869 26939 12872
rect 26881 12863 26939 12869
rect 26970 12860 26976 12872
rect 27028 12900 27034 12912
rect 28626 12900 28632 12912
rect 27028 12872 28632 12900
rect 27028 12860 27034 12872
rect 28626 12860 28632 12872
rect 28684 12860 28690 12912
rect 32309 12903 32367 12909
rect 32309 12869 32321 12903
rect 32355 12900 32367 12903
rect 33134 12900 33140 12912
rect 32355 12872 33140 12900
rect 32355 12869 32367 12872
rect 32309 12863 32367 12869
rect 33134 12860 33140 12872
rect 33192 12900 33198 12912
rect 33873 12903 33931 12909
rect 33873 12900 33885 12903
rect 33192 12872 33885 12900
rect 33192 12860 33198 12872
rect 33873 12869 33885 12872
rect 33919 12900 33931 12903
rect 37826 12900 37832 12912
rect 33919 12872 37832 12900
rect 33919 12869 33931 12872
rect 33873 12863 33931 12869
rect 37826 12860 37832 12872
rect 37884 12860 37890 12912
rect 37967 12903 38025 12909
rect 37967 12869 37979 12903
rect 38013 12900 38025 12903
rect 38470 12900 38476 12912
rect 38013 12872 38476 12900
rect 38013 12869 38025 12872
rect 37967 12863 38025 12869
rect 38470 12860 38476 12872
rect 38528 12860 38534 12912
rect 28353 12835 28411 12841
rect 28353 12801 28365 12835
rect 28399 12832 28411 12835
rect 29273 12835 29331 12841
rect 29273 12832 29285 12835
rect 28399 12804 29285 12832
rect 28399 12801 28411 12804
rect 28353 12795 28411 12801
rect 29273 12801 29285 12804
rect 29319 12832 29331 12835
rect 29454 12832 29460 12844
rect 29319 12804 29460 12832
rect 29319 12801 29331 12804
rect 29273 12795 29331 12801
rect 29454 12792 29460 12804
rect 29512 12792 29518 12844
rect 35802 12832 35808 12844
rect 35715 12804 35808 12832
rect 35802 12792 35808 12804
rect 35860 12832 35866 12844
rect 36449 12835 36507 12841
rect 36449 12832 36461 12835
rect 35860 12804 36461 12832
rect 35860 12792 35866 12804
rect 36449 12801 36461 12804
rect 36495 12801 36507 12835
rect 36449 12795 36507 12801
rect 38378 12792 38384 12844
rect 38436 12832 38442 12844
rect 39209 12835 39267 12841
rect 39209 12832 39221 12835
rect 38436 12804 39221 12832
rect 38436 12792 38442 12804
rect 39209 12801 39221 12804
rect 39255 12801 39267 12835
rect 39209 12795 39267 12801
rect 27154 12724 27160 12776
rect 27212 12764 27218 12776
rect 27617 12767 27675 12773
rect 27617 12764 27629 12767
rect 27212 12736 27629 12764
rect 27212 12724 27218 12736
rect 25914 12699 25972 12705
rect 25914 12665 25926 12699
rect 25960 12665 25972 12699
rect 25914 12659 25972 12665
rect 27448 12640 27476 12736
rect 27617 12733 27629 12736
rect 27663 12733 27675 12767
rect 27617 12727 27675 12733
rect 27798 12724 27804 12776
rect 27856 12764 27862 12776
rect 28169 12767 28227 12773
rect 28169 12764 28181 12767
rect 27856 12736 28181 12764
rect 27856 12724 27862 12736
rect 28169 12733 28181 12736
rect 28215 12764 28227 12767
rect 28718 12764 28724 12776
rect 28215 12736 28724 12764
rect 28215 12733 28227 12736
rect 28169 12727 28227 12733
rect 28718 12724 28724 12736
rect 28776 12724 28782 12776
rect 30466 12724 30472 12776
rect 30524 12764 30530 12776
rect 31018 12764 31024 12776
rect 30524 12736 31024 12764
rect 30524 12724 30530 12736
rect 31018 12724 31024 12736
rect 31076 12724 31082 12776
rect 32582 12724 32588 12776
rect 32640 12764 32646 12776
rect 32861 12767 32919 12773
rect 32861 12764 32873 12767
rect 32640 12736 32873 12764
rect 32640 12724 32646 12736
rect 32861 12733 32873 12736
rect 32907 12733 32919 12767
rect 35342 12764 35348 12776
rect 35303 12736 35348 12764
rect 32861 12727 32919 12733
rect 35342 12724 35348 12736
rect 35400 12724 35406 12776
rect 35526 12764 35532 12776
rect 35487 12736 35532 12764
rect 35526 12724 35532 12736
rect 35584 12724 35590 12776
rect 36668 12767 36726 12773
rect 36668 12733 36680 12767
rect 36714 12733 36726 12767
rect 36668 12727 36726 12733
rect 37896 12767 37954 12773
rect 37896 12733 37908 12767
rect 37942 12764 37954 12767
rect 38194 12764 38200 12776
rect 37942 12736 38200 12764
rect 37942 12733 37954 12736
rect 37896 12727 37954 12733
rect 28626 12696 28632 12708
rect 28539 12668 28632 12696
rect 28626 12656 28632 12668
rect 28684 12696 28690 12708
rect 29089 12699 29147 12705
rect 29089 12696 29101 12699
rect 28684 12668 29101 12696
rect 28684 12656 28690 12668
rect 29089 12665 29101 12668
rect 29135 12696 29147 12699
rect 29635 12699 29693 12705
rect 29635 12696 29647 12699
rect 29135 12668 29647 12696
rect 29135 12665 29147 12668
rect 29089 12659 29147 12665
rect 29635 12665 29647 12668
rect 29681 12696 29693 12699
rect 30926 12696 30932 12708
rect 29681 12668 30932 12696
rect 29681 12665 29693 12668
rect 29635 12659 29693 12665
rect 30926 12656 30932 12668
rect 30984 12696 30990 12708
rect 31383 12699 31441 12705
rect 31383 12696 31395 12699
rect 30984 12668 31395 12696
rect 30984 12656 30990 12668
rect 31383 12665 31395 12668
rect 31429 12696 31441 12699
rect 32398 12696 32404 12708
rect 31429 12668 32404 12696
rect 31429 12665 31441 12668
rect 31383 12659 31441 12665
rect 32398 12656 32404 12668
rect 32456 12656 32462 12708
rect 32766 12696 32772 12708
rect 32727 12668 32772 12696
rect 32766 12656 32772 12668
rect 32824 12656 32830 12708
rect 35434 12656 35440 12708
rect 35492 12696 35498 12708
rect 36683 12696 36711 12727
rect 38194 12724 38200 12736
rect 38252 12724 38258 12776
rect 37093 12699 37151 12705
rect 37093 12696 37105 12699
rect 35492 12668 37105 12696
rect 35492 12656 35498 12668
rect 37093 12665 37105 12668
rect 37139 12665 37151 12699
rect 38930 12696 38936 12708
rect 38891 12668 38936 12696
rect 37093 12659 37151 12665
rect 38930 12656 38936 12668
rect 38988 12656 38994 12708
rect 39025 12699 39083 12705
rect 39025 12665 39037 12699
rect 39071 12665 39083 12699
rect 39025 12659 39083 12665
rect 19242 12628 19248 12640
rect 18340 12600 19248 12628
rect 19242 12588 19248 12600
rect 19300 12628 19306 12640
rect 19613 12631 19671 12637
rect 19613 12628 19625 12631
rect 19300 12600 19625 12628
rect 19300 12588 19306 12600
rect 19613 12597 19625 12600
rect 19659 12597 19671 12631
rect 20438 12628 20444 12640
rect 20399 12600 20444 12628
rect 19613 12591 19671 12597
rect 20438 12588 20444 12600
rect 20496 12588 20502 12640
rect 21818 12628 21824 12640
rect 21779 12600 21824 12628
rect 21818 12588 21824 12600
rect 21876 12588 21882 12640
rect 27430 12628 27436 12640
rect 27391 12600 27436 12628
rect 27430 12588 27436 12600
rect 27488 12588 27494 12640
rect 31938 12628 31944 12640
rect 31899 12600 31944 12628
rect 31938 12588 31944 12600
rect 31996 12588 32002 12640
rect 34698 12628 34704 12640
rect 34659 12600 34704 12628
rect 34698 12588 34704 12600
rect 34756 12588 34762 12640
rect 36173 12631 36231 12637
rect 36173 12597 36185 12631
rect 36219 12628 36231 12631
rect 36538 12628 36544 12640
rect 36219 12600 36544 12628
rect 36219 12597 36231 12600
rect 36173 12591 36231 12597
rect 36538 12588 36544 12600
rect 36596 12588 36602 12640
rect 38749 12631 38807 12637
rect 38749 12597 38761 12631
rect 38795 12628 38807 12631
rect 39040 12628 39068 12659
rect 41690 12628 41696 12640
rect 38795 12600 41696 12628
rect 38795 12597 38807 12600
rect 38749 12591 38807 12597
rect 41690 12588 41696 12600
rect 41748 12588 41754 12640
rect 1104 12538 48852 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 48852 12538
rect 1104 12464 48852 12486
rect 9030 12384 9036 12436
rect 9088 12424 9094 12436
rect 11149 12427 11207 12433
rect 11149 12424 11161 12427
rect 9088 12396 11161 12424
rect 9088 12384 9094 12396
rect 11149 12393 11161 12396
rect 11195 12393 11207 12427
rect 11149 12387 11207 12393
rect 13817 12427 13875 12433
rect 13817 12393 13829 12427
rect 13863 12424 13875 12427
rect 13906 12424 13912 12436
rect 13863 12396 13912 12424
rect 13863 12393 13875 12396
rect 13817 12387 13875 12393
rect 13906 12384 13912 12396
rect 13964 12384 13970 12436
rect 14182 12384 14188 12436
rect 14240 12424 14246 12436
rect 14921 12427 14979 12433
rect 14921 12424 14933 12427
rect 14240 12396 14933 12424
rect 14240 12384 14246 12396
rect 14921 12393 14933 12396
rect 14967 12424 14979 12427
rect 15378 12424 15384 12436
rect 14967 12396 15384 12424
rect 14967 12393 14979 12396
rect 14921 12387 14979 12393
rect 15378 12384 15384 12396
rect 15436 12384 15442 12436
rect 17218 12384 17224 12436
rect 17276 12424 17282 12436
rect 18693 12427 18751 12433
rect 18693 12424 18705 12427
rect 17276 12396 18705 12424
rect 17276 12384 17282 12396
rect 18693 12393 18705 12396
rect 18739 12393 18751 12427
rect 18693 12387 18751 12393
rect 19935 12427 19993 12433
rect 19935 12393 19947 12427
rect 19981 12424 19993 12427
rect 22002 12424 22008 12436
rect 19981 12396 22008 12424
rect 19981 12393 19993 12396
rect 19935 12387 19993 12393
rect 22002 12384 22008 12396
rect 22060 12384 22066 12436
rect 22189 12427 22247 12433
rect 22189 12393 22201 12427
rect 22235 12424 22247 12427
rect 22554 12424 22560 12436
rect 22235 12396 22560 12424
rect 22235 12393 22247 12396
rect 22189 12387 22247 12393
rect 22554 12384 22560 12396
rect 22612 12384 22618 12436
rect 23382 12424 23388 12436
rect 23343 12396 23388 12424
rect 23382 12384 23388 12396
rect 23440 12384 23446 12436
rect 23934 12424 23940 12436
rect 23895 12396 23940 12424
rect 23934 12384 23940 12396
rect 23992 12384 23998 12436
rect 25130 12424 25136 12436
rect 25091 12396 25136 12424
rect 25130 12384 25136 12396
rect 25188 12384 25194 12436
rect 31202 12424 31208 12436
rect 31163 12396 31208 12424
rect 31202 12384 31208 12396
rect 31260 12384 31266 12436
rect 35161 12427 35219 12433
rect 35161 12393 35173 12427
rect 35207 12424 35219 12427
rect 35342 12424 35348 12436
rect 35207 12396 35348 12424
rect 35207 12393 35219 12396
rect 35161 12387 35219 12393
rect 35342 12384 35348 12396
rect 35400 12384 35406 12436
rect 37918 12424 37924 12436
rect 37879 12396 37924 12424
rect 37918 12384 37924 12396
rect 37976 12384 37982 12436
rect 38930 12424 38936 12436
rect 38891 12396 38936 12424
rect 38930 12384 38936 12396
rect 38988 12384 38994 12436
rect 39390 12424 39396 12436
rect 39351 12396 39396 12424
rect 39390 12384 39396 12396
rect 39448 12384 39454 12436
rect 39942 12424 39948 12436
rect 39903 12396 39948 12424
rect 39942 12384 39948 12396
rect 40000 12384 40006 12436
rect 41690 12424 41696 12436
rect 41651 12396 41696 12424
rect 41690 12384 41696 12396
rect 41748 12384 41754 12436
rect 9950 12356 9956 12368
rect 9863 12328 9956 12356
rect 9950 12316 9956 12328
rect 10008 12356 10014 12368
rect 10318 12356 10324 12368
rect 10008 12328 10324 12356
rect 10008 12316 10014 12328
rect 10318 12316 10324 12328
rect 10376 12316 10382 12368
rect 10502 12356 10508 12368
rect 10463 12328 10508 12356
rect 10502 12316 10508 12328
rect 10560 12316 10566 12368
rect 12891 12359 12949 12365
rect 12891 12325 12903 12359
rect 12937 12356 12949 12359
rect 13630 12356 13636 12368
rect 12937 12328 13636 12356
rect 12937 12325 12949 12328
rect 12891 12319 12949 12325
rect 13630 12316 13636 12328
rect 13688 12316 13694 12368
rect 16206 12316 16212 12368
rect 16264 12356 16270 12368
rect 16387 12359 16445 12365
rect 16387 12356 16399 12359
rect 16264 12328 16399 12356
rect 16264 12316 16270 12328
rect 16387 12325 16399 12328
rect 16433 12356 16445 12359
rect 18135 12359 18193 12365
rect 18135 12356 18147 12359
rect 16433 12328 18147 12356
rect 16433 12325 16445 12328
rect 16387 12319 16445 12325
rect 18135 12325 18147 12328
rect 18181 12356 18193 12359
rect 18322 12356 18328 12368
rect 18181 12328 18328 12356
rect 18181 12325 18193 12328
rect 18135 12319 18193 12325
rect 18322 12316 18328 12328
rect 18380 12316 18386 12368
rect 21266 12316 21272 12368
rect 21324 12356 21330 12368
rect 21590 12359 21648 12365
rect 21590 12356 21602 12359
rect 21324 12328 21602 12356
rect 21324 12316 21330 12328
rect 21590 12325 21602 12328
rect 21636 12325 21648 12359
rect 21590 12319 21648 12325
rect 27893 12359 27951 12365
rect 27893 12325 27905 12359
rect 27939 12356 27951 12359
rect 28258 12356 28264 12368
rect 27939 12328 28264 12356
rect 27939 12325 27951 12328
rect 27893 12319 27951 12325
rect 28258 12316 28264 12328
rect 28316 12316 28322 12368
rect 29457 12359 29515 12365
rect 29457 12325 29469 12359
rect 29503 12356 29515 12359
rect 30466 12356 30472 12368
rect 29503 12328 30472 12356
rect 29503 12325 29515 12328
rect 29457 12319 29515 12325
rect 30466 12316 30472 12328
rect 30524 12316 30530 12368
rect 30647 12359 30705 12365
rect 30647 12325 30659 12359
rect 30693 12356 30705 12359
rect 30926 12356 30932 12368
rect 30693 12328 30932 12356
rect 30693 12325 30705 12328
rect 30647 12319 30705 12325
rect 30926 12316 30932 12328
rect 30984 12316 30990 12368
rect 32582 12316 32588 12368
rect 32640 12356 32646 12368
rect 33045 12359 33103 12365
rect 33045 12356 33057 12359
rect 32640 12328 33057 12356
rect 32640 12316 32646 12328
rect 33045 12325 33057 12328
rect 33091 12356 33103 12359
rect 33778 12356 33784 12368
rect 33091 12328 33784 12356
rect 33091 12325 33103 12328
rect 33045 12319 33103 12325
rect 33778 12316 33784 12328
rect 33836 12356 33842 12368
rect 34057 12359 34115 12365
rect 34057 12356 34069 12359
rect 33836 12328 34069 12356
rect 33836 12316 33842 12328
rect 34057 12325 34069 12328
rect 34103 12325 34115 12359
rect 34057 12319 34115 12325
rect 40862 12316 40868 12368
rect 40920 12356 40926 12368
rect 41135 12359 41193 12365
rect 41135 12356 41147 12359
rect 40920 12328 41147 12356
rect 40920 12316 40926 12328
rect 41135 12325 41147 12328
rect 41181 12356 41193 12359
rect 41598 12356 41604 12368
rect 41181 12328 41604 12356
rect 41181 12325 41193 12328
rect 41135 12319 41193 12325
rect 41598 12316 41604 12328
rect 41656 12316 41662 12368
rect 10226 12288 10232 12300
rect 10187 12260 10232 12288
rect 10226 12248 10232 12260
rect 10284 12248 10290 12300
rect 13449 12291 13507 12297
rect 13449 12257 13461 12291
rect 13495 12288 13507 12291
rect 15194 12288 15200 12300
rect 13495 12260 15200 12288
rect 13495 12257 13507 12260
rect 13449 12251 13507 12257
rect 15194 12248 15200 12260
rect 15252 12288 15258 12300
rect 15473 12291 15531 12297
rect 15473 12288 15485 12291
rect 15252 12260 15485 12288
rect 15252 12248 15258 12260
rect 15473 12257 15485 12260
rect 15519 12257 15531 12291
rect 15473 12251 15531 12257
rect 19864 12291 19922 12297
rect 19864 12257 19876 12291
rect 19910 12288 19922 12291
rect 20070 12288 20076 12300
rect 19910 12260 20076 12288
rect 19910 12257 19922 12260
rect 19864 12251 19922 12257
rect 20070 12248 20076 12260
rect 20128 12248 20134 12300
rect 24854 12288 24860 12300
rect 24815 12260 24860 12288
rect 24854 12248 24860 12260
rect 24912 12248 24918 12300
rect 25222 12248 25228 12300
rect 25280 12288 25286 12300
rect 25317 12291 25375 12297
rect 25317 12288 25329 12291
rect 25280 12260 25329 12288
rect 25280 12248 25286 12260
rect 25317 12257 25329 12260
rect 25363 12257 25375 12291
rect 25317 12251 25375 12257
rect 26786 12248 26792 12300
rect 26844 12288 26850 12300
rect 27157 12291 27215 12297
rect 27157 12288 27169 12291
rect 26844 12260 27169 12288
rect 26844 12248 26850 12260
rect 27157 12257 27169 12260
rect 27203 12288 27215 12291
rect 27430 12288 27436 12300
rect 27203 12260 27436 12288
rect 27203 12257 27215 12260
rect 27157 12251 27215 12257
rect 27430 12248 27436 12260
rect 27488 12248 27494 12300
rect 27706 12288 27712 12300
rect 27667 12260 27712 12288
rect 27706 12248 27712 12260
rect 27764 12248 27770 12300
rect 28718 12288 28724 12300
rect 28679 12260 28724 12288
rect 28718 12248 28724 12260
rect 28776 12248 28782 12300
rect 29273 12291 29331 12297
rect 29273 12257 29285 12291
rect 29319 12288 29331 12291
rect 32398 12288 32404 12300
rect 29319 12260 29960 12288
rect 32359 12260 32404 12288
rect 29319 12257 29331 12260
rect 29273 12251 29331 12257
rect 12526 12220 12532 12232
rect 12487 12192 12532 12220
rect 12526 12180 12532 12192
rect 12584 12180 12590 12232
rect 16022 12220 16028 12232
rect 15983 12192 16028 12220
rect 16022 12180 16028 12192
rect 16080 12180 16086 12232
rect 17770 12220 17776 12232
rect 17731 12192 17776 12220
rect 17770 12180 17776 12192
rect 17828 12180 17834 12232
rect 20717 12223 20775 12229
rect 20717 12189 20729 12223
rect 20763 12220 20775 12223
rect 20990 12220 20996 12232
rect 20763 12192 20996 12220
rect 20763 12189 20775 12192
rect 20717 12183 20775 12189
rect 20990 12180 20996 12192
rect 21048 12220 21054 12232
rect 21269 12223 21327 12229
rect 21269 12220 21281 12223
rect 21048 12192 21281 12220
rect 21048 12180 21054 12192
rect 21269 12189 21281 12192
rect 21315 12189 21327 12223
rect 21269 12183 21327 12189
rect 22738 12180 22744 12232
rect 22796 12220 22802 12232
rect 23017 12223 23075 12229
rect 23017 12220 23029 12223
rect 22796 12192 23029 12220
rect 22796 12180 22802 12192
rect 23017 12189 23029 12192
rect 23063 12189 23075 12223
rect 23017 12183 23075 12189
rect 13998 12112 14004 12164
rect 14056 12152 14062 12164
rect 18690 12152 18696 12164
rect 14056 12124 18696 12152
rect 14056 12112 14062 12124
rect 18690 12112 18696 12124
rect 18748 12152 18754 12164
rect 18969 12155 19027 12161
rect 18969 12152 18981 12155
rect 18748 12124 18981 12152
rect 18748 12112 18754 12124
rect 18969 12121 18981 12124
rect 19015 12121 19027 12155
rect 18969 12115 19027 12121
rect 16942 12084 16948 12096
rect 16903 12056 16948 12084
rect 16942 12044 16948 12056
rect 17000 12044 17006 12096
rect 17218 12044 17224 12096
rect 17276 12084 17282 12096
rect 20806 12084 20812 12096
rect 17276 12056 20812 12084
rect 17276 12044 17282 12056
rect 20806 12044 20812 12056
rect 20864 12044 20870 12096
rect 21082 12084 21088 12096
rect 21043 12056 21088 12084
rect 21082 12044 21088 12056
rect 21140 12044 21146 12096
rect 24210 12084 24216 12096
rect 24171 12056 24216 12084
rect 24210 12044 24216 12056
rect 24268 12044 24274 12096
rect 26510 12044 26516 12096
rect 26568 12084 26574 12096
rect 29932 12093 29960 12260
rect 32398 12248 32404 12260
rect 32456 12288 32462 12300
rect 33318 12288 33324 12300
rect 32456 12260 33324 12288
rect 32456 12248 32462 12260
rect 33318 12248 33324 12260
rect 33376 12248 33382 12300
rect 34790 12248 34796 12300
rect 34848 12288 34854 12300
rect 35472 12291 35530 12297
rect 35472 12288 35484 12291
rect 34848 12260 35484 12288
rect 34848 12248 34854 12260
rect 35472 12257 35484 12260
rect 35518 12288 35530 12291
rect 36170 12288 36176 12300
rect 35518 12260 36176 12288
rect 35518 12257 35530 12260
rect 35472 12251 35530 12257
rect 36170 12248 36176 12260
rect 36228 12288 36234 12300
rect 36449 12291 36507 12297
rect 36449 12288 36461 12291
rect 36228 12260 36461 12288
rect 36228 12248 36234 12260
rect 36449 12257 36461 12260
rect 36495 12257 36507 12291
rect 36449 12251 36507 12257
rect 30285 12223 30343 12229
rect 30285 12189 30297 12223
rect 30331 12220 30343 12223
rect 30558 12220 30564 12232
rect 30331 12192 30564 12220
rect 30331 12189 30343 12192
rect 30285 12183 30343 12189
rect 30558 12180 30564 12192
rect 30616 12180 30622 12232
rect 33962 12220 33968 12232
rect 33923 12192 33968 12220
rect 33962 12180 33968 12192
rect 34020 12180 34026 12232
rect 34238 12220 34244 12232
rect 34199 12192 34244 12220
rect 34238 12180 34244 12192
rect 34296 12180 34302 12232
rect 35618 12180 35624 12232
rect 35676 12220 35682 12232
rect 38473 12223 38531 12229
rect 38473 12220 38485 12223
rect 35676 12192 38485 12220
rect 35676 12180 35682 12192
rect 38473 12189 38485 12192
rect 38519 12220 38531 12223
rect 38838 12220 38844 12232
rect 38519 12192 38844 12220
rect 38519 12189 38531 12192
rect 38473 12183 38531 12189
rect 38838 12180 38844 12192
rect 38896 12180 38902 12232
rect 39022 12220 39028 12232
rect 38983 12192 39028 12220
rect 39022 12180 39028 12192
rect 39080 12180 39086 12232
rect 40773 12223 40831 12229
rect 40773 12189 40785 12223
rect 40819 12220 40831 12223
rect 41138 12220 41144 12232
rect 40819 12192 41144 12220
rect 40819 12189 40831 12192
rect 40773 12183 40831 12189
rect 41138 12180 41144 12192
rect 41196 12180 41202 12232
rect 26697 12087 26755 12093
rect 26697 12084 26709 12087
rect 26568 12056 26709 12084
rect 26568 12044 26574 12056
rect 26697 12053 26709 12056
rect 26743 12053 26755 12087
rect 26697 12047 26755 12053
rect 29917 12087 29975 12093
rect 29917 12053 29929 12087
rect 29963 12084 29975 12087
rect 30282 12084 30288 12096
rect 29963 12056 30288 12084
rect 29963 12053 29975 12056
rect 29917 12047 29975 12053
rect 30282 12044 30288 12056
rect 30340 12044 30346 12096
rect 35250 12044 35256 12096
rect 35308 12084 35314 12096
rect 35575 12087 35633 12093
rect 35575 12084 35587 12087
rect 35308 12056 35587 12084
rect 35308 12044 35314 12056
rect 35575 12053 35587 12056
rect 35621 12053 35633 12087
rect 36630 12084 36636 12096
rect 36591 12056 36636 12084
rect 35575 12047 35633 12053
rect 36630 12044 36636 12056
rect 36688 12044 36694 12096
rect 36906 12084 36912 12096
rect 36867 12056 36912 12084
rect 36906 12044 36912 12056
rect 36964 12044 36970 12096
rect 1104 11994 48852 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 48852 11994
rect 1104 11920 48852 11942
rect 9493 11883 9551 11889
rect 9493 11849 9505 11883
rect 9539 11880 9551 11883
rect 10226 11880 10232 11892
rect 9539 11852 10232 11880
rect 9539 11849 9551 11852
rect 9493 11843 9551 11849
rect 10226 11840 10232 11852
rect 10284 11840 10290 11892
rect 15838 11880 15844 11892
rect 15799 11852 15844 11880
rect 15838 11840 15844 11852
rect 15896 11840 15902 11892
rect 16022 11840 16028 11892
rect 16080 11880 16086 11892
rect 16485 11883 16543 11889
rect 16485 11880 16497 11883
rect 16080 11852 16497 11880
rect 16080 11840 16086 11852
rect 16485 11849 16497 11852
rect 16531 11849 16543 11883
rect 16485 11843 16543 11849
rect 16942 11840 16948 11892
rect 17000 11880 17006 11892
rect 17129 11883 17187 11889
rect 17129 11880 17141 11883
rect 17000 11852 17141 11880
rect 17000 11840 17006 11852
rect 17129 11849 17141 11852
rect 17175 11849 17187 11883
rect 17129 11843 17187 11849
rect 17865 11883 17923 11889
rect 17865 11849 17877 11883
rect 17911 11880 17923 11883
rect 18322 11880 18328 11892
rect 17911 11852 18328 11880
rect 17911 11849 17923 11852
rect 17865 11843 17923 11849
rect 18322 11840 18328 11852
rect 18380 11840 18386 11892
rect 19889 11883 19947 11889
rect 19889 11849 19901 11883
rect 19935 11880 19947 11883
rect 20070 11880 20076 11892
rect 19935 11852 20076 11880
rect 19935 11849 19947 11852
rect 19889 11843 19947 11849
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 21266 11840 21272 11892
rect 21324 11880 21330 11892
rect 21453 11883 21511 11889
rect 21453 11880 21465 11883
rect 21324 11852 21465 11880
rect 21324 11840 21330 11852
rect 21453 11849 21465 11852
rect 21499 11849 21511 11883
rect 21453 11843 21511 11849
rect 8662 11772 8668 11824
rect 8720 11812 8726 11824
rect 11241 11815 11299 11821
rect 11241 11812 11253 11815
rect 8720 11784 11253 11812
rect 8720 11772 8726 11784
rect 11241 11781 11253 11784
rect 11287 11781 11299 11815
rect 11241 11775 11299 11781
rect 12253 11815 12311 11821
rect 12253 11781 12265 11815
rect 12299 11812 12311 11815
rect 13630 11812 13636 11824
rect 12299 11784 13636 11812
rect 12299 11781 12311 11784
rect 12253 11775 12311 11781
rect 12268 11744 12296 11775
rect 13630 11772 13636 11784
rect 13688 11812 13694 11824
rect 14829 11815 14887 11821
rect 14829 11812 14841 11815
rect 13688 11784 14841 11812
rect 13688 11772 13694 11784
rect 14829 11781 14841 11784
rect 14875 11812 14887 11815
rect 16206 11812 16212 11824
rect 14875 11784 16212 11812
rect 14875 11781 14887 11784
rect 14829 11775 14887 11781
rect 11808 11716 12296 11744
rect 10318 11676 10324 11688
rect 10279 11648 10324 11676
rect 10318 11636 10324 11648
rect 10376 11636 10382 11688
rect 9861 11611 9919 11617
rect 9861 11577 9873 11611
rect 9907 11608 9919 11611
rect 10229 11611 10287 11617
rect 10229 11608 10241 11611
rect 9907 11580 10241 11608
rect 9907 11577 9919 11580
rect 9861 11571 9919 11577
rect 10229 11577 10241 11580
rect 10275 11608 10287 11611
rect 10502 11608 10508 11620
rect 10275 11580 10508 11608
rect 10275 11577 10287 11580
rect 10229 11571 10287 11577
rect 10502 11568 10508 11580
rect 10560 11608 10566 11620
rect 10683 11611 10741 11617
rect 10683 11608 10695 11611
rect 10560 11580 10695 11608
rect 10560 11568 10566 11580
rect 10683 11577 10695 11580
rect 10729 11608 10741 11611
rect 11808 11608 11836 11716
rect 12526 11704 12532 11756
rect 12584 11744 12590 11756
rect 13173 11747 13231 11753
rect 13173 11744 13185 11747
rect 12584 11716 13185 11744
rect 12584 11704 12590 11716
rect 13173 11713 13185 11716
rect 13219 11744 13231 11747
rect 13817 11747 13875 11753
rect 13817 11744 13829 11747
rect 13219 11716 13829 11744
rect 13219 11713 13231 11716
rect 13173 11707 13231 11713
rect 13817 11713 13829 11716
rect 13863 11713 13875 11747
rect 13817 11707 13875 11713
rect 14921 11747 14979 11753
rect 14921 11713 14933 11747
rect 14967 11744 14979 11747
rect 15010 11744 15016 11756
rect 14967 11716 15016 11744
rect 14967 11713 14979 11716
rect 14921 11707 14979 11713
rect 15010 11704 15016 11716
rect 15068 11704 15074 11756
rect 11885 11679 11943 11685
rect 11885 11645 11897 11679
rect 11931 11676 11943 11679
rect 12710 11676 12716 11688
rect 11931 11648 12716 11676
rect 11931 11645 11943 11648
rect 11885 11639 11943 11645
rect 12710 11636 12716 11648
rect 12768 11636 12774 11688
rect 12802 11636 12808 11688
rect 12860 11676 12866 11688
rect 12897 11679 12955 11685
rect 12897 11676 12909 11679
rect 12860 11648 12909 11676
rect 12860 11636 12866 11648
rect 12897 11645 12909 11648
rect 12943 11676 12955 11679
rect 13449 11679 13507 11685
rect 13449 11676 13461 11679
rect 12943 11648 13461 11676
rect 12943 11645 12955 11648
rect 12897 11639 12955 11645
rect 13449 11645 13461 11648
rect 13495 11645 13507 11679
rect 13449 11639 13507 11645
rect 15257 11617 15285 11784
rect 16206 11772 16212 11784
rect 16264 11772 16270 11824
rect 16390 11772 16396 11824
rect 16448 11812 16454 11824
rect 16807 11815 16865 11821
rect 16807 11812 16819 11815
rect 16448 11784 16819 11812
rect 16448 11772 16454 11784
rect 16807 11781 16819 11784
rect 16853 11781 16865 11815
rect 21082 11812 21088 11824
rect 16807 11775 16865 11781
rect 18892 11784 21088 11812
rect 16736 11679 16794 11685
rect 16736 11645 16748 11679
rect 16782 11676 16794 11679
rect 16942 11676 16948 11688
rect 16782 11648 16948 11676
rect 16782 11645 16794 11648
rect 16736 11639 16794 11645
rect 16942 11636 16948 11648
rect 17000 11636 17006 11688
rect 18892 11685 18920 11784
rect 21082 11772 21088 11784
rect 21140 11772 21146 11824
rect 21468 11812 21496 11843
rect 22922 11840 22928 11892
rect 22980 11880 22986 11892
rect 24581 11883 24639 11889
rect 24581 11880 24593 11883
rect 22980 11852 24593 11880
rect 22980 11840 22986 11852
rect 24581 11849 24593 11852
rect 24627 11849 24639 11883
rect 30926 11880 30932 11892
rect 30887 11852 30932 11880
rect 24581 11843 24639 11849
rect 30926 11840 30932 11852
rect 30984 11840 30990 11892
rect 31481 11883 31539 11889
rect 31481 11849 31493 11883
rect 31527 11880 31539 11883
rect 31938 11880 31944 11892
rect 31527 11852 31944 11880
rect 31527 11849 31539 11852
rect 31481 11843 31539 11849
rect 22554 11812 22560 11824
rect 21468 11784 22560 11812
rect 22554 11772 22560 11784
rect 22612 11812 22618 11824
rect 23017 11815 23075 11821
rect 23017 11812 23029 11815
rect 22612 11784 23029 11812
rect 22612 11772 22618 11784
rect 23017 11781 23029 11784
rect 23063 11812 23075 11815
rect 23293 11815 23351 11821
rect 23293 11812 23305 11815
rect 23063 11784 23305 11812
rect 23063 11781 23075 11784
rect 23017 11775 23075 11781
rect 23293 11781 23305 11784
rect 23339 11812 23351 11815
rect 23382 11812 23388 11824
rect 23339 11784 23388 11812
rect 23339 11781 23351 11784
rect 23293 11775 23351 11781
rect 23382 11772 23388 11784
rect 23440 11772 23446 11824
rect 20990 11744 20996 11756
rect 20951 11716 20996 11744
rect 20990 11704 20996 11716
rect 21048 11704 21054 11756
rect 21913 11747 21971 11753
rect 21913 11713 21925 11747
rect 21959 11744 21971 11747
rect 21959 11716 23060 11744
rect 21959 11713 21971 11716
rect 21913 11707 21971 11713
rect 18509 11679 18567 11685
rect 18509 11645 18521 11679
rect 18555 11676 18567 11679
rect 18877 11679 18935 11685
rect 18877 11676 18889 11679
rect 18555 11648 18889 11676
rect 18555 11645 18567 11648
rect 18509 11639 18567 11645
rect 18877 11645 18889 11648
rect 18923 11645 18935 11679
rect 18877 11639 18935 11645
rect 18966 11636 18972 11688
rect 19024 11676 19030 11688
rect 19061 11679 19119 11685
rect 19061 11676 19073 11679
rect 19024 11648 19073 11676
rect 19024 11636 19030 11648
rect 19061 11645 19073 11648
rect 19107 11645 19119 11679
rect 19061 11639 19119 11645
rect 20349 11679 20407 11685
rect 20349 11645 20361 11679
rect 20395 11676 20407 11679
rect 20438 11676 20444 11688
rect 20395 11648 20444 11676
rect 20395 11645 20407 11648
rect 20349 11639 20407 11645
rect 20438 11636 20444 11648
rect 20496 11676 20502 11688
rect 20717 11679 20775 11685
rect 20717 11676 20729 11679
rect 20496 11648 20729 11676
rect 20496 11636 20502 11648
rect 20717 11645 20729 11648
rect 20763 11645 20775 11679
rect 20717 11639 20775 11645
rect 10729 11580 11836 11608
rect 15242 11611 15300 11617
rect 10729 11577 10741 11580
rect 10683 11571 10741 11577
rect 15242 11577 15254 11611
rect 15288 11577 15300 11611
rect 20732 11608 20760 11639
rect 20806 11636 20812 11688
rect 20864 11676 20870 11688
rect 20901 11679 20959 11685
rect 20901 11676 20913 11679
rect 20864 11648 20913 11676
rect 20864 11636 20870 11648
rect 20901 11645 20913 11648
rect 20947 11645 20959 11679
rect 20901 11639 20959 11645
rect 21928 11608 21956 11707
rect 22296 11685 22324 11716
rect 23032 11688 23060 11716
rect 23566 11704 23572 11756
rect 23624 11744 23630 11756
rect 23661 11747 23719 11753
rect 23661 11744 23673 11747
rect 23624 11716 23673 11744
rect 23624 11704 23630 11716
rect 23661 11713 23673 11716
rect 23707 11744 23719 11747
rect 24210 11744 24216 11756
rect 23707 11716 24216 11744
rect 23707 11713 23719 11716
rect 23661 11707 23719 11713
rect 24210 11704 24216 11716
rect 24268 11704 24274 11756
rect 26510 11744 26516 11756
rect 26471 11716 26516 11744
rect 26510 11704 26516 11716
rect 26568 11704 26574 11756
rect 27433 11747 27491 11753
rect 27433 11713 27445 11747
rect 27479 11744 27491 11747
rect 28350 11744 28356 11756
rect 27479 11716 28356 11744
rect 27479 11713 27491 11716
rect 27433 11707 27491 11713
rect 28350 11704 28356 11716
rect 28408 11704 28414 11756
rect 22281 11679 22339 11685
rect 22281 11645 22293 11679
rect 22327 11645 22339 11679
rect 22462 11676 22468 11688
rect 22423 11648 22468 11676
rect 22281 11639 22339 11645
rect 22462 11636 22468 11648
rect 22520 11636 22526 11688
rect 23014 11636 23020 11688
rect 23072 11676 23078 11688
rect 24854 11676 24860 11688
rect 23072 11648 24860 11676
rect 23072 11636 23078 11648
rect 24854 11636 24860 11648
rect 24912 11676 24918 11688
rect 25593 11679 25651 11685
rect 25593 11676 25605 11679
rect 24912 11648 25605 11676
rect 24912 11636 24918 11648
rect 25593 11645 25605 11648
rect 25639 11676 25651 11679
rect 25777 11679 25835 11685
rect 25777 11676 25789 11679
rect 25639 11648 25789 11676
rect 25639 11645 25651 11648
rect 25593 11639 25651 11645
rect 25777 11645 25789 11648
rect 25823 11645 25835 11679
rect 25777 11639 25835 11645
rect 22738 11608 22744 11620
rect 20732 11580 21956 11608
rect 22699 11580 22744 11608
rect 15242 11571 15300 11577
rect 22738 11568 22744 11580
rect 22796 11568 22802 11620
rect 23293 11611 23351 11617
rect 23293 11577 23305 11611
rect 23339 11608 23351 11611
rect 24023 11611 24081 11617
rect 24023 11608 24035 11611
rect 23339 11580 24035 11608
rect 23339 11577 23351 11580
rect 23293 11571 23351 11577
rect 24023 11577 24035 11580
rect 24069 11608 24081 11611
rect 24670 11608 24676 11620
rect 24069 11580 24676 11608
rect 24069 11577 24081 11580
rect 24023 11571 24081 11577
rect 24670 11568 24676 11580
rect 24728 11568 24734 11620
rect 25792 11608 25820 11639
rect 25866 11636 25872 11688
rect 25924 11676 25930 11688
rect 26237 11679 26295 11685
rect 26237 11676 26249 11679
rect 25924 11648 26249 11676
rect 25924 11636 25930 11648
rect 26237 11645 26249 11648
rect 26283 11645 26295 11679
rect 26237 11639 26295 11645
rect 30101 11679 30159 11685
rect 30101 11645 30113 11679
rect 30147 11645 30159 11679
rect 30282 11676 30288 11688
rect 30243 11648 30288 11676
rect 30101 11639 30159 11645
rect 26786 11608 26792 11620
rect 25792 11580 26792 11608
rect 26786 11568 26792 11580
rect 26844 11568 26850 11620
rect 27249 11611 27307 11617
rect 27249 11577 27261 11611
rect 27295 11608 27307 11611
rect 27522 11608 27528 11620
rect 27295 11580 27528 11608
rect 27295 11577 27307 11580
rect 27249 11571 27307 11577
rect 27522 11568 27528 11580
rect 27580 11568 27586 11620
rect 27890 11568 27896 11620
rect 27948 11608 27954 11620
rect 28077 11611 28135 11617
rect 28077 11608 28089 11611
rect 27948 11580 28089 11608
rect 27948 11568 27954 11580
rect 28077 11577 28089 11580
rect 28123 11577 28135 11611
rect 28077 11571 28135 11577
rect 28258 11568 28264 11620
rect 28316 11608 28322 11620
rect 29733 11611 29791 11617
rect 29733 11608 29745 11611
rect 28316 11580 29745 11608
rect 28316 11568 28322 11580
rect 29733 11577 29745 11580
rect 29779 11608 29791 11611
rect 30116 11608 30144 11639
rect 30282 11636 30288 11648
rect 30340 11636 30346 11688
rect 31655 11685 31683 11852
rect 31938 11840 31944 11852
rect 31996 11840 32002 11892
rect 32125 11883 32183 11889
rect 32125 11849 32137 11883
rect 32171 11880 32183 11883
rect 32398 11880 32404 11892
rect 32171 11852 32404 11880
rect 32171 11849 32183 11852
rect 32125 11843 32183 11849
rect 32398 11840 32404 11852
rect 32456 11840 32462 11892
rect 33962 11880 33968 11892
rect 33106 11852 33968 11880
rect 31711 11815 31769 11821
rect 31711 11781 31723 11815
rect 31757 11812 31769 11815
rect 33106 11812 33134 11852
rect 33962 11840 33968 11852
rect 34020 11880 34026 11892
rect 34241 11883 34299 11889
rect 34241 11880 34253 11883
rect 34020 11852 34253 11880
rect 34020 11840 34026 11852
rect 34241 11849 34253 11852
rect 34287 11849 34299 11883
rect 36170 11880 36176 11892
rect 36131 11852 36176 11880
rect 34241 11843 34299 11849
rect 36170 11840 36176 11852
rect 36228 11840 36234 11892
rect 38286 11880 38292 11892
rect 38247 11852 38292 11880
rect 38286 11840 38292 11852
rect 38344 11840 38350 11892
rect 39390 11840 39396 11892
rect 39448 11880 39454 11892
rect 39577 11883 39635 11889
rect 39577 11880 39589 11883
rect 39448 11852 39589 11880
rect 39448 11840 39454 11852
rect 39577 11849 39589 11852
rect 39623 11880 39635 11883
rect 40862 11880 40868 11892
rect 39623 11852 40868 11880
rect 39623 11849 39635 11852
rect 39577 11843 39635 11849
rect 40862 11840 40868 11852
rect 40920 11840 40926 11892
rect 31757 11784 33134 11812
rect 31757 11781 31769 11784
rect 31711 11775 31769 11781
rect 33778 11772 33784 11824
rect 33836 11812 33842 11824
rect 33873 11815 33931 11821
rect 33873 11812 33885 11815
rect 33836 11784 33885 11812
rect 33836 11772 33842 11784
rect 33873 11781 33885 11784
rect 33919 11781 33931 11815
rect 33873 11775 33931 11781
rect 32674 11744 32680 11756
rect 32635 11716 32680 11744
rect 32674 11704 32680 11716
rect 32732 11704 32738 11756
rect 33321 11747 33379 11753
rect 33321 11713 33333 11747
rect 33367 11744 33379 11747
rect 34238 11744 34244 11756
rect 33367 11716 34244 11744
rect 33367 11713 33379 11716
rect 33321 11707 33379 11713
rect 34238 11704 34244 11716
rect 34296 11704 34302 11756
rect 36725 11747 36783 11753
rect 36725 11713 36737 11747
rect 36771 11744 36783 11747
rect 36906 11744 36912 11756
rect 36771 11716 36912 11744
rect 36771 11713 36783 11716
rect 36725 11707 36783 11713
rect 36906 11704 36912 11716
rect 36964 11704 36970 11756
rect 39022 11704 39028 11756
rect 39080 11744 39086 11756
rect 39209 11747 39267 11753
rect 39209 11744 39221 11747
rect 39080 11716 39221 11744
rect 39080 11704 39086 11716
rect 39209 11713 39221 11716
rect 39255 11744 39267 11747
rect 39853 11747 39911 11753
rect 39853 11744 39865 11747
rect 39255 11716 39865 11744
rect 39255 11713 39267 11716
rect 39209 11707 39267 11713
rect 39853 11713 39865 11716
rect 39899 11713 39911 11747
rect 39853 11707 39911 11713
rect 31640 11679 31698 11685
rect 31640 11645 31652 11679
rect 31686 11645 31698 11679
rect 31640 11639 31698 11645
rect 34701 11679 34759 11685
rect 34701 11645 34713 11679
rect 34747 11676 34759 11679
rect 35529 11679 35587 11685
rect 35529 11676 35541 11679
rect 34747 11648 35541 11676
rect 34747 11645 34759 11648
rect 34701 11639 34759 11645
rect 35529 11645 35541 11648
rect 35575 11676 35587 11679
rect 36630 11676 36636 11688
rect 35575 11648 36636 11676
rect 35575 11645 35587 11648
rect 35529 11639 35587 11645
rect 36630 11636 36636 11648
rect 36688 11636 36694 11688
rect 38286 11636 38292 11688
rect 38344 11676 38350 11688
rect 38473 11679 38531 11685
rect 38473 11676 38485 11679
rect 38344 11648 38485 11676
rect 38344 11636 38350 11648
rect 38473 11645 38485 11648
rect 38519 11645 38531 11679
rect 38473 11639 38531 11645
rect 38838 11636 38844 11688
rect 38896 11676 38902 11688
rect 38933 11679 38991 11685
rect 38933 11676 38945 11679
rect 38896 11648 38945 11676
rect 38896 11636 38902 11648
rect 38933 11645 38945 11648
rect 38979 11645 38991 11679
rect 38933 11639 38991 11645
rect 30374 11608 30380 11620
rect 29779 11580 30380 11608
rect 29779 11577 29791 11580
rect 29733 11571 29791 11577
rect 30374 11568 30380 11580
rect 30432 11568 30438 11620
rect 30558 11608 30564 11620
rect 30519 11580 30564 11608
rect 30558 11568 30564 11580
rect 30616 11568 30622 11620
rect 32493 11611 32551 11617
rect 32493 11577 32505 11611
rect 32539 11608 32551 11611
rect 32766 11608 32772 11620
rect 32539 11580 32772 11608
rect 32539 11577 32551 11580
rect 32493 11571 32551 11577
rect 32766 11568 32772 11580
rect 32824 11568 32830 11620
rect 34330 11568 34336 11620
rect 34388 11608 34394 11620
rect 34885 11611 34943 11617
rect 34885 11608 34897 11611
rect 34388 11580 34897 11608
rect 34388 11568 34394 11580
rect 34885 11577 34897 11580
rect 34931 11577 34943 11611
rect 36538 11608 36544 11620
rect 36451 11580 36544 11608
rect 34885 11571 34943 11577
rect 36538 11568 36544 11580
rect 36596 11608 36602 11620
rect 37087 11611 37145 11617
rect 37087 11608 37099 11611
rect 36596 11580 37099 11608
rect 36596 11568 36602 11580
rect 37087 11577 37099 11580
rect 37133 11608 37145 11611
rect 39390 11608 39396 11620
rect 37133 11580 39396 11608
rect 37133 11577 37145 11580
rect 37087 11571 37145 11577
rect 39390 11568 39396 11580
rect 39448 11568 39454 11620
rect 18506 11500 18512 11552
rect 18564 11540 18570 11552
rect 18693 11543 18751 11549
rect 18693 11540 18705 11543
rect 18564 11512 18705 11540
rect 18564 11500 18570 11512
rect 18693 11509 18705 11512
rect 18739 11509 18751 11543
rect 25222 11540 25228 11552
rect 25183 11512 25228 11540
rect 18693 11503 18751 11509
rect 25222 11500 25228 11512
rect 25280 11500 25286 11552
rect 27982 11500 27988 11552
rect 28040 11540 28046 11552
rect 28353 11543 28411 11549
rect 28353 11540 28365 11543
rect 28040 11512 28365 11540
rect 28040 11500 28046 11512
rect 28353 11509 28365 11512
rect 28399 11509 28411 11543
rect 28718 11540 28724 11552
rect 28679 11512 28724 11540
rect 28353 11503 28411 11509
rect 28718 11500 28724 11512
rect 28776 11500 28782 11552
rect 37642 11540 37648 11552
rect 37603 11512 37648 11540
rect 37642 11500 37648 11512
rect 37700 11500 37706 11552
rect 41138 11540 41144 11552
rect 41099 11512 41144 11540
rect 41138 11500 41144 11512
rect 41196 11500 41202 11552
rect 1104 11450 48852 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 48852 11450
rect 1104 11376 48852 11398
rect 9950 11336 9956 11348
rect 9911 11308 9956 11336
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 10318 11336 10324 11348
rect 10279 11308 10324 11336
rect 10318 11296 10324 11308
rect 10376 11336 10382 11348
rect 11057 11339 11115 11345
rect 11057 11336 11069 11339
rect 10376 11308 11069 11336
rect 10376 11296 10382 11308
rect 11057 11305 11069 11308
rect 11103 11305 11115 11339
rect 11057 11299 11115 11305
rect 11790 11296 11796 11348
rect 11848 11336 11854 11348
rect 12434 11336 12440 11348
rect 11848 11308 12440 11336
rect 11848 11296 11854 11308
rect 12434 11296 12440 11308
rect 12492 11336 12498 11348
rect 13173 11339 13231 11345
rect 13173 11336 13185 11339
rect 12492 11308 13185 11336
rect 12492 11296 12498 11308
rect 13173 11305 13185 11308
rect 13219 11305 13231 11339
rect 15010 11336 15016 11348
rect 14971 11308 15016 11336
rect 13173 11299 13231 11305
rect 15010 11296 15016 11308
rect 15068 11296 15074 11348
rect 16022 11336 16028 11348
rect 15983 11308 16028 11336
rect 16022 11296 16028 11308
rect 16080 11296 16086 11348
rect 17770 11336 17776 11348
rect 17731 11308 17776 11336
rect 17770 11296 17776 11308
rect 17828 11336 17834 11348
rect 17957 11339 18015 11345
rect 17957 11336 17969 11339
rect 17828 11308 17969 11336
rect 17828 11296 17834 11308
rect 17957 11305 17969 11308
rect 18003 11305 18015 11339
rect 17957 11299 18015 11305
rect 18966 11296 18972 11348
rect 19024 11336 19030 11348
rect 19705 11339 19763 11345
rect 19705 11336 19717 11339
rect 19024 11308 19717 11336
rect 19024 11296 19030 11308
rect 19705 11305 19717 11308
rect 19751 11305 19763 11339
rect 19705 11299 19763 11305
rect 22738 11296 22744 11348
rect 22796 11336 22802 11348
rect 23845 11339 23903 11345
rect 23845 11336 23857 11339
rect 22796 11308 23857 11336
rect 22796 11296 22802 11308
rect 23845 11305 23857 11308
rect 23891 11305 23903 11339
rect 23845 11299 23903 11305
rect 24578 11296 24584 11348
rect 24636 11336 24642 11348
rect 24673 11339 24731 11345
rect 24673 11336 24685 11339
rect 24636 11308 24685 11336
rect 24636 11296 24642 11308
rect 24673 11305 24685 11308
rect 24719 11305 24731 11339
rect 26602 11336 26608 11348
rect 26563 11308 26608 11336
rect 24673 11299 24731 11305
rect 26602 11296 26608 11308
rect 26660 11296 26666 11348
rect 27617 11339 27675 11345
rect 27617 11305 27629 11339
rect 27663 11336 27675 11339
rect 27706 11336 27712 11348
rect 27663 11308 27712 11336
rect 27663 11305 27675 11308
rect 27617 11299 27675 11305
rect 27706 11296 27712 11308
rect 27764 11336 27770 11348
rect 28258 11336 28264 11348
rect 27764 11308 28264 11336
rect 27764 11296 27770 11308
rect 28258 11296 28264 11308
rect 28316 11296 28322 11348
rect 30558 11336 30564 11348
rect 30519 11308 30564 11336
rect 30558 11296 30564 11308
rect 30616 11296 30622 11348
rect 32674 11336 32680 11348
rect 32635 11308 32680 11336
rect 32674 11296 32680 11308
rect 32732 11296 32738 11348
rect 35621 11339 35679 11345
rect 35621 11305 35633 11339
rect 35667 11336 35679 11339
rect 36170 11336 36176 11348
rect 35667 11308 36176 11336
rect 35667 11305 35679 11308
rect 35621 11299 35679 11305
rect 36170 11296 36176 11308
rect 36228 11296 36234 11348
rect 40494 11336 40500 11348
rect 39592 11308 40500 11336
rect 9968 11268 9996 11296
rect 9968 11240 10548 11268
rect 10520 11209 10548 11240
rect 11882 11228 11888 11280
rect 11940 11268 11946 11280
rect 12345 11271 12403 11277
rect 12345 11268 12357 11271
rect 11940 11240 12357 11268
rect 11940 11228 11946 11240
rect 12345 11237 12357 11240
rect 12391 11268 12403 11271
rect 17678 11268 17684 11280
rect 12391 11240 17684 11268
rect 12391 11237 12403 11240
rect 12345 11231 12403 11237
rect 17678 11228 17684 11240
rect 17736 11228 17742 11280
rect 19334 11228 19340 11280
rect 19392 11268 19398 11280
rect 19429 11271 19487 11277
rect 19429 11268 19441 11271
rect 19392 11240 19441 11268
rect 19392 11228 19398 11240
rect 19429 11237 19441 11240
rect 19475 11268 19487 11271
rect 20346 11268 20352 11280
rect 19475 11240 20352 11268
rect 19475 11237 19487 11240
rect 19429 11231 19487 11237
rect 20346 11228 20352 11240
rect 20404 11228 20410 11280
rect 20714 11228 20720 11280
rect 20772 11268 20778 11280
rect 20901 11271 20959 11277
rect 20901 11268 20913 11271
rect 20772 11240 20913 11268
rect 20772 11228 20778 11240
rect 20901 11237 20913 11240
rect 20947 11237 20959 11271
rect 23566 11268 23572 11280
rect 23527 11240 23572 11268
rect 20901 11231 20959 11237
rect 23566 11228 23572 11240
rect 23624 11228 23630 11280
rect 24213 11271 24271 11277
rect 24213 11237 24225 11271
rect 24259 11268 24271 11271
rect 24259 11240 24900 11268
rect 24259 11237 24271 11240
rect 24213 11231 24271 11237
rect 10229 11203 10287 11209
rect 10229 11169 10241 11203
rect 10275 11169 10287 11203
rect 10229 11163 10287 11169
rect 10505 11203 10563 11209
rect 10505 11169 10517 11203
rect 10551 11169 10563 11203
rect 12526 11200 12532 11212
rect 12487 11172 12532 11200
rect 10505 11163 10563 11169
rect 10244 11132 10272 11163
rect 12526 11160 12532 11172
rect 12584 11160 12590 11212
rect 12894 11200 12900 11212
rect 12855 11172 12900 11200
rect 12894 11160 12900 11172
rect 12952 11160 12958 11212
rect 13722 11200 13728 11212
rect 13683 11172 13728 11200
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 13814 11160 13820 11212
rect 13872 11200 13878 11212
rect 13909 11203 13967 11209
rect 13909 11200 13921 11203
rect 13872 11172 13921 11200
rect 13872 11160 13878 11172
rect 13909 11169 13921 11172
rect 13955 11169 13967 11203
rect 16206 11200 16212 11212
rect 16167 11172 16212 11200
rect 13909 11163 13967 11169
rect 16206 11160 16212 11172
rect 16264 11160 16270 11212
rect 16393 11203 16451 11209
rect 16393 11169 16405 11203
rect 16439 11169 16451 11203
rect 16393 11163 16451 11169
rect 18141 11203 18199 11209
rect 18141 11169 18153 11203
rect 18187 11200 18199 11203
rect 18230 11200 18236 11212
rect 18187 11172 18236 11200
rect 18187 11169 18199 11172
rect 18141 11163 18199 11169
rect 10318 11132 10324 11144
rect 10244 11104 10324 11132
rect 10318 11092 10324 11104
rect 10376 11092 10382 11144
rect 14274 11132 14280 11144
rect 14235 11104 14280 11132
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 15378 11092 15384 11144
rect 15436 11132 15442 11144
rect 16408 11132 16436 11163
rect 18230 11160 18236 11172
rect 18288 11160 18294 11212
rect 18325 11203 18383 11209
rect 18325 11169 18337 11203
rect 18371 11200 18383 11203
rect 18877 11203 18935 11209
rect 18877 11200 18889 11203
rect 18371 11172 18889 11200
rect 18371 11169 18383 11172
rect 18325 11163 18383 11169
rect 18877 11169 18889 11172
rect 18923 11200 18935 11203
rect 18966 11200 18972 11212
rect 18923 11172 18972 11200
rect 18923 11169 18935 11172
rect 18877 11163 18935 11169
rect 17402 11132 17408 11144
rect 15436 11104 17408 11132
rect 15436 11092 15442 11104
rect 17402 11092 17408 11104
rect 17460 11132 17466 11144
rect 18340 11132 18368 11163
rect 18966 11160 18972 11172
rect 19024 11160 19030 11212
rect 19613 11203 19671 11209
rect 19613 11169 19625 11203
rect 19659 11200 19671 11203
rect 19886 11200 19892 11212
rect 19659 11172 19892 11200
rect 19659 11169 19671 11172
rect 19613 11163 19671 11169
rect 19886 11160 19892 11172
rect 19944 11160 19950 11212
rect 21085 11203 21143 11209
rect 21085 11169 21097 11203
rect 21131 11169 21143 11203
rect 21085 11163 21143 11169
rect 21453 11203 21511 11209
rect 21453 11169 21465 11203
rect 21499 11200 21511 11203
rect 23014 11200 23020 11212
rect 21499 11172 23020 11200
rect 21499 11169 21511 11172
rect 21453 11163 21511 11169
rect 17460 11104 18368 11132
rect 19904 11132 19932 11160
rect 21100 11132 21128 11163
rect 23014 11160 23020 11172
rect 23072 11160 23078 11212
rect 23198 11160 23204 11212
rect 23256 11200 23262 11212
rect 23293 11203 23351 11209
rect 23293 11200 23305 11203
rect 23256 11172 23305 11200
rect 23256 11160 23262 11172
rect 23293 11169 23305 11172
rect 23339 11169 23351 11203
rect 23293 11163 23351 11169
rect 23658 11160 23664 11212
rect 23716 11200 23722 11212
rect 24302 11200 24308 11212
rect 23716 11172 24308 11200
rect 23716 11160 23722 11172
rect 24302 11160 24308 11172
rect 24360 11200 24366 11212
rect 24872 11209 24900 11240
rect 29178 11228 29184 11280
rect 29236 11268 29242 11280
rect 30282 11268 30288 11280
rect 29236 11240 30288 11268
rect 29236 11228 29242 11240
rect 24397 11203 24455 11209
rect 24397 11200 24409 11203
rect 24360 11172 24409 11200
rect 24360 11160 24366 11172
rect 24397 11169 24409 11172
rect 24443 11169 24455 11203
rect 24397 11163 24455 11169
rect 24857 11203 24915 11209
rect 24857 11169 24869 11203
rect 24903 11200 24915 11203
rect 25038 11200 25044 11212
rect 24903 11172 25044 11200
rect 24903 11169 24915 11172
rect 24857 11163 24915 11169
rect 25038 11160 25044 11172
rect 25096 11160 25102 11212
rect 25314 11160 25320 11212
rect 25372 11200 25378 11212
rect 26050 11200 26056 11212
rect 25372 11172 26056 11200
rect 25372 11160 25378 11172
rect 26050 11160 26056 11172
rect 26108 11200 26114 11212
rect 26513 11203 26571 11209
rect 26513 11200 26525 11203
rect 26108 11172 26525 11200
rect 26108 11160 26114 11172
rect 26513 11169 26525 11172
rect 26559 11169 26571 11203
rect 26513 11163 26571 11169
rect 26694 11160 26700 11212
rect 26752 11200 26758 11212
rect 26973 11203 27031 11209
rect 26973 11200 26985 11203
rect 26752 11172 26985 11200
rect 26752 11160 26758 11172
rect 26973 11169 26985 11172
rect 27019 11200 27031 11203
rect 27982 11200 27988 11212
rect 27019 11172 27988 11200
rect 27019 11169 27031 11172
rect 26973 11163 27031 11169
rect 27982 11160 27988 11172
rect 28040 11160 28046 11212
rect 28144 11203 28202 11209
rect 28144 11169 28156 11203
rect 28190 11200 28202 11203
rect 28258 11200 28264 11212
rect 28190 11172 28264 11200
rect 28190 11169 28202 11172
rect 28144 11163 28202 11169
rect 28258 11160 28264 11172
rect 28316 11160 28322 11212
rect 30024 11209 30052 11240
rect 30282 11228 30288 11240
rect 30340 11228 30346 11280
rect 35526 11228 35532 11280
rect 35584 11268 35590 11280
rect 36817 11271 36875 11277
rect 35584 11240 36584 11268
rect 35584 11228 35590 11240
rect 36556 11212 36584 11240
rect 36817 11237 36829 11271
rect 36863 11268 36875 11271
rect 36906 11268 36912 11280
rect 36863 11240 36912 11268
rect 36863 11237 36875 11240
rect 36817 11231 36875 11237
rect 36906 11228 36912 11240
rect 36964 11228 36970 11280
rect 37642 11228 37648 11280
rect 37700 11268 37706 11280
rect 37921 11271 37979 11277
rect 37921 11268 37933 11271
rect 37700 11240 37933 11268
rect 37700 11228 37706 11240
rect 37921 11237 37933 11240
rect 37967 11237 37979 11271
rect 37921 11231 37979 11237
rect 29549 11203 29607 11209
rect 29549 11169 29561 11203
rect 29595 11169 29607 11203
rect 29549 11163 29607 11169
rect 30009 11203 30067 11209
rect 30009 11169 30021 11203
rect 30055 11169 30067 11203
rect 30009 11163 30067 11169
rect 25774 11132 25780 11144
rect 19904 11104 21128 11132
rect 25735 11104 25780 11132
rect 17460 11092 17466 11104
rect 25774 11092 25780 11104
rect 25832 11132 25838 11144
rect 29564 11132 29592 11163
rect 31846 11160 31852 11212
rect 31904 11200 31910 11212
rect 32160 11203 32218 11209
rect 32160 11200 32172 11203
rect 31904 11172 32172 11200
rect 31904 11160 31910 11172
rect 32160 11169 32172 11172
rect 32206 11169 32218 11203
rect 32160 11163 32218 11169
rect 35161 11203 35219 11209
rect 35161 11169 35173 11203
rect 35207 11200 35219 11203
rect 35250 11200 35256 11212
rect 35207 11172 35256 11200
rect 35207 11169 35219 11172
rect 35161 11163 35219 11169
rect 35250 11160 35256 11172
rect 35308 11160 35314 11212
rect 36262 11200 36268 11212
rect 36223 11172 36268 11200
rect 36262 11160 36268 11172
rect 36320 11160 36326 11212
rect 36538 11200 36544 11212
rect 36451 11172 36544 11200
rect 36538 11160 36544 11172
rect 36596 11160 36602 11212
rect 39390 11160 39396 11212
rect 39448 11200 39454 11212
rect 39592 11209 39620 11308
rect 40494 11296 40500 11308
rect 40552 11296 40558 11348
rect 40037 11271 40095 11277
rect 40037 11237 40049 11271
rect 40083 11268 40095 11271
rect 41138 11268 41144 11280
rect 40083 11240 41144 11268
rect 40083 11237 40095 11240
rect 40037 11231 40095 11237
rect 41138 11228 41144 11240
rect 41196 11228 41202 11280
rect 39577 11203 39635 11209
rect 39577 11200 39589 11203
rect 39448 11172 39589 11200
rect 39448 11160 39454 11172
rect 39577 11169 39589 11172
rect 39623 11169 39635 11203
rect 39758 11200 39764 11212
rect 39719 11172 39764 11200
rect 39577 11163 39635 11169
rect 39758 11160 39764 11172
rect 39816 11160 39822 11212
rect 29730 11132 29736 11144
rect 25832 11104 29736 11132
rect 25832 11092 25838 11104
rect 29730 11092 29736 11104
rect 29788 11092 29794 11144
rect 30285 11135 30343 11141
rect 30285 11101 30297 11135
rect 30331 11132 30343 11135
rect 30558 11132 30564 11144
rect 30331 11104 30564 11132
rect 30331 11101 30343 11104
rect 30285 11095 30343 11101
rect 30558 11092 30564 11104
rect 30616 11132 30622 11144
rect 30929 11135 30987 11141
rect 30929 11132 30941 11135
rect 30616 11104 30941 11132
rect 30616 11092 30622 11104
rect 30929 11101 30941 11104
rect 30975 11101 30987 11135
rect 30929 11095 30987 11101
rect 36722 11092 36728 11144
rect 36780 11132 36786 11144
rect 37829 11135 37887 11141
rect 37829 11132 37841 11135
rect 36780 11104 37841 11132
rect 36780 11092 36786 11104
rect 37829 11101 37841 11104
rect 37875 11101 37887 11135
rect 38286 11132 38292 11144
rect 38247 11104 38292 11132
rect 37829 11095 37887 11101
rect 38286 11092 38292 11104
rect 38344 11092 38350 11144
rect 15746 11024 15752 11076
rect 15804 11064 15810 11076
rect 22005 11067 22063 11073
rect 22005 11064 22017 11067
rect 15804 11036 22017 11064
rect 15804 11024 15810 11036
rect 22005 11033 22017 11036
rect 22051 11064 22063 11067
rect 22462 11064 22468 11076
rect 22051 11036 22468 11064
rect 22051 11033 22063 11036
rect 22005 11027 22063 11033
rect 22462 11024 22468 11036
rect 22520 11024 22526 11076
rect 27246 11024 27252 11076
rect 27304 11064 27310 11076
rect 28215 11067 28273 11073
rect 28215 11064 28227 11067
rect 27304 11036 28227 11064
rect 27304 11024 27310 11036
rect 28215 11033 28227 11036
rect 28261 11033 28273 11067
rect 28215 11027 28273 11033
rect 16206 10956 16212 11008
rect 16264 10996 16270 11008
rect 17126 10996 17132 11008
rect 16264 10968 17132 10996
rect 16264 10956 16270 10968
rect 17126 10956 17132 10968
rect 17184 10996 17190 11008
rect 20533 10999 20591 11005
rect 20533 10996 20545 10999
rect 17184 10968 20545 10996
rect 17184 10956 17190 10968
rect 20533 10965 20545 10968
rect 20579 10996 20591 10999
rect 20806 10996 20812 11008
rect 20579 10968 20812 10996
rect 20579 10965 20591 10968
rect 20533 10959 20591 10965
rect 20806 10956 20812 10968
rect 20864 10956 20870 11008
rect 22649 10999 22707 11005
rect 22649 10965 22661 10999
rect 22695 10996 22707 10999
rect 22830 10996 22836 11008
rect 22695 10968 22836 10996
rect 22695 10965 22707 10968
rect 22649 10959 22707 10965
rect 22830 10956 22836 10968
rect 22888 10956 22894 11008
rect 27985 10999 28043 11005
rect 27985 10965 27997 10999
rect 28031 10996 28043 10999
rect 28350 10996 28356 11008
rect 28031 10968 28356 10996
rect 28031 10965 28043 10968
rect 27985 10959 28043 10965
rect 28350 10956 28356 10968
rect 28408 10956 28414 11008
rect 29270 10996 29276 11008
rect 29231 10968 29276 10996
rect 29270 10956 29276 10968
rect 29328 10956 29334 11008
rect 32263 10999 32321 11005
rect 32263 10965 32275 10999
rect 32309 10996 32321 10999
rect 32490 10996 32496 11008
rect 32309 10968 32496 10996
rect 32309 10965 32321 10968
rect 32263 10959 32321 10965
rect 32490 10956 32496 10968
rect 32548 10956 32554 11008
rect 34698 10956 34704 11008
rect 34756 10996 34762 11008
rect 34793 10999 34851 11005
rect 34793 10996 34805 10999
rect 34756 10968 34805 10996
rect 34756 10956 34762 10968
rect 34793 10965 34805 10968
rect 34839 10965 34851 10999
rect 34793 10959 34851 10965
rect 1104 10906 48852 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 48852 10906
rect 1104 10832 48852 10854
rect 10778 10792 10784 10804
rect 10739 10764 10784 10792
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 11882 10792 11888 10804
rect 11843 10764 11888 10792
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 12710 10792 12716 10804
rect 12671 10764 12716 10792
rect 12710 10752 12716 10764
rect 12768 10752 12774 10804
rect 14553 10795 14611 10801
rect 14553 10761 14565 10795
rect 14599 10792 14611 10795
rect 14642 10792 14648 10804
rect 14599 10764 14648 10792
rect 14599 10761 14611 10764
rect 14553 10755 14611 10761
rect 14642 10752 14648 10764
rect 14700 10752 14706 10804
rect 14921 10795 14979 10801
rect 14921 10761 14933 10795
rect 14967 10792 14979 10795
rect 18414 10792 18420 10804
rect 14967 10764 18420 10792
rect 14967 10761 14979 10764
rect 14921 10755 14979 10761
rect 18414 10752 18420 10764
rect 18472 10792 18478 10804
rect 18601 10795 18659 10801
rect 18601 10792 18613 10795
rect 18472 10764 18613 10792
rect 18472 10752 18478 10764
rect 18601 10761 18613 10764
rect 18647 10761 18659 10795
rect 19058 10792 19064 10804
rect 19019 10764 19064 10792
rect 18601 10755 18659 10761
rect 14660 10724 14688 10752
rect 16850 10724 16856 10736
rect 14660 10696 16856 10724
rect 16850 10684 16856 10696
rect 16908 10684 16914 10736
rect 17126 10724 17132 10736
rect 17087 10696 17132 10724
rect 17126 10684 17132 10696
rect 17184 10684 17190 10736
rect 17402 10724 17408 10736
rect 17363 10696 17408 10724
rect 17402 10684 17408 10696
rect 17460 10724 17466 10736
rect 17773 10727 17831 10733
rect 17773 10724 17785 10727
rect 17460 10696 17785 10724
rect 17460 10684 17466 10696
rect 17773 10693 17785 10696
rect 17819 10693 17831 10727
rect 17773 10687 17831 10693
rect 9674 10656 9680 10668
rect 9635 10628 9680 10656
rect 9674 10616 9680 10628
rect 9732 10616 9738 10668
rect 13630 10616 13636 10668
rect 13688 10656 13694 10668
rect 15562 10656 15568 10668
rect 13688 10628 15332 10656
rect 15475 10628 15568 10656
rect 13688 10616 13694 10628
rect 9309 10591 9367 10597
rect 9309 10557 9321 10591
rect 9355 10588 9367 10591
rect 10045 10591 10103 10597
rect 10045 10588 10057 10591
rect 9355 10560 10057 10588
rect 9355 10557 9367 10560
rect 9309 10551 9367 10557
rect 10045 10557 10057 10560
rect 10091 10588 10103 10591
rect 10686 10588 10692 10600
rect 10091 10560 10692 10588
rect 10091 10557 10103 10560
rect 10045 10551 10103 10557
rect 10686 10548 10692 10560
rect 10744 10588 10750 10600
rect 12434 10588 12440 10600
rect 10744 10560 11468 10588
rect 12395 10560 12440 10588
rect 10744 10548 10750 10560
rect 9033 10523 9091 10529
rect 9033 10489 9045 10523
rect 9079 10520 9091 10523
rect 9125 10523 9183 10529
rect 9125 10520 9137 10523
rect 9079 10492 9137 10520
rect 9079 10489 9091 10492
rect 9033 10483 9091 10489
rect 9125 10489 9137 10492
rect 9171 10520 9183 10523
rect 9766 10520 9772 10532
rect 9171 10492 9772 10520
rect 9171 10489 9183 10492
rect 9125 10483 9183 10489
rect 9766 10480 9772 10492
rect 9824 10480 9830 10532
rect 10413 10523 10471 10529
rect 10413 10489 10425 10523
rect 10459 10520 10471 10523
rect 10502 10520 10508 10532
rect 10459 10492 10508 10520
rect 10459 10489 10471 10492
rect 10413 10483 10471 10489
rect 10502 10480 10508 10492
rect 10560 10480 10566 10532
rect 11440 10529 11468 10560
rect 12434 10548 12440 10560
rect 12492 10548 12498 10600
rect 12621 10591 12679 10597
rect 12621 10557 12633 10591
rect 12667 10588 12679 10591
rect 13357 10591 13415 10597
rect 13357 10588 13369 10591
rect 12667 10560 13369 10588
rect 12667 10557 12679 10560
rect 12621 10551 12679 10557
rect 13357 10557 13369 10560
rect 13403 10588 13415 10591
rect 14461 10591 14519 10597
rect 14461 10588 14473 10591
rect 13403 10560 14473 10588
rect 13403 10557 13415 10560
rect 13357 10551 13415 10557
rect 14461 10557 14473 10560
rect 14507 10588 14519 10591
rect 14507 10560 15240 10588
rect 14507 10557 14519 10560
rect 14461 10551 14519 10557
rect 11425 10523 11483 10529
rect 11425 10489 11437 10523
rect 11471 10520 11483 10523
rect 12253 10523 12311 10529
rect 12253 10520 12265 10523
rect 11471 10492 12265 10520
rect 11471 10489 11483 10492
rect 11425 10483 11483 10489
rect 12253 10489 12265 10492
rect 12299 10520 12311 10523
rect 12526 10520 12532 10532
rect 12299 10492 12532 10520
rect 12299 10489 12311 10492
rect 12253 10483 12311 10489
rect 12526 10480 12532 10492
rect 12584 10520 12590 10532
rect 12636 10520 12664 10551
rect 13722 10520 13728 10532
rect 12584 10492 12664 10520
rect 13509 10492 13728 10520
rect 12584 10480 12590 10492
rect 9214 10412 9220 10464
rect 9272 10452 9278 10464
rect 12710 10452 12716 10464
rect 9272 10424 12716 10452
rect 9272 10412 9278 10424
rect 12710 10412 12716 10424
rect 12768 10452 12774 10464
rect 13509 10452 13537 10492
rect 13722 10480 13728 10492
rect 13780 10520 13786 10532
rect 14093 10523 14151 10529
rect 14093 10520 14105 10523
rect 13780 10492 14105 10520
rect 13780 10480 13786 10492
rect 14093 10489 14105 10492
rect 14139 10489 14151 10523
rect 14274 10520 14280 10532
rect 14187 10492 14280 10520
rect 14093 10483 14151 10489
rect 14274 10480 14280 10492
rect 14332 10520 14338 10532
rect 14921 10523 14979 10529
rect 14921 10520 14933 10523
rect 14332 10492 14933 10520
rect 14332 10480 14338 10492
rect 14921 10489 14933 10492
rect 14967 10489 14979 10523
rect 14921 10483 14979 10489
rect 15212 10464 15240 10560
rect 15304 10520 15332 10628
rect 15562 10616 15568 10628
rect 15620 10656 15626 10668
rect 16117 10659 16175 10665
rect 16117 10656 16129 10659
rect 15620 10628 16129 10656
rect 15620 10616 15626 10628
rect 16117 10625 16129 10628
rect 16163 10625 16175 10659
rect 16117 10619 16175 10625
rect 16761 10659 16819 10665
rect 16761 10625 16773 10659
rect 16807 10656 16819 10659
rect 17678 10656 17684 10668
rect 16807 10628 17684 10656
rect 16807 10625 16819 10628
rect 16761 10619 16819 10625
rect 17678 10616 17684 10628
rect 17736 10616 17742 10668
rect 15654 10548 15660 10600
rect 15712 10588 15718 10600
rect 16025 10591 16083 10597
rect 16025 10588 16037 10591
rect 15712 10560 16037 10588
rect 15712 10548 15718 10560
rect 16025 10557 16037 10560
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 16301 10591 16359 10597
rect 16301 10557 16313 10591
rect 16347 10557 16359 10591
rect 18616 10588 18644 10755
rect 19058 10752 19064 10764
rect 19116 10752 19122 10804
rect 20714 10752 20720 10804
rect 20772 10792 20778 10804
rect 21821 10795 21879 10801
rect 21821 10792 21833 10795
rect 20772 10764 21833 10792
rect 20772 10752 20778 10764
rect 21821 10761 21833 10764
rect 21867 10761 21879 10795
rect 23014 10792 23020 10804
rect 22975 10764 23020 10792
rect 21821 10755 21879 10761
rect 23014 10752 23020 10764
rect 23072 10752 23078 10804
rect 24302 10792 24308 10804
rect 24263 10764 24308 10792
rect 24302 10752 24308 10764
rect 24360 10752 24366 10804
rect 27525 10795 27583 10801
rect 27525 10761 27537 10795
rect 27571 10792 27583 10795
rect 28169 10795 28227 10801
rect 28169 10792 28181 10795
rect 27571 10764 28181 10792
rect 27571 10761 27583 10764
rect 27525 10755 27583 10761
rect 28169 10761 28181 10764
rect 28215 10792 28227 10795
rect 28258 10792 28264 10804
rect 28215 10764 28264 10792
rect 28215 10761 28227 10764
rect 28169 10755 28227 10761
rect 28258 10752 28264 10764
rect 28316 10752 28322 10804
rect 28350 10752 28356 10804
rect 28408 10792 28414 10804
rect 29411 10795 29469 10801
rect 29411 10792 29423 10795
rect 28408 10764 29423 10792
rect 28408 10752 28414 10764
rect 29411 10761 29423 10764
rect 29457 10761 29469 10795
rect 29730 10792 29736 10804
rect 29691 10764 29736 10792
rect 29411 10755 29469 10761
rect 29730 10752 29736 10764
rect 29788 10752 29794 10804
rect 30469 10795 30527 10801
rect 30469 10761 30481 10795
rect 30515 10792 30527 10795
rect 30926 10792 30932 10804
rect 30515 10764 30932 10792
rect 30515 10761 30527 10764
rect 30469 10755 30527 10761
rect 30926 10752 30932 10764
rect 30984 10752 30990 10804
rect 34333 10795 34391 10801
rect 34333 10761 34345 10795
rect 34379 10792 34391 10795
rect 35250 10792 35256 10804
rect 34379 10764 35256 10792
rect 34379 10761 34391 10764
rect 34333 10755 34391 10761
rect 35250 10752 35256 10764
rect 35308 10752 35314 10804
rect 36173 10795 36231 10801
rect 36173 10761 36185 10795
rect 36219 10792 36231 10795
rect 36262 10792 36268 10804
rect 36219 10764 36268 10792
rect 36219 10761 36231 10764
rect 36173 10755 36231 10761
rect 36262 10752 36268 10764
rect 36320 10752 36326 10804
rect 36538 10792 36544 10804
rect 36499 10764 36544 10792
rect 36538 10752 36544 10764
rect 36596 10752 36602 10804
rect 36722 10752 36728 10804
rect 36780 10792 36786 10804
rect 37277 10795 37335 10801
rect 37277 10792 37289 10795
rect 36780 10764 37289 10792
rect 36780 10752 36786 10764
rect 37277 10761 37289 10764
rect 37323 10761 37335 10795
rect 37277 10755 37335 10761
rect 37642 10752 37648 10804
rect 37700 10792 37706 10804
rect 38289 10795 38347 10801
rect 38289 10792 38301 10795
rect 37700 10764 38301 10792
rect 37700 10752 37706 10764
rect 38289 10761 38301 10764
rect 38335 10761 38347 10795
rect 39390 10792 39396 10804
rect 39351 10764 39396 10792
rect 38289 10755 38347 10761
rect 39390 10752 39396 10764
rect 39448 10752 39454 10804
rect 27982 10684 27988 10736
rect 28040 10724 28046 10736
rect 28997 10727 29055 10733
rect 28997 10724 29009 10727
rect 28040 10696 29009 10724
rect 28040 10684 28046 10696
rect 28997 10693 29009 10696
rect 29043 10724 29055 10727
rect 29178 10724 29184 10736
rect 29043 10696 29184 10724
rect 29043 10693 29055 10696
rect 28997 10687 29055 10693
rect 29178 10684 29184 10696
rect 29236 10684 29242 10736
rect 34698 10724 34704 10736
rect 34659 10696 34704 10724
rect 34698 10684 34704 10696
rect 34756 10684 34762 10736
rect 37734 10684 37740 10736
rect 37792 10724 37798 10736
rect 37921 10727 37979 10733
rect 37921 10724 37933 10727
rect 37792 10696 37933 10724
rect 37792 10684 37798 10696
rect 37921 10693 37933 10696
rect 37967 10724 37979 10727
rect 38838 10724 38844 10736
rect 37967 10696 38844 10724
rect 37967 10693 37979 10696
rect 37921 10687 37979 10693
rect 38838 10684 38844 10696
rect 38896 10684 38902 10736
rect 38930 10684 38936 10736
rect 38988 10724 38994 10736
rect 39669 10727 39727 10733
rect 39669 10724 39681 10727
rect 38988 10696 39681 10724
rect 38988 10684 38994 10696
rect 39669 10693 39681 10696
rect 39715 10724 39727 10727
rect 39758 10724 39764 10736
rect 39715 10696 39764 10724
rect 39715 10693 39727 10696
rect 39669 10687 39727 10693
rect 39758 10684 39764 10696
rect 39816 10684 39822 10736
rect 22281 10659 22339 10665
rect 22281 10656 22293 10659
rect 21376 10628 22293 10656
rect 18785 10591 18843 10597
rect 18785 10588 18797 10591
rect 18616 10560 18797 10588
rect 16301 10551 16359 10557
rect 18785 10557 18797 10560
rect 18831 10557 18843 10591
rect 18785 10551 18843 10557
rect 18969 10591 19027 10597
rect 18969 10557 18981 10591
rect 19015 10588 19027 10591
rect 20809 10591 20867 10597
rect 19015 10560 19472 10588
rect 19015 10557 19027 10560
rect 18969 10551 19027 10557
rect 15933 10523 15991 10529
rect 15933 10520 15945 10523
rect 15304 10492 15945 10520
rect 15933 10489 15945 10492
rect 15979 10520 15991 10523
rect 16316 10520 16344 10551
rect 15979 10492 16344 10520
rect 15979 10489 15991 10492
rect 15933 10483 15991 10489
rect 19444 10464 19472 10560
rect 20809 10557 20821 10591
rect 20855 10557 20867 10591
rect 20809 10551 20867 10557
rect 19886 10480 19892 10532
rect 19944 10520 19950 10532
rect 19981 10523 20039 10529
rect 19981 10520 19993 10523
rect 19944 10492 19993 10520
rect 19944 10480 19950 10492
rect 19981 10489 19993 10492
rect 20027 10520 20039 10523
rect 20625 10523 20683 10529
rect 20625 10520 20637 10523
rect 20027 10492 20637 10520
rect 20027 10489 20039 10492
rect 19981 10483 20039 10489
rect 20625 10489 20637 10492
rect 20671 10489 20683 10523
rect 20824 10520 20852 10551
rect 20898 10548 20904 10600
rect 20956 10588 20962 10600
rect 21376 10597 21404 10628
rect 22281 10625 22293 10628
rect 22327 10625 22339 10659
rect 26602 10656 26608 10668
rect 26563 10628 26608 10656
rect 22281 10619 22339 10625
rect 26602 10616 26608 10628
rect 26660 10616 26666 10668
rect 30558 10656 30564 10668
rect 30519 10628 30564 10656
rect 30558 10616 30564 10628
rect 30616 10616 30622 10668
rect 32493 10659 32551 10665
rect 32493 10625 32505 10659
rect 32539 10656 32551 10659
rect 33502 10656 33508 10668
rect 32539 10628 33508 10656
rect 32539 10625 32551 10628
rect 32493 10619 32551 10625
rect 33502 10616 33508 10628
rect 33560 10616 33566 10668
rect 21361 10591 21419 10597
rect 21361 10588 21373 10591
rect 20956 10560 21373 10588
rect 20956 10548 20962 10560
rect 21361 10557 21373 10560
rect 21407 10557 21419 10591
rect 21361 10551 21419 10557
rect 22624 10591 22682 10597
rect 22624 10557 22636 10591
rect 22670 10588 22682 10591
rect 22830 10588 22836 10600
rect 22670 10560 22836 10588
rect 22670 10557 22682 10560
rect 22624 10551 22682 10557
rect 22830 10548 22836 10560
rect 22888 10548 22894 10600
rect 23566 10588 23572 10600
rect 23527 10560 23572 10588
rect 23566 10548 23572 10560
rect 23624 10548 23630 10600
rect 24854 10588 24860 10600
rect 24815 10560 24860 10588
rect 24854 10548 24860 10560
rect 24912 10548 24918 10600
rect 25777 10591 25835 10597
rect 25777 10557 25789 10591
rect 25823 10588 25835 10591
rect 29270 10588 29276 10600
rect 29328 10597 29334 10600
rect 29328 10591 29366 10597
rect 25823 10560 29276 10588
rect 25823 10557 25835 10560
rect 25777 10551 25835 10557
rect 29270 10548 29276 10560
rect 29354 10557 29366 10591
rect 29328 10551 29366 10557
rect 37528 10591 37586 10597
rect 37528 10557 37540 10591
rect 37574 10588 37586 10591
rect 37752 10588 37780 10684
rect 37574 10560 37780 10588
rect 37574 10557 37586 10560
rect 37528 10551 37586 10557
rect 29328 10548 29334 10551
rect 20990 10520 20996 10532
rect 20824 10492 20996 10520
rect 20625 10483 20683 10489
rect 20990 10480 20996 10492
rect 21048 10480 21054 10532
rect 21542 10520 21548 10532
rect 21503 10492 21548 10520
rect 21542 10480 21548 10492
rect 21600 10480 21606 10532
rect 23290 10480 23296 10532
rect 23348 10520 23354 10532
rect 23799 10523 23857 10529
rect 23799 10520 23811 10523
rect 23348 10492 23811 10520
rect 23348 10480 23354 10492
rect 23799 10489 23811 10492
rect 23845 10489 23857 10523
rect 23799 10483 23857 10489
rect 24670 10480 24676 10532
rect 24728 10520 24734 10532
rect 24765 10523 24823 10529
rect 24765 10520 24777 10523
rect 24728 10492 24777 10520
rect 24728 10480 24734 10492
rect 24765 10489 24777 10492
rect 24811 10520 24823 10523
rect 25219 10523 25277 10529
rect 25219 10520 25231 10523
rect 24811 10492 25231 10520
rect 24811 10489 24823 10492
rect 24765 10483 24823 10489
rect 25219 10489 25231 10492
rect 25265 10520 25277 10523
rect 26513 10523 26571 10529
rect 26513 10520 26525 10523
rect 25265 10492 26525 10520
rect 25265 10489 25277 10492
rect 25219 10483 25277 10489
rect 26513 10489 26525 10492
rect 26559 10520 26571 10523
rect 26967 10523 27025 10529
rect 26967 10520 26979 10523
rect 26559 10492 26979 10520
rect 26559 10489 26571 10492
rect 26513 10483 26571 10489
rect 26967 10489 26979 10492
rect 27013 10489 27025 10523
rect 26967 10483 27025 10489
rect 32309 10523 32367 10529
rect 32309 10489 32321 10523
rect 32355 10520 32367 10523
rect 32582 10520 32588 10532
rect 32355 10492 32588 10520
rect 32355 10489 32367 10492
rect 32309 10483 32367 10489
rect 32582 10480 32588 10492
rect 32640 10480 32646 10532
rect 33134 10480 33140 10532
rect 33192 10520 33198 10532
rect 34974 10520 34980 10532
rect 33192 10492 34980 10520
rect 33192 10480 33198 10492
rect 34974 10480 34980 10492
rect 35032 10480 35038 10532
rect 35069 10523 35127 10529
rect 35069 10489 35081 10523
rect 35115 10489 35127 10523
rect 35069 10483 35127 10489
rect 35621 10523 35679 10529
rect 35621 10489 35633 10523
rect 35667 10520 35679 10523
rect 36170 10520 36176 10532
rect 35667 10492 36176 10520
rect 35667 10489 35679 10492
rect 35621 10483 35679 10489
rect 12768 10424 13537 10452
rect 12768 10412 12774 10424
rect 13814 10412 13820 10464
rect 13872 10452 13878 10464
rect 15194 10452 15200 10464
rect 13872 10424 13917 10452
rect 15155 10424 15200 10452
rect 13872 10412 13878 10424
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 18322 10452 18328 10464
rect 18283 10424 18328 10452
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 19426 10412 19432 10464
rect 19484 10452 19490 10464
rect 19613 10455 19671 10461
rect 19613 10452 19625 10455
rect 19484 10424 19625 10452
rect 19484 10412 19490 10424
rect 19613 10421 19625 10424
rect 19659 10421 19671 10455
rect 19613 10415 19671 10421
rect 22695 10455 22753 10461
rect 22695 10421 22707 10455
rect 22741 10452 22753 10455
rect 22922 10452 22928 10464
rect 22741 10424 22928 10452
rect 22741 10421 22753 10424
rect 22695 10415 22753 10421
rect 22922 10412 22928 10424
rect 22980 10412 22986 10464
rect 23198 10412 23204 10464
rect 23256 10452 23262 10464
rect 23385 10455 23443 10461
rect 23385 10452 23397 10455
rect 23256 10424 23397 10452
rect 23256 10412 23262 10424
rect 23385 10421 23397 10424
rect 23431 10421 23443 10455
rect 26050 10452 26056 10464
rect 26011 10424 26056 10452
rect 23385 10415 23443 10421
rect 26050 10412 26056 10424
rect 26108 10412 26114 10464
rect 30926 10452 30932 10464
rect 30887 10424 30932 10452
rect 30926 10412 30932 10424
rect 30984 10412 30990 10464
rect 31478 10452 31484 10464
rect 31439 10424 31484 10452
rect 31478 10412 31484 10424
rect 31536 10412 31542 10464
rect 31846 10452 31852 10464
rect 31807 10424 31852 10452
rect 31846 10412 31852 10424
rect 31904 10412 31910 10464
rect 33502 10452 33508 10464
rect 33463 10424 33508 10452
rect 33502 10412 33508 10424
rect 33560 10412 33566 10464
rect 34698 10412 34704 10464
rect 34756 10452 34762 10464
rect 35084 10452 35112 10483
rect 36170 10480 36176 10492
rect 36228 10480 36234 10532
rect 34756 10424 35112 10452
rect 37599 10455 37657 10461
rect 34756 10412 34762 10424
rect 37599 10421 37611 10455
rect 37645 10452 37657 10455
rect 37826 10452 37832 10464
rect 37645 10424 37832 10452
rect 37645 10421 37657 10424
rect 37599 10415 37657 10421
rect 37826 10412 37832 10424
rect 37884 10412 37890 10464
rect 1104 10362 48852 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 48852 10362
rect 1104 10288 48852 10310
rect 10137 10251 10195 10257
rect 10137 10217 10149 10251
rect 10183 10248 10195 10251
rect 10318 10248 10324 10260
rect 10183 10220 10324 10248
rect 10183 10217 10195 10220
rect 10137 10211 10195 10217
rect 10318 10208 10324 10220
rect 10376 10248 10382 10260
rect 10781 10251 10839 10257
rect 10781 10248 10793 10251
rect 10376 10220 10793 10248
rect 10376 10208 10382 10220
rect 10781 10217 10793 10220
rect 10827 10217 10839 10251
rect 10781 10211 10839 10217
rect 12161 10251 12219 10257
rect 12161 10217 12173 10251
rect 12207 10217 12219 10251
rect 12161 10211 12219 10217
rect 10505 10183 10563 10189
rect 10505 10149 10517 10183
rect 10551 10180 10563 10183
rect 10594 10180 10600 10192
rect 10551 10152 10600 10180
rect 10551 10149 10563 10152
rect 10505 10143 10563 10149
rect 10594 10140 10600 10152
rect 10652 10180 10658 10192
rect 11238 10180 11244 10192
rect 10652 10152 11244 10180
rect 10652 10140 10658 10152
rect 11238 10140 11244 10152
rect 11296 10180 11302 10192
rect 12176 10180 12204 10211
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 13725 10251 13783 10257
rect 13725 10248 13737 10251
rect 12492 10220 13737 10248
rect 12492 10208 12498 10220
rect 13725 10217 13737 10220
rect 13771 10217 13783 10251
rect 14274 10248 14280 10260
rect 14235 10220 14280 10248
rect 13725 10211 13783 10217
rect 14274 10208 14280 10220
rect 14332 10208 14338 10260
rect 19334 10248 19340 10260
rect 19295 10220 19340 10248
rect 19334 10208 19340 10220
rect 19392 10208 19398 10260
rect 21223 10251 21281 10257
rect 21223 10217 21235 10251
rect 21269 10248 21281 10251
rect 22278 10248 22284 10260
rect 21269 10220 22284 10248
rect 21269 10217 21281 10220
rect 21223 10211 21281 10217
rect 22278 10208 22284 10220
rect 22336 10208 22342 10260
rect 22465 10251 22523 10257
rect 22465 10217 22477 10251
rect 22511 10248 22523 10251
rect 22554 10248 22560 10260
rect 22511 10220 22560 10248
rect 22511 10217 22523 10220
rect 22465 10211 22523 10217
rect 22554 10208 22560 10220
rect 22612 10208 22618 10260
rect 23017 10251 23075 10257
rect 23017 10217 23029 10251
rect 23063 10248 23075 10251
rect 23566 10248 23572 10260
rect 23063 10220 23572 10248
rect 23063 10217 23075 10220
rect 23017 10211 23075 10217
rect 23566 10208 23572 10220
rect 23624 10248 23630 10260
rect 23661 10251 23719 10257
rect 23661 10248 23673 10251
rect 23624 10220 23673 10248
rect 23624 10208 23630 10220
rect 23661 10217 23673 10220
rect 23707 10217 23719 10251
rect 23661 10211 23719 10217
rect 26329 10251 26387 10257
rect 26329 10217 26341 10251
rect 26375 10248 26387 10251
rect 26602 10248 26608 10260
rect 26375 10220 26608 10248
rect 26375 10217 26387 10220
rect 26329 10211 26387 10217
rect 26602 10208 26608 10220
rect 26660 10208 26666 10260
rect 31205 10251 31263 10257
rect 27356 10220 30788 10248
rect 27356 10192 27384 10220
rect 11296 10152 12204 10180
rect 13096 10152 13538 10180
rect 11296 10140 11302 10152
rect 10686 10112 10692 10124
rect 10647 10084 10692 10112
rect 10686 10072 10692 10084
rect 10744 10072 10750 10124
rect 11882 10112 11888 10124
rect 11843 10084 11888 10112
rect 11882 10072 11888 10084
rect 11940 10072 11946 10124
rect 12070 10115 12128 10121
rect 12070 10081 12082 10115
rect 12116 10112 12128 10115
rect 12158 10112 12164 10124
rect 12116 10084 12164 10112
rect 12116 10081 12128 10084
rect 12070 10075 12128 10081
rect 12158 10072 12164 10084
rect 12216 10112 12222 10124
rect 13096 10112 13124 10152
rect 13510 10124 13538 10152
rect 14550 10140 14556 10192
rect 14608 10180 14614 10192
rect 16114 10180 16120 10192
rect 14608 10152 16120 10180
rect 14608 10140 14614 10152
rect 16114 10140 16120 10152
rect 16172 10140 16178 10192
rect 17678 10140 17684 10192
rect 17736 10180 17742 10192
rect 18049 10183 18107 10189
rect 18049 10180 18061 10183
rect 17736 10152 18061 10180
rect 17736 10140 17742 10152
rect 18049 10149 18061 10152
rect 18095 10149 18107 10183
rect 18049 10143 18107 10149
rect 18322 10140 18328 10192
rect 18380 10180 18386 10192
rect 18601 10183 18659 10189
rect 18601 10180 18613 10183
rect 18380 10152 18613 10180
rect 18380 10140 18386 10152
rect 18601 10149 18613 10152
rect 18647 10180 18659 10183
rect 18647 10152 21956 10180
rect 18647 10149 18659 10152
rect 18601 10143 18659 10149
rect 13262 10112 13268 10124
rect 12216 10084 13124 10112
rect 13223 10084 13268 10112
rect 12216 10072 12222 10084
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 13492 10112 13498 10124
rect 13453 10084 13498 10112
rect 13492 10072 13498 10084
rect 13550 10072 13556 10124
rect 16853 10115 16911 10121
rect 16853 10081 16865 10115
rect 16899 10112 16911 10115
rect 17494 10112 17500 10124
rect 16899 10084 17500 10112
rect 16899 10081 16911 10084
rect 16853 10075 16911 10081
rect 17494 10072 17500 10084
rect 17552 10112 17558 10124
rect 18230 10112 18236 10124
rect 17552 10084 18236 10112
rect 17552 10072 17558 10084
rect 18230 10072 18236 10084
rect 18288 10072 18294 10124
rect 19426 10112 19432 10124
rect 19387 10084 19432 10112
rect 19426 10072 19432 10084
rect 19484 10072 19490 10124
rect 19610 10112 19616 10124
rect 19571 10084 19616 10112
rect 19610 10072 19616 10084
rect 19668 10072 19674 10124
rect 21152 10115 21210 10121
rect 21152 10081 21164 10115
rect 21198 10112 21210 10115
rect 21450 10112 21456 10124
rect 21198 10084 21456 10112
rect 21198 10081 21210 10084
rect 21152 10075 21210 10081
rect 21450 10072 21456 10084
rect 21508 10112 21514 10124
rect 21818 10112 21824 10124
rect 21508 10084 21824 10112
rect 21508 10072 21514 10084
rect 21818 10072 21824 10084
rect 21876 10072 21882 10124
rect 21928 10112 21956 10152
rect 23474 10140 23480 10192
rect 23532 10180 23538 10192
rect 23532 10152 24808 10180
rect 23532 10140 23538 10152
rect 23198 10112 23204 10124
rect 21928 10084 23204 10112
rect 23198 10072 23204 10084
rect 23256 10072 23262 10124
rect 24302 10112 24308 10124
rect 24263 10084 24308 10112
rect 24302 10072 24308 10084
rect 24360 10072 24366 10124
rect 24780 10121 24808 10152
rect 24854 10140 24860 10192
rect 24912 10180 24918 10192
rect 25041 10183 25099 10189
rect 25041 10180 25053 10183
rect 24912 10152 25053 10180
rect 24912 10140 24918 10152
rect 25041 10149 25053 10152
rect 25087 10180 25099 10183
rect 25317 10183 25375 10189
rect 25317 10180 25329 10183
rect 25087 10152 25329 10180
rect 25087 10149 25099 10152
rect 25041 10143 25099 10149
rect 25317 10149 25329 10152
rect 25363 10149 25375 10183
rect 27246 10180 27252 10192
rect 27207 10152 27252 10180
rect 25317 10143 25375 10149
rect 27246 10140 27252 10152
rect 27304 10140 27310 10192
rect 27338 10140 27344 10192
rect 27396 10180 27402 10192
rect 27890 10180 27896 10192
rect 27396 10152 27489 10180
rect 27851 10152 27896 10180
rect 27396 10140 27402 10152
rect 27890 10140 27896 10152
rect 27948 10140 27954 10192
rect 30647 10183 30705 10189
rect 30647 10149 30659 10183
rect 30693 10149 30705 10183
rect 30760 10180 30788 10220
rect 31205 10217 31217 10251
rect 31251 10248 31263 10251
rect 31846 10248 31852 10260
rect 31251 10220 31852 10248
rect 31251 10217 31263 10220
rect 31205 10211 31263 10217
rect 31846 10208 31852 10220
rect 31904 10208 31910 10260
rect 31956 10220 32628 10248
rect 31956 10180 31984 10220
rect 32490 10180 32496 10192
rect 30760 10152 31984 10180
rect 32451 10152 32496 10180
rect 30647 10143 30705 10149
rect 24765 10115 24823 10121
rect 24765 10081 24777 10115
rect 24811 10081 24823 10115
rect 24765 10075 24823 10081
rect 28813 10115 28871 10121
rect 28813 10081 28825 10115
rect 28859 10081 28871 10115
rect 29178 10112 29184 10124
rect 29139 10084 29184 10112
rect 28813 10075 28871 10081
rect 15194 10004 15200 10056
rect 15252 10044 15258 10056
rect 15749 10047 15807 10053
rect 15749 10044 15761 10047
rect 15252 10016 15761 10044
rect 15252 10004 15258 10016
rect 15749 10013 15761 10016
rect 15795 10044 15807 10047
rect 16022 10044 16028 10056
rect 15795 10016 16028 10044
rect 15795 10013 15807 10016
rect 15749 10007 15807 10013
rect 16022 10004 16028 10016
rect 16080 10044 16086 10056
rect 16209 10047 16267 10053
rect 16209 10044 16221 10047
rect 16080 10016 16221 10044
rect 16080 10004 16086 10016
rect 16209 10013 16221 10016
rect 16255 10013 16267 10047
rect 19444 10044 19472 10072
rect 20257 10047 20315 10053
rect 20257 10044 20269 10047
rect 19444 10016 20269 10044
rect 16209 10007 16267 10013
rect 20257 10013 20269 10016
rect 20303 10013 20315 10047
rect 22094 10044 22100 10056
rect 22055 10016 22100 10044
rect 20257 10007 20315 10013
rect 22094 10004 22100 10016
rect 22152 10004 22158 10056
rect 10502 9936 10508 9988
rect 10560 9976 10566 9988
rect 13173 9979 13231 9985
rect 10560 9948 12848 9976
rect 10560 9936 10566 9948
rect 10870 9868 10876 9920
rect 10928 9908 10934 9920
rect 11333 9911 11391 9917
rect 11333 9908 11345 9911
rect 10928 9880 11345 9908
rect 10928 9868 10934 9880
rect 11333 9877 11345 9880
rect 11379 9877 11391 9911
rect 11333 9871 11391 9877
rect 11882 9868 11888 9920
rect 11940 9908 11946 9920
rect 12618 9908 12624 9920
rect 11940 9880 12624 9908
rect 11940 9868 11946 9880
rect 12618 9868 12624 9880
rect 12676 9908 12682 9920
rect 12713 9911 12771 9917
rect 12713 9908 12725 9911
rect 12676 9880 12725 9908
rect 12676 9868 12682 9880
rect 12713 9877 12725 9880
rect 12759 9877 12771 9911
rect 12820 9908 12848 9948
rect 13173 9945 13185 9979
rect 13219 9976 13231 9979
rect 13357 9979 13415 9985
rect 13357 9976 13369 9979
rect 13219 9948 13369 9976
rect 13219 9945 13231 9948
rect 13173 9939 13231 9945
rect 13357 9945 13369 9948
rect 13403 9976 13415 9979
rect 15562 9976 15568 9988
rect 13403 9948 15568 9976
rect 13403 9945 13415 9948
rect 13357 9939 13415 9945
rect 15562 9936 15568 9948
rect 15620 9936 15626 9988
rect 20990 9936 20996 9988
rect 21048 9976 21054 9988
rect 21545 9979 21603 9985
rect 21545 9976 21557 9979
rect 21048 9948 21557 9976
rect 21048 9936 21054 9948
rect 21545 9945 21557 9948
rect 21591 9976 21603 9979
rect 21726 9976 21732 9988
rect 21591 9948 21732 9976
rect 21591 9945 21603 9948
rect 21545 9939 21603 9945
rect 21726 9936 21732 9948
rect 21784 9936 21790 9988
rect 22922 9936 22928 9988
rect 22980 9976 22986 9988
rect 23382 9976 23388 9988
rect 22980 9948 23388 9976
rect 22980 9936 22986 9948
rect 23382 9936 23388 9948
rect 23440 9976 23446 9988
rect 24121 9979 24179 9985
rect 24121 9976 24133 9979
rect 23440 9948 24133 9976
rect 23440 9936 23446 9948
rect 24121 9945 24133 9948
rect 24167 9945 24179 9979
rect 24121 9939 24179 9945
rect 25222 9936 25228 9988
rect 25280 9976 25286 9988
rect 28718 9976 28724 9988
rect 25280 9948 28724 9976
rect 25280 9936 25286 9948
rect 28718 9936 28724 9948
rect 28776 9976 28782 9988
rect 28828 9976 28856 10075
rect 29178 10072 29184 10084
rect 29236 10072 29242 10124
rect 30662 10112 30690 10143
rect 32490 10140 32496 10152
rect 32548 10140 32554 10192
rect 32600 10189 32628 10220
rect 34974 10208 34980 10260
rect 35032 10248 35038 10260
rect 35529 10251 35587 10257
rect 35529 10248 35541 10251
rect 35032 10220 35541 10248
rect 35032 10208 35038 10220
rect 35529 10217 35541 10220
rect 35575 10217 35587 10251
rect 35529 10211 35587 10217
rect 32585 10183 32643 10189
rect 32585 10149 32597 10183
rect 32631 10180 32643 10183
rect 32766 10180 32772 10192
rect 32631 10152 32772 10180
rect 32631 10149 32643 10152
rect 32585 10143 32643 10149
rect 32766 10140 32772 10152
rect 32824 10140 32830 10192
rect 33134 10140 33140 10192
rect 33192 10180 33198 10192
rect 34057 10183 34115 10189
rect 33192 10152 33237 10180
rect 33192 10140 33198 10152
rect 34057 10149 34069 10183
rect 34103 10180 34115 10183
rect 34238 10180 34244 10192
rect 34103 10152 34244 10180
rect 34103 10149 34115 10152
rect 34057 10143 34115 10149
rect 34238 10140 34244 10152
rect 34296 10140 34302 10192
rect 34330 10140 34336 10192
rect 34388 10180 34394 10192
rect 35158 10180 35164 10192
rect 34388 10152 34433 10180
rect 35119 10152 35164 10180
rect 34388 10140 34394 10152
rect 35158 10140 35164 10152
rect 35216 10140 35222 10192
rect 36262 10180 36268 10192
rect 36175 10152 36268 10180
rect 36262 10140 36268 10152
rect 36320 10180 36326 10192
rect 37737 10183 37795 10189
rect 37737 10180 37749 10183
rect 36320 10152 37749 10180
rect 36320 10140 36326 10152
rect 37737 10149 37749 10152
rect 37783 10149 37795 10183
rect 37737 10143 37795 10149
rect 30926 10112 30932 10124
rect 30662 10084 30932 10112
rect 30926 10072 30932 10084
rect 30984 10072 30990 10124
rect 37826 10112 37832 10124
rect 37787 10084 37832 10112
rect 37826 10072 37832 10084
rect 37884 10072 37890 10124
rect 29457 10047 29515 10053
rect 29457 10013 29469 10047
rect 29503 10044 29515 10047
rect 30285 10047 30343 10053
rect 30285 10044 30297 10047
rect 29503 10016 30297 10044
rect 29503 10013 29515 10016
rect 29457 10007 29515 10013
rect 30285 10013 30297 10016
rect 30331 10044 30343 10047
rect 31202 10044 31208 10056
rect 30331 10016 31208 10044
rect 30331 10013 30343 10016
rect 30285 10007 30343 10013
rect 31202 10004 31208 10016
rect 31260 10004 31266 10056
rect 34238 10044 34244 10056
rect 34199 10016 34244 10044
rect 34238 10004 34244 10016
rect 34296 10004 34302 10056
rect 34885 10047 34943 10053
rect 34885 10013 34897 10047
rect 34931 10044 34943 10047
rect 36170 10044 36176 10056
rect 34931 10016 36176 10044
rect 34931 10013 34943 10016
rect 34885 10007 34943 10013
rect 36170 10004 36176 10016
rect 36228 10004 36234 10056
rect 36814 10044 36820 10056
rect 36775 10016 36820 10044
rect 36814 10004 36820 10016
rect 36872 10004 36878 10056
rect 28776 9948 28856 9976
rect 28776 9936 28782 9948
rect 14182 9908 14188 9920
rect 12820 9880 14188 9908
rect 12713 9871 12771 9877
rect 14182 9868 14188 9880
rect 14240 9868 14246 9920
rect 15654 9868 15660 9920
rect 15712 9908 15718 9920
rect 16025 9911 16083 9917
rect 16025 9908 16037 9911
rect 15712 9880 16037 9908
rect 15712 9868 15718 9880
rect 16025 9877 16037 9880
rect 16071 9877 16083 9911
rect 16025 9871 16083 9877
rect 19705 9911 19763 9917
rect 19705 9877 19717 9911
rect 19751 9908 19763 9911
rect 21082 9908 21088 9920
rect 19751 9880 21088 9908
rect 19751 9877 19763 9880
rect 19705 9871 19763 9877
rect 21082 9868 21088 9880
rect 21140 9868 21146 9920
rect 21910 9908 21916 9920
rect 21871 9880 21916 9908
rect 21910 9868 21916 9880
rect 21968 9868 21974 9920
rect 26602 9868 26608 9920
rect 26660 9908 26666 9920
rect 26697 9911 26755 9917
rect 26697 9908 26709 9911
rect 26660 9880 26709 9908
rect 26660 9868 26666 9880
rect 26697 9877 26709 9880
rect 26743 9877 26755 9911
rect 26697 9871 26755 9877
rect 1104 9818 48852 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 48852 9818
rect 1104 9744 48852 9766
rect 8386 9664 8392 9716
rect 8444 9704 8450 9716
rect 8481 9707 8539 9713
rect 8481 9704 8493 9707
rect 8444 9676 8493 9704
rect 8444 9664 8450 9676
rect 8481 9673 8493 9676
rect 8527 9673 8539 9707
rect 8481 9667 8539 9673
rect 10505 9707 10563 9713
rect 10505 9673 10517 9707
rect 10551 9704 10563 9707
rect 10686 9704 10692 9716
rect 10551 9676 10692 9704
rect 10551 9673 10563 9676
rect 10505 9667 10563 9673
rect 10686 9664 10692 9676
rect 10744 9664 10750 9716
rect 14829 9707 14887 9713
rect 14829 9673 14841 9707
rect 14875 9704 14887 9707
rect 15194 9704 15200 9716
rect 14875 9676 15200 9704
rect 14875 9673 14887 9676
rect 14829 9667 14887 9673
rect 13630 9636 13636 9648
rect 13591 9608 13636 9636
rect 13630 9596 13636 9608
rect 13688 9596 13694 9648
rect 8757 9571 8815 9577
rect 8757 9537 8769 9571
rect 8803 9568 8815 9571
rect 13725 9571 13783 9577
rect 8803 9540 11376 9568
rect 8803 9537 8815 9540
rect 8757 9531 8815 9537
rect 8272 9503 8330 9509
rect 8272 9469 8284 9503
rect 8318 9500 8330 9503
rect 8772 9500 8800 9531
rect 8318 9472 8800 9500
rect 9401 9503 9459 9509
rect 8318 9469 8330 9472
rect 8272 9463 8330 9469
rect 9401 9469 9413 9503
rect 9447 9500 9459 9503
rect 10045 9503 10103 9509
rect 10045 9500 10057 9503
rect 9447 9472 10057 9500
rect 9447 9469 9459 9472
rect 9401 9463 9459 9469
rect 9125 9435 9183 9441
rect 9125 9401 9137 9435
rect 9171 9432 9183 9435
rect 9214 9432 9220 9444
rect 9171 9404 9220 9432
rect 9171 9401 9183 9404
rect 9125 9395 9183 9401
rect 9214 9392 9220 9404
rect 9272 9392 9278 9444
rect 9766 9432 9772 9444
rect 9727 9404 9772 9432
rect 9766 9392 9772 9404
rect 9824 9392 9830 9444
rect 9876 9364 9904 9472
rect 10045 9469 10057 9472
rect 10091 9469 10103 9503
rect 10045 9463 10103 9469
rect 11348 9444 11376 9540
rect 13725 9537 13737 9571
rect 13771 9568 13783 9571
rect 14844 9568 14872 9667
rect 15194 9664 15200 9676
rect 15252 9664 15258 9716
rect 17037 9707 17095 9713
rect 17037 9704 17049 9707
rect 15810 9676 17049 9704
rect 15654 9596 15660 9648
rect 15712 9636 15718 9648
rect 15810 9645 15838 9676
rect 17037 9673 17049 9676
rect 17083 9673 17095 9707
rect 17037 9667 17095 9673
rect 17497 9707 17555 9713
rect 17497 9673 17509 9707
rect 17543 9704 17555 9707
rect 17678 9704 17684 9716
rect 17543 9676 17684 9704
rect 17543 9673 17555 9676
rect 17497 9667 17555 9673
rect 17678 9664 17684 9676
rect 17736 9664 17742 9716
rect 18046 9664 18052 9716
rect 18104 9704 18110 9716
rect 18325 9707 18383 9713
rect 18325 9704 18337 9707
rect 18104 9676 18337 9704
rect 18104 9664 18110 9676
rect 18325 9673 18337 9676
rect 18371 9673 18383 9707
rect 20898 9704 20904 9716
rect 20859 9676 20904 9704
rect 18325 9667 18383 9673
rect 20898 9664 20904 9676
rect 20956 9664 20962 9716
rect 21269 9707 21327 9713
rect 21269 9673 21281 9707
rect 21315 9704 21327 9707
rect 21726 9704 21732 9716
rect 21315 9676 21732 9704
rect 21315 9673 21327 9676
rect 21269 9667 21327 9673
rect 21726 9664 21732 9676
rect 21784 9704 21790 9716
rect 22554 9704 22560 9716
rect 21784 9676 22560 9704
rect 21784 9664 21790 9676
rect 22554 9664 22560 9676
rect 22612 9664 22618 9716
rect 24302 9664 24308 9716
rect 24360 9704 24366 9716
rect 25133 9707 25191 9713
rect 25133 9704 25145 9707
rect 24360 9676 25145 9704
rect 24360 9664 24366 9676
rect 25133 9673 25145 9676
rect 25179 9673 25191 9707
rect 25133 9667 25191 9673
rect 27249 9707 27307 9713
rect 27249 9673 27261 9707
rect 27295 9704 27307 9707
rect 27338 9704 27344 9716
rect 27295 9676 27344 9704
rect 27295 9673 27307 9676
rect 27249 9667 27307 9673
rect 27338 9664 27344 9676
rect 27396 9664 27402 9716
rect 28718 9704 28724 9716
rect 28679 9676 28724 9704
rect 28718 9664 28724 9676
rect 28776 9664 28782 9716
rect 29549 9707 29607 9713
rect 29549 9673 29561 9707
rect 29595 9704 29607 9707
rect 30282 9704 30288 9716
rect 29595 9676 30288 9704
rect 29595 9673 29607 9676
rect 29549 9667 29607 9673
rect 15795 9639 15853 9645
rect 15795 9636 15807 9639
rect 15712 9608 15807 9636
rect 15712 9596 15718 9608
rect 15795 9605 15807 9608
rect 15841 9605 15853 9639
rect 15930 9636 15936 9648
rect 15891 9608 15936 9636
rect 15795 9599 15853 9605
rect 15930 9596 15936 9608
rect 15988 9596 15994 9648
rect 16114 9636 16120 9648
rect 16075 9608 16120 9636
rect 16114 9596 16120 9608
rect 16172 9636 16178 9648
rect 16172 9608 19840 9636
rect 16172 9596 16178 9608
rect 13771 9540 14872 9568
rect 15672 9540 15884 9568
rect 13771 9537 13783 9540
rect 13725 9531 13783 9537
rect 13504 9503 13562 9509
rect 13504 9469 13516 9503
rect 13550 9469 13562 9503
rect 14090 9500 14096 9512
rect 14003 9472 14096 9500
rect 13504 9463 13562 9469
rect 9950 9392 9956 9444
rect 10008 9432 10014 9444
rect 10689 9435 10747 9441
rect 10689 9432 10701 9435
rect 10008 9404 10701 9432
rect 10008 9392 10014 9404
rect 10689 9401 10701 9404
rect 10735 9401 10747 9435
rect 10689 9395 10747 9401
rect 10781 9435 10839 9441
rect 10781 9401 10793 9435
rect 10827 9432 10839 9435
rect 10870 9432 10876 9444
rect 10827 9404 10876 9432
rect 10827 9401 10839 9404
rect 10781 9395 10839 9401
rect 10870 9392 10876 9404
rect 10928 9392 10934 9444
rect 11330 9432 11336 9444
rect 11291 9404 11336 9432
rect 11330 9392 11336 9404
rect 11388 9392 11394 9444
rect 13354 9432 13360 9444
rect 13315 9404 13360 9432
rect 13354 9392 13360 9404
rect 13412 9392 13418 9444
rect 11885 9367 11943 9373
rect 11885 9364 11897 9367
rect 9876 9336 11897 9364
rect 11885 9333 11897 9336
rect 11931 9364 11943 9367
rect 12066 9364 12072 9376
rect 11931 9336 12072 9364
rect 11931 9333 11943 9336
rect 11885 9327 11943 9333
rect 12066 9324 12072 9336
rect 12124 9324 12130 9376
rect 12897 9367 12955 9373
rect 12897 9333 12909 9367
rect 12943 9364 12955 9367
rect 13262 9364 13268 9376
rect 12943 9336 13268 9364
rect 12943 9333 12955 9336
rect 12897 9327 12955 9333
rect 13262 9324 13268 9336
rect 13320 9364 13326 9376
rect 13519 9364 13547 9463
rect 14090 9460 14096 9472
rect 14148 9500 14154 9512
rect 15672 9500 15700 9540
rect 14148 9472 15700 9500
rect 14148 9460 14154 9472
rect 15657 9435 15715 9441
rect 15657 9401 15669 9435
rect 15703 9401 15715 9435
rect 15856 9432 15884 9540
rect 16022 9528 16028 9580
rect 16080 9568 16086 9580
rect 18874 9568 18880 9580
rect 16080 9540 16125 9568
rect 18064 9540 18880 9568
rect 16080 9528 16086 9540
rect 16666 9460 16672 9512
rect 16724 9500 16730 9512
rect 18064 9509 18092 9540
rect 18874 9528 18880 9540
rect 18932 9528 18938 9580
rect 19812 9568 19840 9608
rect 20254 9568 20260 9580
rect 19812 9540 20260 9568
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 16724 9472 18061 9500
rect 16724 9460 16730 9472
rect 18049 9469 18061 9472
rect 18095 9469 18107 9503
rect 18230 9500 18236 9512
rect 18191 9472 18236 9500
rect 18049 9463 18107 9469
rect 18230 9460 18236 9472
rect 18288 9500 18294 9512
rect 19812 9509 19840 9540
rect 20254 9528 20260 9540
rect 20312 9528 20318 9580
rect 20533 9571 20591 9577
rect 20533 9537 20545 9571
rect 20579 9568 20591 9571
rect 21361 9571 21419 9577
rect 21361 9568 21373 9571
rect 20579 9540 21373 9568
rect 20579 9537 20591 9540
rect 20533 9531 20591 9537
rect 21361 9537 21373 9540
rect 21407 9568 21419 9571
rect 21910 9568 21916 9580
rect 21407 9540 21916 9568
rect 21407 9537 21419 9540
rect 21361 9531 21419 9537
rect 21910 9528 21916 9540
rect 21968 9528 21974 9580
rect 23382 9528 23388 9580
rect 23440 9568 23446 9580
rect 24213 9571 24271 9577
rect 24213 9568 24225 9571
rect 23440 9540 24225 9568
rect 23440 9528 23446 9540
rect 24213 9537 24225 9540
rect 24259 9537 24271 9571
rect 28353 9571 28411 9577
rect 28353 9568 28365 9571
rect 24213 9531 24271 9537
rect 26620 9540 28365 9568
rect 26620 9512 26648 9540
rect 28353 9537 28365 9540
rect 28399 9537 28411 9571
rect 28353 9531 28411 9537
rect 19797 9503 19855 9509
rect 18288 9472 19334 9500
rect 18288 9460 18294 9472
rect 19306 9432 19334 9472
rect 19797 9469 19809 9503
rect 19843 9469 19855 9503
rect 19797 9463 19855 9469
rect 19978 9460 19984 9512
rect 20036 9500 20042 9512
rect 20349 9503 20407 9509
rect 20349 9500 20361 9503
rect 20036 9472 20361 9500
rect 20036 9460 20042 9472
rect 20349 9469 20361 9472
rect 20395 9500 20407 9503
rect 20898 9500 20904 9512
rect 20395 9472 20904 9500
rect 20395 9469 20407 9472
rect 20349 9463 20407 9469
rect 20898 9460 20904 9472
rect 20956 9460 20962 9512
rect 23106 9500 23112 9512
rect 21238 9472 23112 9500
rect 19521 9435 19579 9441
rect 19521 9432 19533 9435
rect 15856 9404 19012 9432
rect 19306 9404 19533 9432
rect 15657 9395 15715 9401
rect 13320 9336 13547 9364
rect 13320 9324 13326 9336
rect 14090 9324 14096 9376
rect 14148 9364 14154 9376
rect 14369 9367 14427 9373
rect 14369 9364 14381 9367
rect 14148 9336 14381 9364
rect 14148 9324 14154 9336
rect 14369 9333 14381 9336
rect 14415 9333 14427 9367
rect 15102 9364 15108 9376
rect 15063 9336 15108 9364
rect 14369 9327 14427 9333
rect 15102 9324 15108 9336
rect 15160 9324 15166 9376
rect 15470 9364 15476 9376
rect 15431 9336 15476 9364
rect 15470 9324 15476 9336
rect 15528 9364 15534 9376
rect 15672 9364 15700 9395
rect 15528 9336 15700 9364
rect 15528 9324 15534 9336
rect 15930 9324 15936 9376
rect 15988 9364 15994 9376
rect 16669 9367 16727 9373
rect 16669 9364 16681 9367
rect 15988 9336 16681 9364
rect 15988 9324 15994 9336
rect 16669 9333 16681 9336
rect 16715 9364 16727 9367
rect 17773 9367 17831 9373
rect 17773 9364 17785 9367
rect 16715 9336 17785 9364
rect 16715 9333 16727 9336
rect 16669 9327 16727 9333
rect 17773 9333 17785 9336
rect 17819 9364 17831 9367
rect 18230 9364 18236 9376
rect 17819 9336 18236 9364
rect 17819 9333 17831 9336
rect 17773 9327 17831 9333
rect 18230 9324 18236 9336
rect 18288 9364 18294 9376
rect 18877 9367 18935 9373
rect 18877 9364 18889 9367
rect 18288 9336 18889 9364
rect 18288 9324 18294 9336
rect 18877 9333 18889 9336
rect 18923 9333 18935 9367
rect 18984 9364 19012 9404
rect 19521 9401 19533 9404
rect 19567 9432 19579 9435
rect 19610 9432 19616 9444
rect 19567 9404 19616 9432
rect 19567 9401 19579 9404
rect 19521 9395 19579 9401
rect 19610 9392 19616 9404
rect 19668 9432 19674 9444
rect 21238 9432 21266 9472
rect 23106 9460 23112 9472
rect 23164 9460 23170 9512
rect 25958 9500 25964 9512
rect 25919 9472 25964 9500
rect 25958 9460 25964 9472
rect 26016 9500 26022 9512
rect 26145 9503 26203 9509
rect 26145 9500 26157 9503
rect 26016 9472 26157 9500
rect 26016 9460 26022 9472
rect 26145 9469 26157 9472
rect 26191 9469 26203 9503
rect 26602 9500 26608 9512
rect 26563 9472 26608 9500
rect 26145 9463 26203 9469
rect 26602 9460 26608 9472
rect 26660 9460 26666 9512
rect 27744 9503 27802 9509
rect 27744 9500 27756 9503
rect 27632 9472 27756 9500
rect 19668 9404 21266 9432
rect 19668 9392 19674 9404
rect 22094 9392 22100 9444
rect 22152 9432 22158 9444
rect 22925 9435 22983 9441
rect 22925 9432 22937 9435
rect 22152 9404 22937 9432
rect 22152 9392 22158 9404
rect 22925 9401 22937 9404
rect 22971 9401 22983 9435
rect 22925 9395 22983 9401
rect 24305 9435 24363 9441
rect 24305 9401 24317 9435
rect 24351 9401 24363 9435
rect 24854 9432 24860 9444
rect 24815 9404 24860 9432
rect 24305 9395 24363 9401
rect 20990 9364 20996 9376
rect 18984 9336 20996 9364
rect 18877 9327 18935 9333
rect 20990 9324 20996 9336
rect 21048 9324 21054 9376
rect 21726 9364 21732 9376
rect 21687 9336 21732 9364
rect 21726 9324 21732 9336
rect 21784 9324 21790 9376
rect 21818 9324 21824 9376
rect 21876 9364 21882 9376
rect 22281 9367 22339 9373
rect 22281 9364 22293 9367
rect 21876 9336 22293 9364
rect 21876 9324 21882 9336
rect 22281 9333 22293 9336
rect 22327 9333 22339 9367
rect 22281 9327 22339 9333
rect 23474 9324 23480 9376
rect 23532 9364 23538 9376
rect 24029 9367 24087 9373
rect 23532 9336 23577 9364
rect 23532 9324 23538 9336
rect 24029 9333 24041 9367
rect 24075 9364 24087 9367
rect 24320 9364 24348 9395
rect 24854 9392 24860 9404
rect 24912 9392 24918 9444
rect 26878 9432 26884 9444
rect 26839 9404 26884 9432
rect 26878 9392 26884 9404
rect 26936 9392 26942 9444
rect 27632 9376 27660 9472
rect 27744 9469 27756 9472
rect 27790 9469 27802 9503
rect 29638 9500 29644 9512
rect 29599 9472 29644 9500
rect 27744 9463 27802 9469
rect 29638 9460 29644 9472
rect 29696 9460 29702 9512
rect 30018 9441 30046 9676
rect 30282 9664 30288 9676
rect 30340 9704 30346 9716
rect 30926 9704 30932 9716
rect 30340 9676 30932 9704
rect 30340 9664 30346 9676
rect 30926 9664 30932 9676
rect 30984 9664 30990 9716
rect 31202 9704 31208 9716
rect 31163 9676 31208 9704
rect 31202 9664 31208 9676
rect 31260 9664 31266 9716
rect 33502 9664 33508 9716
rect 33560 9704 33566 9716
rect 33919 9707 33977 9713
rect 33919 9704 33931 9707
rect 33560 9676 33931 9704
rect 33560 9664 33566 9676
rect 33919 9673 33931 9676
rect 33965 9673 33977 9707
rect 34330 9704 34336 9716
rect 34291 9676 34336 9704
rect 33919 9667 33977 9673
rect 34330 9664 34336 9676
rect 34388 9704 34394 9716
rect 34609 9707 34667 9713
rect 34609 9704 34621 9707
rect 34388 9676 34621 9704
rect 34388 9664 34394 9676
rect 34609 9673 34621 9676
rect 34655 9673 34667 9707
rect 34609 9667 34667 9673
rect 32490 9596 32496 9648
rect 32548 9636 32554 9648
rect 33597 9639 33655 9645
rect 33597 9636 33609 9639
rect 32548 9608 33609 9636
rect 32548 9596 32554 9608
rect 33597 9605 33609 9608
rect 33643 9605 33655 9639
rect 33597 9599 33655 9605
rect 31478 9528 31484 9580
rect 31536 9568 31542 9580
rect 31536 9540 33859 9568
rect 31536 9528 31542 9540
rect 33831 9512 33859 9540
rect 33778 9500 33784 9512
rect 33836 9509 33859 9512
rect 33836 9503 33874 9509
rect 33726 9472 33784 9500
rect 33778 9460 33784 9472
rect 33862 9469 33874 9503
rect 33836 9463 33874 9469
rect 33836 9460 33842 9463
rect 30003 9435 30061 9441
rect 30003 9401 30015 9435
rect 30049 9401 30061 9435
rect 30003 9395 30061 9401
rect 31757 9435 31815 9441
rect 31757 9401 31769 9435
rect 31803 9432 31815 9435
rect 32122 9432 32128 9444
rect 31803 9404 32128 9432
rect 31803 9401 31815 9404
rect 31757 9395 31815 9401
rect 32122 9392 32128 9404
rect 32180 9432 32186 9444
rect 32309 9435 32367 9441
rect 32309 9432 32321 9435
rect 32180 9404 32321 9432
rect 32180 9392 32186 9404
rect 32309 9401 32321 9404
rect 32355 9401 32367 9435
rect 32309 9395 32367 9401
rect 32401 9435 32459 9441
rect 32401 9401 32413 9435
rect 32447 9432 32459 9435
rect 32766 9432 32772 9444
rect 32447 9404 32772 9432
rect 32447 9401 32459 9404
rect 32401 9395 32459 9401
rect 24394 9364 24400 9376
rect 24075 9336 24400 9364
rect 24075 9333 24087 9336
rect 24029 9327 24087 9333
rect 24394 9324 24400 9336
rect 24452 9364 24458 9376
rect 25866 9364 25872 9376
rect 24452 9336 25872 9364
rect 24452 9324 24458 9336
rect 25866 9324 25872 9336
rect 25924 9324 25930 9376
rect 27614 9364 27620 9376
rect 27575 9336 27620 9364
rect 27614 9324 27620 9336
rect 27672 9324 27678 9376
rect 27847 9367 27905 9373
rect 27847 9333 27859 9367
rect 27893 9364 27905 9367
rect 27982 9364 27988 9376
rect 27893 9336 27988 9364
rect 27893 9333 27905 9336
rect 27847 9327 27905 9333
rect 27982 9324 27988 9336
rect 28040 9324 28046 9376
rect 30558 9364 30564 9376
rect 30519 9336 30564 9364
rect 30558 9324 30564 9336
rect 30616 9324 30622 9376
rect 32033 9367 32091 9373
rect 32033 9333 32045 9367
rect 32079 9364 32091 9367
rect 32416 9364 32444 9395
rect 32766 9392 32772 9404
rect 32824 9392 32830 9444
rect 32950 9432 32956 9444
rect 32911 9404 32956 9432
rect 32950 9392 32956 9404
rect 33008 9392 33014 9444
rect 34624 9432 34652 9667
rect 36170 9664 36176 9716
rect 36228 9704 36234 9716
rect 36449 9707 36507 9713
rect 36449 9704 36461 9707
rect 36228 9676 36461 9704
rect 36228 9664 36234 9676
rect 36449 9673 36461 9676
rect 36495 9673 36507 9707
rect 36449 9667 36507 9673
rect 37826 9664 37832 9716
rect 37884 9704 37890 9716
rect 38289 9707 38347 9713
rect 38289 9704 38301 9707
rect 37884 9676 38301 9704
rect 37884 9664 37890 9676
rect 38289 9673 38301 9676
rect 38335 9673 38347 9707
rect 38289 9667 38347 9673
rect 39025 9639 39083 9645
rect 39025 9605 39037 9639
rect 39071 9605 39083 9639
rect 39025 9599 39083 9605
rect 34977 9571 35035 9577
rect 34977 9537 34989 9571
rect 35023 9568 35035 9571
rect 35250 9568 35256 9580
rect 35023 9540 35256 9568
rect 35023 9537 35035 9540
rect 34977 9531 35035 9537
rect 35250 9528 35256 9540
rect 35308 9528 35314 9580
rect 36173 9571 36231 9577
rect 36173 9537 36185 9571
rect 36219 9568 36231 9571
rect 36262 9568 36268 9580
rect 36219 9540 36268 9568
rect 36219 9537 36231 9540
rect 36173 9531 36231 9537
rect 36262 9528 36268 9540
rect 36320 9528 36326 9580
rect 39040 9568 39068 9599
rect 37936 9540 39068 9568
rect 37936 9509 37964 9540
rect 37185 9503 37243 9509
rect 37185 9469 37197 9503
rect 37231 9500 37243 9503
rect 37921 9503 37979 9509
rect 37921 9500 37933 9503
rect 37231 9472 37933 9500
rect 37231 9469 37243 9472
rect 37185 9463 37243 9469
rect 37921 9469 37933 9472
rect 37967 9469 37979 9503
rect 38838 9500 38844 9512
rect 38799 9472 38844 9500
rect 37921 9463 37979 9469
rect 38838 9460 38844 9472
rect 38896 9500 38902 9512
rect 39301 9503 39359 9509
rect 39301 9500 39313 9503
rect 38896 9472 39313 9500
rect 38896 9460 38902 9472
rect 39301 9469 39313 9472
rect 39347 9469 39359 9503
rect 39301 9463 39359 9469
rect 34698 9432 34704 9444
rect 34611 9404 34704 9432
rect 34698 9392 34704 9404
rect 34756 9432 34762 9444
rect 35066 9432 35072 9444
rect 34756 9404 35072 9432
rect 34756 9392 34762 9404
rect 35066 9392 35072 9404
rect 35124 9392 35130 9444
rect 35158 9392 35164 9444
rect 35216 9432 35222 9444
rect 35621 9435 35679 9441
rect 35621 9432 35633 9435
rect 35216 9404 35633 9432
rect 35216 9392 35222 9404
rect 35621 9401 35633 9404
rect 35667 9432 35679 9435
rect 37826 9432 37832 9444
rect 35667 9404 37832 9432
rect 35667 9401 35679 9404
rect 35621 9395 35679 9401
rect 37826 9392 37832 9404
rect 37884 9392 37890 9444
rect 32079 9336 32444 9364
rect 32784 9364 32812 9392
rect 33229 9367 33287 9373
rect 33229 9364 33241 9367
rect 32784 9336 33241 9364
rect 32079 9333 32091 9336
rect 32033 9327 32091 9333
rect 33229 9333 33241 9336
rect 33275 9333 33287 9367
rect 33229 9327 33287 9333
rect 37737 9367 37795 9373
rect 37737 9333 37749 9367
rect 37783 9364 37795 9367
rect 37918 9364 37924 9376
rect 37783 9336 37924 9364
rect 37783 9333 37795 9336
rect 37737 9327 37795 9333
rect 37918 9324 37924 9336
rect 37976 9324 37982 9376
rect 1104 9274 48852 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 48852 9274
rect 1104 9200 48852 9222
rect 8711 9163 8769 9169
rect 8711 9129 8723 9163
rect 8757 9160 8769 9163
rect 9950 9160 9956 9172
rect 8757 9132 9956 9160
rect 8757 9129 8769 9132
rect 8711 9123 8769 9129
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 10965 9163 11023 9169
rect 10965 9160 10977 9163
rect 10928 9132 10977 9160
rect 10928 9120 10934 9132
rect 10965 9129 10977 9132
rect 11011 9129 11023 9163
rect 11238 9160 11244 9172
rect 11199 9132 11244 9160
rect 10965 9123 11023 9129
rect 11238 9120 11244 9132
rect 11296 9120 11302 9172
rect 18874 9160 18880 9172
rect 18835 9132 18880 9160
rect 18874 9120 18880 9132
rect 18932 9120 18938 9172
rect 20254 9160 20260 9172
rect 20215 9132 20260 9160
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 21450 9160 21456 9172
rect 21411 9132 21456 9160
rect 21450 9120 21456 9132
rect 21508 9120 21514 9172
rect 21818 9160 21824 9172
rect 21779 9132 21824 9160
rect 21818 9120 21824 9132
rect 21876 9120 21882 9172
rect 22830 9160 22836 9172
rect 22791 9132 22836 9160
rect 22830 9120 22836 9132
rect 22888 9120 22894 9172
rect 27154 9160 27160 9172
rect 27115 9132 27160 9160
rect 27154 9120 27160 9132
rect 27212 9120 27218 9172
rect 27246 9120 27252 9172
rect 27304 9160 27310 9172
rect 27985 9163 28043 9169
rect 27985 9160 27997 9163
rect 27304 9132 27997 9160
rect 27304 9120 27310 9132
rect 27985 9129 27997 9132
rect 28031 9129 28043 9163
rect 33778 9160 33784 9172
rect 33739 9132 33784 9160
rect 27985 9123 28043 9129
rect 33778 9120 33784 9132
rect 33836 9120 33842 9172
rect 34238 9160 34244 9172
rect 34151 9132 34244 9160
rect 9858 9052 9864 9104
rect 9916 9092 9922 9104
rect 10366 9095 10424 9101
rect 10366 9092 10378 9095
rect 9916 9064 10378 9092
rect 9916 9052 9922 9064
rect 10366 9061 10378 9064
rect 10412 9061 10424 9095
rect 13998 9092 14004 9104
rect 10366 9055 10424 9061
rect 12084 9064 13768 9092
rect 13959 9064 14004 9092
rect 12084 9036 12112 9064
rect 13740 9036 13768 9064
rect 13998 9052 14004 9064
rect 14056 9052 14062 9104
rect 17862 9052 17868 9104
rect 17920 9092 17926 9104
rect 18049 9095 18107 9101
rect 18049 9092 18061 9095
rect 17920 9064 18061 9092
rect 17920 9052 17926 9064
rect 18049 9061 18061 9064
rect 18095 9092 18107 9095
rect 19334 9092 19340 9104
rect 18095 9064 19340 9092
rect 18095 9061 18107 9064
rect 18049 9055 18107 9061
rect 19334 9052 19340 9064
rect 19392 9052 19398 9104
rect 19978 9092 19984 9104
rect 19939 9064 19984 9092
rect 19978 9052 19984 9064
rect 20036 9052 20042 9104
rect 8640 9027 8698 9033
rect 8640 8993 8652 9027
rect 8686 9024 8698 9027
rect 8754 9024 8760 9036
rect 8686 8996 8760 9024
rect 8686 8993 8698 8996
rect 8640 8987 8698 8993
rect 8754 8984 8760 8996
rect 8812 8984 8818 9036
rect 11882 9024 11888 9036
rect 11843 8996 11888 9024
rect 11882 8984 11888 8996
rect 11940 8984 11946 9036
rect 12066 8984 12072 9036
rect 12124 9024 12130 9036
rect 13262 9024 13268 9036
rect 12124 8996 12217 9024
rect 13223 8996 13268 9024
rect 12124 8984 12130 8996
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 13541 9027 13599 9033
rect 13541 8993 13553 9027
rect 13587 9024 13599 9027
rect 13630 9024 13636 9036
rect 13587 8996 13636 9024
rect 13587 8993 13599 8996
rect 13541 8987 13599 8993
rect 10042 8956 10048 8968
rect 10003 8928 10048 8956
rect 10042 8916 10048 8928
rect 10100 8916 10106 8968
rect 13354 8956 13360 8968
rect 12728 8928 13360 8956
rect 8570 8848 8576 8900
rect 8628 8888 8634 8900
rect 12728 8897 12756 8928
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 12713 8891 12771 8897
rect 12713 8888 12725 8891
rect 8628 8860 12725 8888
rect 8628 8848 8634 8860
rect 12713 8857 12725 8860
rect 12759 8857 12771 8891
rect 12713 8851 12771 8857
rect 10410 8780 10416 8832
rect 10468 8820 10474 8832
rect 12161 8823 12219 8829
rect 12161 8820 12173 8823
rect 10468 8792 12173 8820
rect 10468 8780 10474 8792
rect 12161 8789 12173 8792
rect 12207 8820 12219 8823
rect 12618 8820 12624 8832
rect 12207 8792 12624 8820
rect 12207 8789 12219 8792
rect 12161 8783 12219 8789
rect 12618 8780 12624 8792
rect 12676 8780 12682 8832
rect 13170 8820 13176 8832
rect 13131 8792 13176 8820
rect 13170 8780 13176 8792
rect 13228 8820 13234 8832
rect 13556 8820 13584 8987
rect 13630 8984 13636 8996
rect 13688 8984 13694 9036
rect 13722 8984 13728 9036
rect 13780 9024 13786 9036
rect 15654 9024 15660 9036
rect 13780 8996 15660 9024
rect 13780 8984 13786 8996
rect 15654 8984 15660 8996
rect 15712 8984 15718 9036
rect 15838 8984 15844 9036
rect 15896 9033 15902 9036
rect 15896 9027 15945 9033
rect 15896 8993 15899 9027
rect 15933 8993 15945 9027
rect 18230 9024 18236 9036
rect 18191 8996 18236 9024
rect 15896 8987 15945 8993
rect 15896 8984 15902 8987
rect 18230 8984 18236 8996
rect 18288 8984 18294 9036
rect 19150 8984 19156 9036
rect 19208 9024 19214 9036
rect 19429 9027 19487 9033
rect 19429 9024 19441 9027
rect 19208 8996 19441 9024
rect 19208 8984 19214 8996
rect 19429 8993 19441 8996
rect 19475 8993 19487 9027
rect 19429 8987 19487 8993
rect 19613 9027 19671 9033
rect 19613 8993 19625 9027
rect 19659 9024 19671 9027
rect 19886 9024 19892 9036
rect 19659 8996 19892 9024
rect 19659 8993 19671 8996
rect 19613 8987 19671 8993
rect 19886 8984 19892 8996
rect 19944 8984 19950 9036
rect 20968 9027 21026 9033
rect 20968 8993 20980 9027
rect 21014 9024 21026 9027
rect 21836 9024 21864 9120
rect 22278 9101 22284 9104
rect 22275 9092 22284 9101
rect 22191 9064 22284 9092
rect 22275 9055 22284 9064
rect 22336 9092 22342 9104
rect 22554 9092 22560 9104
rect 22336 9064 22560 9092
rect 22278 9052 22284 9055
rect 22336 9052 22342 9064
rect 22554 9052 22560 9064
rect 22612 9052 22618 9104
rect 24302 9092 24308 9104
rect 24263 9064 24308 9092
rect 24302 9052 24308 9064
rect 24360 9052 24366 9104
rect 29365 9095 29423 9101
rect 29365 9061 29377 9095
rect 29411 9092 29423 9095
rect 29638 9092 29644 9104
rect 29411 9064 29644 9092
rect 29411 9061 29423 9064
rect 29365 9055 29423 9061
rect 29638 9052 29644 9064
rect 29696 9052 29702 9104
rect 32309 9095 32367 9101
rect 32309 9061 32321 9095
rect 32355 9092 32367 9095
rect 32582 9092 32588 9104
rect 32355 9064 32588 9092
rect 32355 9061 32367 9064
rect 32309 9055 32367 9061
rect 32582 9052 32588 9064
rect 32640 9052 32646 9104
rect 32861 9095 32919 9101
rect 32861 9061 32873 9095
rect 32907 9092 32919 9095
rect 32950 9092 32956 9104
rect 32907 9064 32956 9092
rect 32907 9061 32919 9064
rect 32861 9055 32919 9061
rect 32950 9052 32956 9064
rect 33008 9092 33014 9104
rect 34164 9101 34192 9132
rect 34238 9120 34244 9132
rect 34296 9160 34302 9172
rect 34606 9160 34612 9172
rect 34296 9132 34612 9160
rect 34296 9120 34302 9132
rect 34606 9120 34612 9132
rect 34664 9120 34670 9172
rect 34149 9095 34207 9101
rect 33008 9064 33134 9092
rect 33008 9052 33014 9064
rect 21014 8996 21864 9024
rect 26789 9027 26847 9033
rect 21014 8993 21026 8996
rect 20968 8987 21026 8993
rect 26789 8993 26801 9027
rect 26835 9024 26847 9027
rect 26878 9024 26884 9036
rect 26835 8996 26884 9024
rect 26835 8993 26847 8996
rect 26789 8987 26847 8993
rect 26878 8984 26884 8996
rect 26936 8984 26942 9036
rect 26970 8984 26976 9036
rect 27028 9024 27034 9036
rect 28626 9024 28632 9036
rect 27028 8996 28632 9024
rect 27028 8984 27034 8996
rect 28626 8984 28632 8996
rect 28684 8984 28690 9036
rect 28994 8984 29000 9036
rect 29052 9024 29058 9036
rect 29089 9027 29147 9033
rect 29089 9024 29101 9027
rect 29052 8996 29101 9024
rect 29052 8984 29058 8996
rect 29089 8993 29101 8996
rect 29135 8993 29147 9027
rect 29089 8987 29147 8993
rect 30193 9027 30251 9033
rect 30193 8993 30205 9027
rect 30239 8993 30251 9027
rect 30650 9024 30656 9036
rect 30611 8996 30656 9024
rect 30193 8987 30251 8993
rect 14182 8916 14188 8968
rect 14240 8956 14246 8968
rect 16117 8959 16175 8965
rect 16117 8956 16129 8959
rect 14240 8928 16129 8956
rect 14240 8916 14246 8928
rect 16117 8925 16129 8928
rect 16163 8956 16175 8959
rect 16574 8956 16580 8968
rect 16163 8928 16580 8956
rect 16163 8925 16175 8928
rect 16117 8919 16175 8925
rect 16574 8916 16580 8928
rect 16632 8916 16638 8968
rect 21542 8916 21548 8968
rect 21600 8956 21606 8968
rect 21913 8959 21971 8965
rect 21913 8956 21925 8959
rect 21600 8928 21925 8956
rect 21600 8916 21606 8928
rect 21913 8925 21925 8928
rect 21959 8956 21971 8959
rect 22554 8956 22560 8968
rect 21959 8928 22560 8956
rect 21959 8925 21971 8928
rect 21913 8919 21971 8925
rect 22554 8916 22560 8928
rect 22612 8916 22618 8968
rect 24210 8956 24216 8968
rect 23446 8928 24216 8956
rect 15749 8891 15807 8897
rect 15749 8857 15761 8891
rect 15795 8857 15807 8891
rect 15749 8851 15807 8857
rect 21039 8891 21097 8897
rect 21039 8857 21051 8891
rect 21085 8888 21097 8891
rect 23446 8888 23474 8928
rect 24210 8916 24216 8928
rect 24268 8916 24274 8968
rect 24857 8959 24915 8965
rect 24857 8925 24869 8959
rect 24903 8956 24915 8959
rect 24946 8956 24952 8968
rect 24903 8928 24952 8956
rect 24903 8925 24915 8928
rect 24857 8919 24915 8925
rect 24946 8916 24952 8928
rect 25004 8916 25010 8968
rect 28718 8916 28724 8968
rect 28776 8956 28782 8968
rect 29914 8956 29920 8968
rect 28776 8928 29920 8956
rect 28776 8916 28782 8928
rect 29914 8916 29920 8928
rect 29972 8956 29978 8968
rect 30208 8956 30236 8987
rect 30650 8984 30656 8996
rect 30708 8984 30714 9036
rect 30926 8956 30932 8968
rect 29972 8928 30236 8956
rect 30887 8928 30932 8956
rect 29972 8916 29978 8928
rect 30926 8916 30932 8928
rect 30984 8916 30990 8968
rect 31754 8916 31760 8968
rect 31812 8956 31818 8968
rect 32217 8959 32275 8965
rect 32217 8956 32229 8959
rect 31812 8928 32229 8956
rect 31812 8916 31818 8928
rect 32217 8925 32229 8928
rect 32263 8925 32275 8959
rect 33106 8956 33134 9064
rect 34149 9061 34161 9095
rect 34195 9061 34207 9095
rect 34149 9055 34207 9061
rect 35066 9052 35072 9104
rect 35124 9092 35130 9104
rect 35713 9095 35771 9101
rect 35713 9092 35725 9095
rect 35124 9064 35725 9092
rect 35124 9052 35130 9064
rect 35713 9061 35725 9064
rect 35759 9061 35771 9095
rect 37918 9092 37924 9104
rect 37879 9064 37924 9092
rect 35713 9055 35771 9061
rect 37918 9052 37924 9064
rect 37976 9052 37982 9104
rect 34701 9027 34759 9033
rect 34701 8993 34713 9027
rect 34747 9024 34759 9027
rect 35158 9024 35164 9036
rect 34747 8996 35164 9024
rect 34747 8993 34759 8996
rect 34701 8987 34759 8993
rect 35158 8984 35164 8996
rect 35216 8984 35222 9036
rect 34054 8956 34060 8968
rect 33106 8928 34060 8956
rect 32217 8919 32275 8925
rect 34054 8916 34060 8928
rect 34112 8916 34118 8968
rect 35621 8959 35679 8965
rect 35621 8925 35633 8959
rect 35667 8925 35679 8959
rect 35621 8919 35679 8925
rect 21085 8860 23474 8888
rect 21085 8857 21097 8860
rect 21039 8851 21097 8857
rect 13228 8792 13584 8820
rect 13228 8780 13234 8792
rect 14274 8780 14280 8832
rect 14332 8820 14338 8832
rect 15473 8823 15531 8829
rect 15473 8820 15485 8823
rect 14332 8792 15485 8820
rect 14332 8780 14338 8792
rect 15473 8789 15485 8792
rect 15519 8820 15531 8823
rect 15562 8820 15568 8832
rect 15519 8792 15568 8820
rect 15519 8789 15531 8792
rect 15473 8783 15531 8789
rect 15562 8780 15568 8792
rect 15620 8820 15626 8832
rect 15764 8820 15792 8851
rect 35526 8848 35532 8900
rect 35584 8888 35590 8900
rect 35636 8888 35664 8919
rect 35802 8916 35808 8968
rect 35860 8956 35866 8968
rect 35897 8959 35955 8965
rect 35897 8956 35909 8959
rect 35860 8928 35909 8956
rect 35860 8916 35866 8928
rect 35897 8925 35909 8928
rect 35943 8925 35955 8959
rect 37826 8956 37832 8968
rect 37787 8928 37832 8956
rect 35897 8919 35955 8925
rect 37826 8916 37832 8928
rect 37884 8916 37890 8968
rect 38102 8956 38108 8968
rect 38063 8928 38108 8956
rect 38102 8916 38108 8928
rect 38160 8916 38166 8968
rect 35584 8860 35664 8888
rect 35584 8848 35590 8860
rect 15620 8792 15792 8820
rect 15620 8780 15626 8792
rect 16022 8780 16028 8832
rect 16080 8820 16086 8832
rect 18325 8823 18383 8829
rect 18325 8820 18337 8823
rect 16080 8792 18337 8820
rect 16080 8780 16086 8792
rect 18325 8789 18337 8792
rect 18371 8789 18383 8823
rect 18325 8783 18383 8789
rect 23934 8780 23940 8832
rect 23992 8820 23998 8832
rect 26145 8823 26203 8829
rect 26145 8820 26157 8823
rect 23992 8792 26157 8820
rect 23992 8780 23998 8792
rect 26145 8789 26157 8792
rect 26191 8820 26203 8823
rect 26602 8820 26608 8832
rect 26191 8792 26608 8820
rect 26191 8789 26203 8792
rect 26145 8783 26203 8789
rect 26602 8780 26608 8792
rect 26660 8780 26666 8832
rect 27709 8823 27767 8829
rect 27709 8789 27721 8823
rect 27755 8820 27767 8823
rect 27890 8820 27896 8832
rect 27755 8792 27896 8820
rect 27755 8789 27767 8792
rect 27709 8783 27767 8789
rect 27890 8780 27896 8792
rect 27948 8780 27954 8832
rect 34790 8780 34796 8832
rect 34848 8820 34854 8832
rect 34977 8823 35035 8829
rect 34977 8820 34989 8823
rect 34848 8792 34989 8820
rect 34848 8780 34854 8792
rect 34977 8789 34989 8792
rect 35023 8789 35035 8823
rect 36538 8820 36544 8832
rect 36499 8792 36544 8820
rect 34977 8783 35035 8789
rect 36538 8780 36544 8792
rect 36596 8780 36602 8832
rect 1104 8730 48852 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 48852 8730
rect 1104 8656 48852 8678
rect 8665 8619 8723 8625
rect 8665 8585 8677 8619
rect 8711 8616 8723 8619
rect 8754 8616 8760 8628
rect 8711 8588 8760 8616
rect 8711 8585 8723 8588
rect 8665 8579 8723 8585
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 11609 8619 11667 8625
rect 11609 8585 11621 8619
rect 11655 8616 11667 8619
rect 12066 8616 12072 8628
rect 11655 8588 12072 8616
rect 11655 8585 11667 8588
rect 11609 8579 11667 8585
rect 12066 8576 12072 8588
rect 12124 8576 12130 8628
rect 13354 8576 13360 8628
rect 13412 8616 13418 8628
rect 14274 8616 14280 8628
rect 13412 8588 14280 8616
rect 13412 8576 13418 8588
rect 14274 8576 14280 8588
rect 14332 8576 14338 8628
rect 17862 8616 17868 8628
rect 17823 8588 17868 8616
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 19150 8576 19156 8628
rect 19208 8616 19214 8628
rect 19981 8619 20039 8625
rect 19981 8616 19993 8619
rect 19208 8588 19993 8616
rect 19208 8576 19214 8588
rect 19981 8585 19993 8588
rect 20027 8616 20039 8619
rect 20530 8616 20536 8628
rect 20027 8588 20536 8616
rect 20027 8585 20039 8588
rect 19981 8579 20039 8585
rect 20530 8576 20536 8588
rect 20588 8576 20594 8628
rect 20717 8619 20775 8625
rect 20717 8585 20729 8619
rect 20763 8616 20775 8619
rect 20898 8616 20904 8628
rect 20763 8588 20904 8616
rect 20763 8585 20775 8588
rect 20717 8579 20775 8585
rect 20898 8576 20904 8588
rect 20956 8576 20962 8628
rect 22278 8616 22284 8628
rect 22239 8588 22284 8616
rect 22278 8576 22284 8588
rect 22336 8576 22342 8628
rect 22554 8616 22560 8628
rect 22515 8588 22560 8616
rect 22554 8576 22560 8588
rect 22612 8576 22618 8628
rect 24210 8576 24216 8628
rect 24268 8616 24274 8628
rect 25133 8619 25191 8625
rect 25133 8616 25145 8619
rect 24268 8588 25145 8616
rect 24268 8576 24274 8588
rect 25133 8585 25145 8588
rect 25179 8585 25191 8619
rect 25133 8579 25191 8585
rect 25593 8619 25651 8625
rect 25593 8585 25605 8619
rect 25639 8616 25651 8619
rect 25866 8616 25872 8628
rect 25639 8588 25872 8616
rect 25639 8585 25651 8588
rect 25593 8579 25651 8585
rect 25866 8576 25872 8588
rect 25924 8616 25930 8628
rect 27338 8616 27344 8628
rect 25924 8588 27344 8616
rect 25924 8576 25930 8588
rect 27338 8576 27344 8588
rect 27396 8616 27402 8628
rect 27433 8619 27491 8625
rect 27433 8616 27445 8619
rect 27396 8588 27445 8616
rect 27396 8576 27402 8588
rect 27433 8585 27445 8588
rect 27479 8585 27491 8619
rect 28626 8616 28632 8628
rect 28587 8588 28632 8616
rect 27433 8579 27491 8585
rect 28626 8576 28632 8588
rect 28684 8576 28690 8628
rect 29914 8616 29920 8628
rect 29875 8588 29920 8616
rect 29914 8576 29920 8588
rect 29972 8576 29978 8628
rect 30282 8616 30288 8628
rect 30243 8588 30288 8616
rect 30282 8576 30288 8588
rect 30340 8576 30346 8628
rect 31754 8616 31760 8628
rect 31715 8588 31760 8616
rect 31754 8576 31760 8588
rect 31812 8576 31818 8628
rect 32582 8576 32588 8628
rect 32640 8616 32646 8628
rect 32677 8619 32735 8625
rect 32677 8616 32689 8619
rect 32640 8588 32689 8616
rect 32640 8576 32646 8588
rect 32677 8585 32689 8588
rect 32723 8585 32735 8619
rect 34238 8616 34244 8628
rect 34199 8588 34244 8616
rect 32677 8579 32735 8585
rect 34238 8576 34244 8588
rect 34296 8576 34302 8628
rect 34698 8616 34704 8628
rect 34659 8588 34704 8616
rect 34698 8576 34704 8588
rect 34756 8616 34762 8628
rect 35897 8619 35955 8625
rect 35897 8616 35909 8619
rect 34756 8588 35909 8616
rect 34756 8576 34762 8588
rect 35897 8585 35909 8588
rect 35943 8585 35955 8619
rect 36262 8616 36268 8628
rect 36223 8588 36268 8616
rect 35897 8579 35955 8585
rect 36262 8576 36268 8588
rect 36320 8576 36326 8628
rect 37826 8576 37832 8628
rect 37884 8616 37890 8628
rect 38841 8619 38899 8625
rect 38841 8616 38853 8619
rect 37884 8588 38853 8616
rect 37884 8576 37890 8588
rect 38841 8585 38853 8588
rect 38887 8585 38899 8619
rect 38841 8579 38899 8585
rect 15654 8508 15660 8560
rect 15712 8548 15718 8560
rect 16025 8551 16083 8557
rect 16025 8548 16037 8551
rect 15712 8520 16037 8548
rect 15712 8508 15718 8520
rect 16025 8517 16037 8520
rect 16071 8548 16083 8551
rect 16206 8548 16212 8560
rect 16071 8520 16212 8548
rect 16071 8517 16083 8520
rect 16025 8511 16083 8517
rect 16206 8508 16212 8520
rect 16264 8548 16270 8560
rect 16945 8551 17003 8557
rect 16945 8548 16957 8551
rect 16264 8520 16957 8548
rect 16264 8508 16270 8520
rect 16945 8517 16957 8520
rect 16991 8548 17003 8551
rect 17313 8551 17371 8557
rect 17313 8548 17325 8551
rect 16991 8520 17325 8548
rect 16991 8517 17003 8520
rect 16945 8511 17003 8517
rect 17313 8517 17325 8520
rect 17359 8517 17371 8551
rect 17313 8511 17371 8517
rect 9585 8483 9643 8489
rect 9585 8449 9597 8483
rect 9631 8480 9643 8483
rect 12805 8483 12863 8489
rect 9631 8452 10548 8480
rect 9631 8449 9643 8452
rect 9585 8443 9643 8449
rect 10520 8424 10548 8452
rect 12805 8449 12817 8483
rect 12851 8480 12863 8483
rect 13170 8480 13176 8492
rect 12851 8452 13176 8480
rect 12851 8449 12863 8452
rect 12805 8443 12863 8449
rect 13170 8440 13176 8452
rect 13228 8480 13234 8492
rect 13265 8483 13323 8489
rect 13265 8480 13277 8483
rect 13228 8452 13277 8480
rect 13228 8440 13234 8452
rect 13265 8449 13277 8452
rect 13311 8480 13323 8483
rect 15013 8483 15071 8489
rect 15013 8480 15025 8483
rect 13311 8452 15025 8480
rect 13311 8449 13323 8452
rect 13265 8443 13323 8449
rect 15013 8449 15025 8452
rect 15059 8480 15071 8483
rect 15102 8480 15108 8492
rect 15059 8452 15108 8480
rect 15059 8449 15071 8452
rect 15013 8443 15071 8449
rect 15102 8440 15108 8452
rect 15160 8480 15166 8492
rect 15381 8483 15439 8489
rect 15381 8480 15393 8483
rect 15160 8452 15393 8480
rect 15160 8440 15166 8452
rect 15381 8449 15393 8452
rect 15427 8480 15439 8483
rect 15838 8480 15844 8492
rect 15427 8452 15844 8480
rect 15427 8449 15439 8452
rect 15381 8443 15439 8449
rect 15838 8440 15844 8452
rect 15896 8480 15902 8492
rect 16666 8480 16672 8492
rect 15896 8452 16252 8480
rect 16627 8452 16672 8480
rect 15896 8440 15902 8452
rect 10321 8415 10379 8421
rect 10321 8381 10333 8415
rect 10367 8381 10379 8415
rect 10502 8412 10508 8424
rect 10415 8384 10508 8412
rect 10321 8375 10379 8381
rect 9217 8347 9275 8353
rect 9217 8313 9229 8347
rect 9263 8344 9275 8347
rect 10336 8344 10364 8375
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 13538 8372 13544 8424
rect 13596 8412 13602 8424
rect 13909 8415 13967 8421
rect 13909 8412 13921 8415
rect 13596 8384 13921 8412
rect 13596 8372 13602 8384
rect 13909 8381 13921 8384
rect 13955 8412 13967 8415
rect 14090 8412 14096 8424
rect 13955 8384 14096 8412
rect 13955 8381 13967 8384
rect 13909 8375 13967 8381
rect 14090 8372 14096 8384
rect 14148 8372 14154 8424
rect 16224 8421 16252 8452
rect 16666 8440 16672 8452
rect 16724 8440 16730 8492
rect 20916 8480 20944 8576
rect 23477 8551 23535 8557
rect 23477 8517 23489 8551
rect 23523 8548 23535 8551
rect 24302 8548 24308 8560
rect 23523 8520 24308 8548
rect 23523 8517 23535 8520
rect 23477 8511 23535 8517
rect 24302 8508 24308 8520
rect 24360 8508 24366 8560
rect 26881 8551 26939 8557
rect 26881 8517 26893 8551
rect 26927 8548 26939 8551
rect 27154 8548 27160 8560
rect 26927 8520 27160 8548
rect 26927 8517 26939 8520
rect 26881 8511 26939 8517
rect 27154 8508 27160 8520
rect 27212 8508 27218 8560
rect 33873 8551 33931 8557
rect 33873 8517 33885 8551
rect 33919 8548 33931 8551
rect 35802 8548 35808 8560
rect 33919 8520 35808 8548
rect 33919 8517 33931 8520
rect 33873 8511 33931 8517
rect 35802 8508 35808 8520
rect 35860 8508 35866 8560
rect 21358 8480 21364 8492
rect 20916 8452 21364 8480
rect 21358 8440 21364 8452
rect 21416 8480 21422 8492
rect 21913 8483 21971 8489
rect 21416 8452 21680 8480
rect 21416 8440 21422 8452
rect 15933 8415 15991 8421
rect 15933 8381 15945 8415
rect 15979 8381 15991 8415
rect 15933 8375 15991 8381
rect 16209 8415 16267 8421
rect 16209 8381 16221 8415
rect 16255 8381 16267 8415
rect 18782 8412 18788 8424
rect 18743 8384 18788 8412
rect 16209 8375 16267 8381
rect 10410 8344 10416 8356
rect 9263 8316 10088 8344
rect 10336 8316 10416 8344
rect 9263 8313 9275 8316
rect 9217 8307 9275 8313
rect 10060 8288 10088 8316
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 11882 8304 11888 8356
rect 11940 8344 11946 8356
rect 11977 8347 12035 8353
rect 11977 8344 11989 8347
rect 11940 8316 11989 8344
rect 11940 8304 11946 8316
rect 11977 8313 11989 8316
rect 12023 8344 12035 8347
rect 12023 8316 13814 8344
rect 12023 8313 12035 8316
rect 11977 8307 12035 8313
rect 9858 8276 9864 8288
rect 9819 8248 9864 8276
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 10042 8236 10048 8288
rect 10100 8276 10106 8288
rect 10137 8279 10195 8285
rect 10137 8276 10149 8279
rect 10100 8248 10149 8276
rect 10100 8236 10106 8248
rect 10137 8245 10149 8248
rect 10183 8245 10195 8279
rect 10137 8239 10195 8245
rect 13173 8279 13231 8285
rect 13173 8245 13185 8279
rect 13219 8276 13231 8279
rect 13262 8276 13268 8288
rect 13219 8248 13268 8276
rect 13219 8245 13231 8248
rect 13173 8239 13231 8245
rect 13262 8236 13268 8248
rect 13320 8276 13326 8288
rect 13630 8276 13636 8288
rect 13320 8248 13636 8276
rect 13320 8236 13326 8248
rect 13630 8236 13636 8248
rect 13688 8236 13694 8288
rect 13786 8276 13814 8316
rect 15470 8276 15476 8288
rect 13786 8248 15476 8276
rect 15470 8236 15476 8248
rect 15528 8276 15534 8288
rect 15841 8279 15899 8285
rect 15841 8276 15853 8279
rect 15528 8248 15853 8276
rect 15528 8236 15534 8248
rect 15841 8245 15853 8248
rect 15887 8276 15899 8279
rect 15948 8276 15976 8375
rect 18782 8372 18788 8384
rect 18840 8372 18846 8424
rect 18966 8412 18972 8424
rect 18927 8384 18972 8412
rect 18966 8372 18972 8384
rect 19024 8372 19030 8424
rect 20438 8372 20444 8424
rect 20496 8412 20502 8424
rect 20993 8415 21051 8421
rect 20993 8412 21005 8415
rect 20496 8384 21005 8412
rect 20496 8372 20502 8384
rect 20993 8381 21005 8384
rect 21039 8412 21051 8415
rect 21177 8415 21235 8421
rect 21177 8412 21189 8415
rect 21039 8384 21189 8412
rect 21039 8381 21051 8384
rect 20993 8375 21051 8381
rect 21177 8381 21189 8384
rect 21223 8412 21235 8415
rect 21266 8412 21272 8424
rect 21223 8384 21272 8412
rect 21223 8381 21235 8384
rect 21177 8375 21235 8381
rect 21266 8372 21272 8384
rect 21324 8372 21330 8424
rect 21652 8421 21680 8452
rect 21913 8449 21925 8483
rect 21959 8480 21971 8483
rect 22094 8480 22100 8492
rect 21959 8452 22100 8480
rect 21959 8449 21971 8452
rect 21913 8443 21971 8449
rect 22094 8440 22100 8452
rect 22152 8440 22158 8492
rect 23290 8440 23296 8492
rect 23348 8480 23354 8492
rect 24026 8480 24032 8492
rect 23348 8452 24032 8480
rect 23348 8440 23354 8452
rect 24026 8440 24032 8452
rect 24084 8480 24090 8492
rect 24213 8483 24271 8489
rect 24213 8480 24225 8483
rect 24084 8452 24225 8480
rect 24084 8440 24090 8452
rect 24213 8449 24225 8452
rect 24259 8449 24271 8483
rect 28350 8480 28356 8492
rect 28311 8452 28356 8480
rect 24213 8443 24271 8449
rect 28350 8440 28356 8452
rect 28408 8440 28414 8492
rect 32122 8440 32128 8492
rect 32180 8480 32186 8492
rect 32355 8483 32413 8489
rect 32355 8480 32367 8483
rect 32180 8452 32367 8480
rect 32180 8440 32186 8452
rect 32355 8449 32367 8452
rect 32401 8449 32413 8483
rect 32355 8443 32413 8449
rect 33134 8440 33140 8492
rect 33192 8480 33198 8492
rect 33321 8483 33379 8489
rect 33321 8480 33333 8483
rect 33192 8452 33333 8480
rect 33192 8440 33198 8452
rect 33321 8449 33333 8452
rect 33367 8449 33379 8483
rect 34974 8480 34980 8492
rect 34935 8452 34980 8480
rect 33321 8443 33379 8449
rect 34974 8440 34980 8452
rect 35032 8440 35038 8492
rect 35250 8480 35256 8492
rect 35211 8452 35256 8480
rect 35250 8440 35256 8452
rect 35308 8480 35314 8492
rect 36538 8480 36544 8492
rect 35308 8452 36544 8480
rect 35308 8440 35314 8452
rect 36538 8440 36544 8452
rect 36596 8440 36602 8492
rect 37182 8480 37188 8492
rect 37095 8452 37188 8480
rect 37182 8440 37188 8452
rect 37240 8480 37246 8492
rect 38102 8480 38108 8492
rect 37240 8452 38108 8480
rect 37240 8440 37246 8452
rect 38102 8440 38108 8452
rect 38160 8440 38166 8492
rect 21637 8415 21695 8421
rect 21637 8381 21649 8415
rect 21683 8412 21695 8415
rect 23474 8412 23480 8424
rect 21683 8384 23480 8412
rect 21683 8381 21695 8384
rect 21637 8375 21695 8381
rect 23474 8372 23480 8384
rect 23532 8412 23538 8424
rect 23934 8412 23940 8424
rect 23532 8384 23940 8412
rect 23532 8372 23538 8384
rect 23934 8372 23940 8384
rect 23992 8372 23998 8424
rect 30469 8415 30527 8421
rect 30469 8412 30481 8415
rect 29564 8384 30481 8412
rect 18230 8304 18236 8356
rect 18288 8344 18294 8356
rect 18325 8347 18383 8353
rect 18325 8344 18337 8347
rect 18288 8316 18337 8344
rect 18288 8304 18294 8316
rect 18325 8313 18337 8316
rect 18371 8344 18383 8347
rect 18693 8347 18751 8353
rect 18693 8344 18705 8347
rect 18371 8316 18705 8344
rect 18371 8313 18383 8316
rect 18325 8307 18383 8313
rect 18693 8313 18705 8316
rect 18739 8344 18751 8347
rect 18984 8344 19012 8372
rect 18739 8316 19012 8344
rect 19705 8347 19763 8353
rect 18739 8313 18751 8316
rect 18693 8307 18751 8313
rect 19705 8313 19717 8347
rect 19751 8344 19763 8347
rect 19886 8344 19892 8356
rect 19751 8316 19892 8344
rect 19751 8313 19763 8316
rect 19705 8307 19763 8313
rect 19886 8304 19892 8316
rect 19944 8304 19950 8356
rect 24029 8347 24087 8353
rect 24029 8313 24041 8347
rect 24075 8344 24087 8347
rect 24302 8344 24308 8356
rect 24075 8316 24308 8344
rect 24075 8313 24087 8316
rect 24029 8307 24087 8313
rect 24302 8304 24308 8316
rect 24360 8304 24366 8356
rect 24854 8344 24860 8356
rect 24815 8316 24860 8344
rect 24854 8304 24860 8316
rect 24912 8304 24918 8356
rect 25777 8347 25835 8353
rect 25777 8313 25789 8347
rect 25823 8313 25835 8347
rect 25777 8307 25835 8313
rect 16114 8276 16120 8288
rect 15887 8248 16120 8276
rect 15887 8245 15899 8248
rect 15841 8239 15899 8245
rect 16114 8236 16120 8248
rect 16172 8236 16178 8288
rect 19058 8276 19064 8288
rect 19019 8248 19064 8276
rect 19058 8236 19064 8248
rect 19116 8236 19122 8288
rect 24320 8276 24348 8304
rect 25130 8276 25136 8288
rect 24320 8248 25136 8276
rect 25130 8236 25136 8248
rect 25188 8236 25194 8288
rect 25682 8236 25688 8288
rect 25740 8276 25746 8288
rect 25792 8276 25820 8307
rect 25866 8304 25872 8356
rect 25924 8344 25930 8356
rect 26421 8347 26479 8353
rect 25924 8316 25969 8344
rect 25924 8304 25930 8316
rect 26421 8313 26433 8347
rect 26467 8344 26479 8347
rect 27246 8344 27252 8356
rect 26467 8316 27252 8344
rect 26467 8313 26479 8316
rect 26421 8307 26479 8313
rect 27246 8304 27252 8316
rect 27304 8304 27310 8356
rect 27706 8344 27712 8356
rect 27667 8316 27712 8344
rect 27706 8304 27712 8316
rect 27764 8304 27770 8356
rect 27801 8347 27859 8353
rect 27801 8313 27813 8347
rect 27847 8313 27859 8347
rect 27801 8307 27859 8313
rect 25740 8248 25820 8276
rect 25740 8236 25746 8248
rect 27338 8236 27344 8288
rect 27396 8276 27402 8288
rect 27816 8276 27844 8307
rect 29564 8288 29592 8384
rect 30469 8381 30481 8384
rect 30515 8381 30527 8415
rect 30469 8375 30527 8381
rect 31389 8415 31447 8421
rect 31389 8381 31401 8415
rect 31435 8412 31447 8415
rect 32033 8415 32091 8421
rect 32033 8412 32045 8415
rect 31435 8384 32045 8412
rect 31435 8381 31447 8384
rect 31389 8375 31447 8381
rect 32033 8381 32045 8384
rect 32079 8412 32091 8415
rect 32252 8415 32310 8421
rect 32252 8412 32264 8415
rect 32079 8384 32264 8412
rect 32079 8381 32091 8384
rect 32033 8375 32091 8381
rect 32252 8381 32264 8384
rect 32298 8381 32310 8415
rect 38010 8412 38016 8424
rect 37971 8384 38016 8412
rect 32252 8375 32310 8381
rect 38010 8372 38016 8384
rect 38068 8412 38074 8424
rect 38470 8412 38476 8424
rect 38068 8384 38476 8412
rect 38068 8372 38074 8384
rect 38470 8372 38476 8384
rect 38528 8372 38534 8424
rect 30282 8304 30288 8356
rect 30340 8344 30346 8356
rect 30790 8347 30848 8353
rect 30790 8344 30802 8347
rect 30340 8316 30802 8344
rect 30340 8304 30346 8316
rect 30790 8313 30802 8316
rect 30836 8344 30848 8347
rect 31662 8344 31668 8356
rect 30836 8316 31668 8344
rect 30836 8313 30848 8316
rect 30790 8307 30848 8313
rect 31662 8304 31668 8316
rect 31720 8304 31726 8356
rect 33137 8347 33195 8353
rect 33137 8313 33149 8347
rect 33183 8344 33195 8347
rect 33413 8347 33471 8353
rect 33413 8344 33425 8347
rect 33183 8316 33425 8344
rect 33183 8313 33195 8316
rect 33137 8307 33195 8313
rect 33413 8313 33425 8316
rect 33459 8344 33471 8347
rect 34238 8344 34244 8356
rect 33459 8316 34244 8344
rect 33459 8313 33471 8316
rect 33413 8307 33471 8313
rect 34238 8304 34244 8316
rect 34296 8304 34302 8356
rect 34698 8304 34704 8356
rect 34756 8344 34762 8356
rect 35069 8347 35127 8353
rect 35069 8344 35081 8347
rect 34756 8316 35081 8344
rect 34756 8304 34762 8316
rect 35069 8313 35081 8316
rect 35115 8313 35127 8347
rect 35069 8307 35127 8313
rect 36262 8304 36268 8356
rect 36320 8344 36326 8356
rect 36633 8347 36691 8353
rect 36633 8344 36645 8347
rect 36320 8316 36645 8344
rect 36320 8304 36326 8316
rect 36633 8313 36645 8316
rect 36679 8313 36691 8347
rect 36633 8307 36691 8313
rect 28994 8276 29000 8288
rect 27396 8248 27844 8276
rect 28955 8248 29000 8276
rect 27396 8236 27402 8248
rect 28994 8236 29000 8248
rect 29052 8236 29058 8288
rect 29546 8276 29552 8288
rect 29507 8248 29552 8276
rect 29546 8236 29552 8248
rect 29604 8236 29610 8288
rect 36354 8236 36360 8288
rect 36412 8276 36418 8288
rect 37737 8279 37795 8285
rect 37737 8276 37749 8279
rect 36412 8248 37749 8276
rect 36412 8236 36418 8248
rect 37737 8245 37749 8248
rect 37783 8276 37795 8279
rect 37918 8276 37924 8288
rect 37783 8248 37924 8276
rect 37783 8245 37795 8248
rect 37737 8239 37795 8245
rect 37918 8236 37924 8248
rect 37976 8236 37982 8288
rect 38194 8276 38200 8288
rect 38155 8248 38200 8276
rect 38194 8236 38200 8248
rect 38252 8236 38258 8288
rect 1104 8186 48852 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 48852 8186
rect 1104 8112 48852 8134
rect 13357 8075 13415 8081
rect 13357 8041 13369 8075
rect 13403 8072 13415 8075
rect 13538 8072 13544 8084
rect 13403 8044 13544 8072
rect 13403 8041 13415 8044
rect 13357 8035 13415 8041
rect 13538 8032 13544 8044
rect 13596 8032 13602 8084
rect 13722 8072 13728 8084
rect 13648 8044 13728 8072
rect 10594 8004 10600 8016
rect 10555 7976 10600 8004
rect 10594 7964 10600 7976
rect 10652 7964 10658 8016
rect 12158 8004 12164 8016
rect 12119 7976 12164 8004
rect 12158 7964 12164 7976
rect 12216 7964 12222 8016
rect 13648 8013 13676 8044
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 17494 8072 17500 8084
rect 17455 8044 17500 8072
rect 17494 8032 17500 8044
rect 17552 8032 17558 8084
rect 18782 8072 18788 8084
rect 18743 8044 18788 8072
rect 18782 8032 18788 8044
rect 18840 8072 18846 8084
rect 24026 8072 24032 8084
rect 18840 8044 19472 8072
rect 23987 8044 24032 8072
rect 18840 8032 18846 8044
rect 19444 8016 19472 8044
rect 24026 8032 24032 8044
rect 24084 8032 24090 8084
rect 26050 8072 26056 8084
rect 24320 8044 26056 8072
rect 13633 8007 13691 8013
rect 13633 7973 13645 8007
rect 13679 7973 13691 8007
rect 13633 7967 13691 7973
rect 16577 8007 16635 8013
rect 16577 7973 16589 8007
rect 16623 8004 16635 8007
rect 17126 8004 17132 8016
rect 16623 7976 17132 8004
rect 16623 7973 16635 7976
rect 16577 7967 16635 7973
rect 17126 7964 17132 7976
rect 17184 7964 17190 8016
rect 19426 8004 19432 8016
rect 19339 7976 19432 8004
rect 19426 7964 19432 7976
rect 19484 7964 19490 8016
rect 19981 8007 20039 8013
rect 19981 7973 19993 8007
rect 20027 8004 20039 8007
rect 21450 8004 21456 8016
rect 20027 7976 21456 8004
rect 20027 7973 20039 7976
rect 19981 7967 20039 7973
rect 21450 7964 21456 7976
rect 21508 8004 21514 8016
rect 23014 8004 23020 8016
rect 21508 7976 22416 8004
rect 22927 7976 23020 8004
rect 21508 7964 21514 7976
rect 13722 7936 13728 7948
rect 13683 7908 13728 7936
rect 13722 7896 13728 7908
rect 13780 7896 13786 7948
rect 15838 7936 15844 7948
rect 15799 7908 15844 7936
rect 15838 7896 15844 7908
rect 15896 7896 15902 7948
rect 17402 7936 17408 7948
rect 17363 7908 17408 7936
rect 17402 7896 17408 7908
rect 17460 7896 17466 7948
rect 17862 7896 17868 7948
rect 17920 7936 17926 7948
rect 17957 7939 18015 7945
rect 17957 7936 17969 7939
rect 17920 7908 17969 7936
rect 17920 7896 17926 7908
rect 17957 7905 17969 7908
rect 18003 7936 18015 7939
rect 19058 7936 19064 7948
rect 18003 7908 19064 7936
rect 18003 7905 18015 7908
rect 17957 7899 18015 7905
rect 19058 7896 19064 7908
rect 19116 7896 19122 7948
rect 19610 7936 19616 7948
rect 19571 7908 19616 7936
rect 19610 7896 19616 7908
rect 19668 7936 19674 7948
rect 19886 7936 19892 7948
rect 19668 7908 19892 7936
rect 19668 7896 19674 7908
rect 19886 7896 19892 7908
rect 19944 7896 19950 7948
rect 21082 7936 21088 7948
rect 21043 7908 21088 7936
rect 21082 7896 21088 7908
rect 21140 7896 21146 7948
rect 21358 7936 21364 7948
rect 21319 7908 21364 7936
rect 21358 7896 21364 7908
rect 21416 7896 21422 7948
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7868 8631 7871
rect 10505 7871 10563 7877
rect 10505 7868 10517 7871
rect 8619 7840 10517 7868
rect 8619 7837 8631 7840
rect 8573 7831 8631 7837
rect 10505 7837 10517 7840
rect 10551 7868 10563 7871
rect 11146 7868 11152 7880
rect 10551 7840 11152 7868
rect 10551 7837 10563 7840
rect 10505 7831 10563 7837
rect 11146 7828 11152 7840
rect 11204 7828 11210 7880
rect 12066 7868 12072 7880
rect 12027 7840 12072 7868
rect 12066 7828 12072 7840
rect 12124 7828 12130 7880
rect 12345 7871 12403 7877
rect 12345 7837 12357 7871
rect 12391 7837 12403 7871
rect 16206 7868 16212 7880
rect 16167 7840 16212 7868
rect 12345 7831 12403 7837
rect 11057 7803 11115 7809
rect 11057 7769 11069 7803
rect 11103 7800 11115 7803
rect 11330 7800 11336 7812
rect 11103 7772 11336 7800
rect 11103 7769 11115 7772
rect 11057 7763 11115 7769
rect 11330 7760 11336 7772
rect 11388 7800 11394 7812
rect 12360 7800 12388 7831
rect 16206 7828 16212 7840
rect 16264 7828 16270 7880
rect 21637 7871 21695 7877
rect 21637 7837 21649 7871
rect 21683 7868 21695 7871
rect 21818 7868 21824 7880
rect 21683 7840 21824 7868
rect 21683 7837 21695 7840
rect 21637 7831 21695 7837
rect 21818 7828 21824 7840
rect 21876 7868 21882 7880
rect 21913 7871 21971 7877
rect 21913 7868 21925 7871
rect 21876 7840 21925 7868
rect 21876 7828 21882 7840
rect 21913 7837 21925 7840
rect 21959 7837 21971 7871
rect 22388 7868 22416 7976
rect 22940 7945 22968 7976
rect 23014 7964 23020 7976
rect 23072 8004 23078 8016
rect 24320 8004 24348 8044
rect 26050 8032 26056 8044
rect 26108 8032 26114 8084
rect 26329 8075 26387 8081
rect 26329 8041 26341 8075
rect 26375 8072 26387 8075
rect 26878 8072 26884 8084
rect 26375 8044 26884 8072
rect 26375 8041 26387 8044
rect 26329 8035 26387 8041
rect 26878 8032 26884 8044
rect 26936 8032 26942 8084
rect 27706 8072 27712 8084
rect 27667 8044 27712 8072
rect 27706 8032 27712 8044
rect 27764 8072 27770 8084
rect 28215 8075 28273 8081
rect 28215 8072 28227 8075
rect 27764 8044 28227 8072
rect 27764 8032 27770 8044
rect 28215 8041 28227 8044
rect 28261 8041 28273 8075
rect 29546 8072 29552 8084
rect 29507 8044 29552 8072
rect 28215 8035 28273 8041
rect 29546 8032 29552 8044
rect 29604 8032 29610 8084
rect 31067 8075 31125 8081
rect 31067 8041 31079 8075
rect 31113 8072 31125 8075
rect 31754 8072 31760 8084
rect 31113 8044 31760 8072
rect 31113 8041 31125 8044
rect 31067 8035 31125 8041
rect 31754 8032 31760 8044
rect 31812 8032 31818 8084
rect 32214 8072 32220 8084
rect 32175 8044 32220 8072
rect 32214 8032 32220 8044
rect 32272 8032 32278 8084
rect 34054 8072 34060 8084
rect 34015 8044 34060 8072
rect 34054 8032 34060 8044
rect 34112 8032 34118 8084
rect 35526 8072 35532 8084
rect 35487 8044 35532 8072
rect 35526 8032 35532 8044
rect 35584 8032 35590 8084
rect 35989 8075 36047 8081
rect 35989 8041 36001 8075
rect 36035 8072 36047 8075
rect 36354 8072 36360 8084
rect 36035 8044 36360 8072
rect 36035 8041 36047 8044
rect 35989 8035 36047 8041
rect 36354 8032 36360 8044
rect 36412 8072 36418 8084
rect 37182 8072 37188 8084
rect 36412 8044 37188 8072
rect 36412 8032 36418 8044
rect 37182 8032 37188 8044
rect 37240 8032 37246 8084
rect 23072 7976 24348 8004
rect 23072 7964 23078 7976
rect 24394 7964 24400 8016
rect 24452 8004 24458 8016
rect 24946 8004 24952 8016
rect 24452 7976 24497 8004
rect 24907 7976 24952 8004
rect 24452 7964 24458 7976
rect 24946 7964 24952 7976
rect 25004 7964 25010 8016
rect 25130 7964 25136 8016
rect 25188 8004 25194 8016
rect 26418 8004 26424 8016
rect 25188 7976 26424 8004
rect 25188 7964 25194 7976
rect 26418 7964 26424 7976
rect 26476 8004 26482 8016
rect 26697 8007 26755 8013
rect 26697 8004 26709 8007
rect 26476 7976 26709 8004
rect 26476 7964 26482 7976
rect 26697 7973 26709 7976
rect 26743 8004 26755 8007
rect 27522 8004 27528 8016
rect 26743 7976 27528 8004
rect 26743 7973 26755 7976
rect 26697 7967 26755 7973
rect 27522 7964 27528 7976
rect 27580 7964 27586 8016
rect 28994 7964 29000 8016
rect 29052 8004 29058 8016
rect 29052 7976 29776 8004
rect 29052 7964 29058 7976
rect 22925 7939 22983 7945
rect 22925 7905 22937 7939
rect 22971 7905 22983 7939
rect 22925 7899 22983 7905
rect 23109 7939 23167 7945
rect 23109 7905 23121 7939
rect 23155 7905 23167 7939
rect 23109 7899 23167 7905
rect 22830 7868 22836 7880
rect 22388 7840 22836 7868
rect 21913 7831 21971 7837
rect 22830 7828 22836 7840
rect 22888 7868 22894 7880
rect 23124 7868 23152 7899
rect 27890 7896 27896 7948
rect 27948 7936 27954 7948
rect 28112 7939 28170 7945
rect 28112 7936 28124 7939
rect 27948 7908 28124 7936
rect 27948 7896 27954 7908
rect 28112 7905 28124 7908
rect 28158 7905 28170 7939
rect 28112 7899 28170 7905
rect 28258 7896 28264 7948
rect 28316 7936 28322 7948
rect 29273 7939 29331 7945
rect 29273 7936 29285 7939
rect 28316 7908 29285 7936
rect 28316 7896 28322 7908
rect 29273 7905 29285 7908
rect 29319 7936 29331 7939
rect 29454 7936 29460 7948
rect 29319 7908 29460 7936
rect 29319 7905 29331 7908
rect 29273 7899 29331 7905
rect 29454 7896 29460 7908
rect 29512 7896 29518 7948
rect 29748 7945 29776 7976
rect 33134 7964 33140 8016
rect 33192 8004 33198 8016
rect 33229 8007 33287 8013
rect 33229 8004 33241 8007
rect 33192 7976 33241 8004
rect 33192 7964 33198 7976
rect 33229 7973 33241 7976
rect 33275 7973 33287 8007
rect 33229 7967 33287 7973
rect 34238 7964 34244 8016
rect 34296 8004 34302 8016
rect 34333 8007 34391 8013
rect 34333 8004 34345 8007
rect 34296 7976 34345 8004
rect 34296 7964 34302 7976
rect 34333 7973 34345 7976
rect 34379 7973 34391 8007
rect 34333 7967 34391 7973
rect 34885 8007 34943 8013
rect 34885 7973 34897 8007
rect 34931 8004 34943 8007
rect 35250 8004 35256 8016
rect 34931 7976 35256 8004
rect 34931 7973 34943 7976
rect 34885 7967 34943 7973
rect 35250 7964 35256 7976
rect 35308 7964 35314 8016
rect 36262 8004 36268 8016
rect 36223 7976 36268 8004
rect 36262 7964 36268 7976
rect 36320 7964 36326 8016
rect 36814 8004 36820 8016
rect 36775 7976 36820 8004
rect 36814 7964 36820 7976
rect 36872 7964 36878 8016
rect 37918 8004 37924 8016
rect 37879 7976 37924 8004
rect 37918 7964 37924 7976
rect 37976 7964 37982 8016
rect 29733 7939 29791 7945
rect 29733 7905 29745 7939
rect 29779 7905 29791 7939
rect 29733 7899 29791 7905
rect 30558 7896 30564 7948
rect 30616 7936 30622 7948
rect 30964 7939 31022 7945
rect 30964 7936 30976 7939
rect 30616 7908 30976 7936
rect 30616 7896 30622 7908
rect 30964 7905 30976 7908
rect 31010 7936 31022 7939
rect 31389 7939 31447 7945
rect 31389 7936 31401 7939
rect 31010 7908 31401 7936
rect 31010 7905 31022 7908
rect 30964 7899 31022 7905
rect 31389 7905 31401 7908
rect 31435 7905 31447 7939
rect 32122 7936 32128 7948
rect 32083 7908 32128 7936
rect 31389 7899 31447 7905
rect 32122 7896 32128 7908
rect 32180 7896 32186 7948
rect 32585 7939 32643 7945
rect 32585 7905 32597 7939
rect 32631 7905 32643 7939
rect 32585 7899 32643 7905
rect 23382 7868 23388 7880
rect 22888 7840 23152 7868
rect 23343 7840 23388 7868
rect 22888 7828 22894 7840
rect 23382 7828 23388 7840
rect 23440 7828 23446 7880
rect 24302 7868 24308 7880
rect 24263 7840 24308 7868
rect 24302 7828 24308 7840
rect 24360 7828 24366 7880
rect 26602 7868 26608 7880
rect 26563 7840 26608 7868
rect 26602 7828 26608 7840
rect 26660 7828 26666 7880
rect 27246 7868 27252 7880
rect 27207 7840 27252 7868
rect 27246 7828 27252 7840
rect 27304 7828 27310 7880
rect 32600 7868 32628 7899
rect 33134 7868 33140 7880
rect 30668 7840 33140 7868
rect 15930 7800 15936 7812
rect 11388 7772 12388 7800
rect 15580 7772 15936 7800
rect 11388 7760 11394 7772
rect 15580 7744 15608 7772
rect 15930 7760 15936 7772
rect 15988 7809 15994 7812
rect 15988 7803 16037 7809
rect 15988 7769 15991 7803
rect 16025 7769 16037 7803
rect 15988 7763 16037 7769
rect 15988 7760 15994 7763
rect 25038 7760 25044 7812
rect 25096 7800 25102 7812
rect 30285 7803 30343 7809
rect 30285 7800 30297 7803
rect 25096 7772 30297 7800
rect 25096 7760 25102 7772
rect 30285 7769 30297 7772
rect 30331 7800 30343 7803
rect 30558 7800 30564 7812
rect 30331 7772 30564 7800
rect 30331 7769 30343 7772
rect 30285 7763 30343 7769
rect 30558 7760 30564 7772
rect 30616 7800 30622 7812
rect 30668 7809 30696 7840
rect 33134 7828 33140 7840
rect 33192 7828 33198 7880
rect 34241 7871 34299 7877
rect 34241 7837 34253 7871
rect 34287 7868 34299 7871
rect 34514 7868 34520 7880
rect 34287 7840 34520 7868
rect 34287 7837 34299 7840
rect 34241 7831 34299 7837
rect 34514 7828 34520 7840
rect 34572 7828 34578 7880
rect 35802 7828 35808 7880
rect 35860 7868 35866 7880
rect 36170 7868 36176 7880
rect 35860 7840 36176 7868
rect 35860 7828 35866 7840
rect 36170 7828 36176 7840
rect 36228 7828 36234 7880
rect 36832 7868 36860 7964
rect 38470 7896 38476 7948
rect 38528 7936 38534 7948
rect 39298 7936 39304 7948
rect 39356 7945 39362 7948
rect 39356 7939 39394 7945
rect 38528 7908 39304 7936
rect 38528 7896 38534 7908
rect 39298 7896 39304 7908
rect 39382 7905 39394 7939
rect 39356 7899 39394 7905
rect 39356 7896 39362 7899
rect 37826 7868 37832 7880
rect 36832 7840 37832 7868
rect 37826 7828 37832 7840
rect 37884 7828 37890 7880
rect 38102 7868 38108 7880
rect 38063 7840 38108 7868
rect 38102 7828 38108 7840
rect 38160 7828 38166 7880
rect 30653 7803 30711 7809
rect 30653 7800 30665 7803
rect 30616 7772 30665 7800
rect 30616 7760 30622 7772
rect 30653 7769 30665 7772
rect 30699 7769 30711 7803
rect 30653 7763 30711 7769
rect 10137 7735 10195 7741
rect 10137 7701 10149 7735
rect 10183 7732 10195 7735
rect 10410 7732 10416 7744
rect 10183 7704 10416 7732
rect 10183 7701 10195 7704
rect 10137 7695 10195 7701
rect 10410 7692 10416 7704
rect 10468 7692 10474 7744
rect 15562 7732 15568 7744
rect 15523 7704 15568 7732
rect 15562 7692 15568 7704
rect 15620 7692 15626 7744
rect 16114 7692 16120 7744
rect 16172 7732 16178 7744
rect 16942 7732 16948 7744
rect 16172 7704 16217 7732
rect 16903 7704 16948 7732
rect 16172 7692 16178 7704
rect 16942 7692 16948 7704
rect 17000 7692 17006 7744
rect 23658 7732 23664 7744
rect 23619 7704 23664 7732
rect 23658 7692 23664 7704
rect 23716 7692 23722 7744
rect 25682 7732 25688 7744
rect 25643 7704 25688 7732
rect 25682 7692 25688 7704
rect 25740 7692 25746 7744
rect 38470 7692 38476 7744
rect 38528 7732 38534 7744
rect 39439 7735 39497 7741
rect 39439 7732 39451 7735
rect 38528 7704 39451 7732
rect 38528 7692 38534 7704
rect 39439 7701 39451 7704
rect 39485 7701 39497 7735
rect 39439 7695 39497 7701
rect 1104 7642 48852 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 48852 7642
rect 1104 7568 48852 7590
rect 9858 7528 9864 7540
rect 9819 7500 9864 7528
rect 9858 7488 9864 7500
rect 9916 7488 9922 7540
rect 10594 7488 10600 7540
rect 10652 7528 10658 7540
rect 10873 7531 10931 7537
rect 10873 7528 10885 7531
rect 10652 7500 10885 7528
rect 10652 7488 10658 7500
rect 10873 7497 10885 7500
rect 10919 7497 10931 7531
rect 11146 7528 11152 7540
rect 11107 7500 11152 7528
rect 10873 7491 10931 7497
rect 11146 7488 11152 7500
rect 11204 7488 11210 7540
rect 14274 7488 14280 7540
rect 14332 7528 14338 7540
rect 15470 7537 15476 7540
rect 14369 7531 14427 7537
rect 14369 7528 14381 7531
rect 14332 7500 14381 7528
rect 14332 7488 14338 7500
rect 14369 7497 14381 7500
rect 14415 7497 14427 7531
rect 14369 7491 14427 7497
rect 15454 7531 15476 7537
rect 15454 7497 15466 7531
rect 15454 7491 15476 7497
rect 9493 7463 9551 7469
rect 9493 7460 9505 7463
rect 8772 7432 9505 7460
rect 8481 7327 8539 7333
rect 8481 7293 8493 7327
rect 8527 7324 8539 7327
rect 8570 7324 8576 7336
rect 8527 7296 8576 7324
rect 8527 7293 8539 7296
rect 8481 7287 8539 7293
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 8772 7333 8800 7432
rect 9493 7429 9505 7432
rect 9539 7460 9551 7463
rect 11885 7463 11943 7469
rect 9539 7432 11514 7460
rect 9539 7429 9551 7432
rect 9493 7423 9551 7429
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7392 9183 7395
rect 10226 7392 10232 7404
rect 9171 7364 10232 7392
rect 9171 7361 9183 7364
rect 9125 7355 9183 7361
rect 10226 7352 10232 7364
rect 10284 7352 10290 7404
rect 11486 7392 11514 7432
rect 11885 7429 11897 7463
rect 11931 7460 11943 7463
rect 12158 7460 12164 7472
rect 11931 7432 12164 7460
rect 11931 7429 11943 7432
rect 11885 7423 11943 7429
rect 12158 7420 12164 7432
rect 12216 7460 12222 7472
rect 13357 7463 13415 7469
rect 13357 7460 13369 7463
rect 12216 7432 13369 7460
rect 12216 7420 12222 7432
rect 13357 7429 13369 7432
rect 13403 7429 13415 7463
rect 14384 7460 14412 7491
rect 15470 7488 15476 7491
rect 15528 7488 15534 7540
rect 15746 7528 15752 7540
rect 15707 7500 15752 7528
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 17083 7531 17141 7537
rect 17083 7497 17095 7531
rect 17129 7528 17141 7531
rect 17954 7528 17960 7540
rect 17129 7500 17960 7528
rect 17129 7497 17141 7500
rect 17083 7491 17141 7497
rect 17954 7488 17960 7500
rect 18012 7488 18018 7540
rect 20717 7531 20775 7537
rect 20717 7497 20729 7531
rect 20763 7528 20775 7531
rect 21174 7528 21180 7540
rect 20763 7500 21180 7528
rect 20763 7497 20775 7500
rect 20717 7491 20775 7497
rect 21174 7488 21180 7500
rect 21232 7528 21238 7540
rect 21358 7528 21364 7540
rect 21232 7500 21364 7528
rect 21232 7488 21238 7500
rect 21358 7488 21364 7500
rect 21416 7488 21422 7540
rect 21729 7531 21787 7537
rect 21729 7497 21741 7531
rect 21775 7528 21787 7531
rect 22278 7528 22284 7540
rect 21775 7500 22284 7528
rect 21775 7497 21787 7500
rect 21729 7491 21787 7497
rect 22278 7488 22284 7500
rect 22336 7488 22342 7540
rect 23014 7528 23020 7540
rect 22975 7500 23020 7528
rect 23014 7488 23020 7500
rect 23072 7488 23078 7540
rect 24302 7528 24308 7540
rect 23124 7500 24308 7528
rect 14734 7460 14740 7472
rect 14384 7432 14740 7460
rect 13357 7423 13415 7429
rect 14734 7420 14740 7432
rect 14792 7460 14798 7472
rect 15565 7463 15623 7469
rect 15565 7460 15577 7463
rect 14792 7432 15577 7460
rect 14792 7420 14798 7432
rect 15565 7429 15577 7432
rect 15611 7429 15623 7463
rect 17402 7460 17408 7472
rect 17363 7432 17408 7460
rect 15565 7423 15623 7429
rect 17402 7420 17408 7432
rect 17460 7420 17466 7472
rect 17862 7460 17868 7472
rect 17823 7432 17868 7460
rect 17862 7420 17868 7432
rect 17920 7420 17926 7472
rect 19610 7460 19616 7472
rect 19523 7432 19616 7460
rect 13541 7395 13599 7401
rect 13541 7392 13553 7395
rect 11486 7364 13553 7392
rect 13541 7361 13553 7364
rect 13587 7392 13599 7395
rect 13722 7392 13728 7404
rect 13587 7364 13728 7392
rect 13587 7361 13599 7364
rect 13541 7355 13599 7361
rect 13722 7352 13728 7364
rect 13780 7392 13786 7404
rect 15105 7395 15163 7401
rect 15105 7392 15117 7395
rect 13780 7364 15117 7392
rect 13780 7352 13786 7364
rect 15105 7361 15117 7364
rect 15151 7392 15163 7395
rect 15657 7395 15715 7401
rect 15657 7392 15669 7395
rect 15151 7364 15669 7392
rect 15151 7361 15163 7364
rect 15105 7355 15163 7361
rect 15657 7361 15669 7364
rect 15703 7361 15715 7395
rect 15657 7355 15715 7361
rect 18877 7395 18935 7401
rect 18877 7361 18889 7395
rect 18923 7392 18935 7395
rect 19536 7392 19564 7432
rect 19610 7420 19616 7432
rect 19668 7460 19674 7472
rect 20947 7463 21005 7469
rect 19668 7432 20116 7460
rect 19668 7420 19674 7432
rect 18923 7364 19564 7392
rect 18923 7361 18935 7364
rect 18877 7355 18935 7361
rect 8757 7327 8815 7333
rect 8757 7293 8769 7327
rect 8803 7293 8815 7327
rect 9950 7324 9956 7336
rect 9911 7296 9956 7324
rect 8757 7287 8815 7293
rect 9950 7284 9956 7296
rect 10008 7284 10014 7336
rect 12434 7324 12440 7336
rect 12395 7296 12440 7324
rect 12434 7284 12440 7296
rect 12492 7324 12498 7336
rect 14001 7327 14059 7333
rect 14001 7324 14013 7327
rect 12492 7296 14013 7324
rect 12492 7284 12498 7296
rect 14001 7293 14013 7296
rect 14047 7293 14059 7327
rect 14001 7287 14059 7293
rect 14090 7284 14096 7336
rect 14148 7324 14154 7336
rect 14829 7327 14887 7333
rect 14829 7324 14841 7327
rect 14148 7296 14841 7324
rect 14148 7284 14154 7296
rect 14829 7293 14841 7296
rect 14875 7324 14887 7327
rect 15289 7327 15347 7333
rect 15289 7324 15301 7327
rect 14875 7296 15301 7324
rect 14875 7293 14887 7296
rect 14829 7287 14887 7293
rect 15289 7293 15301 7296
rect 15335 7324 15347 7327
rect 15838 7324 15844 7336
rect 15335 7296 15844 7324
rect 15335 7293 15347 7296
rect 15289 7287 15347 7293
rect 15838 7284 15844 7296
rect 15896 7324 15902 7336
rect 16853 7327 16911 7333
rect 15896 7296 16804 7324
rect 15896 7284 15902 7296
rect 9858 7216 9864 7268
rect 9916 7256 9922 7268
rect 10274 7259 10332 7265
rect 10274 7256 10286 7259
rect 9916 7228 10286 7256
rect 9916 7216 9922 7228
rect 10274 7225 10286 7228
rect 10320 7256 10332 7259
rect 10778 7256 10784 7268
rect 10320 7228 10784 7256
rect 10320 7225 10332 7228
rect 10274 7219 10332 7225
rect 10778 7216 10784 7228
rect 10836 7256 10842 7268
rect 12161 7259 12219 7265
rect 12161 7256 12173 7259
rect 10836 7228 12173 7256
rect 10836 7216 10842 7228
rect 12161 7225 12173 7228
rect 12207 7256 12219 7259
rect 12758 7259 12816 7265
rect 12758 7256 12770 7259
rect 12207 7228 12770 7256
rect 12207 7225 12219 7228
rect 12161 7219 12219 7225
rect 12758 7225 12770 7228
rect 12804 7225 12816 7259
rect 12758 7219 12816 7225
rect 15746 7216 15752 7268
rect 15804 7256 15810 7268
rect 16114 7256 16120 7268
rect 15804 7228 16120 7256
rect 15804 7216 15810 7228
rect 16114 7216 16120 7228
rect 16172 7256 16178 7268
rect 16301 7259 16359 7265
rect 16301 7256 16313 7259
rect 16172 7228 16313 7256
rect 16172 7216 16178 7228
rect 16301 7225 16313 7228
rect 16347 7225 16359 7259
rect 16301 7219 16359 7225
rect 13262 7148 13268 7200
rect 13320 7188 13326 7200
rect 16776 7197 16804 7296
rect 16853 7293 16865 7327
rect 16899 7324 16911 7327
rect 16942 7324 16948 7336
rect 16899 7296 16948 7324
rect 16899 7293 16911 7296
rect 16853 7287 16911 7293
rect 16942 7284 16948 7296
rect 17000 7284 17006 7336
rect 19536 7333 19564 7364
rect 19521 7327 19579 7333
rect 19521 7293 19533 7327
rect 19567 7293 19579 7327
rect 19521 7287 19579 7293
rect 18966 7216 18972 7268
rect 19024 7256 19030 7268
rect 20088 7265 20116 7432
rect 20947 7429 20959 7463
rect 20993 7460 21005 7463
rect 23124 7460 23152 7500
rect 24302 7488 24308 7500
rect 24360 7488 24366 7540
rect 24394 7488 24400 7540
rect 24452 7528 24458 7540
rect 24857 7531 24915 7537
rect 24857 7528 24869 7531
rect 24452 7500 24869 7528
rect 24452 7488 24458 7500
rect 24857 7497 24869 7500
rect 24903 7497 24915 7531
rect 24857 7491 24915 7497
rect 26329 7531 26387 7537
rect 26329 7497 26341 7531
rect 26375 7528 26387 7531
rect 26418 7528 26424 7540
rect 26375 7500 26424 7528
rect 26375 7497 26387 7500
rect 26329 7491 26387 7497
rect 26418 7488 26424 7500
rect 26476 7488 26482 7540
rect 26697 7531 26755 7537
rect 26697 7497 26709 7531
rect 26743 7528 26755 7531
rect 27154 7528 27160 7540
rect 26743 7500 27160 7528
rect 26743 7497 26755 7500
rect 26697 7491 26755 7497
rect 27154 7488 27160 7500
rect 27212 7488 27218 7540
rect 27614 7488 27620 7540
rect 27672 7528 27678 7540
rect 27709 7531 27767 7537
rect 27709 7528 27721 7531
rect 27672 7500 27721 7528
rect 27672 7488 27678 7500
rect 27709 7497 27721 7500
rect 27755 7497 27767 7531
rect 27709 7491 27767 7497
rect 27890 7488 27896 7540
rect 27948 7528 27954 7540
rect 28353 7531 28411 7537
rect 28353 7528 28365 7531
rect 27948 7500 28365 7528
rect 27948 7488 27954 7500
rect 28353 7497 28365 7500
rect 28399 7497 28411 7531
rect 29454 7528 29460 7540
rect 29415 7500 29460 7528
rect 28353 7491 28411 7497
rect 29454 7488 29460 7500
rect 29512 7488 29518 7540
rect 29730 7488 29736 7540
rect 29788 7528 29794 7540
rect 31297 7531 31355 7537
rect 31297 7528 31309 7531
rect 29788 7500 31309 7528
rect 29788 7488 29794 7500
rect 31297 7497 31309 7500
rect 31343 7528 31355 7531
rect 32122 7528 32128 7540
rect 31343 7500 32128 7528
rect 31343 7497 31355 7500
rect 31297 7491 31355 7497
rect 32122 7488 32128 7500
rect 32180 7488 32186 7540
rect 33134 7488 33140 7540
rect 33192 7528 33198 7540
rect 33410 7528 33416 7540
rect 33192 7500 33416 7528
rect 33192 7488 33198 7500
rect 33410 7488 33416 7500
rect 33468 7488 33474 7540
rect 33505 7531 33563 7537
rect 33505 7497 33517 7531
rect 33551 7528 33563 7531
rect 33594 7528 33600 7540
rect 33551 7500 33600 7528
rect 33551 7497 33563 7500
rect 33505 7491 33563 7497
rect 33594 7488 33600 7500
rect 33652 7488 33658 7540
rect 34238 7528 34244 7540
rect 34199 7500 34244 7528
rect 34238 7488 34244 7500
rect 34296 7488 34302 7540
rect 36081 7531 36139 7537
rect 36081 7497 36093 7531
rect 36127 7528 36139 7531
rect 36262 7528 36268 7540
rect 36127 7500 36268 7528
rect 36127 7497 36139 7500
rect 36081 7491 36139 7497
rect 36262 7488 36268 7500
rect 36320 7488 36326 7540
rect 37826 7488 37832 7540
rect 37884 7528 37890 7540
rect 38749 7531 38807 7537
rect 38749 7528 38761 7531
rect 37884 7500 38761 7528
rect 37884 7488 37890 7500
rect 38749 7497 38761 7500
rect 38795 7497 38807 7531
rect 39298 7528 39304 7540
rect 39259 7500 39304 7528
rect 38749 7491 38807 7497
rect 39298 7488 39304 7500
rect 39356 7488 39362 7540
rect 20993 7432 23152 7460
rect 23477 7463 23535 7469
rect 20993 7429 21005 7432
rect 20947 7423 21005 7429
rect 23477 7429 23489 7463
rect 23523 7460 23535 7463
rect 23750 7460 23756 7472
rect 23523 7432 23756 7460
rect 23523 7429 23535 7432
rect 23477 7423 23535 7429
rect 23750 7420 23756 7432
rect 23808 7420 23814 7472
rect 25547 7463 25605 7469
rect 25547 7429 25559 7463
rect 25593 7460 25605 7463
rect 26602 7460 26608 7472
rect 25593 7432 26608 7460
rect 25593 7429 25605 7432
rect 25547 7423 25605 7429
rect 26602 7420 26608 7432
rect 26660 7460 26666 7472
rect 27985 7463 28043 7469
rect 27985 7460 27997 7463
rect 26660 7432 27997 7460
rect 26660 7420 26666 7432
rect 27985 7429 27997 7432
rect 28031 7429 28043 7463
rect 27985 7423 28043 7429
rect 28810 7420 28816 7472
rect 28868 7460 28874 7472
rect 29917 7463 29975 7469
rect 29917 7460 29929 7463
rect 28868 7432 29929 7460
rect 28868 7420 28874 7432
rect 29917 7429 29929 7432
rect 29963 7429 29975 7463
rect 31662 7460 31668 7472
rect 31623 7432 31668 7460
rect 29917 7423 29975 7429
rect 21082 7352 21088 7404
rect 21140 7392 21146 7404
rect 21361 7395 21419 7401
rect 21361 7392 21373 7395
rect 21140 7364 21373 7392
rect 21140 7352 21146 7364
rect 21361 7361 21373 7364
rect 21407 7392 21419 7395
rect 21634 7392 21640 7404
rect 21407 7364 21640 7392
rect 21407 7361 21419 7364
rect 21361 7355 21419 7361
rect 21634 7352 21640 7364
rect 21692 7352 21698 7404
rect 21818 7392 21824 7404
rect 21779 7364 21824 7392
rect 21818 7352 21824 7364
rect 21876 7352 21882 7404
rect 23658 7392 23664 7404
rect 23619 7364 23664 7392
rect 23658 7352 23664 7364
rect 23716 7352 23722 7404
rect 20806 7324 20812 7336
rect 20767 7296 20812 7324
rect 20806 7284 20812 7296
rect 20864 7284 20870 7336
rect 22741 7327 22799 7333
rect 22741 7293 22753 7327
rect 22787 7324 22799 7327
rect 24486 7324 24492 7336
rect 22787 7296 24492 7324
rect 22787 7293 22799 7296
rect 22741 7287 22799 7293
rect 24486 7284 24492 7296
rect 24544 7284 24550 7336
rect 24581 7327 24639 7333
rect 24581 7293 24593 7327
rect 24627 7324 24639 7327
rect 25444 7327 25502 7333
rect 25444 7324 25456 7327
rect 24627 7296 25456 7324
rect 24627 7293 24639 7296
rect 24581 7287 24639 7293
rect 25444 7293 25456 7296
rect 25490 7324 25502 7327
rect 25869 7327 25927 7333
rect 25869 7324 25881 7327
rect 25490 7296 25881 7324
rect 25490 7293 25502 7296
rect 25444 7287 25502 7293
rect 25869 7293 25881 7296
rect 25915 7293 25927 7327
rect 26786 7324 26792 7336
rect 26747 7296 26792 7324
rect 25869 7287 25927 7293
rect 26786 7284 26792 7296
rect 26844 7284 26850 7336
rect 29932 7324 29960 7423
rect 31662 7420 31668 7432
rect 31720 7420 31726 7472
rect 32769 7463 32827 7469
rect 32769 7429 32781 7463
rect 32815 7460 32827 7463
rect 35802 7460 35808 7472
rect 32815 7432 35808 7460
rect 32815 7429 32827 7432
rect 32769 7423 32827 7429
rect 35802 7420 35808 7432
rect 35860 7420 35866 7472
rect 36817 7463 36875 7469
rect 36817 7429 36829 7463
rect 36863 7460 36875 7463
rect 37274 7460 37280 7472
rect 36863 7432 37280 7460
rect 36863 7429 36875 7432
rect 36817 7423 36875 7429
rect 37274 7420 37280 7432
rect 37332 7460 37338 7472
rect 38102 7460 38108 7472
rect 37332 7432 38108 7460
rect 37332 7420 37338 7432
rect 38102 7420 38108 7432
rect 38160 7420 38166 7472
rect 36265 7395 36323 7401
rect 36265 7361 36277 7395
rect 36311 7392 36323 7395
rect 36354 7392 36360 7404
rect 36311 7364 36360 7392
rect 36311 7361 36323 7364
rect 36265 7355 36323 7361
rect 36354 7352 36360 7364
rect 36412 7352 36418 7404
rect 37645 7395 37703 7401
rect 37645 7361 37657 7395
rect 37691 7392 37703 7395
rect 37737 7395 37795 7401
rect 37737 7392 37749 7395
rect 37691 7364 37749 7392
rect 37691 7361 37703 7364
rect 37645 7355 37703 7361
rect 37737 7361 37749 7364
rect 37783 7392 37795 7395
rect 37918 7392 37924 7404
rect 37783 7364 37924 7392
rect 37783 7361 37795 7364
rect 37737 7355 37795 7361
rect 37918 7352 37924 7364
rect 37976 7352 37982 7404
rect 30101 7327 30159 7333
rect 30101 7324 30113 7327
rect 29932 7296 30113 7324
rect 30101 7293 30113 7296
rect 30147 7293 30159 7327
rect 30558 7324 30564 7336
rect 30519 7296 30564 7324
rect 30101 7287 30159 7293
rect 30558 7284 30564 7296
rect 30616 7284 30622 7336
rect 31846 7324 31852 7336
rect 31807 7296 31852 7324
rect 31846 7284 31852 7296
rect 31904 7284 31910 7336
rect 33594 7324 33600 7336
rect 33555 7296 33600 7324
rect 33594 7284 33600 7296
rect 33652 7324 33658 7336
rect 34920 7327 34978 7333
rect 34920 7324 34932 7327
rect 33652 7296 34932 7324
rect 33652 7284 33658 7296
rect 34920 7293 34932 7296
rect 34966 7324 34978 7327
rect 35345 7327 35403 7333
rect 35345 7324 35357 7327
rect 34966 7296 35357 7324
rect 34966 7293 34978 7296
rect 34920 7287 34978 7293
rect 35345 7293 35357 7296
rect 35391 7293 35403 7327
rect 35345 7287 35403 7293
rect 37277 7327 37335 7333
rect 37277 7293 37289 7327
rect 37323 7324 37335 7327
rect 38194 7324 38200 7336
rect 37323 7296 38200 7324
rect 37323 7293 37335 7296
rect 37277 7287 37335 7293
rect 38194 7284 38200 7296
rect 38252 7284 38258 7336
rect 20073 7259 20131 7265
rect 19024 7228 19472 7256
rect 19024 7216 19030 7228
rect 13541 7191 13599 7197
rect 13541 7188 13553 7191
rect 13320 7160 13553 7188
rect 13320 7148 13326 7160
rect 13541 7157 13553 7160
rect 13587 7188 13599 7191
rect 13633 7191 13691 7197
rect 13633 7188 13645 7191
rect 13587 7160 13645 7188
rect 13587 7157 13599 7160
rect 13541 7151 13599 7157
rect 13633 7157 13645 7160
rect 13679 7157 13691 7191
rect 13633 7151 13691 7157
rect 16761 7191 16819 7197
rect 16761 7157 16773 7191
rect 16807 7188 16819 7191
rect 19334 7188 19340 7200
rect 16807 7160 19340 7188
rect 16807 7157 16819 7160
rect 16761 7151 16819 7157
rect 19334 7148 19340 7160
rect 19392 7148 19398 7200
rect 19444 7197 19472 7228
rect 20073 7225 20085 7259
rect 20119 7256 20131 7259
rect 20119 7228 23474 7256
rect 20119 7225 20131 7228
rect 20073 7219 20131 7225
rect 19429 7191 19487 7197
rect 19429 7157 19441 7191
rect 19475 7188 19487 7191
rect 19978 7188 19984 7200
rect 19475 7160 19984 7188
rect 19475 7157 19487 7160
rect 19429 7151 19487 7157
rect 19978 7148 19984 7160
rect 20036 7188 20042 7200
rect 21542 7188 21548 7200
rect 20036 7160 21548 7188
rect 20036 7148 20042 7160
rect 21542 7148 21548 7160
rect 21600 7148 21606 7200
rect 22189 7191 22247 7197
rect 22189 7157 22201 7191
rect 22235 7188 22247 7191
rect 22278 7188 22284 7200
rect 22235 7160 22284 7188
rect 22235 7157 22247 7160
rect 22189 7151 22247 7157
rect 22278 7148 22284 7160
rect 22336 7148 22342 7200
rect 23446 7188 23474 7228
rect 23750 7216 23756 7268
rect 23808 7256 23814 7268
rect 24023 7259 24081 7265
rect 24023 7256 24035 7259
rect 23808 7228 24035 7256
rect 23808 7216 23814 7228
rect 24023 7225 24035 7228
rect 24069 7256 24081 7259
rect 27042 7259 27100 7265
rect 27042 7256 27054 7259
rect 24069 7228 27054 7256
rect 24069 7225 24081 7228
rect 24023 7219 24081 7225
rect 27042 7225 27054 7228
rect 27088 7256 27100 7259
rect 27154 7256 27160 7268
rect 27088 7228 27160 7256
rect 27088 7225 27100 7228
rect 27042 7219 27100 7225
rect 27154 7216 27160 7228
rect 27212 7216 27218 7268
rect 30834 7256 30840 7268
rect 30795 7228 30840 7256
rect 30834 7216 30840 7228
rect 30892 7216 30898 7268
rect 31662 7216 31668 7268
rect 31720 7256 31726 7268
rect 32170 7259 32228 7265
rect 32170 7256 32182 7259
rect 31720 7228 32182 7256
rect 31720 7216 31726 7228
rect 32170 7225 32182 7228
rect 32216 7256 32228 7259
rect 32490 7256 32496 7268
rect 32216 7228 32496 7256
rect 32216 7225 32228 7228
rect 32170 7219 32228 7225
rect 32490 7216 32496 7228
rect 32548 7216 32554 7268
rect 36354 7216 36360 7268
rect 36412 7256 36418 7268
rect 36412 7228 36457 7256
rect 36412 7216 36418 7228
rect 26326 7188 26332 7200
rect 23446 7160 26332 7188
rect 26326 7148 26332 7160
rect 26384 7148 26390 7200
rect 26694 7148 26700 7200
rect 26752 7188 26758 7200
rect 28994 7188 29000 7200
rect 26752 7160 29000 7188
rect 26752 7148 26758 7160
rect 28994 7148 29000 7160
rect 29052 7148 29058 7200
rect 33778 7188 33784 7200
rect 33739 7160 33784 7188
rect 33778 7148 33784 7160
rect 33836 7148 33842 7200
rect 34514 7188 34520 7200
rect 34475 7160 34520 7188
rect 34514 7148 34520 7160
rect 34572 7148 34578 7200
rect 34606 7148 34612 7200
rect 34664 7188 34670 7200
rect 35023 7191 35081 7197
rect 35023 7188 35035 7191
rect 34664 7160 35035 7188
rect 34664 7148 34670 7160
rect 35023 7157 35035 7160
rect 35069 7157 35081 7191
rect 35023 7151 35081 7157
rect 1104 7098 48852 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 48852 7098
rect 1104 7024 48852 7046
rect 9493 6987 9551 6993
rect 9493 6953 9505 6987
rect 9539 6984 9551 6987
rect 9950 6984 9956 6996
rect 9539 6956 9956 6984
rect 9539 6953 9551 6956
rect 9493 6947 9551 6953
rect 9950 6944 9956 6956
rect 10008 6984 10014 6996
rect 10045 6987 10103 6993
rect 10045 6984 10057 6987
rect 10008 6956 10057 6984
rect 10008 6944 10014 6956
rect 10045 6953 10057 6956
rect 10091 6953 10103 6987
rect 10045 6947 10103 6953
rect 10594 6944 10600 6996
rect 10652 6984 10658 6996
rect 10965 6987 11023 6993
rect 10965 6984 10977 6987
rect 10652 6956 10977 6984
rect 10652 6944 10658 6956
rect 10965 6953 10977 6956
rect 11011 6953 11023 6987
rect 10965 6947 11023 6953
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 12529 6987 12587 6993
rect 12529 6984 12541 6987
rect 12492 6956 12541 6984
rect 12492 6944 12498 6956
rect 12529 6953 12541 6956
rect 12575 6953 12587 6987
rect 12529 6947 12587 6953
rect 14139 6987 14197 6993
rect 14139 6953 14151 6987
rect 14185 6984 14197 6987
rect 14366 6984 14372 6996
rect 14185 6956 14372 6984
rect 14185 6953 14197 6956
rect 14139 6947 14197 6953
rect 14366 6944 14372 6956
rect 14424 6944 14430 6996
rect 15562 6944 15568 6996
rect 15620 6984 15626 6996
rect 16025 6987 16083 6993
rect 16025 6984 16037 6987
rect 15620 6956 16037 6984
rect 15620 6944 15626 6956
rect 16025 6953 16037 6956
rect 16071 6953 16083 6987
rect 16025 6947 16083 6953
rect 16206 6944 16212 6996
rect 16264 6984 16270 6996
rect 16393 6987 16451 6993
rect 16393 6984 16405 6987
rect 16264 6956 16405 6984
rect 16264 6944 16270 6956
rect 16393 6953 16405 6956
rect 16439 6953 16451 6987
rect 16393 6947 16451 6953
rect 17497 6987 17555 6993
rect 17497 6953 17509 6987
rect 17543 6984 17555 6987
rect 19426 6984 19432 6996
rect 17543 6956 18552 6984
rect 19387 6956 19432 6984
rect 17543 6953 17555 6956
rect 17497 6947 17555 6953
rect 18524 6928 18552 6956
rect 19426 6944 19432 6956
rect 19484 6944 19490 6996
rect 22830 6944 22836 6996
rect 22888 6984 22894 6996
rect 22925 6987 22983 6993
rect 22925 6984 22937 6987
rect 22888 6956 22937 6984
rect 22888 6944 22894 6956
rect 22925 6953 22937 6956
rect 22971 6953 22983 6987
rect 22925 6947 22983 6953
rect 23658 6944 23664 6996
rect 23716 6984 23722 6996
rect 23753 6987 23811 6993
rect 23753 6984 23765 6987
rect 23716 6956 23765 6984
rect 23716 6944 23722 6956
rect 23753 6953 23765 6956
rect 23799 6953 23811 6987
rect 23753 6947 23811 6953
rect 24302 6944 24308 6996
rect 24360 6984 24366 6996
rect 24489 6987 24547 6993
rect 24489 6984 24501 6987
rect 24360 6956 24501 6984
rect 24360 6944 24366 6956
rect 24489 6953 24501 6956
rect 24535 6953 24547 6987
rect 24489 6947 24547 6953
rect 25179 6987 25237 6993
rect 25179 6953 25191 6987
rect 25225 6984 25237 6987
rect 25682 6984 25688 6996
rect 25225 6956 25688 6984
rect 25225 6953 25237 6956
rect 25179 6947 25237 6953
rect 25682 6944 25688 6956
rect 25740 6944 25746 6996
rect 26329 6987 26387 6993
rect 26329 6953 26341 6987
rect 26375 6984 26387 6987
rect 26605 6987 26663 6993
rect 26605 6984 26617 6987
rect 26375 6956 26617 6984
rect 26375 6953 26387 6956
rect 26329 6947 26387 6953
rect 26605 6953 26617 6956
rect 26651 6984 26663 6987
rect 26786 6984 26792 6996
rect 26651 6956 26792 6984
rect 26651 6953 26663 6956
rect 26605 6947 26663 6953
rect 26786 6944 26792 6956
rect 26844 6944 26850 6996
rect 27709 6987 27767 6993
rect 27709 6953 27721 6987
rect 27755 6984 27767 6987
rect 27982 6984 27988 6996
rect 27755 6956 27988 6984
rect 27755 6953 27767 6956
rect 27709 6947 27767 6953
rect 27982 6944 27988 6956
rect 28040 6944 28046 6996
rect 30282 6984 30288 6996
rect 30243 6956 30288 6984
rect 30282 6944 30288 6956
rect 30340 6944 30346 6996
rect 31294 6984 31300 6996
rect 31207 6956 31300 6984
rect 31294 6944 31300 6956
rect 31352 6984 31358 6996
rect 32214 6984 32220 6996
rect 31352 6956 32220 6984
rect 31352 6944 31358 6956
rect 32214 6944 32220 6956
rect 32272 6944 32278 6996
rect 32490 6984 32496 6996
rect 32451 6956 32496 6984
rect 32490 6944 32496 6956
rect 32548 6944 32554 6996
rect 33045 6987 33103 6993
rect 33045 6953 33057 6987
rect 33091 6984 33103 6987
rect 33091 6956 34871 6984
rect 33091 6953 33103 6956
rect 33045 6947 33103 6953
rect 16482 6876 16488 6928
rect 16540 6916 16546 6928
rect 16898 6919 16956 6925
rect 16898 6916 16910 6919
rect 16540 6888 16910 6916
rect 16540 6876 16546 6888
rect 16898 6885 16910 6888
rect 16944 6885 16956 6919
rect 16898 6879 16956 6885
rect 17862 6876 17868 6928
rect 17920 6916 17926 6928
rect 18049 6919 18107 6925
rect 18049 6916 18061 6919
rect 17920 6888 18061 6916
rect 17920 6876 17926 6888
rect 18049 6885 18061 6888
rect 18095 6885 18107 6919
rect 18506 6916 18512 6928
rect 18419 6888 18512 6916
rect 18049 6879 18107 6885
rect 18506 6876 18512 6888
rect 18564 6876 18570 6928
rect 22091 6919 22149 6925
rect 22091 6885 22103 6919
rect 22137 6916 22149 6919
rect 22278 6916 22284 6928
rect 22137 6888 22284 6916
rect 22137 6885 22149 6888
rect 22091 6879 22149 6885
rect 22278 6876 22284 6888
rect 22336 6876 22342 6928
rect 28813 6919 28871 6925
rect 28813 6885 28825 6919
rect 28859 6916 28871 6919
rect 28902 6916 28908 6928
rect 28859 6888 28908 6916
rect 28859 6885 28871 6888
rect 28813 6879 28871 6885
rect 28902 6876 28908 6888
rect 28960 6876 28966 6928
rect 34057 6919 34115 6925
rect 34057 6885 34069 6919
rect 34103 6916 34115 6919
rect 34330 6916 34336 6928
rect 34103 6888 34336 6916
rect 34103 6885 34115 6888
rect 34057 6879 34115 6885
rect 34330 6876 34336 6888
rect 34388 6876 34394 6928
rect 10226 6848 10232 6860
rect 10187 6820 10232 6848
rect 10226 6808 10232 6820
rect 10284 6808 10290 6860
rect 10502 6848 10508 6860
rect 10463 6820 10508 6848
rect 10502 6808 10508 6820
rect 10560 6808 10566 6860
rect 12710 6848 12716 6860
rect 12671 6820 12716 6848
rect 12710 6808 12716 6820
rect 12768 6808 12774 6860
rect 12897 6851 12955 6857
rect 12897 6817 12909 6851
rect 12943 6817 12955 6851
rect 12897 6811 12955 6817
rect 10520 6780 10548 6808
rect 12526 6780 12532 6792
rect 10520 6752 12532 6780
rect 12526 6740 12532 6752
rect 12584 6780 12590 6792
rect 12912 6780 12940 6811
rect 13630 6808 13636 6860
rect 13688 6848 13694 6860
rect 14036 6851 14094 6857
rect 14036 6848 14048 6851
rect 13688 6820 14048 6848
rect 13688 6808 13694 6820
rect 14036 6817 14048 6820
rect 14082 6817 14094 6851
rect 14036 6811 14094 6817
rect 15565 6851 15623 6857
rect 15565 6817 15577 6851
rect 15611 6848 15623 6851
rect 15611 6820 18276 6848
rect 15611 6817 15623 6820
rect 15565 6811 15623 6817
rect 16022 6780 16028 6792
rect 12584 6752 16028 6780
rect 12584 6740 12590 6752
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 16574 6780 16580 6792
rect 16535 6752 16580 6780
rect 16574 6740 16580 6752
rect 16632 6740 16638 6792
rect 18248 6780 18276 6820
rect 20806 6808 20812 6860
rect 20864 6848 20870 6860
rect 21177 6851 21235 6857
rect 21177 6848 21189 6851
rect 20864 6820 21189 6848
rect 20864 6808 20870 6820
rect 21177 6817 21189 6820
rect 21223 6848 21235 6851
rect 22649 6851 22707 6857
rect 22649 6848 22661 6851
rect 21223 6820 22661 6848
rect 21223 6817 21235 6820
rect 21177 6811 21235 6817
rect 22649 6817 22661 6820
rect 22695 6817 22707 6851
rect 22649 6811 22707 6817
rect 23474 6808 23480 6860
rect 23532 6848 23538 6860
rect 23934 6848 23940 6860
rect 23532 6820 23577 6848
rect 23895 6820 23940 6848
rect 23532 6808 23538 6820
rect 23934 6808 23940 6820
rect 23992 6808 23998 6860
rect 24486 6808 24492 6860
rect 24544 6848 24550 6860
rect 25076 6851 25134 6857
rect 25076 6848 25088 6851
rect 24544 6820 25088 6848
rect 24544 6808 24550 6820
rect 25076 6817 25088 6820
rect 25122 6848 25134 6851
rect 25498 6848 25504 6860
rect 25122 6820 25504 6848
rect 25122 6817 25134 6820
rect 25076 6811 25134 6817
rect 25498 6808 25504 6820
rect 25556 6808 25562 6860
rect 26510 6848 26516 6860
rect 26471 6820 26516 6848
rect 26510 6808 26516 6820
rect 26568 6808 26574 6860
rect 26694 6808 26700 6860
rect 26752 6848 26758 6860
rect 26973 6851 27031 6857
rect 26973 6848 26985 6851
rect 26752 6820 26985 6848
rect 26752 6808 26758 6820
rect 26973 6817 26985 6820
rect 27019 6817 27031 6851
rect 26973 6811 27031 6817
rect 29454 6808 29460 6860
rect 29512 6848 29518 6860
rect 30190 6848 30196 6860
rect 29512 6820 30196 6848
rect 29512 6808 29518 6820
rect 30190 6808 30196 6820
rect 30248 6808 30254 6860
rect 30558 6808 30564 6860
rect 30616 6848 30622 6860
rect 30653 6851 30711 6857
rect 30653 6848 30665 6851
rect 30616 6820 30665 6848
rect 30616 6808 30622 6820
rect 30653 6817 30665 6820
rect 30699 6817 30711 6851
rect 30653 6811 30711 6817
rect 30834 6808 30840 6860
rect 30892 6848 30898 6860
rect 31938 6848 31944 6860
rect 30892 6820 31944 6848
rect 30892 6808 30898 6820
rect 31938 6808 31944 6820
rect 31996 6848 32002 6860
rect 32125 6851 32183 6857
rect 32125 6848 32137 6851
rect 31996 6820 32137 6848
rect 31996 6808 32002 6820
rect 32125 6817 32137 6820
rect 32171 6817 32183 6851
rect 34843 6848 34871 6956
rect 36170 6944 36176 6996
rect 36228 6984 36234 6996
rect 37001 6987 37059 6993
rect 37001 6984 37013 6987
rect 36228 6956 37013 6984
rect 36228 6944 36234 6956
rect 37001 6953 37013 6956
rect 37047 6953 37059 6987
rect 37001 6947 37059 6953
rect 35802 6876 35808 6928
rect 35860 6916 35866 6928
rect 36357 6919 36415 6925
rect 36357 6916 36369 6919
rect 35860 6888 36369 6916
rect 35860 6876 35866 6888
rect 36357 6885 36369 6888
rect 36403 6916 36415 6919
rect 36906 6916 36912 6928
rect 36403 6888 36912 6916
rect 36403 6885 36415 6888
rect 36357 6879 36415 6885
rect 36906 6876 36912 6888
rect 36964 6876 36970 6928
rect 35472 6851 35530 6857
rect 35472 6848 35484 6851
rect 34843 6820 35484 6848
rect 32125 6811 32183 6817
rect 35472 6817 35484 6820
rect 35518 6848 35530 6851
rect 35894 6848 35900 6860
rect 35518 6820 35900 6848
rect 35518 6817 35530 6820
rect 35472 6811 35530 6817
rect 35894 6808 35900 6820
rect 35952 6808 35958 6860
rect 38381 6851 38439 6857
rect 38381 6817 38393 6851
rect 38427 6848 38439 6851
rect 38470 6848 38476 6860
rect 38427 6820 38476 6848
rect 38427 6817 38439 6820
rect 38381 6811 38439 6817
rect 38470 6808 38476 6820
rect 38528 6808 38534 6860
rect 18417 6783 18475 6789
rect 18417 6780 18429 6783
rect 18248 6752 18429 6780
rect 18417 6749 18429 6752
rect 18463 6780 18475 6783
rect 19058 6780 19064 6792
rect 18463 6752 19064 6780
rect 18463 6749 18475 6752
rect 18417 6743 18475 6749
rect 19058 6740 19064 6752
rect 19116 6740 19122 6792
rect 21729 6783 21787 6789
rect 21729 6749 21741 6783
rect 21775 6749 21787 6783
rect 28718 6780 28724 6792
rect 28679 6752 28724 6780
rect 21729 6743 21787 6749
rect 16942 6672 16948 6724
rect 17000 6712 17006 6724
rect 18969 6715 19027 6721
rect 18969 6712 18981 6715
rect 17000 6684 18981 6712
rect 17000 6672 17006 6684
rect 18969 6681 18981 6684
rect 19015 6681 19027 6715
rect 18969 6675 19027 6681
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 11977 6647 12035 6653
rect 11977 6644 11989 6647
rect 11296 6616 11989 6644
rect 11296 6604 11302 6616
rect 11977 6613 11989 6616
rect 12023 6644 12035 6647
rect 12066 6644 12072 6656
rect 12023 6616 12072 6644
rect 12023 6613 12035 6616
rect 11977 6607 12035 6613
rect 12066 6604 12072 6616
rect 12124 6604 12130 6656
rect 21358 6604 21364 6656
rect 21416 6644 21422 6656
rect 21545 6647 21603 6653
rect 21545 6644 21557 6647
rect 21416 6616 21557 6644
rect 21416 6604 21422 6616
rect 21545 6613 21557 6616
rect 21591 6644 21603 6647
rect 21744 6644 21772 6743
rect 28718 6740 28724 6752
rect 28776 6740 28782 6792
rect 29365 6783 29423 6789
rect 29365 6749 29377 6783
rect 29411 6780 29423 6783
rect 30006 6780 30012 6792
rect 29411 6752 30012 6780
rect 29411 6749 29423 6752
rect 29365 6743 29423 6749
rect 30006 6740 30012 6752
rect 30064 6740 30070 6792
rect 33781 6783 33839 6789
rect 33781 6749 33793 6783
rect 33827 6780 33839 6783
rect 33965 6783 34023 6789
rect 33965 6780 33977 6783
rect 33827 6752 33977 6780
rect 33827 6749 33839 6752
rect 33781 6743 33839 6749
rect 33965 6749 33977 6752
rect 34011 6780 34023 6783
rect 35575 6783 35633 6789
rect 35575 6780 35587 6783
rect 34011 6752 35587 6780
rect 34011 6749 34023 6752
rect 33965 6743 34023 6749
rect 35575 6749 35587 6752
rect 35621 6749 35633 6783
rect 35575 6743 35633 6749
rect 36265 6783 36323 6789
rect 36265 6749 36277 6783
rect 36311 6780 36323 6783
rect 36354 6780 36360 6792
rect 36311 6752 36360 6780
rect 36311 6749 36323 6752
rect 36265 6743 36323 6749
rect 36354 6740 36360 6752
rect 36412 6780 36418 6792
rect 37737 6783 37795 6789
rect 37737 6780 37749 6783
rect 36412 6752 37749 6780
rect 36412 6740 36418 6752
rect 37737 6749 37749 6752
rect 37783 6749 37795 6783
rect 37737 6743 37795 6749
rect 34054 6672 34060 6724
rect 34112 6712 34118 6724
rect 34517 6715 34575 6721
rect 34517 6712 34529 6715
rect 34112 6684 34529 6712
rect 34112 6672 34118 6684
rect 34517 6681 34529 6684
rect 34563 6681 34575 6715
rect 36587 6715 36645 6721
rect 36587 6712 36599 6715
rect 34517 6675 34575 6681
rect 35820 6684 36599 6712
rect 29638 6644 29644 6656
rect 21591 6616 21772 6644
rect 29599 6616 29644 6644
rect 21591 6613 21603 6616
rect 21545 6607 21603 6613
rect 29638 6604 29644 6616
rect 29696 6604 29702 6656
rect 31846 6604 31852 6656
rect 31904 6644 31910 6656
rect 31941 6647 31999 6653
rect 31941 6644 31953 6647
rect 31904 6616 31953 6644
rect 31904 6604 31910 6616
rect 31941 6613 31953 6616
rect 31987 6644 31999 6647
rect 32766 6644 32772 6656
rect 31987 6616 32772 6644
rect 31987 6613 31999 6616
rect 31941 6607 31999 6613
rect 32766 6604 32772 6616
rect 32824 6604 32830 6656
rect 33318 6604 33324 6656
rect 33376 6644 33382 6656
rect 35820 6644 35848 6684
rect 36587 6681 36599 6684
rect 36633 6681 36645 6715
rect 36587 6675 36645 6681
rect 33376 6616 35848 6644
rect 33376 6604 33382 6616
rect 1104 6554 48852 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 48852 6554
rect 1104 6480 48852 6502
rect 9309 6443 9367 6449
rect 9309 6409 9321 6443
rect 9355 6440 9367 6443
rect 10502 6440 10508 6452
rect 9355 6412 10508 6440
rect 9355 6409 9367 6412
rect 9309 6403 9367 6409
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6440 12311 6443
rect 12710 6440 12716 6452
rect 12299 6412 12716 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 14734 6440 14740 6452
rect 14695 6412 14740 6440
rect 14734 6400 14740 6412
rect 14792 6400 14798 6452
rect 19058 6440 19064 6452
rect 19019 6412 19064 6440
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 21821 6443 21879 6449
rect 21821 6409 21833 6443
rect 21867 6440 21879 6443
rect 22278 6440 22284 6452
rect 21867 6412 22284 6440
rect 21867 6409 21879 6412
rect 21821 6403 21879 6409
rect 22278 6400 22284 6412
rect 22336 6400 22342 6452
rect 23474 6400 23480 6452
rect 23532 6440 23538 6452
rect 23845 6443 23903 6449
rect 23845 6440 23857 6443
rect 23532 6412 23857 6440
rect 23532 6400 23538 6412
rect 23845 6409 23857 6412
rect 23891 6409 23903 6443
rect 25498 6440 25504 6452
rect 25459 6412 25504 6440
rect 23845 6403 23903 6409
rect 25498 6400 25504 6412
rect 25556 6400 25562 6452
rect 25958 6440 25964 6452
rect 25919 6412 25964 6440
rect 25958 6400 25964 6412
rect 26016 6400 26022 6452
rect 27522 6440 27528 6452
rect 27483 6412 27528 6440
rect 27522 6400 27528 6412
rect 27580 6400 27586 6452
rect 30190 6400 30196 6452
rect 30248 6440 30254 6452
rect 30285 6443 30343 6449
rect 30285 6440 30297 6443
rect 30248 6412 30297 6440
rect 30248 6400 30254 6412
rect 30285 6409 30297 6412
rect 30331 6409 30343 6443
rect 30834 6440 30840 6452
rect 30747 6412 30840 6440
rect 30285 6403 30343 6409
rect 30834 6400 30840 6412
rect 30892 6440 30898 6452
rect 31662 6440 31668 6452
rect 30892 6412 31668 6440
rect 30892 6400 30898 6412
rect 10045 6375 10103 6381
rect 10045 6341 10057 6375
rect 10091 6372 10103 6375
rect 10226 6372 10232 6384
rect 10091 6344 10232 6372
rect 10091 6341 10103 6344
rect 10045 6335 10103 6341
rect 10226 6332 10232 6344
rect 10284 6372 10290 6384
rect 15378 6372 15384 6384
rect 10284 6344 15384 6372
rect 10284 6332 10290 6344
rect 10428 6245 10456 6344
rect 15378 6332 15384 6344
rect 15436 6372 15442 6384
rect 15841 6375 15899 6381
rect 15841 6372 15853 6375
rect 15436 6344 15853 6372
rect 15436 6332 15442 6344
rect 15841 6341 15853 6344
rect 15887 6341 15899 6375
rect 15841 6335 15899 6341
rect 12529 6307 12587 6313
rect 12529 6273 12541 6307
rect 12575 6304 12587 6307
rect 12802 6304 12808 6316
rect 12575 6276 12808 6304
rect 12575 6273 12587 6276
rect 12529 6267 12587 6273
rect 12802 6264 12808 6276
rect 12860 6264 12866 6316
rect 10413 6239 10471 6245
rect 10413 6205 10425 6239
rect 10459 6205 10471 6239
rect 10413 6199 10471 6205
rect 10597 6239 10655 6245
rect 10597 6205 10609 6239
rect 10643 6205 10655 6239
rect 14553 6239 14611 6245
rect 14553 6236 14565 6239
rect 10597 6199 10655 6205
rect 14384 6208 14565 6236
rect 9677 6171 9735 6177
rect 9677 6137 9689 6171
rect 9723 6168 9735 6171
rect 10612 6168 10640 6199
rect 10686 6168 10692 6180
rect 9723 6140 10692 6168
rect 9723 6137 9735 6140
rect 9677 6131 9735 6137
rect 10686 6128 10692 6140
rect 10744 6128 10750 6180
rect 10870 6168 10876 6180
rect 10831 6140 10876 6168
rect 10870 6128 10876 6140
rect 10928 6128 10934 6180
rect 12621 6171 12679 6177
rect 11808 6140 12480 6168
rect 11808 6112 11836 6140
rect 11790 6100 11796 6112
rect 11751 6072 11796 6100
rect 11790 6060 11796 6072
rect 11848 6060 11854 6112
rect 12452 6100 12480 6140
rect 12621 6137 12633 6171
rect 12667 6137 12679 6171
rect 12621 6131 12679 6137
rect 13173 6171 13231 6177
rect 13173 6137 13185 6171
rect 13219 6168 13231 6171
rect 13630 6168 13636 6180
rect 13219 6140 13636 6168
rect 13219 6137 13231 6140
rect 13173 6131 13231 6137
rect 12636 6100 12664 6131
rect 13630 6128 13636 6140
rect 13688 6168 13694 6180
rect 13909 6171 13967 6177
rect 13909 6168 13921 6171
rect 13688 6140 13921 6168
rect 13688 6128 13694 6140
rect 13909 6137 13921 6140
rect 13955 6137 13967 6171
rect 13909 6131 13967 6137
rect 14384 6112 14412 6208
rect 14553 6205 14565 6208
rect 14599 6236 14611 6239
rect 15746 6236 15752 6248
rect 14599 6208 15752 6236
rect 14599 6205 14611 6208
rect 14553 6199 14611 6205
rect 15746 6196 15752 6208
rect 15804 6196 15810 6248
rect 15856 6236 15884 6335
rect 16850 6332 16856 6384
rect 16908 6372 16914 6384
rect 20441 6375 20499 6381
rect 20441 6372 20453 6375
rect 16908 6344 20453 6372
rect 16908 6332 16914 6344
rect 20441 6341 20453 6344
rect 20487 6341 20499 6375
rect 20441 6335 20499 6341
rect 16574 6264 16580 6316
rect 16632 6304 16638 6316
rect 16761 6307 16819 6313
rect 16761 6304 16773 6307
rect 16632 6276 16773 6304
rect 16632 6264 16638 6276
rect 16761 6273 16773 6276
rect 16807 6304 16819 6307
rect 17405 6307 17463 6313
rect 17405 6304 17417 6307
rect 16807 6276 17417 6304
rect 16807 6273 16819 6276
rect 16761 6267 16819 6273
rect 17405 6273 17417 6276
rect 17451 6273 17463 6307
rect 17405 6267 17463 6273
rect 17862 6264 17868 6316
rect 17920 6304 17926 6316
rect 17920 6276 18552 6304
rect 17920 6264 17926 6276
rect 16025 6239 16083 6245
rect 16025 6236 16037 6239
rect 15856 6208 16037 6236
rect 16025 6205 16037 6208
rect 16071 6205 16083 6239
rect 16025 6199 16083 6205
rect 16485 6239 16543 6245
rect 16485 6205 16497 6239
rect 16531 6236 16543 6239
rect 17880 6236 17908 6264
rect 18524 6245 18552 6276
rect 16531 6208 17908 6236
rect 18049 6239 18107 6245
rect 16531 6205 16543 6208
rect 16485 6199 16543 6205
rect 18049 6205 18061 6239
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 18509 6239 18567 6245
rect 18509 6205 18521 6239
rect 18555 6205 18567 6239
rect 18509 6199 18567 6205
rect 19664 6239 19722 6245
rect 19664 6205 19676 6239
rect 19710 6236 19722 6239
rect 20162 6236 20168 6248
rect 19710 6208 20168 6236
rect 19710 6205 19722 6208
rect 19664 6199 19722 6205
rect 15565 6171 15623 6177
rect 15565 6137 15577 6171
rect 15611 6168 15623 6171
rect 16500 6168 16528 6199
rect 18064 6168 18092 6199
rect 20162 6196 20168 6208
rect 20220 6196 20226 6248
rect 20456 6236 20484 6335
rect 23566 6332 23572 6384
rect 23624 6372 23630 6384
rect 24305 6375 24363 6381
rect 24305 6372 24317 6375
rect 23624 6344 24317 6372
rect 23624 6332 23630 6344
rect 24305 6341 24317 6344
rect 24351 6372 24363 6375
rect 26510 6372 26516 6384
rect 24351 6344 26516 6372
rect 24351 6341 24363 6344
rect 24305 6335 24363 6341
rect 21358 6304 21364 6316
rect 21319 6276 21364 6304
rect 21358 6264 21364 6276
rect 21416 6264 21422 6316
rect 23477 6307 23535 6313
rect 23477 6273 23489 6307
rect 23523 6304 23535 6307
rect 23934 6304 23940 6316
rect 23523 6276 23940 6304
rect 23523 6273 23535 6276
rect 23477 6267 23535 6273
rect 23934 6264 23940 6276
rect 23992 6264 23998 6316
rect 20625 6239 20683 6245
rect 20625 6236 20637 6239
rect 20456 6208 20637 6236
rect 20625 6205 20637 6208
rect 20671 6236 20683 6239
rect 20898 6236 20904 6248
rect 20671 6208 20904 6236
rect 20671 6205 20683 6208
rect 20625 6199 20683 6205
rect 20898 6196 20904 6208
rect 20956 6196 20962 6248
rect 21174 6236 21180 6248
rect 21135 6208 21180 6236
rect 21174 6196 21180 6208
rect 21232 6196 21238 6248
rect 21542 6196 21548 6248
rect 21600 6236 21606 6248
rect 22373 6239 22431 6245
rect 22373 6236 22385 6239
rect 21600 6208 22385 6236
rect 21600 6196 21606 6208
rect 22373 6205 22385 6208
rect 22419 6236 22431 6239
rect 23017 6239 23075 6245
rect 23017 6236 23029 6239
rect 22419 6208 23029 6236
rect 22419 6205 22431 6208
rect 22373 6199 22431 6205
rect 23017 6205 23029 6208
rect 23063 6205 23075 6239
rect 24320 6236 24348 6335
rect 26510 6332 26516 6344
rect 26568 6372 26574 6384
rect 27065 6375 27123 6381
rect 27065 6372 27077 6375
rect 26568 6344 27077 6372
rect 26568 6332 26574 6344
rect 27065 6341 27077 6344
rect 27111 6341 27123 6375
rect 27065 6335 27123 6341
rect 27709 6307 27767 6313
rect 27709 6273 27721 6307
rect 27755 6304 27767 6307
rect 27982 6304 27988 6316
rect 27755 6276 27988 6304
rect 27755 6273 27767 6276
rect 27709 6267 27767 6273
rect 27982 6264 27988 6276
rect 28040 6264 28046 6316
rect 28350 6304 28356 6316
rect 28311 6276 28356 6304
rect 28350 6264 28356 6276
rect 28408 6264 28414 6316
rect 29365 6307 29423 6313
rect 29365 6273 29377 6307
rect 29411 6304 29423 6307
rect 29638 6304 29644 6316
rect 29411 6276 29644 6304
rect 29411 6273 29423 6276
rect 29365 6267 29423 6273
rect 29638 6264 29644 6276
rect 29696 6264 29702 6316
rect 30929 6307 30987 6313
rect 30929 6273 30941 6307
rect 30975 6304 30987 6307
rect 31294 6304 31300 6316
rect 30975 6276 31300 6304
rect 30975 6273 30987 6276
rect 30929 6267 30987 6273
rect 31294 6264 31300 6276
rect 31352 6264 31358 6316
rect 24489 6239 24547 6245
rect 24489 6236 24501 6239
rect 24320 6208 24501 6236
rect 23017 6199 23075 6205
rect 24489 6205 24501 6208
rect 24535 6205 24547 6239
rect 24489 6199 24547 6205
rect 24762 6196 24768 6248
rect 24820 6236 24826 6248
rect 25038 6236 25044 6248
rect 24820 6208 25044 6236
rect 24820 6196 24826 6208
rect 25038 6196 25044 6208
rect 25096 6196 25102 6248
rect 25958 6196 25964 6248
rect 26016 6236 26022 6248
rect 26053 6239 26111 6245
rect 26053 6236 26065 6239
rect 26016 6208 26065 6236
rect 26016 6196 26022 6208
rect 26053 6205 26065 6208
rect 26099 6205 26111 6239
rect 26510 6236 26516 6248
rect 26471 6208 26516 6236
rect 26053 6199 26111 6205
rect 26510 6196 26516 6208
rect 26568 6196 26574 6248
rect 26786 6236 26792 6248
rect 26747 6208 26792 6236
rect 26786 6196 26792 6208
rect 26844 6196 26850 6248
rect 15611 6140 16528 6168
rect 17880 6140 18092 6168
rect 19751 6171 19809 6177
rect 15611 6137 15623 6140
rect 15565 6131 15623 6137
rect 17880 6112 17908 6140
rect 19751 6137 19763 6171
rect 19797 6168 19809 6171
rect 19886 6168 19892 6180
rect 19797 6140 19892 6168
rect 19797 6137 19809 6140
rect 19751 6131 19809 6137
rect 19886 6128 19892 6140
rect 19944 6128 19950 6180
rect 20530 6128 20536 6180
rect 20588 6168 20594 6180
rect 22186 6168 22192 6180
rect 20588 6140 22192 6168
rect 20588 6128 20594 6140
rect 22186 6128 22192 6140
rect 22244 6128 22250 6180
rect 25225 6171 25283 6177
rect 25225 6137 25237 6171
rect 25271 6168 25283 6171
rect 26970 6168 26976 6180
rect 25271 6140 26976 6168
rect 25271 6137 25283 6140
rect 25225 6131 25283 6137
rect 26970 6128 26976 6140
rect 27028 6128 27034 6180
rect 27522 6128 27528 6180
rect 27580 6168 27586 6180
rect 27801 6171 27859 6177
rect 27801 6168 27813 6171
rect 27580 6140 27813 6168
rect 27580 6128 27586 6140
rect 27801 6137 27813 6140
rect 27847 6137 27859 6171
rect 27801 6131 27859 6137
rect 29454 6128 29460 6180
rect 29512 6168 29518 6180
rect 30006 6168 30012 6180
rect 29512 6140 29557 6168
rect 29967 6140 30012 6168
rect 29512 6128 29518 6140
rect 30006 6128 30012 6140
rect 30064 6128 30070 6180
rect 31291 6171 31349 6177
rect 31291 6137 31303 6171
rect 31337 6168 31349 6171
rect 31398 6168 31426 6412
rect 31662 6400 31668 6412
rect 31720 6440 31726 6452
rect 32125 6443 32183 6449
rect 32125 6440 32137 6443
rect 31720 6412 32137 6440
rect 31720 6400 31726 6412
rect 32125 6409 32137 6412
rect 32171 6409 32183 6443
rect 32125 6403 32183 6409
rect 33778 6400 33784 6452
rect 33836 6440 33842 6452
rect 34609 6443 34667 6449
rect 34609 6440 34621 6443
rect 33836 6412 34621 6440
rect 33836 6400 33842 6412
rect 34609 6409 34621 6412
rect 34655 6409 34667 6443
rect 35894 6440 35900 6452
rect 35855 6412 35900 6440
rect 34609 6403 34667 6409
rect 32769 6307 32827 6313
rect 32769 6273 32781 6307
rect 32815 6304 32827 6307
rect 33318 6304 33324 6316
rect 32815 6276 33324 6304
rect 32815 6273 32827 6276
rect 32769 6267 32827 6273
rect 33318 6264 33324 6276
rect 33376 6264 33382 6316
rect 34624 6236 34652 6403
rect 35894 6400 35900 6412
rect 35952 6400 35958 6452
rect 36906 6440 36912 6452
rect 36867 6412 36912 6440
rect 36906 6400 36912 6412
rect 36964 6400 36970 6452
rect 37274 6440 37280 6452
rect 37235 6412 37280 6440
rect 37274 6400 37280 6412
rect 37332 6400 37338 6452
rect 38013 6443 38071 6449
rect 38013 6409 38025 6443
rect 38059 6440 38071 6443
rect 38470 6440 38476 6452
rect 38059 6412 38476 6440
rect 38059 6409 38071 6412
rect 38013 6403 38071 6409
rect 38470 6400 38476 6412
rect 38528 6400 38534 6452
rect 34977 6239 35035 6245
rect 34977 6236 34989 6239
rect 34624 6208 34989 6236
rect 34977 6205 34989 6208
rect 35023 6205 35035 6239
rect 34977 6199 35035 6205
rect 36516 6239 36574 6245
rect 36516 6205 36528 6239
rect 36562 6236 36574 6239
rect 37274 6236 37280 6248
rect 36562 6208 37280 6236
rect 36562 6205 36574 6208
rect 36516 6199 36574 6205
rect 37274 6196 37280 6208
rect 37332 6196 37338 6248
rect 37528 6239 37586 6245
rect 37528 6205 37540 6239
rect 37574 6236 37586 6239
rect 38286 6236 38292 6248
rect 37574 6208 38292 6236
rect 37574 6205 37586 6208
rect 37528 6199 37586 6205
rect 38286 6196 38292 6208
rect 38344 6196 38350 6248
rect 31337 6140 31426 6168
rect 33413 6171 33471 6177
rect 31337 6137 31349 6140
rect 31291 6131 31349 6137
rect 33413 6137 33425 6171
rect 33459 6137 33471 6171
rect 33413 6131 33471 6137
rect 33965 6171 34023 6177
rect 33965 6137 33977 6171
rect 34011 6168 34023 6171
rect 34054 6168 34060 6180
rect 34011 6140 34060 6168
rect 34011 6137 34023 6140
rect 33965 6131 34023 6137
rect 14366 6100 14372 6112
rect 12452 6072 12664 6100
rect 14327 6072 14372 6100
rect 14366 6060 14372 6072
rect 14424 6060 14430 6112
rect 16482 6060 16488 6112
rect 16540 6100 16546 6112
rect 17037 6103 17095 6109
rect 17037 6100 17049 6103
rect 16540 6072 17049 6100
rect 16540 6060 16546 6072
rect 17037 6069 17049 6072
rect 17083 6069 17095 6103
rect 17862 6100 17868 6112
rect 17823 6072 17868 6100
rect 17037 6063 17095 6069
rect 17862 6060 17868 6072
rect 17920 6060 17926 6112
rect 18138 6100 18144 6112
rect 18099 6072 18144 6100
rect 18138 6060 18144 6072
rect 18196 6060 18202 6112
rect 22462 6100 22468 6112
rect 22423 6072 22468 6100
rect 22462 6060 22468 6072
rect 22520 6060 22526 6112
rect 28721 6103 28779 6109
rect 28721 6069 28733 6103
rect 28767 6100 28779 6103
rect 28902 6100 28908 6112
rect 28767 6072 28908 6100
rect 28767 6069 28779 6072
rect 28721 6063 28779 6069
rect 28902 6060 28908 6072
rect 28960 6060 28966 6112
rect 29089 6103 29147 6109
rect 29089 6069 29101 6103
rect 29135 6100 29147 6103
rect 29472 6100 29500 6128
rect 31846 6100 31852 6112
rect 29135 6072 29500 6100
rect 31807 6072 31852 6100
rect 29135 6069 29147 6072
rect 29089 6063 29147 6069
rect 31846 6060 31852 6072
rect 31904 6060 31910 6112
rect 33134 6060 33140 6112
rect 33192 6100 33198 6112
rect 33428 6100 33456 6131
rect 34054 6128 34060 6140
rect 34112 6128 34118 6180
rect 34885 6171 34943 6177
rect 34885 6137 34897 6171
rect 34931 6137 34943 6171
rect 34885 6131 34943 6137
rect 34330 6100 34336 6112
rect 33192 6072 33456 6100
rect 34291 6072 34336 6100
rect 33192 6060 33198 6072
rect 34330 6060 34336 6072
rect 34388 6100 34394 6112
rect 34900 6100 34928 6131
rect 34388 6072 34928 6100
rect 34388 6060 34394 6072
rect 35250 6060 35256 6112
rect 35308 6100 35314 6112
rect 36587 6103 36645 6109
rect 36587 6100 36599 6103
rect 35308 6072 36599 6100
rect 35308 6060 35314 6072
rect 36587 6069 36599 6072
rect 36633 6069 36645 6103
rect 36587 6063 36645 6069
rect 37599 6103 37657 6109
rect 37599 6069 37611 6103
rect 37645 6100 37657 6103
rect 37826 6100 37832 6112
rect 37645 6072 37832 6100
rect 37645 6069 37657 6072
rect 37599 6063 37657 6069
rect 37826 6060 37832 6072
rect 37884 6060 37890 6112
rect 1104 6010 48852 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 48852 6010
rect 1104 5936 48852 5958
rect 10226 5896 10232 5908
rect 10187 5868 10232 5896
rect 10226 5856 10232 5868
rect 10284 5856 10290 5908
rect 10778 5856 10784 5908
rect 10836 5896 10842 5908
rect 10873 5899 10931 5905
rect 10873 5896 10885 5899
rect 10836 5868 10885 5896
rect 10836 5856 10842 5868
rect 10873 5865 10885 5868
rect 10919 5865 10931 5899
rect 12526 5896 12532 5908
rect 12487 5868 12532 5896
rect 10873 5859 10931 5865
rect 12526 5856 12532 5868
rect 12584 5856 12590 5908
rect 13078 5896 13084 5908
rect 13039 5868 13084 5896
rect 13078 5856 13084 5868
rect 13136 5856 13142 5908
rect 17402 5896 17408 5908
rect 15856 5868 17408 5896
rect 12710 5720 12716 5772
rect 12768 5760 12774 5772
rect 12989 5763 13047 5769
rect 12989 5760 13001 5763
rect 12768 5732 13001 5760
rect 12768 5720 12774 5732
rect 12989 5729 13001 5732
rect 13035 5729 13047 5763
rect 12989 5723 13047 5729
rect 10505 5695 10563 5701
rect 10505 5661 10517 5695
rect 10551 5692 10563 5695
rect 10870 5692 10876 5704
rect 10551 5664 10876 5692
rect 10551 5661 10563 5664
rect 10505 5655 10563 5661
rect 10870 5652 10876 5664
rect 10928 5692 10934 5704
rect 11330 5692 11336 5704
rect 10928 5664 11336 5692
rect 10928 5652 10934 5664
rect 11330 5652 11336 5664
rect 11388 5652 11394 5704
rect 13004 5692 13032 5723
rect 13170 5720 13176 5772
rect 13228 5760 13234 5772
rect 13449 5763 13507 5769
rect 13449 5760 13461 5763
rect 13228 5732 13461 5760
rect 13228 5720 13234 5732
rect 13449 5729 13461 5732
rect 13495 5729 13507 5763
rect 13449 5723 13507 5729
rect 15746 5720 15752 5772
rect 15804 5760 15810 5772
rect 15856 5769 15884 5868
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 18138 5896 18144 5908
rect 18099 5868 18144 5896
rect 18138 5856 18144 5868
rect 18196 5856 18202 5908
rect 18506 5896 18512 5908
rect 18467 5868 18512 5896
rect 18506 5856 18512 5868
rect 18564 5856 18570 5908
rect 20990 5896 20996 5908
rect 20951 5868 20996 5896
rect 20990 5856 20996 5868
rect 21048 5856 21054 5908
rect 22186 5896 22192 5908
rect 22147 5868 22192 5896
rect 22186 5856 22192 5868
rect 22244 5856 22250 5908
rect 23934 5856 23940 5908
rect 23992 5896 23998 5908
rect 26694 5896 26700 5908
rect 23992 5868 26700 5896
rect 23992 5856 23998 5868
rect 26694 5856 26700 5868
rect 26752 5856 26758 5908
rect 28626 5856 28632 5908
rect 28684 5896 28690 5908
rect 28684 5868 30420 5896
rect 28684 5856 28690 5868
rect 17310 5828 17316 5840
rect 17271 5800 17316 5828
rect 17310 5788 17316 5800
rect 17368 5788 17374 5840
rect 18874 5828 18880 5840
rect 18835 5800 18880 5828
rect 18874 5788 18880 5800
rect 18932 5788 18938 5840
rect 20717 5831 20775 5837
rect 20717 5797 20729 5831
rect 20763 5828 20775 5831
rect 21174 5828 21180 5840
rect 20763 5800 21180 5828
rect 20763 5797 20775 5800
rect 20717 5791 20775 5797
rect 21174 5788 21180 5800
rect 21232 5788 21238 5840
rect 22830 5828 22836 5840
rect 22743 5800 22836 5828
rect 15841 5763 15899 5769
rect 15841 5760 15853 5763
rect 15804 5732 15853 5760
rect 15804 5720 15810 5732
rect 15841 5729 15853 5732
rect 15887 5729 15899 5763
rect 16114 5760 16120 5772
rect 16075 5732 16120 5760
rect 15841 5723 15899 5729
rect 16114 5720 16120 5732
rect 16172 5720 16178 5772
rect 20898 5760 20904 5772
rect 20859 5732 20904 5760
rect 20898 5720 20904 5732
rect 20956 5720 20962 5772
rect 21450 5760 21456 5772
rect 21411 5732 21456 5760
rect 21450 5720 21456 5732
rect 21508 5720 21514 5772
rect 22756 5769 22784 5800
rect 22830 5788 22836 5800
rect 22888 5828 22894 5840
rect 23474 5828 23480 5840
rect 22888 5800 23480 5828
rect 22888 5788 22894 5800
rect 23474 5788 23480 5800
rect 23532 5788 23538 5840
rect 24581 5831 24639 5837
rect 24581 5797 24593 5831
rect 24627 5828 24639 5831
rect 24762 5828 24768 5840
rect 24627 5800 24768 5828
rect 24627 5797 24639 5800
rect 24581 5791 24639 5797
rect 22741 5763 22799 5769
rect 22741 5729 22753 5763
rect 22787 5729 22799 5763
rect 22922 5760 22928 5772
rect 22883 5732 22928 5760
rect 22741 5723 22799 5729
rect 22922 5720 22928 5732
rect 22980 5760 22986 5772
rect 24596 5760 24624 5791
rect 24762 5788 24768 5800
rect 24820 5788 24826 5840
rect 24857 5831 24915 5837
rect 24857 5797 24869 5831
rect 24903 5828 24915 5831
rect 25038 5828 25044 5840
rect 24903 5800 25044 5828
rect 24903 5797 24915 5800
rect 24857 5791 24915 5797
rect 25038 5788 25044 5800
rect 25096 5788 25102 5840
rect 27154 5788 27160 5840
rect 27212 5828 27218 5840
rect 27386 5831 27444 5837
rect 27386 5828 27398 5831
rect 27212 5800 27398 5828
rect 27212 5788 27218 5800
rect 27386 5797 27398 5800
rect 27432 5828 27444 5831
rect 27522 5828 27528 5840
rect 27432 5800 27528 5828
rect 27432 5797 27444 5800
rect 27386 5791 27444 5797
rect 27522 5788 27528 5800
rect 27580 5788 27586 5840
rect 29822 5837 29828 5840
rect 29819 5828 29828 5837
rect 29783 5800 29828 5828
rect 29819 5791 29828 5800
rect 29822 5788 29828 5791
rect 29880 5788 29886 5840
rect 22980 5732 24624 5760
rect 22980 5720 22986 5732
rect 26970 5720 26976 5772
rect 27028 5760 27034 5772
rect 27065 5763 27123 5769
rect 27065 5760 27077 5763
rect 27028 5732 27077 5760
rect 27028 5720 27034 5732
rect 27065 5729 27077 5732
rect 27111 5729 27123 5763
rect 27065 5723 27123 5729
rect 29457 5763 29515 5769
rect 29457 5729 29469 5763
rect 29503 5760 29515 5763
rect 30282 5760 30288 5772
rect 29503 5732 30288 5760
rect 29503 5729 29515 5732
rect 29457 5723 29515 5729
rect 30282 5720 30288 5732
rect 30340 5720 30346 5772
rect 30392 5760 30420 5868
rect 30926 5856 30932 5908
rect 30984 5896 30990 5908
rect 31021 5899 31079 5905
rect 31021 5896 31033 5899
rect 30984 5868 31033 5896
rect 30984 5856 30990 5868
rect 31021 5865 31033 5868
rect 31067 5865 31079 5899
rect 31938 5896 31944 5908
rect 31899 5868 31944 5896
rect 31021 5859 31079 5865
rect 31938 5856 31944 5868
rect 31996 5856 32002 5908
rect 32030 5856 32036 5908
rect 32088 5896 32094 5908
rect 32217 5899 32275 5905
rect 32217 5896 32229 5899
rect 32088 5868 32229 5896
rect 32088 5856 32094 5868
rect 32217 5865 32229 5868
rect 32263 5865 32275 5899
rect 32217 5859 32275 5865
rect 33229 5899 33287 5905
rect 33229 5865 33241 5899
rect 33275 5896 33287 5899
rect 33410 5896 33416 5908
rect 33275 5868 33416 5896
rect 33275 5865 33287 5868
rect 33229 5859 33287 5865
rect 33410 5856 33416 5868
rect 33468 5856 33474 5908
rect 30745 5831 30803 5837
rect 30745 5797 30757 5831
rect 30791 5828 30803 5831
rect 30791 5800 32628 5828
rect 30791 5797 30803 5800
rect 30745 5791 30803 5797
rect 32122 5760 32128 5772
rect 30392 5732 32128 5760
rect 32122 5720 32128 5732
rect 32180 5720 32186 5772
rect 32600 5769 32628 5800
rect 33134 5788 33140 5840
rect 33192 5828 33198 5840
rect 33781 5831 33839 5837
rect 33781 5828 33793 5831
rect 33192 5800 33793 5828
rect 33192 5788 33198 5800
rect 33781 5797 33793 5800
rect 33827 5797 33839 5831
rect 33781 5791 33839 5797
rect 35805 5831 35863 5837
rect 35805 5797 35817 5831
rect 35851 5828 35863 5831
rect 36078 5828 36084 5840
rect 35851 5800 36084 5828
rect 35851 5797 35863 5800
rect 35805 5791 35863 5797
rect 36078 5788 36084 5800
rect 36136 5788 36142 5840
rect 36354 5828 36360 5840
rect 36315 5800 36360 5828
rect 36354 5788 36360 5800
rect 36412 5788 36418 5840
rect 32585 5763 32643 5769
rect 32585 5729 32597 5763
rect 32631 5760 32643 5763
rect 33410 5760 33416 5772
rect 32631 5732 33416 5760
rect 32631 5729 32643 5732
rect 32585 5723 32643 5729
rect 33410 5720 33416 5732
rect 33468 5720 33474 5772
rect 34146 5720 34152 5772
rect 34204 5760 34210 5772
rect 34425 5763 34483 5769
rect 34425 5760 34437 5763
rect 34204 5732 34437 5760
rect 34204 5720 34210 5732
rect 34425 5729 34437 5732
rect 34471 5760 34483 5763
rect 34606 5760 34612 5772
rect 34471 5732 34612 5760
rect 34471 5729 34483 5732
rect 34425 5723 34483 5729
rect 34606 5720 34612 5732
rect 34664 5720 34670 5772
rect 37645 5763 37703 5769
rect 37645 5729 37657 5763
rect 37691 5760 37703 5763
rect 37826 5760 37832 5772
rect 37691 5732 37832 5760
rect 37691 5729 37703 5732
rect 37645 5723 37703 5729
rect 37826 5720 37832 5732
rect 37884 5720 37890 5772
rect 15764 5692 15792 5720
rect 16206 5692 16212 5704
rect 13004 5664 15792 5692
rect 16167 5664 16212 5692
rect 16206 5652 16212 5664
rect 16264 5652 16270 5704
rect 16850 5652 16856 5704
rect 16908 5692 16914 5704
rect 17221 5695 17279 5701
rect 17221 5692 17233 5695
rect 16908 5664 17233 5692
rect 16908 5652 16914 5664
rect 17221 5661 17233 5664
rect 17267 5661 17279 5695
rect 17221 5655 17279 5661
rect 17497 5695 17555 5701
rect 17497 5661 17509 5695
rect 17543 5661 17555 5695
rect 18782 5692 18788 5704
rect 18743 5664 18788 5692
rect 17497 5655 17555 5661
rect 16942 5584 16948 5636
rect 17000 5624 17006 5636
rect 17512 5624 17540 5655
rect 18782 5652 18788 5664
rect 18840 5652 18846 5704
rect 19061 5695 19119 5701
rect 19061 5661 19073 5695
rect 19107 5661 19119 5695
rect 23106 5692 23112 5704
rect 23067 5664 23112 5692
rect 19061 5655 19119 5661
rect 19076 5624 19104 5655
rect 23106 5652 23112 5664
rect 23164 5652 23170 5704
rect 24118 5652 24124 5704
rect 24176 5692 24182 5704
rect 24765 5695 24823 5701
rect 24765 5692 24777 5695
rect 24176 5664 24777 5692
rect 24176 5652 24182 5664
rect 24765 5661 24777 5664
rect 24811 5661 24823 5695
rect 24765 5655 24823 5661
rect 25409 5695 25467 5701
rect 25409 5661 25421 5695
rect 25455 5692 25467 5695
rect 28718 5692 28724 5704
rect 25455 5664 28724 5692
rect 25455 5661 25467 5664
rect 25409 5655 25467 5661
rect 28718 5652 28724 5664
rect 28776 5692 28782 5704
rect 30098 5692 30104 5704
rect 28776 5664 30104 5692
rect 28776 5652 28782 5664
rect 30098 5652 30104 5664
rect 30156 5652 30162 5704
rect 30190 5652 30196 5704
rect 30248 5692 30254 5704
rect 35434 5692 35440 5704
rect 30248 5664 35440 5692
rect 30248 5652 30254 5664
rect 35434 5652 35440 5664
rect 35492 5652 35498 5704
rect 35713 5695 35771 5701
rect 35713 5661 35725 5695
rect 35759 5692 35771 5695
rect 36906 5692 36912 5704
rect 35759 5664 36912 5692
rect 35759 5661 35771 5664
rect 35713 5655 35771 5661
rect 36906 5652 36912 5664
rect 36964 5652 36970 5704
rect 17000 5596 19104 5624
rect 17000 5584 17006 5596
rect 30006 5584 30012 5636
rect 30064 5624 30070 5636
rect 36170 5624 36176 5636
rect 30064 5596 36176 5624
rect 30064 5584 30070 5596
rect 36170 5584 36176 5596
rect 36228 5584 36234 5636
rect 11422 5556 11428 5568
rect 11383 5528 11428 5556
rect 11422 5516 11428 5528
rect 11480 5516 11486 5568
rect 12802 5556 12808 5568
rect 12763 5528 12808 5556
rect 12802 5516 12808 5528
rect 12860 5516 12866 5568
rect 24762 5516 24768 5568
rect 24820 5556 24826 5568
rect 26053 5559 26111 5565
rect 26053 5556 26065 5559
rect 24820 5528 26065 5556
rect 24820 5516 24826 5528
rect 26053 5525 26065 5528
rect 26099 5556 26111 5559
rect 26510 5556 26516 5568
rect 26099 5528 26516 5556
rect 26099 5525 26111 5528
rect 26053 5519 26111 5525
rect 26510 5516 26516 5528
rect 26568 5516 26574 5568
rect 27154 5516 27160 5568
rect 27212 5556 27218 5568
rect 27985 5559 28043 5565
rect 27985 5556 27997 5559
rect 27212 5528 27997 5556
rect 27212 5516 27218 5528
rect 27985 5525 27997 5528
rect 28031 5525 28043 5559
rect 29362 5556 29368 5568
rect 29323 5528 29368 5556
rect 27985 5519 28043 5525
rect 29362 5516 29368 5528
rect 29420 5516 29426 5568
rect 29546 5516 29552 5568
rect 29604 5556 29610 5568
rect 30377 5559 30435 5565
rect 30377 5556 30389 5559
rect 29604 5528 30389 5556
rect 29604 5516 29610 5528
rect 30377 5525 30389 5528
rect 30423 5525 30435 5559
rect 30377 5519 30435 5525
rect 36538 5516 36544 5568
rect 36596 5556 36602 5568
rect 37875 5559 37933 5565
rect 37875 5556 37887 5559
rect 36596 5528 37887 5556
rect 36596 5516 36602 5528
rect 37875 5525 37887 5528
rect 37921 5525 37933 5559
rect 37875 5519 37933 5525
rect 1104 5466 48852 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 48852 5466
rect 1104 5392 48852 5414
rect 10137 5355 10195 5361
rect 10137 5321 10149 5355
rect 10183 5352 10195 5355
rect 10505 5355 10563 5361
rect 10505 5352 10517 5355
rect 10183 5324 10517 5352
rect 10183 5321 10195 5324
rect 10137 5315 10195 5321
rect 10505 5321 10517 5324
rect 10551 5352 10563 5355
rect 10778 5352 10784 5364
rect 10551 5324 10784 5352
rect 10551 5321 10563 5324
rect 10505 5315 10563 5321
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 11517 5355 11575 5361
rect 11517 5321 11529 5355
rect 11563 5352 11575 5355
rect 11790 5352 11796 5364
rect 11563 5324 11796 5352
rect 11563 5321 11575 5324
rect 11517 5315 11575 5321
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 12710 5352 12716 5364
rect 12671 5324 12716 5352
rect 12710 5312 12716 5324
rect 12768 5312 12774 5364
rect 15378 5352 15384 5364
rect 15339 5324 15384 5352
rect 15378 5312 15384 5324
rect 15436 5312 15442 5364
rect 16850 5352 16856 5364
rect 16811 5324 16856 5352
rect 16850 5312 16856 5324
rect 16908 5312 16914 5364
rect 17221 5355 17279 5361
rect 17221 5321 17233 5355
rect 17267 5352 17279 5355
rect 17310 5352 17316 5364
rect 17267 5324 17316 5352
rect 17267 5321 17279 5324
rect 17221 5315 17279 5321
rect 17310 5312 17316 5324
rect 17368 5312 17374 5364
rect 18874 5312 18880 5364
rect 18932 5352 18938 5364
rect 18969 5355 19027 5361
rect 18969 5352 18981 5355
rect 18932 5324 18981 5352
rect 18932 5312 18938 5324
rect 18969 5321 18981 5324
rect 19015 5352 19027 5355
rect 19245 5355 19303 5361
rect 19245 5352 19257 5355
rect 19015 5324 19257 5352
rect 19015 5321 19027 5324
rect 18969 5315 19027 5321
rect 19245 5321 19257 5324
rect 19291 5321 19303 5355
rect 19245 5315 19303 5321
rect 20165 5355 20223 5361
rect 20165 5321 20177 5355
rect 20211 5352 20223 5355
rect 20254 5352 20260 5364
rect 20211 5324 20260 5352
rect 20211 5321 20223 5324
rect 20165 5315 20223 5321
rect 20254 5312 20260 5324
rect 20312 5312 20318 5364
rect 20898 5312 20904 5364
rect 20956 5352 20962 5364
rect 21269 5355 21327 5361
rect 21269 5352 21281 5355
rect 20956 5324 21281 5352
rect 20956 5312 20962 5324
rect 21269 5321 21281 5324
rect 21315 5321 21327 5355
rect 22830 5352 22836 5364
rect 22791 5324 22836 5352
rect 21269 5315 21327 5321
rect 22830 5312 22836 5324
rect 22888 5312 22894 5364
rect 22922 5312 22928 5364
rect 22980 5352 22986 5364
rect 23201 5355 23259 5361
rect 23201 5352 23213 5355
rect 22980 5324 23213 5352
rect 22980 5312 22986 5324
rect 23201 5321 23213 5324
rect 23247 5321 23259 5355
rect 23201 5315 23259 5321
rect 23382 5312 23388 5364
rect 23440 5352 23446 5364
rect 24118 5352 24124 5364
rect 23440 5312 23474 5352
rect 24079 5324 24124 5352
rect 24118 5312 24124 5324
rect 24176 5312 24182 5364
rect 26970 5312 26976 5364
rect 27028 5352 27034 5364
rect 27893 5355 27951 5361
rect 27893 5352 27905 5355
rect 27028 5324 27905 5352
rect 27028 5312 27034 5324
rect 27893 5321 27905 5324
rect 27939 5321 27951 5355
rect 27893 5315 27951 5321
rect 29822 5312 29828 5364
rect 29880 5352 29886 5364
rect 30285 5355 30343 5361
rect 30285 5352 30297 5355
rect 29880 5324 30297 5352
rect 29880 5312 29886 5324
rect 30285 5321 30297 5324
rect 30331 5352 30343 5355
rect 30834 5352 30840 5364
rect 30331 5324 30840 5352
rect 30331 5321 30343 5324
rect 30285 5315 30343 5321
rect 30834 5312 30840 5324
rect 30892 5312 30898 5364
rect 32122 5352 32128 5364
rect 32083 5324 32128 5352
rect 32122 5312 32128 5324
rect 32180 5312 32186 5364
rect 34146 5352 34152 5364
rect 34107 5324 34152 5352
rect 34146 5312 34152 5324
rect 34204 5312 34210 5364
rect 36906 5352 36912 5364
rect 36867 5324 36912 5352
rect 36906 5312 36912 5324
rect 36964 5312 36970 5364
rect 37826 5312 37832 5364
rect 37884 5352 37890 5364
rect 37921 5355 37979 5361
rect 37921 5352 37933 5355
rect 37884 5324 37933 5352
rect 37884 5312 37890 5324
rect 37921 5321 37933 5324
rect 37967 5352 37979 5355
rect 38289 5355 38347 5361
rect 38289 5352 38301 5355
rect 37967 5324 38301 5352
rect 37967 5321 37979 5324
rect 37921 5315 37979 5321
rect 38289 5321 38301 5324
rect 38335 5321 38347 5355
rect 38289 5315 38347 5321
rect 10796 5284 10824 5312
rect 12989 5287 13047 5293
rect 12989 5284 13001 5287
rect 10796 5256 13001 5284
rect 12989 5253 13001 5256
rect 13035 5253 13047 5287
rect 12989 5247 13047 5253
rect 10594 5148 10600 5160
rect 10507 5120 10600 5148
rect 10594 5108 10600 5120
rect 10652 5148 10658 5160
rect 11793 5151 11851 5157
rect 11793 5148 11805 5151
rect 10652 5120 11805 5148
rect 10652 5108 10658 5120
rect 11793 5117 11805 5120
rect 11839 5117 11851 5151
rect 11793 5111 11851 5117
rect 10778 5040 10784 5092
rect 10836 5080 10842 5092
rect 10918 5083 10976 5089
rect 10918 5080 10930 5083
rect 10836 5052 10930 5080
rect 10836 5040 10842 5052
rect 10918 5049 10930 5052
rect 10964 5049 10976 5083
rect 13004 5080 13032 5247
rect 13078 5176 13084 5228
rect 13136 5216 13142 5228
rect 13173 5219 13231 5225
rect 13173 5216 13185 5219
rect 13136 5188 13185 5216
rect 13136 5176 13142 5188
rect 13173 5185 13185 5188
rect 13219 5216 13231 5219
rect 14369 5219 14427 5225
rect 14369 5216 14381 5219
rect 13219 5188 14381 5216
rect 13219 5185 13231 5188
rect 13173 5179 13231 5185
rect 14369 5185 14381 5188
rect 14415 5185 14427 5219
rect 14369 5179 14427 5185
rect 16482 5176 16488 5228
rect 16540 5216 16546 5228
rect 17773 5219 17831 5225
rect 17773 5216 17785 5219
rect 16540 5188 17785 5216
rect 16540 5176 16546 5188
rect 17773 5185 17785 5188
rect 17819 5185 17831 5219
rect 17773 5179 17831 5185
rect 18049 5219 18107 5225
rect 18049 5185 18061 5219
rect 18095 5216 18107 5219
rect 18138 5216 18144 5228
rect 18095 5188 18144 5216
rect 18095 5185 18107 5188
rect 18049 5179 18107 5185
rect 15378 5108 15384 5160
rect 15436 5148 15442 5160
rect 15565 5151 15623 5157
rect 15565 5148 15577 5151
rect 15436 5120 15577 5148
rect 15436 5108 15442 5120
rect 15565 5117 15577 5120
rect 15611 5117 15623 5151
rect 16114 5148 16120 5160
rect 16075 5120 16120 5148
rect 15565 5111 15623 5117
rect 16114 5108 16120 5120
rect 16172 5108 16178 5160
rect 13494 5083 13552 5089
rect 13494 5080 13506 5083
rect 13004 5052 13506 5080
rect 10918 5043 10976 5049
rect 13494 5049 13506 5052
rect 13540 5080 13552 5083
rect 15010 5080 15016 5092
rect 13540 5052 15016 5080
rect 13540 5049 13552 5052
rect 13494 5043 13552 5049
rect 15010 5040 15016 5052
rect 15068 5040 15074 5092
rect 15105 5083 15163 5089
rect 15105 5049 15117 5083
rect 15151 5080 15163 5083
rect 16132 5080 16160 5108
rect 15151 5052 16160 5080
rect 17788 5080 17816 5179
rect 18138 5176 18144 5188
rect 18196 5176 18202 5228
rect 22554 5216 22560 5228
rect 22388 5188 22560 5216
rect 20254 5148 20260 5160
rect 20215 5120 20260 5148
rect 20254 5108 20260 5120
rect 20312 5108 20318 5160
rect 20346 5108 20352 5160
rect 20404 5148 20410 5160
rect 20809 5151 20867 5157
rect 20809 5148 20821 5151
rect 20404 5120 20821 5148
rect 20404 5108 20410 5120
rect 20809 5117 20821 5120
rect 20855 5148 20867 5151
rect 21450 5148 21456 5160
rect 20855 5120 21456 5148
rect 20855 5117 20867 5120
rect 20809 5111 20867 5117
rect 21450 5108 21456 5120
rect 21508 5108 21514 5160
rect 21634 5108 21640 5160
rect 21692 5148 21698 5160
rect 22388 5157 22416 5188
rect 22554 5176 22560 5188
rect 22612 5216 22618 5228
rect 22940 5216 22968 5312
rect 23446 5284 23474 5312
rect 25777 5287 25835 5293
rect 25777 5284 25789 5287
rect 23446 5256 25789 5284
rect 25777 5253 25789 5256
rect 25823 5253 25835 5287
rect 25777 5247 25835 5253
rect 26237 5287 26295 5293
rect 26237 5253 26249 5287
rect 26283 5284 26295 5287
rect 26694 5284 26700 5296
rect 26283 5256 26700 5284
rect 26283 5253 26295 5256
rect 26237 5247 26295 5253
rect 25792 5216 25820 5247
rect 26694 5244 26700 5256
rect 26752 5284 26758 5296
rect 27522 5284 27528 5296
rect 26752 5256 27528 5284
rect 26752 5244 26758 5256
rect 27522 5244 27528 5256
rect 27580 5284 27586 5296
rect 31849 5287 31907 5293
rect 27580 5256 28994 5284
rect 27580 5244 27586 5256
rect 26329 5219 26387 5225
rect 26329 5216 26341 5219
rect 22612 5188 22968 5216
rect 23446 5188 25728 5216
rect 25792 5188 26341 5216
rect 22612 5176 22618 5188
rect 21729 5151 21787 5157
rect 21729 5148 21741 5151
rect 21692 5120 21741 5148
rect 21692 5108 21698 5120
rect 21729 5117 21741 5120
rect 21775 5148 21787 5151
rect 21821 5151 21879 5157
rect 21821 5148 21833 5151
rect 21775 5120 21833 5148
rect 21775 5117 21787 5120
rect 21729 5111 21787 5117
rect 21821 5117 21833 5120
rect 21867 5117 21879 5151
rect 21821 5111 21879 5117
rect 22373 5151 22431 5157
rect 22373 5117 22385 5151
rect 22419 5117 22431 5151
rect 22373 5111 22431 5117
rect 22830 5108 22836 5160
rect 22888 5148 22894 5160
rect 23446 5148 23474 5188
rect 24578 5148 24584 5160
rect 22888 5120 23474 5148
rect 24539 5120 24584 5148
rect 22888 5108 22894 5120
rect 24578 5108 24584 5120
rect 24636 5108 24642 5160
rect 25700 5148 25728 5188
rect 26329 5185 26341 5188
rect 26375 5185 26387 5219
rect 28966 5216 28994 5256
rect 31849 5253 31861 5287
rect 31895 5284 31907 5287
rect 34609 5287 34667 5293
rect 34609 5284 34621 5287
rect 31895 5256 34621 5284
rect 31895 5253 31907 5256
rect 31849 5247 31907 5253
rect 34609 5253 34621 5256
rect 34655 5253 34667 5287
rect 34609 5247 34667 5253
rect 29086 5216 29092 5228
rect 28966 5188 29092 5216
rect 26329 5179 26387 5185
rect 29086 5176 29092 5188
rect 29144 5176 29150 5228
rect 29822 5216 29828 5228
rect 29783 5188 29828 5216
rect 29822 5176 29828 5188
rect 29880 5176 29886 5228
rect 30926 5216 30932 5228
rect 30887 5188 30932 5216
rect 30926 5176 30932 5188
rect 30984 5176 30990 5228
rect 28112 5151 28170 5157
rect 28112 5148 28124 5151
rect 25700 5120 28124 5148
rect 28112 5117 28124 5120
rect 28158 5148 28170 5151
rect 28537 5151 28595 5157
rect 28537 5148 28549 5151
rect 28158 5120 28549 5148
rect 28158 5117 28170 5120
rect 28112 5111 28170 5117
rect 28537 5117 28549 5120
rect 28583 5117 28595 5151
rect 28537 5111 28595 5117
rect 30374 5108 30380 5160
rect 30432 5148 30438 5160
rect 32585 5151 32643 5157
rect 32585 5148 32597 5151
rect 30432 5120 32597 5148
rect 30432 5108 30438 5120
rect 32585 5117 32597 5120
rect 32631 5148 32643 5151
rect 32677 5151 32735 5157
rect 32677 5148 32689 5151
rect 32631 5120 32689 5148
rect 32631 5117 32643 5120
rect 32585 5111 32643 5117
rect 32677 5117 32689 5120
rect 32723 5117 32735 5151
rect 32677 5111 32735 5117
rect 33229 5151 33287 5157
rect 33229 5117 33241 5151
rect 33275 5148 33287 5151
rect 33410 5148 33416 5160
rect 33275 5120 33416 5148
rect 33275 5117 33287 5120
rect 33229 5111 33287 5117
rect 33410 5108 33416 5120
rect 33468 5148 33474 5160
rect 33689 5151 33747 5157
rect 33689 5148 33701 5151
rect 33468 5120 33701 5148
rect 33468 5108 33474 5120
rect 33689 5117 33701 5120
rect 33735 5117 33747 5151
rect 34624 5148 34652 5247
rect 34920 5151 34978 5157
rect 34920 5148 34932 5151
rect 34624 5120 34932 5148
rect 33689 5111 33747 5117
rect 34920 5117 34932 5120
rect 34966 5117 34978 5151
rect 36538 5148 36544 5160
rect 36499 5120 36544 5148
rect 34920 5111 34978 5117
rect 36538 5108 36544 5120
rect 36596 5108 36602 5160
rect 37461 5151 37519 5157
rect 37461 5117 37473 5151
rect 37507 5148 37519 5151
rect 37826 5148 37832 5160
rect 37507 5120 37832 5148
rect 37507 5117 37519 5120
rect 37461 5111 37519 5117
rect 37826 5108 37832 5120
rect 37884 5108 37890 5160
rect 18370 5083 18428 5089
rect 18370 5080 18382 5083
rect 17788 5052 18382 5080
rect 15151 5049 15163 5052
rect 15105 5043 15163 5049
rect 18370 5049 18382 5052
rect 18416 5080 18428 5083
rect 20714 5080 20720 5092
rect 18416 5052 20720 5080
rect 18416 5049 18428 5052
rect 18370 5043 18428 5049
rect 20714 5040 20720 5052
rect 20772 5040 20778 5092
rect 20993 5083 21051 5089
rect 20993 5049 21005 5083
rect 21039 5080 21051 5083
rect 21174 5080 21180 5092
rect 21039 5052 21180 5080
rect 21039 5049 21051 5052
rect 20993 5043 21051 5049
rect 21174 5040 21180 5052
rect 21232 5040 21238 5092
rect 22557 5083 22615 5089
rect 22557 5049 22569 5083
rect 22603 5080 22615 5083
rect 23658 5080 23664 5092
rect 22603 5052 23664 5080
rect 22603 5049 22615 5052
rect 22557 5043 22615 5049
rect 23658 5040 23664 5052
rect 23716 5040 23722 5092
rect 24486 5080 24492 5092
rect 24399 5052 24492 5080
rect 24486 5040 24492 5052
rect 24544 5080 24550 5092
rect 26694 5089 26700 5092
rect 24943 5083 25001 5089
rect 24943 5080 24955 5083
rect 24544 5052 24955 5080
rect 24544 5040 24550 5052
rect 24943 5049 24955 5052
rect 24989 5080 25001 5083
rect 26691 5080 26700 5089
rect 24989 5052 26700 5080
rect 24989 5049 25001 5052
rect 24943 5043 25001 5049
rect 26691 5043 26700 5052
rect 26694 5040 26700 5043
rect 26752 5040 26758 5092
rect 28810 5040 28816 5092
rect 28868 5080 28874 5092
rect 29362 5080 29368 5092
rect 28868 5052 29368 5080
rect 28868 5040 28874 5052
rect 29362 5040 29368 5052
rect 29420 5040 29426 5092
rect 29457 5083 29515 5089
rect 29457 5049 29469 5083
rect 29503 5080 29515 5083
rect 31018 5080 31024 5092
rect 29503 5052 31024 5080
rect 29503 5049 29515 5052
rect 29457 5043 29515 5049
rect 9582 5012 9588 5024
rect 9543 4984 9588 5012
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 14090 5012 14096 5024
rect 14051 4984 14096 5012
rect 14090 4972 14096 4984
rect 14148 4972 14154 5024
rect 15654 5012 15660 5024
rect 15615 4984 15660 5012
rect 15654 4972 15660 4984
rect 15712 4972 15718 5024
rect 25498 5012 25504 5024
rect 25459 4984 25504 5012
rect 25498 4972 25504 4984
rect 25556 4972 25562 5024
rect 26510 4972 26516 5024
rect 26568 5012 26574 5024
rect 27249 5015 27307 5021
rect 27249 5012 27261 5015
rect 26568 4984 27261 5012
rect 26568 4972 26574 4984
rect 27249 4981 27261 4984
rect 27295 4981 27307 5015
rect 27249 4975 27307 4981
rect 28215 5015 28273 5021
rect 28215 4981 28227 5015
rect 28261 5012 28273 5015
rect 28442 5012 28448 5024
rect 28261 4984 28448 5012
rect 28261 4981 28273 4984
rect 28215 4975 28273 4981
rect 28442 4972 28448 4984
rect 28500 4972 28506 5024
rect 28902 4972 28908 5024
rect 28960 5012 28966 5024
rect 29089 5015 29147 5021
rect 29089 5012 29101 5015
rect 28960 4984 29101 5012
rect 28960 4972 28966 4984
rect 29089 4981 29101 4984
rect 29135 5012 29147 5015
rect 29472 5012 29500 5043
rect 31018 5040 31024 5052
rect 31076 5040 31082 5092
rect 31250 5083 31308 5089
rect 31250 5049 31262 5083
rect 31296 5049 31308 5083
rect 36630 5080 36636 5092
rect 36591 5052 36636 5080
rect 31250 5043 31308 5049
rect 29135 4984 29500 5012
rect 29135 4981 29147 4984
rect 29089 4975 29147 4981
rect 30834 4972 30840 5024
rect 30892 5012 30898 5024
rect 31265 5012 31293 5043
rect 36630 5040 36636 5052
rect 36688 5040 36694 5092
rect 32766 5012 32772 5024
rect 30892 4984 31293 5012
rect 32727 4984 32772 5012
rect 30892 4972 30898 4984
rect 32766 4972 32772 4984
rect 32824 4972 32830 5024
rect 34238 4972 34244 5024
rect 34296 5012 34302 5024
rect 35023 5015 35081 5021
rect 35023 5012 35035 5015
rect 34296 4984 35035 5012
rect 34296 4972 34302 4984
rect 35023 4981 35035 4984
rect 35069 4981 35081 5015
rect 35023 4975 35081 4981
rect 35713 5015 35771 5021
rect 35713 4981 35725 5015
rect 35759 5012 35771 5015
rect 36078 5012 36084 5024
rect 35759 4984 36084 5012
rect 35759 4981 35771 4984
rect 35713 4975 35771 4981
rect 36078 4972 36084 4984
rect 36136 4972 36142 5024
rect 37642 5012 37648 5024
rect 37603 4984 37648 5012
rect 37642 4972 37648 4984
rect 37700 4972 37706 5024
rect 1104 4922 48852 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 48852 4922
rect 1104 4848 48852 4870
rect 10594 4808 10600 4820
rect 10555 4780 10600 4808
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 11330 4808 11336 4820
rect 11291 4780 11336 4808
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 12023 4811 12081 4817
rect 12023 4777 12035 4811
rect 12069 4808 12081 4811
rect 12802 4808 12808 4820
rect 12069 4780 12808 4808
rect 12069 4777 12081 4780
rect 12023 4771 12081 4777
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 15657 4811 15715 4817
rect 15657 4777 15669 4811
rect 15703 4808 15715 4811
rect 15746 4808 15752 4820
rect 15703 4780 15752 4808
rect 15703 4777 15715 4780
rect 15657 4771 15715 4777
rect 15746 4768 15752 4780
rect 15804 4768 15810 4820
rect 16025 4811 16083 4817
rect 16025 4777 16037 4811
rect 16071 4808 16083 4811
rect 16114 4808 16120 4820
rect 16071 4780 16120 4808
rect 16071 4777 16083 4780
rect 16025 4771 16083 4777
rect 16114 4768 16120 4780
rect 16172 4808 16178 4820
rect 17037 4811 17095 4817
rect 16172 4780 16620 4808
rect 16172 4768 16178 4780
rect 12434 4740 12440 4752
rect 12395 4712 12440 4740
rect 12434 4700 12440 4712
rect 12492 4700 12498 4752
rect 13449 4743 13507 4749
rect 13449 4709 13461 4743
rect 13495 4740 13507 4743
rect 14090 4740 14096 4752
rect 13495 4712 14096 4740
rect 13495 4709 13507 4712
rect 13449 4703 13507 4709
rect 14090 4700 14096 4712
rect 14148 4740 14154 4752
rect 14645 4743 14703 4749
rect 14645 4740 14657 4743
rect 14148 4712 14657 4740
rect 14148 4700 14154 4712
rect 14645 4709 14657 4712
rect 14691 4709 14703 4743
rect 14645 4703 14703 4709
rect 15010 4700 15016 4752
rect 15068 4740 15074 4752
rect 16482 4749 16488 4752
rect 16438 4743 16488 4749
rect 16438 4740 16450 4743
rect 15068 4712 16450 4740
rect 15068 4700 15074 4712
rect 16438 4709 16450 4712
rect 16484 4709 16488 4743
rect 16438 4703 16488 4709
rect 16482 4700 16488 4703
rect 16540 4700 16546 4752
rect 16592 4740 16620 4780
rect 17037 4777 17049 4811
rect 17083 4808 17095 4811
rect 17310 4808 17316 4820
rect 17083 4780 17316 4808
rect 17083 4777 17095 4780
rect 17037 4771 17095 4777
rect 17310 4768 17316 4780
rect 17368 4768 17374 4820
rect 18782 4768 18788 4820
rect 18840 4808 18846 4820
rect 18877 4811 18935 4817
rect 18877 4808 18889 4811
rect 18840 4780 18889 4808
rect 18840 4768 18846 4780
rect 18877 4777 18889 4780
rect 18923 4777 18935 4811
rect 20346 4808 20352 4820
rect 20307 4780 20352 4808
rect 18877 4771 18935 4777
rect 20346 4768 20352 4780
rect 20404 4808 20410 4820
rect 21085 4811 21143 4817
rect 21085 4808 21097 4811
rect 20404 4780 21097 4808
rect 20404 4768 20410 4780
rect 21085 4777 21097 4780
rect 21131 4777 21143 4811
rect 22554 4808 22560 4820
rect 22515 4780 22560 4808
rect 21085 4771 21143 4777
rect 22554 4768 22560 4780
rect 22612 4768 22618 4820
rect 24397 4811 24455 4817
rect 24397 4777 24409 4811
rect 24443 4808 24455 4811
rect 24578 4808 24584 4820
rect 24443 4780 24584 4808
rect 24443 4777 24455 4780
rect 24397 4771 24455 4777
rect 24578 4768 24584 4780
rect 24636 4768 24642 4820
rect 26786 4768 26792 4820
rect 26844 4808 26850 4820
rect 27525 4811 27583 4817
rect 27525 4808 27537 4811
rect 26844 4780 27537 4808
rect 26844 4768 26850 4780
rect 27525 4777 27537 4780
rect 27571 4777 27583 4811
rect 30282 4808 30288 4820
rect 30243 4780 30288 4808
rect 27525 4771 27583 4777
rect 30282 4768 30288 4780
rect 30340 4768 30346 4820
rect 35989 4811 36047 4817
rect 35989 4777 36001 4811
rect 36035 4808 36047 4811
rect 36538 4808 36544 4820
rect 36035 4780 36544 4808
rect 36035 4777 36047 4780
rect 35989 4771 36047 4777
rect 36538 4768 36544 4780
rect 36596 4768 36602 4820
rect 17586 4740 17592 4752
rect 16592 4712 17592 4740
rect 17586 4700 17592 4712
rect 17644 4740 17650 4752
rect 22462 4740 22468 4752
rect 17644 4712 22468 4740
rect 17644 4700 17650 4712
rect 10502 4672 10508 4684
rect 10463 4644 10508 4672
rect 10502 4632 10508 4644
rect 10560 4632 10566 4684
rect 10686 4632 10692 4684
rect 10744 4672 10750 4684
rect 10781 4675 10839 4681
rect 10781 4672 10793 4675
rect 10744 4644 10793 4672
rect 10744 4632 10750 4644
rect 10781 4641 10793 4644
rect 10827 4641 10839 4675
rect 10781 4635 10839 4641
rect 11952 4675 12010 4681
rect 11952 4641 11964 4675
rect 11998 4672 12010 4675
rect 12452 4672 12480 4700
rect 11998 4644 12480 4672
rect 11998 4641 12010 4644
rect 11952 4635 12010 4641
rect 10796 4604 10824 4635
rect 16022 4632 16028 4684
rect 16080 4672 16086 4684
rect 16117 4675 16175 4681
rect 16117 4672 16129 4675
rect 16080 4644 16129 4672
rect 16080 4632 16086 4644
rect 16117 4641 16129 4644
rect 16163 4672 16175 4675
rect 17494 4672 17500 4684
rect 16163 4644 17500 4672
rect 16163 4641 16175 4644
rect 16117 4635 16175 4641
rect 17494 4632 17500 4644
rect 17552 4632 17558 4684
rect 17862 4672 17868 4684
rect 17823 4644 17868 4672
rect 17862 4632 17868 4644
rect 17920 4632 17926 4684
rect 18432 4681 18460 4712
rect 22462 4700 22468 4712
rect 22520 4700 22526 4752
rect 18417 4675 18475 4681
rect 18417 4641 18429 4675
rect 18463 4641 18475 4675
rect 18417 4635 18475 4641
rect 19429 4675 19487 4681
rect 19429 4641 19441 4675
rect 19475 4641 19487 4675
rect 19429 4635 19487 4641
rect 12989 4607 13047 4613
rect 12989 4604 13001 4607
rect 10796 4576 13001 4604
rect 12989 4573 13001 4576
rect 13035 4604 13047 4607
rect 13170 4604 13176 4616
rect 13035 4576 13176 4604
rect 13035 4573 13047 4576
rect 12989 4567 13047 4573
rect 13170 4564 13176 4576
rect 13228 4564 13234 4616
rect 13354 4604 13360 4616
rect 13315 4576 13360 4604
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 13630 4604 13636 4616
rect 13591 4576 13636 4604
rect 13630 4564 13636 4576
rect 13688 4564 13694 4616
rect 18506 4604 18512 4616
rect 18467 4576 18512 4604
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 19444 4604 19472 4635
rect 19518 4632 19524 4684
rect 19576 4672 19582 4684
rect 19613 4675 19671 4681
rect 19613 4672 19625 4675
rect 19576 4644 19625 4672
rect 19576 4632 19582 4644
rect 19613 4641 19625 4644
rect 19659 4672 19671 4675
rect 19978 4672 19984 4684
rect 19659 4644 19984 4672
rect 19659 4641 19671 4644
rect 19613 4635 19671 4641
rect 19978 4632 19984 4644
rect 20036 4632 20042 4684
rect 21266 4632 21272 4684
rect 21324 4672 21330 4684
rect 21453 4675 21511 4681
rect 21453 4672 21465 4675
rect 21324 4644 21465 4672
rect 21324 4632 21330 4644
rect 21453 4641 21465 4644
rect 21499 4641 21511 4675
rect 21453 4635 21511 4641
rect 22005 4675 22063 4681
rect 22005 4641 22017 4675
rect 22051 4672 22063 4675
rect 22572 4672 22600 4768
rect 23471 4743 23529 4749
rect 23471 4709 23483 4743
rect 23517 4740 23529 4743
rect 24486 4740 24492 4752
rect 23517 4712 24492 4740
rect 23517 4709 23529 4712
rect 23471 4703 23529 4709
rect 24486 4700 24492 4712
rect 24544 4700 24550 4752
rect 24765 4743 24823 4749
rect 24765 4709 24777 4743
rect 24811 4740 24823 4743
rect 25038 4740 25044 4752
rect 24811 4712 25044 4740
rect 24811 4709 24823 4712
rect 24765 4703 24823 4709
rect 25038 4700 25044 4712
rect 25096 4700 25102 4752
rect 26697 4743 26755 4749
rect 26697 4709 26709 4743
rect 26743 4740 26755 4743
rect 27062 4740 27068 4752
rect 26743 4712 27068 4740
rect 26743 4709 26755 4712
rect 26697 4703 26755 4709
rect 27062 4700 27068 4712
rect 27120 4700 27126 4752
rect 29086 4700 29092 4752
rect 29144 4740 29150 4752
rect 29451 4743 29509 4749
rect 29451 4740 29463 4743
rect 29144 4712 29463 4740
rect 29144 4700 29150 4712
rect 29451 4709 29463 4712
rect 29497 4740 29509 4743
rect 30834 4740 30840 4752
rect 29497 4712 30840 4740
rect 29497 4709 29509 4712
rect 29451 4703 29509 4709
rect 30834 4700 30840 4712
rect 30892 4700 30898 4752
rect 32214 4700 32220 4752
rect 32272 4740 32278 4752
rect 32585 4743 32643 4749
rect 32585 4740 32597 4743
rect 32272 4712 32597 4740
rect 32272 4700 32278 4712
rect 32585 4709 32597 4712
rect 32631 4740 32643 4743
rect 33134 4740 33140 4752
rect 32631 4712 33140 4740
rect 32631 4709 32643 4712
rect 32585 4703 32643 4709
rect 33134 4700 33140 4712
rect 33192 4700 33198 4752
rect 34146 4740 34152 4752
rect 34107 4712 34152 4740
rect 34146 4700 34152 4712
rect 34204 4700 34210 4752
rect 36078 4740 36084 4752
rect 36039 4712 36084 4740
rect 36078 4700 36084 4712
rect 36136 4700 36142 4752
rect 23106 4672 23112 4684
rect 22051 4644 22600 4672
rect 23067 4644 23112 4672
rect 22051 4641 22063 4644
rect 22005 4635 22063 4641
rect 23106 4632 23112 4644
rect 23164 4632 23170 4684
rect 28166 4681 28172 4684
rect 28144 4675 28172 4681
rect 28144 4672 28156 4675
rect 28079 4644 28156 4672
rect 28144 4641 28156 4644
rect 28224 4672 28230 4684
rect 29546 4672 29552 4684
rect 28224 4644 29552 4672
rect 28144 4635 28172 4641
rect 28166 4632 28172 4635
rect 28224 4632 28230 4644
rect 29546 4632 29552 4644
rect 29604 4632 29610 4684
rect 30374 4632 30380 4684
rect 30432 4672 30438 4684
rect 31088 4675 31146 4681
rect 31088 4672 31100 4675
rect 30432 4644 31100 4672
rect 30432 4632 30438 4644
rect 31088 4641 31100 4644
rect 31134 4672 31146 4675
rect 31846 4672 31852 4684
rect 31134 4644 31852 4672
rect 31134 4641 31146 4644
rect 31088 4635 31146 4641
rect 31846 4632 31852 4644
rect 31904 4632 31910 4684
rect 35986 4632 35992 4684
rect 36044 4672 36050 4684
rect 36725 4675 36783 4681
rect 36725 4672 36737 4675
rect 36044 4644 36737 4672
rect 36044 4632 36050 4644
rect 36725 4641 36737 4644
rect 36771 4672 36783 4675
rect 37642 4672 37648 4684
rect 36771 4644 37648 4672
rect 36771 4641 36783 4644
rect 36725 4635 36783 4641
rect 37642 4632 37648 4644
rect 37700 4632 37706 4684
rect 20622 4604 20628 4616
rect 19444 4576 20628 4604
rect 20622 4564 20628 4576
rect 20680 4564 20686 4616
rect 22186 4604 22192 4616
rect 22147 4576 22192 4604
rect 22186 4564 22192 4576
rect 22244 4564 22250 4616
rect 24949 4607 25007 4613
rect 24949 4573 24961 4607
rect 24995 4604 25007 4607
rect 25222 4604 25228 4616
rect 24995 4576 25228 4604
rect 24995 4573 25007 4576
rect 24949 4567 25007 4573
rect 25222 4564 25228 4576
rect 25280 4564 25286 4616
rect 26602 4604 26608 4616
rect 26563 4576 26608 4604
rect 26602 4564 26608 4576
rect 26660 4564 26666 4616
rect 27249 4607 27307 4613
rect 27249 4573 27261 4607
rect 27295 4604 27307 4607
rect 27338 4604 27344 4616
rect 27295 4576 27344 4604
rect 27295 4573 27307 4576
rect 27249 4567 27307 4573
rect 27338 4564 27344 4576
rect 27396 4564 27402 4616
rect 28997 4607 29055 4613
rect 28997 4573 29009 4607
rect 29043 4604 29055 4607
rect 29089 4607 29147 4613
rect 29089 4604 29101 4607
rect 29043 4576 29101 4604
rect 29043 4573 29055 4576
rect 28997 4567 29055 4573
rect 29089 4573 29101 4576
rect 29135 4604 29147 4607
rect 32030 4604 32036 4616
rect 29135 4576 32036 4604
rect 29135 4573 29147 4576
rect 29089 4567 29147 4573
rect 32030 4564 32036 4576
rect 32088 4564 32094 4616
rect 32493 4607 32551 4613
rect 32493 4573 32505 4607
rect 32539 4604 32551 4607
rect 33502 4604 33508 4616
rect 32539 4576 33508 4604
rect 32539 4573 32551 4576
rect 32493 4567 32551 4573
rect 33502 4564 33508 4576
rect 33560 4564 33566 4616
rect 34054 4604 34060 4616
rect 33967 4576 34060 4604
rect 34054 4564 34060 4576
rect 34112 4604 34118 4616
rect 34698 4604 34704 4616
rect 34112 4576 34704 4604
rect 34112 4564 34118 4576
rect 34698 4564 34704 4576
rect 34756 4564 34762 4616
rect 13188 4536 13216 4564
rect 25501 4539 25559 4545
rect 13188 4508 18092 4536
rect 13722 4428 13728 4480
rect 13780 4468 13786 4480
rect 14277 4471 14335 4477
rect 14277 4468 14289 4471
rect 13780 4440 14289 4468
rect 13780 4428 13786 4440
rect 14277 4437 14289 4440
rect 14323 4437 14335 4471
rect 15102 4468 15108 4480
rect 15063 4440 15108 4468
rect 14277 4431 14335 4437
rect 15102 4428 15108 4440
rect 15160 4428 15166 4480
rect 17770 4468 17776 4480
rect 17731 4440 17776 4468
rect 17770 4428 17776 4440
rect 17828 4428 17834 4480
rect 18064 4468 18092 4508
rect 25501 4505 25513 4539
rect 25547 4536 25559 4539
rect 25590 4536 25596 4548
rect 25547 4508 25596 4536
rect 25547 4505 25559 4508
rect 25501 4499 25559 4505
rect 25590 4496 25596 4508
rect 25648 4536 25654 4548
rect 29638 4536 29644 4548
rect 25648 4508 29644 4536
rect 25648 4496 25654 4508
rect 29638 4496 29644 4508
rect 29696 4496 29702 4548
rect 33042 4536 33048 4548
rect 33003 4508 33048 4536
rect 33042 4496 33048 4508
rect 33100 4496 33106 4548
rect 34606 4536 34612 4548
rect 34567 4508 34612 4536
rect 34606 4496 34612 4508
rect 34664 4496 34670 4548
rect 19705 4471 19763 4477
rect 19705 4468 19717 4471
rect 18064 4440 19717 4468
rect 19705 4437 19717 4440
rect 19751 4437 19763 4471
rect 22922 4468 22928 4480
rect 22835 4440 22928 4468
rect 19705 4431 19763 4437
rect 22922 4428 22928 4440
rect 22980 4468 22986 4480
rect 24029 4471 24087 4477
rect 24029 4468 24041 4471
rect 22980 4440 24041 4468
rect 22980 4428 22986 4440
rect 24029 4437 24041 4440
rect 24075 4437 24087 4471
rect 24029 4431 24087 4437
rect 28215 4471 28273 4477
rect 28215 4437 28227 4471
rect 28261 4468 28273 4471
rect 28626 4468 28632 4480
rect 28261 4440 28632 4468
rect 28261 4437 28273 4440
rect 28215 4431 28273 4437
rect 28626 4428 28632 4440
rect 28684 4428 28690 4480
rect 30006 4468 30012 4480
rect 29967 4440 30012 4468
rect 30006 4428 30012 4440
rect 30064 4428 30070 4480
rect 30926 4468 30932 4480
rect 30887 4440 30932 4468
rect 30926 4428 30932 4440
rect 30984 4428 30990 4480
rect 31159 4471 31217 4477
rect 31159 4437 31171 4471
rect 31205 4468 31217 4471
rect 32490 4468 32496 4480
rect 31205 4440 32496 4468
rect 31205 4437 31217 4440
rect 31159 4431 31217 4437
rect 32490 4428 32496 4440
rect 32548 4428 32554 4480
rect 34790 4428 34796 4480
rect 34848 4468 34854 4480
rect 34977 4471 35035 4477
rect 34977 4468 34989 4471
rect 34848 4440 34989 4468
rect 34848 4428 34854 4440
rect 34977 4437 34989 4440
rect 35023 4437 35035 4471
rect 34977 4431 35035 4437
rect 35894 4428 35900 4480
rect 35952 4468 35958 4480
rect 38013 4471 38071 4477
rect 38013 4468 38025 4471
rect 35952 4440 38025 4468
rect 35952 4428 35958 4440
rect 38013 4437 38025 4440
rect 38059 4468 38071 4471
rect 38102 4468 38108 4480
rect 38059 4440 38108 4468
rect 38059 4437 38071 4440
rect 38013 4431 38071 4437
rect 38102 4428 38108 4440
rect 38160 4428 38166 4480
rect 1104 4378 48852 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 48852 4378
rect 1104 4304 48852 4326
rect 10045 4267 10103 4273
rect 10045 4233 10057 4267
rect 10091 4264 10103 4267
rect 10686 4264 10692 4276
rect 10091 4236 10692 4264
rect 10091 4233 10103 4236
rect 10045 4227 10103 4233
rect 10686 4224 10692 4236
rect 10744 4224 10750 4276
rect 12253 4267 12311 4273
rect 12253 4233 12265 4267
rect 12299 4264 12311 4267
rect 12342 4264 12348 4276
rect 12299 4236 12348 4264
rect 12299 4233 12311 4236
rect 12253 4227 12311 4233
rect 12342 4224 12348 4236
rect 12400 4264 12406 4276
rect 14366 4264 14372 4276
rect 12400 4236 14372 4264
rect 12400 4224 12406 4236
rect 14366 4224 14372 4236
rect 14424 4264 14430 4276
rect 15746 4264 15752 4276
rect 14424 4236 15752 4264
rect 14424 4224 14430 4236
rect 15746 4224 15752 4236
rect 15804 4224 15810 4276
rect 16482 4264 16488 4276
rect 16443 4236 16488 4264
rect 16482 4224 16488 4236
rect 16540 4224 16546 4276
rect 16850 4224 16856 4276
rect 16908 4264 16914 4276
rect 17083 4267 17141 4273
rect 17083 4264 17095 4267
rect 16908 4236 17095 4264
rect 16908 4224 16914 4236
rect 17083 4233 17095 4236
rect 17129 4233 17141 4267
rect 17083 4227 17141 4233
rect 17497 4267 17555 4273
rect 17497 4233 17509 4267
rect 17543 4264 17555 4267
rect 17586 4264 17592 4276
rect 17543 4236 17592 4264
rect 17543 4233 17555 4236
rect 17497 4227 17555 4233
rect 17586 4224 17592 4236
rect 17644 4224 17650 4276
rect 17862 4264 17868 4276
rect 17823 4236 17868 4264
rect 17862 4224 17868 4236
rect 17920 4224 17926 4276
rect 19518 4264 19524 4276
rect 19479 4236 19524 4264
rect 19518 4224 19524 4236
rect 19576 4224 19582 4276
rect 20165 4267 20223 4273
rect 20165 4233 20177 4267
rect 20211 4264 20223 4267
rect 20622 4264 20628 4276
rect 20211 4236 20628 4264
rect 20211 4233 20223 4236
rect 20165 4227 20223 4233
rect 20622 4224 20628 4236
rect 20680 4224 20686 4276
rect 21266 4224 21272 4276
rect 21324 4264 21330 4276
rect 22005 4267 22063 4273
rect 22005 4264 22017 4267
rect 21324 4236 22017 4264
rect 21324 4224 21330 4236
rect 22005 4233 22017 4236
rect 22051 4233 22063 4267
rect 22005 4227 22063 4233
rect 22465 4267 22523 4273
rect 22465 4233 22477 4267
rect 22511 4264 22523 4267
rect 22554 4264 22560 4276
rect 22511 4236 22560 4264
rect 22511 4233 22523 4236
rect 22465 4227 22523 4233
rect 22554 4224 22560 4236
rect 22612 4224 22618 4276
rect 25406 4224 25412 4276
rect 25464 4264 25470 4276
rect 28629 4267 28687 4273
rect 28629 4264 28641 4267
rect 25464 4236 28641 4264
rect 25464 4224 25470 4236
rect 28629 4233 28641 4236
rect 28675 4264 28687 4267
rect 28813 4267 28871 4273
rect 28813 4264 28825 4267
rect 28675 4236 28825 4264
rect 28675 4233 28687 4236
rect 28629 4227 28687 4233
rect 28813 4233 28825 4236
rect 28859 4233 28871 4267
rect 30374 4264 30380 4276
rect 30335 4236 30380 4264
rect 28813 4227 28871 4233
rect 30374 4224 30380 4236
rect 30432 4224 30438 4276
rect 30745 4267 30803 4273
rect 30745 4233 30757 4267
rect 30791 4264 30803 4267
rect 31018 4264 31024 4276
rect 30791 4236 31024 4264
rect 30791 4233 30803 4236
rect 30745 4227 30803 4233
rect 31018 4224 31024 4236
rect 31076 4264 31082 4276
rect 33318 4264 33324 4276
rect 31076 4236 33324 4264
rect 31076 4224 31082 4236
rect 33318 4224 33324 4236
rect 33376 4224 33382 4276
rect 33502 4224 33508 4276
rect 33560 4264 33566 4276
rect 34238 4264 34244 4276
rect 33560 4236 34244 4264
rect 33560 4224 33566 4236
rect 34238 4224 34244 4236
rect 34296 4224 34302 4276
rect 35986 4264 35992 4276
rect 35947 4236 35992 4264
rect 35986 4224 35992 4236
rect 36044 4224 36050 4276
rect 36630 4224 36636 4276
rect 36688 4264 36694 4276
rect 37829 4267 37887 4273
rect 37829 4264 37841 4267
rect 36688 4236 37841 4264
rect 36688 4224 36694 4236
rect 37829 4233 37841 4236
rect 37875 4264 37887 4267
rect 38194 4264 38200 4276
rect 37875 4236 38200 4264
rect 37875 4233 37887 4236
rect 37829 4227 37887 4233
rect 38194 4224 38200 4236
rect 38252 4224 38258 4276
rect 10413 4199 10471 4205
rect 10413 4165 10425 4199
rect 10459 4196 10471 4199
rect 10502 4196 10508 4208
rect 10459 4168 10508 4196
rect 10459 4165 10471 4168
rect 10413 4159 10471 4165
rect 10502 4156 10508 4168
rect 10560 4156 10566 4208
rect 11425 4199 11483 4205
rect 11425 4165 11437 4199
rect 11471 4196 11483 4199
rect 13630 4196 13636 4208
rect 11471 4168 13636 4196
rect 11471 4165 11483 4168
rect 11425 4159 11483 4165
rect 13630 4156 13636 4168
rect 13688 4156 13694 4208
rect 26694 4196 26700 4208
rect 26655 4168 26700 4196
rect 26694 4156 26700 4168
rect 26752 4156 26758 4208
rect 28166 4196 28172 4208
rect 28127 4168 28172 4196
rect 28166 4156 28172 4168
rect 28224 4156 28230 4208
rect 29086 4196 29092 4208
rect 29047 4168 29092 4196
rect 29086 4156 29092 4168
rect 29144 4156 29150 4208
rect 32214 4196 32220 4208
rect 32175 4168 32220 4196
rect 32214 4156 32220 4168
rect 32272 4156 32278 4208
rect 33042 4196 33048 4208
rect 32324 4168 32628 4196
rect 33003 4168 33048 4196
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 10873 4131 10931 4137
rect 10873 4128 10885 4131
rect 9640 4100 10885 4128
rect 9640 4088 9646 4100
rect 10873 4097 10885 4100
rect 10919 4128 10931 4131
rect 11793 4131 11851 4137
rect 11793 4128 11805 4131
rect 10919 4100 11805 4128
rect 10919 4097 10931 4100
rect 10873 4091 10931 4097
rect 11793 4097 11805 4100
rect 11839 4097 11851 4131
rect 11793 4091 11851 4097
rect 12710 4088 12716 4140
rect 12768 4128 12774 4140
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12768 4100 12909 4128
rect 12768 4088 12774 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 14182 4128 14188 4140
rect 14143 4100 14188 4128
rect 12897 4091 12955 4097
rect 14182 4088 14188 4100
rect 14240 4088 14246 4140
rect 18414 4128 18420 4140
rect 18375 4100 18420 4128
rect 18414 4088 18420 4100
rect 18472 4088 18478 4140
rect 18782 4088 18788 4140
rect 18840 4128 18846 4140
rect 19751 4131 19809 4137
rect 19751 4128 19763 4131
rect 18840 4100 19763 4128
rect 18840 4088 18846 4100
rect 19751 4097 19763 4100
rect 19797 4097 19809 4131
rect 19751 4091 19809 4097
rect 20809 4131 20867 4137
rect 20809 4097 20821 4131
rect 20855 4128 20867 4131
rect 20990 4128 20996 4140
rect 20855 4100 20996 4128
rect 20855 4097 20867 4100
rect 20809 4091 20867 4097
rect 20990 4088 20996 4100
rect 21048 4088 21054 4140
rect 26786 4128 26792 4140
rect 26747 4100 26792 4128
rect 26786 4088 26792 4100
rect 26844 4088 26850 4140
rect 28813 4131 28871 4137
rect 28813 4097 28825 4131
rect 28859 4128 28871 4131
rect 29365 4131 29423 4137
rect 29365 4128 29377 4131
rect 28859 4100 29377 4128
rect 28859 4097 28871 4100
rect 28813 4091 28871 4097
rect 29365 4097 29377 4100
rect 29411 4097 29423 4131
rect 29365 4091 29423 4097
rect 29822 4088 29828 4140
rect 29880 4128 29886 4140
rect 30009 4131 30067 4137
rect 30009 4128 30021 4131
rect 29880 4100 30021 4128
rect 29880 4088 29886 4100
rect 30009 4097 30021 4100
rect 30055 4128 30067 4131
rect 32324 4128 32352 4168
rect 32490 4128 32496 4140
rect 30055 4100 32352 4128
rect 32451 4100 32496 4128
rect 30055 4097 30067 4100
rect 30009 4091 30067 4097
rect 32490 4088 32496 4100
rect 32548 4088 32554 4140
rect 32600 4128 32628 4168
rect 33042 4156 33048 4168
rect 33100 4156 33106 4208
rect 36354 4156 36360 4208
rect 36412 4196 36418 4208
rect 36412 4168 38424 4196
rect 36412 4156 36418 4168
rect 34790 4128 34796 4140
rect 32600 4100 34796 4128
rect 34790 4088 34796 4100
rect 34848 4128 34854 4140
rect 34977 4131 35035 4137
rect 34977 4128 34989 4131
rect 34848 4100 34989 4128
rect 34848 4088 34854 4100
rect 34977 4097 34989 4100
rect 35023 4097 35035 4131
rect 34977 4091 35035 4097
rect 35621 4131 35679 4137
rect 35621 4097 35633 4131
rect 35667 4128 35679 4131
rect 35894 4128 35900 4140
rect 35667 4100 35900 4128
rect 35667 4097 35679 4100
rect 35621 4091 35679 4097
rect 35894 4088 35900 4100
rect 35952 4088 35958 4140
rect 36262 4088 36268 4140
rect 36320 4128 36326 4140
rect 36541 4131 36599 4137
rect 36541 4128 36553 4131
rect 36320 4100 36553 4128
rect 36320 4088 36326 4100
rect 36541 4097 36553 4100
rect 36587 4097 36599 4131
rect 36814 4128 36820 4140
rect 36775 4100 36820 4128
rect 36541 4091 36599 4097
rect 36814 4088 36820 4100
rect 36872 4088 36878 4140
rect 38102 4128 38108 4140
rect 38063 4100 38108 4128
rect 38102 4088 38108 4100
rect 38160 4088 38166 4140
rect 38396 4137 38424 4168
rect 38381 4131 38439 4137
rect 38381 4128 38393 4131
rect 38359 4100 38393 4128
rect 38381 4097 38393 4100
rect 38427 4097 38439 4131
rect 38381 4091 38439 4097
rect 12342 4020 12348 4072
rect 12400 4060 12406 4072
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 12400 4032 12449 4060
rect 12400 4020 12406 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 12618 4060 12624 4072
rect 12579 4032 12624 4060
rect 12437 4023 12495 4029
rect 12618 4020 12624 4032
rect 12676 4060 12682 4072
rect 13262 4060 13268 4072
rect 12676 4032 13268 4060
rect 12676 4020 12682 4032
rect 13262 4020 13268 4032
rect 13320 4020 13326 4072
rect 13817 4063 13875 4069
rect 13817 4029 13829 4063
rect 13863 4029 13875 4063
rect 13817 4023 13875 4029
rect 10965 3995 11023 4001
rect 10965 3961 10977 3995
rect 11011 3992 11023 3995
rect 11330 3992 11336 4004
rect 11011 3964 11336 3992
rect 11011 3961 11023 3964
rect 10965 3955 11023 3961
rect 11330 3952 11336 3964
rect 11388 3952 11394 4004
rect 13630 3924 13636 3936
rect 13591 3896 13636 3924
rect 13630 3884 13636 3896
rect 13688 3924 13694 3936
rect 13832 3924 13860 4023
rect 15470 4020 15476 4072
rect 15528 4060 15534 4072
rect 15657 4063 15715 4069
rect 15657 4060 15669 4063
rect 15528 4032 15669 4060
rect 15528 4020 15534 4032
rect 15657 4029 15669 4032
rect 15703 4029 15715 4063
rect 16980 4063 17038 4069
rect 16980 4060 16992 4063
rect 15657 4023 15715 4029
rect 16776 4032 16992 4060
rect 14550 3952 14556 4004
rect 14608 3952 14614 4004
rect 16114 3924 16120 3936
rect 13688 3896 13860 3924
rect 16075 3896 16120 3924
rect 13688 3884 13694 3896
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 16574 3884 16580 3936
rect 16632 3924 16638 3936
rect 16776 3933 16804 4032
rect 16980 4029 16992 4032
rect 17026 4029 17038 4063
rect 19648 4063 19706 4069
rect 19648 4060 19660 4063
rect 16980 4023 17038 4029
rect 19076 4032 19660 4060
rect 17770 3952 17776 4004
rect 17828 3992 17834 4004
rect 18141 3995 18199 4001
rect 18141 3992 18153 3995
rect 17828 3964 18153 3992
rect 17828 3952 17834 3964
rect 18141 3961 18153 3964
rect 18187 3961 18199 3995
rect 18141 3955 18199 3961
rect 18230 3952 18236 4004
rect 18288 3992 18294 4004
rect 18288 3964 18333 3992
rect 18288 3952 18294 3964
rect 16761 3927 16819 3933
rect 16761 3924 16773 3927
rect 16632 3896 16773 3924
rect 16632 3884 16638 3896
rect 16761 3893 16773 3896
rect 16807 3893 16819 3927
rect 16761 3887 16819 3893
rect 18874 3884 18880 3936
rect 18932 3924 18938 3936
rect 19076 3933 19104 4032
rect 19648 4029 19660 4032
rect 19694 4060 19706 4063
rect 19886 4060 19892 4072
rect 19694 4032 19892 4060
rect 19694 4029 19706 4032
rect 19648 4023 19706 4029
rect 19886 4020 19892 4032
rect 19944 4020 19950 4072
rect 22624 4063 22682 4069
rect 22624 4029 22636 4063
rect 22670 4060 22682 4063
rect 22922 4060 22928 4072
rect 22670 4032 22928 4060
rect 22670 4029 22682 4032
rect 22624 4023 22682 4029
rect 22922 4020 22928 4032
rect 22980 4020 22986 4072
rect 23658 4060 23664 4072
rect 23619 4032 23664 4060
rect 23658 4020 23664 4032
rect 23716 4020 23722 4072
rect 25498 4020 25504 4072
rect 25556 4060 25562 4072
rect 25628 4063 25686 4069
rect 25628 4060 25640 4063
rect 25556 4032 25640 4060
rect 25556 4020 25562 4032
rect 25628 4029 25640 4032
rect 25674 4029 25686 4063
rect 25628 4023 25686 4029
rect 19150 3952 19156 4004
rect 19208 3992 19214 4004
rect 20530 3992 20536 4004
rect 19208 3964 20536 3992
rect 19208 3952 19214 3964
rect 20530 3952 20536 3964
rect 20588 3952 20594 4004
rect 20714 3992 20720 4004
rect 20675 3964 20720 3992
rect 20714 3952 20720 3964
rect 20772 3992 20778 4004
rect 21130 3995 21188 4001
rect 21130 3992 21142 3995
rect 20772 3964 21142 3992
rect 20772 3952 20778 3964
rect 21130 3961 21142 3964
rect 21176 3961 21188 3995
rect 21130 3955 21188 3961
rect 23201 3995 23259 4001
rect 23201 3961 23213 3995
rect 23247 3992 23259 3995
rect 23842 3992 23848 4004
rect 23247 3964 23848 3992
rect 23247 3961 23259 3964
rect 23201 3955 23259 3961
rect 23842 3952 23848 3964
rect 23900 3992 23906 4004
rect 24023 3995 24081 4001
rect 24023 3992 24035 3995
rect 23900 3964 24035 3992
rect 23900 3952 23906 3964
rect 24023 3961 24035 3964
rect 24069 3992 24081 3995
rect 24486 3992 24492 4004
rect 24069 3964 24492 3992
rect 24069 3961 24081 3964
rect 24023 3955 24081 3961
rect 24486 3952 24492 3964
rect 24544 3952 24550 4004
rect 26694 3952 26700 4004
rect 26752 3992 26758 4004
rect 27151 3995 27209 4001
rect 27151 3992 27163 3995
rect 26752 3964 27163 3992
rect 26752 3952 26758 3964
rect 27151 3961 27163 3964
rect 27197 3961 27209 3995
rect 27151 3955 27209 3961
rect 27338 3952 27344 4004
rect 27396 3992 27402 4004
rect 29454 3992 29460 4004
rect 27396 3964 28523 3992
rect 29415 3964 29460 3992
rect 27396 3952 27402 3964
rect 19061 3927 19119 3933
rect 19061 3924 19073 3927
rect 18932 3896 19073 3924
rect 18932 3884 18938 3896
rect 19061 3893 19073 3896
rect 19107 3893 19119 3927
rect 21726 3924 21732 3936
rect 21687 3896 21732 3924
rect 19061 3887 19119 3893
rect 21726 3884 21732 3896
rect 21784 3884 21790 3936
rect 22695 3927 22753 3933
rect 22695 3893 22707 3927
rect 22741 3924 22753 3927
rect 23290 3924 23296 3936
rect 22741 3896 23296 3924
rect 22741 3893 22753 3896
rect 22695 3887 22753 3893
rect 23290 3884 23296 3896
rect 23348 3884 23354 3936
rect 24578 3924 24584 3936
rect 24539 3896 24584 3924
rect 24578 3884 24584 3896
rect 24636 3884 24642 3936
rect 24949 3927 25007 3933
rect 24949 3893 24961 3927
rect 24995 3924 25007 3927
rect 25038 3924 25044 3936
rect 24995 3896 25044 3924
rect 24995 3893 25007 3896
rect 24949 3887 25007 3893
rect 25038 3884 25044 3896
rect 25096 3884 25102 3936
rect 25222 3924 25228 3936
rect 25183 3896 25228 3924
rect 25222 3884 25228 3896
rect 25280 3884 25286 3936
rect 25731 3927 25789 3933
rect 25731 3893 25743 3927
rect 25777 3924 25789 3927
rect 26050 3924 26056 3936
rect 25777 3896 26056 3924
rect 25777 3893 25789 3896
rect 25731 3887 25789 3893
rect 26050 3884 26056 3896
rect 26108 3884 26114 3936
rect 26329 3927 26387 3933
rect 26329 3893 26341 3927
rect 26375 3924 26387 3927
rect 27062 3924 27068 3936
rect 26375 3896 27068 3924
rect 26375 3893 26387 3896
rect 26329 3887 26387 3893
rect 27062 3884 27068 3896
rect 27120 3884 27126 3936
rect 27709 3927 27767 3933
rect 27709 3893 27721 3927
rect 27755 3924 27767 3927
rect 28258 3924 28264 3936
rect 27755 3896 28264 3924
rect 27755 3893 27767 3896
rect 27709 3887 27767 3893
rect 28258 3884 28264 3896
rect 28316 3884 28322 3936
rect 28495 3924 28523 3964
rect 29454 3952 29460 3964
rect 29512 3952 29518 4004
rect 30926 3992 30932 4004
rect 30839 3964 30932 3992
rect 30926 3952 30932 3964
rect 30984 3952 30990 4004
rect 31018 3952 31024 4004
rect 31076 3992 31082 4004
rect 31573 3995 31631 4001
rect 31076 3964 31121 3992
rect 31076 3952 31082 3964
rect 31573 3961 31585 3995
rect 31619 3992 31631 3995
rect 32306 3992 32312 4004
rect 31619 3964 32312 3992
rect 31619 3961 31631 3964
rect 31573 3955 31631 3961
rect 32306 3952 32312 3964
rect 32364 3952 32370 4004
rect 32585 3995 32643 4001
rect 32585 3961 32597 3995
rect 32631 3992 32643 3995
rect 34330 3992 34336 4004
rect 32631 3964 34336 3992
rect 32631 3961 32643 3964
rect 32585 3955 32643 3961
rect 30944 3924 30972 3952
rect 31938 3924 31944 3936
rect 28495 3896 30972 3924
rect 31851 3896 31944 3924
rect 31938 3884 31944 3896
rect 31996 3924 32002 3936
rect 32600 3924 32628 3955
rect 34330 3952 34336 3964
rect 34388 3952 34394 4004
rect 34701 3995 34759 4001
rect 34701 3961 34713 3995
rect 34747 3992 34759 3995
rect 35066 3992 35072 4004
rect 34747 3964 35072 3992
rect 34747 3961 34759 3964
rect 34701 3955 34759 3961
rect 35066 3952 35072 3964
rect 35124 3952 35130 4004
rect 36633 3995 36691 4001
rect 36633 3961 36645 3995
rect 36679 3961 36691 3995
rect 36633 3955 36691 3961
rect 31996 3896 32628 3924
rect 31996 3884 32002 3896
rect 33318 3884 33324 3936
rect 33376 3924 33382 3936
rect 33965 3927 34023 3933
rect 33965 3924 33977 3927
rect 33376 3896 33977 3924
rect 33376 3884 33382 3896
rect 33965 3893 33977 3896
rect 34011 3924 34023 3927
rect 34146 3924 34152 3936
rect 34011 3896 34152 3924
rect 34011 3893 34023 3896
rect 33965 3887 34023 3893
rect 34146 3884 34152 3896
rect 34204 3884 34210 3936
rect 36354 3924 36360 3936
rect 36315 3896 36360 3924
rect 36354 3884 36360 3896
rect 36412 3924 36418 3936
rect 36648 3924 36676 3955
rect 38194 3952 38200 4004
rect 38252 3992 38258 4004
rect 38252 3964 38297 3992
rect 38252 3952 38258 3964
rect 36412 3896 36676 3924
rect 36412 3884 36418 3896
rect 1104 3834 48852 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 48852 3834
rect 1104 3760 48852 3782
rect 11011 3723 11069 3729
rect 11011 3689 11023 3723
rect 11057 3720 11069 3723
rect 11238 3720 11244 3732
rect 11057 3692 11244 3720
rect 11057 3689 11069 3692
rect 11011 3683 11069 3689
rect 11238 3680 11244 3692
rect 11296 3680 11302 3732
rect 11422 3720 11428 3732
rect 11383 3692 11428 3720
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 14550 3720 14556 3732
rect 13372 3692 14556 3720
rect 13372 3624 13400 3692
rect 14550 3680 14556 3692
rect 14608 3680 14614 3732
rect 16022 3720 16028 3732
rect 15983 3692 16028 3720
rect 16022 3680 16028 3692
rect 16080 3680 16086 3732
rect 16482 3680 16488 3732
rect 16540 3720 16546 3732
rect 16577 3723 16635 3729
rect 16577 3720 16589 3723
rect 16540 3692 16589 3720
rect 16540 3680 16546 3692
rect 16577 3689 16589 3692
rect 16623 3689 16635 3723
rect 16577 3683 16635 3689
rect 17129 3723 17187 3729
rect 17129 3689 17141 3723
rect 17175 3720 17187 3723
rect 17865 3723 17923 3729
rect 17865 3720 17877 3723
rect 17175 3692 17877 3720
rect 17175 3689 17187 3692
rect 17129 3683 17187 3689
rect 17865 3689 17877 3692
rect 17911 3720 17923 3723
rect 18230 3720 18236 3732
rect 17911 3692 18236 3720
rect 17911 3689 17923 3692
rect 17865 3683 17923 3689
rect 18230 3680 18236 3692
rect 18288 3680 18294 3732
rect 20717 3723 20775 3729
rect 20717 3689 20729 3723
rect 20763 3720 20775 3723
rect 20990 3720 20996 3732
rect 20763 3692 20996 3720
rect 20763 3689 20775 3692
rect 20717 3683 20775 3689
rect 20990 3680 20996 3692
rect 21048 3680 21054 3732
rect 23658 3680 23664 3732
rect 23716 3720 23722 3732
rect 24121 3723 24179 3729
rect 24121 3720 24133 3723
rect 23716 3692 24133 3720
rect 23716 3680 23722 3692
rect 24121 3689 24133 3692
rect 24167 3689 24179 3723
rect 24121 3683 24179 3689
rect 25498 3680 25504 3732
rect 25556 3720 25562 3732
rect 25869 3723 25927 3729
rect 25869 3720 25881 3723
rect 25556 3692 25881 3720
rect 25556 3680 25562 3692
rect 25869 3689 25881 3692
rect 25915 3689 25927 3723
rect 26602 3720 26608 3732
rect 26561 3692 26608 3720
rect 25869 3683 25927 3689
rect 26602 3680 26608 3692
rect 26660 3729 26666 3732
rect 26660 3723 26709 3729
rect 26660 3689 26663 3723
rect 26697 3720 26709 3723
rect 26973 3723 27031 3729
rect 26973 3720 26985 3723
rect 26697 3692 26985 3720
rect 26697 3689 26709 3692
rect 26660 3683 26709 3689
rect 26973 3689 26985 3692
rect 27019 3689 27031 3723
rect 26973 3683 27031 3689
rect 26660 3680 26666 3683
rect 28626 3680 28632 3732
rect 28684 3720 28690 3732
rect 29733 3723 29791 3729
rect 28684 3692 29500 3720
rect 28684 3680 28690 3692
rect 18138 3652 18144 3664
rect 18099 3624 18144 3652
rect 18138 3612 18144 3624
rect 18196 3612 18202 3664
rect 22646 3612 22652 3664
rect 22704 3652 22710 3664
rect 22919 3655 22977 3661
rect 22919 3652 22931 3655
rect 22704 3624 22931 3652
rect 22704 3612 22710 3624
rect 22919 3621 22931 3624
rect 22965 3652 22977 3655
rect 23842 3652 23848 3664
rect 22965 3624 23848 3652
rect 22965 3621 22977 3624
rect 22919 3615 22977 3621
rect 23842 3612 23848 3624
rect 23900 3612 23906 3664
rect 25038 3652 25044 3664
rect 24999 3624 25044 3652
rect 25038 3612 25044 3624
rect 25096 3612 25102 3664
rect 25593 3655 25651 3661
rect 25593 3621 25605 3655
rect 25639 3652 25651 3655
rect 27338 3652 27344 3664
rect 25639 3624 27344 3652
rect 25639 3621 25651 3624
rect 25593 3615 25651 3621
rect 27338 3612 27344 3624
rect 27396 3612 27402 3664
rect 28166 3652 28172 3664
rect 28127 3624 28172 3652
rect 28166 3612 28172 3624
rect 28224 3612 28230 3664
rect 28721 3655 28779 3661
rect 28721 3621 28733 3655
rect 28767 3652 28779 3655
rect 28810 3652 28816 3664
rect 28767 3624 28816 3652
rect 28767 3621 28779 3624
rect 28721 3615 28779 3621
rect 28810 3612 28816 3624
rect 28868 3612 28874 3664
rect 29472 3652 29500 3692
rect 29733 3689 29745 3723
rect 29779 3720 29791 3723
rect 30006 3720 30012 3732
rect 29779 3692 30012 3720
rect 29779 3689 29791 3692
rect 29733 3683 29791 3689
rect 30006 3680 30012 3692
rect 30064 3680 30070 3732
rect 30377 3723 30435 3729
rect 30377 3689 30389 3723
rect 30423 3720 30435 3723
rect 32030 3720 32036 3732
rect 30423 3692 32036 3720
rect 30423 3689 30435 3692
rect 30377 3683 30435 3689
rect 32030 3680 32036 3692
rect 32088 3720 32094 3732
rect 32088 3692 32352 3720
rect 32088 3680 32094 3692
rect 30558 3652 30564 3664
rect 29472 3624 30564 3652
rect 30558 3612 30564 3624
rect 30616 3612 30622 3664
rect 30653 3655 30711 3661
rect 30653 3621 30665 3655
rect 30699 3652 30711 3655
rect 30742 3652 30748 3664
rect 30699 3624 30748 3652
rect 30699 3621 30711 3624
rect 30653 3615 30711 3621
rect 30742 3612 30748 3624
rect 30800 3652 30806 3664
rect 32214 3652 32220 3664
rect 30800 3624 32220 3652
rect 30800 3612 30806 3624
rect 32214 3612 32220 3624
rect 32272 3612 32278 3664
rect 32324 3661 32352 3692
rect 32490 3680 32496 3732
rect 32548 3720 32554 3732
rect 33137 3723 33195 3729
rect 33137 3720 33149 3723
rect 32548 3692 33149 3720
rect 32548 3680 32554 3692
rect 33137 3689 33149 3692
rect 33183 3689 33195 3723
rect 34698 3720 34704 3732
rect 34659 3692 34704 3720
rect 33137 3683 33195 3689
rect 34698 3680 34704 3692
rect 34756 3680 34762 3732
rect 36262 3680 36268 3732
rect 36320 3720 36326 3732
rect 36541 3723 36599 3729
rect 36541 3720 36553 3723
rect 36320 3692 36553 3720
rect 36320 3680 36326 3692
rect 36541 3689 36553 3692
rect 36587 3689 36599 3723
rect 36541 3683 36599 3689
rect 32309 3655 32367 3661
rect 32309 3621 32321 3655
rect 32355 3652 32367 3655
rect 32355 3624 32904 3652
rect 32355 3621 32367 3624
rect 32309 3615 32367 3621
rect 10940 3587 10998 3593
rect 10940 3553 10952 3587
rect 10986 3584 10998 3587
rect 11514 3584 11520 3596
rect 10986 3556 11520 3584
rect 10986 3553 10998 3556
rect 10940 3547 10998 3553
rect 11514 3544 11520 3556
rect 11572 3544 11578 3596
rect 13722 3584 13728 3596
rect 13683 3556 13728 3584
rect 13722 3544 13728 3556
rect 13780 3544 13786 3596
rect 19150 3544 19156 3596
rect 19208 3584 19214 3596
rect 19556 3587 19614 3593
rect 19556 3584 19568 3587
rect 19208 3556 19568 3584
rect 19208 3544 19214 3556
rect 19556 3553 19568 3556
rect 19602 3584 19614 3587
rect 19886 3584 19892 3596
rect 19602 3556 19892 3584
rect 19602 3553 19614 3556
rect 19556 3547 19614 3553
rect 19886 3544 19892 3556
rect 19944 3544 19950 3596
rect 20898 3584 20904 3596
rect 20859 3556 20904 3584
rect 20898 3544 20904 3556
rect 20956 3544 20962 3596
rect 21358 3584 21364 3596
rect 21319 3556 21364 3584
rect 21358 3544 21364 3556
rect 21416 3544 21422 3596
rect 22186 3544 22192 3596
rect 22244 3584 22250 3596
rect 22557 3587 22615 3593
rect 22557 3584 22569 3587
rect 22244 3556 22569 3584
rect 22244 3544 22250 3556
rect 22557 3553 22569 3556
rect 22603 3553 22615 3587
rect 26418 3584 26424 3596
rect 26379 3556 26424 3584
rect 22557 3547 22615 3553
rect 26418 3544 26424 3556
rect 26476 3544 26482 3596
rect 29365 3587 29423 3593
rect 29365 3553 29377 3587
rect 29411 3584 29423 3587
rect 29454 3584 29460 3596
rect 29411 3556 29460 3584
rect 29411 3553 29423 3556
rect 29365 3547 29423 3553
rect 29454 3544 29460 3556
rect 29512 3584 29518 3596
rect 30377 3587 30435 3593
rect 30377 3584 30389 3587
rect 29512 3556 30389 3584
rect 29512 3544 29518 3556
rect 30377 3553 30389 3556
rect 30423 3553 30435 3587
rect 32876 3584 32904 3624
rect 33042 3612 33048 3664
rect 33100 3652 33106 3664
rect 33502 3652 33508 3664
rect 33100 3624 33508 3652
rect 33100 3612 33106 3624
rect 33502 3612 33508 3624
rect 33560 3612 33566 3664
rect 33870 3652 33876 3664
rect 33612 3624 33876 3652
rect 33612 3584 33640 3624
rect 33870 3612 33876 3624
rect 33928 3612 33934 3664
rect 35066 3612 35072 3664
rect 35124 3652 35130 3664
rect 35250 3652 35256 3664
rect 35124 3624 35256 3652
rect 35124 3612 35130 3624
rect 35250 3612 35256 3624
rect 35308 3652 35314 3664
rect 35529 3655 35587 3661
rect 35529 3652 35541 3655
rect 35308 3624 35541 3652
rect 35308 3612 35314 3624
rect 35529 3621 35541 3624
rect 35575 3621 35587 3655
rect 35529 3615 35587 3621
rect 32876 3556 33640 3584
rect 30377 3547 30435 3553
rect 35434 3544 35440 3596
rect 35492 3584 35498 3596
rect 35621 3587 35679 3593
rect 35621 3584 35633 3587
rect 35492 3556 35633 3584
rect 35492 3544 35498 3556
rect 35621 3553 35633 3556
rect 35667 3553 35679 3587
rect 37734 3584 37740 3596
rect 37695 3556 37740 3584
rect 35621 3547 35679 3553
rect 37734 3544 37740 3556
rect 37792 3544 37798 3596
rect 11882 3516 11888 3528
rect 11843 3488 11888 3516
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 12253 3519 12311 3525
rect 12253 3485 12265 3519
rect 12299 3516 12311 3519
rect 12434 3516 12440 3528
rect 12299 3488 12440 3516
rect 12299 3485 12311 3488
rect 12253 3479 12311 3485
rect 12434 3476 12440 3488
rect 12492 3476 12498 3528
rect 16206 3516 16212 3528
rect 16119 3488 16212 3516
rect 16206 3476 16212 3488
rect 16264 3516 16270 3528
rect 16758 3516 16764 3528
rect 16264 3488 16764 3516
rect 16264 3476 16270 3488
rect 16758 3476 16764 3488
rect 16816 3476 16822 3528
rect 18049 3519 18107 3525
rect 18049 3485 18061 3519
rect 18095 3516 18107 3519
rect 18230 3516 18236 3528
rect 18095 3488 18236 3516
rect 18095 3485 18107 3488
rect 18049 3479 18107 3485
rect 18230 3476 18236 3488
rect 18288 3476 18294 3528
rect 18325 3519 18383 3525
rect 18325 3485 18337 3519
rect 18371 3516 18383 3519
rect 18414 3516 18420 3528
rect 18371 3488 18420 3516
rect 18371 3485 18383 3488
rect 18325 3479 18383 3485
rect 13354 3408 13360 3460
rect 13412 3448 13418 3460
rect 14829 3451 14887 3457
rect 14829 3448 14841 3451
rect 13412 3420 14841 3448
rect 13412 3408 13418 3420
rect 14829 3417 14841 3420
rect 14875 3417 14887 3451
rect 14829 3411 14887 3417
rect 15562 3408 15568 3460
rect 15620 3448 15626 3460
rect 18340 3448 18368 3479
rect 18414 3476 18420 3488
rect 18472 3476 18478 3528
rect 21450 3516 21456 3528
rect 21411 3488 21456 3516
rect 21450 3476 21456 3488
rect 21508 3476 21514 3528
rect 24949 3519 25007 3525
rect 24949 3485 24961 3519
rect 24995 3516 25007 3519
rect 26050 3516 26056 3528
rect 24995 3488 26056 3516
rect 24995 3485 25007 3488
rect 24949 3479 25007 3485
rect 26050 3476 26056 3488
rect 26108 3476 26114 3528
rect 26970 3476 26976 3528
rect 27028 3516 27034 3528
rect 28077 3519 28135 3525
rect 28077 3516 28089 3519
rect 27028 3488 28089 3516
rect 27028 3476 27034 3488
rect 28077 3485 28089 3488
rect 28123 3516 28135 3519
rect 28994 3516 29000 3528
rect 28123 3488 29000 3516
rect 28123 3485 28135 3488
rect 28077 3479 28135 3485
rect 28994 3476 29000 3488
rect 29052 3476 29058 3528
rect 31202 3516 31208 3528
rect 31115 3488 31208 3516
rect 31202 3476 31208 3488
rect 31260 3516 31266 3528
rect 32214 3516 32220 3528
rect 31260 3488 32220 3516
rect 31260 3476 31266 3488
rect 32214 3476 32220 3488
rect 32272 3476 32278 3528
rect 32306 3476 32312 3528
rect 32364 3516 32370 3528
rect 32493 3519 32551 3525
rect 32493 3516 32505 3519
rect 32364 3488 32505 3516
rect 32364 3476 32370 3488
rect 32493 3485 32505 3488
rect 32539 3516 32551 3519
rect 32539 3488 33134 3516
rect 32539 3485 32551 3488
rect 32493 3479 32551 3485
rect 15620 3420 18368 3448
rect 15620 3408 15626 3420
rect 21174 3408 21180 3460
rect 21232 3448 21238 3460
rect 21913 3451 21971 3457
rect 21913 3448 21925 3451
rect 21232 3420 21925 3448
rect 21232 3408 21238 3420
rect 21913 3417 21925 3420
rect 21959 3417 21971 3451
rect 33106 3448 33134 3488
rect 33502 3476 33508 3528
rect 33560 3516 33566 3528
rect 33778 3516 33784 3528
rect 33560 3488 33784 3516
rect 33560 3476 33566 3488
rect 33778 3476 33784 3488
rect 33836 3476 33842 3528
rect 37093 3519 37151 3525
rect 37093 3516 37105 3519
rect 34256 3488 37105 3516
rect 34256 3448 34284 3488
rect 37093 3485 37105 3488
rect 37139 3516 37151 3519
rect 37182 3516 37188 3528
rect 37139 3488 37188 3516
rect 37139 3485 37151 3488
rect 37093 3479 37151 3485
rect 37182 3476 37188 3488
rect 37240 3476 37246 3528
rect 33106 3420 34284 3448
rect 21913 3411 21971 3417
rect 34330 3408 34336 3460
rect 34388 3448 34394 3460
rect 34606 3448 34612 3460
rect 34388 3420 34612 3448
rect 34388 3408 34394 3420
rect 34606 3408 34612 3420
rect 34664 3408 34670 3460
rect 1670 3340 1676 3392
rect 1728 3380 1734 3392
rect 9217 3383 9275 3389
rect 9217 3380 9229 3383
rect 1728 3352 9229 3380
rect 1728 3340 1734 3352
rect 9217 3349 9229 3352
rect 9263 3380 9275 3383
rect 9950 3380 9956 3392
rect 9263 3352 9956 3380
rect 9263 3349 9275 3352
rect 9217 3343 9275 3349
rect 9950 3340 9956 3352
rect 10008 3340 10014 3392
rect 11514 3340 11520 3392
rect 11572 3380 11578 3392
rect 11701 3383 11759 3389
rect 11701 3380 11713 3383
rect 11572 3352 11713 3380
rect 11572 3340 11578 3352
rect 11701 3349 11713 3352
rect 11747 3349 11759 3383
rect 14182 3380 14188 3392
rect 14143 3352 14188 3380
rect 11701 3343 11759 3349
rect 14182 3340 14188 3352
rect 14240 3340 14246 3392
rect 14274 3340 14280 3392
rect 14332 3380 14338 3392
rect 18874 3380 18880 3392
rect 14332 3352 18880 3380
rect 14332 3340 14338 3352
rect 18874 3340 18880 3352
rect 18932 3340 18938 3392
rect 18966 3340 18972 3392
rect 19024 3380 19030 3392
rect 19061 3383 19119 3389
rect 19061 3380 19073 3383
rect 19024 3352 19073 3380
rect 19024 3340 19030 3352
rect 19061 3349 19073 3352
rect 19107 3380 19119 3383
rect 19659 3383 19717 3389
rect 19659 3380 19671 3383
rect 19107 3352 19671 3380
rect 19107 3349 19119 3352
rect 19061 3343 19119 3349
rect 19659 3349 19671 3352
rect 19705 3349 19717 3383
rect 19659 3343 19717 3349
rect 23474 3340 23480 3392
rect 23532 3380 23538 3392
rect 24762 3380 24768 3392
rect 23532 3352 23577 3380
rect 24723 3352 24768 3380
rect 23532 3340 23538 3352
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 27706 3380 27712 3392
rect 27667 3352 27712 3380
rect 27706 3340 27712 3352
rect 27764 3340 27770 3392
rect 36170 3340 36176 3392
rect 36228 3380 36234 3392
rect 37921 3383 37979 3389
rect 37921 3380 37933 3383
rect 36228 3352 37933 3380
rect 36228 3340 36234 3352
rect 37921 3349 37933 3352
rect 37967 3349 37979 3383
rect 37921 3343 37979 3349
rect 1104 3290 48852 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 48852 3290
rect 1104 3216 48852 3238
rect 8662 3176 8668 3188
rect 8623 3148 8668 3176
rect 8662 3136 8668 3148
rect 8720 3136 8726 3188
rect 11514 3176 11520 3188
rect 11475 3148 11520 3176
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 12943 3179 13001 3185
rect 12943 3145 12955 3179
rect 12989 3176 13001 3179
rect 13354 3176 13360 3188
rect 12989 3148 13360 3176
rect 12989 3145 13001 3148
rect 12943 3139 13001 3145
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 13722 3136 13728 3188
rect 13780 3176 13786 3188
rect 15470 3176 15476 3188
rect 13780 3148 15476 3176
rect 13780 3136 13786 3148
rect 15470 3136 15476 3148
rect 15528 3176 15534 3188
rect 16117 3179 16175 3185
rect 15528 3148 15700 3176
rect 15528 3136 15534 3148
rect 8680 3040 8708 3136
rect 9585 3043 9643 3049
rect 9585 3040 9597 3043
rect 8680 3012 9597 3040
rect 9585 3009 9597 3012
rect 9631 3009 9643 3043
rect 9585 3003 9643 3009
rect 11882 3000 11888 3052
rect 11940 3040 11946 3052
rect 13630 3040 13636 3052
rect 11940 3012 13636 3040
rect 11940 3000 11946 3012
rect 13630 3000 13636 3012
rect 13688 3040 13694 3052
rect 13817 3043 13875 3049
rect 13817 3040 13829 3043
rect 13688 3012 13829 3040
rect 13688 3000 13694 3012
rect 13817 3009 13829 3012
rect 13863 3009 13875 3043
rect 13817 3003 13875 3009
rect 9217 2975 9275 2981
rect 9217 2972 9229 2975
rect 9048 2944 9229 2972
rect 9048 2848 9076 2944
rect 9217 2941 9229 2944
rect 9263 2941 9275 2975
rect 9217 2935 9275 2941
rect 10870 2932 10876 2984
rect 10928 2972 10934 2984
rect 11057 2975 11115 2981
rect 11057 2972 11069 2975
rect 10928 2944 11069 2972
rect 10928 2932 10934 2944
rect 11057 2941 11069 2944
rect 11103 2972 11115 2975
rect 12621 2975 12679 2981
rect 12621 2972 12633 2975
rect 11103 2944 12633 2972
rect 11103 2941 11115 2944
rect 11057 2935 11115 2941
rect 12621 2941 12633 2944
rect 12667 2972 12679 2975
rect 12710 2972 12716 2984
rect 12667 2944 12716 2972
rect 12667 2941 12679 2944
rect 12621 2935 12679 2941
rect 12710 2932 12716 2944
rect 12768 2932 12774 2984
rect 12805 2975 12863 2981
rect 12805 2941 12817 2975
rect 12851 2972 12863 2975
rect 12894 2972 12900 2984
rect 12851 2944 12900 2972
rect 12851 2941 12863 2944
rect 12805 2935 12863 2941
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 14185 2975 14243 2981
rect 14185 2941 14197 2975
rect 14231 2972 14243 2975
rect 14274 2972 14280 2984
rect 14231 2944 14280 2972
rect 14231 2941 14243 2944
rect 14185 2935 14243 2941
rect 14274 2932 14280 2944
rect 14332 2932 14338 2984
rect 15672 2981 15700 3148
rect 16117 3145 16129 3179
rect 16163 3176 16175 3179
rect 16574 3176 16580 3188
rect 16163 3148 16580 3176
rect 16163 3145 16175 3148
rect 16117 3139 16175 3145
rect 16574 3136 16580 3148
rect 16632 3136 16638 3188
rect 16758 3176 16764 3188
rect 16719 3148 16764 3176
rect 16758 3136 16764 3148
rect 16816 3136 16822 3188
rect 17083 3179 17141 3185
rect 17083 3145 17095 3179
rect 17129 3176 17141 3179
rect 17770 3176 17776 3188
rect 17129 3148 17776 3176
rect 17129 3145 17141 3148
rect 17083 3139 17141 3145
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 17865 3179 17923 3185
rect 17865 3145 17877 3179
rect 17911 3176 17923 3179
rect 18138 3176 18144 3188
rect 17911 3148 18144 3176
rect 17911 3145 17923 3148
rect 17865 3139 17923 3145
rect 18138 3136 18144 3148
rect 18196 3136 18202 3188
rect 19886 3176 19892 3188
rect 19847 3148 19892 3176
rect 19886 3136 19892 3148
rect 19944 3136 19950 3188
rect 20717 3179 20775 3185
rect 20717 3145 20729 3179
rect 20763 3176 20775 3179
rect 20898 3176 20904 3188
rect 20763 3148 20904 3176
rect 20763 3145 20775 3148
rect 20717 3139 20775 3145
rect 20898 3136 20904 3148
rect 20956 3136 20962 3188
rect 22186 3136 22192 3188
rect 22244 3176 22250 3188
rect 22925 3179 22983 3185
rect 22925 3176 22937 3179
rect 22244 3148 22937 3176
rect 22244 3136 22250 3148
rect 22925 3145 22937 3148
rect 22971 3145 22983 3179
rect 22925 3139 22983 3145
rect 23106 3136 23112 3188
rect 23164 3176 23170 3188
rect 23293 3179 23351 3185
rect 23293 3176 23305 3179
rect 23164 3148 23305 3176
rect 23164 3136 23170 3148
rect 23293 3145 23305 3148
rect 23339 3145 23351 3179
rect 23293 3139 23351 3145
rect 23799 3179 23857 3185
rect 23799 3145 23811 3179
rect 23845 3176 23857 3179
rect 24026 3176 24032 3188
rect 23845 3148 24032 3176
rect 23845 3145 23857 3148
rect 23799 3139 23857 3145
rect 24026 3136 24032 3148
rect 24084 3136 24090 3188
rect 26050 3176 26056 3188
rect 26011 3148 26056 3176
rect 26050 3136 26056 3148
rect 26108 3136 26114 3188
rect 26510 3176 26516 3188
rect 26471 3148 26516 3176
rect 26510 3136 26516 3148
rect 26568 3136 26574 3188
rect 26743 3179 26801 3185
rect 26743 3145 26755 3179
rect 26789 3176 26801 3179
rect 26970 3176 26976 3188
rect 26789 3148 26976 3176
rect 26789 3145 26801 3148
rect 26743 3139 26801 3145
rect 26970 3136 26976 3148
rect 27028 3136 27034 3188
rect 27154 3176 27160 3188
rect 27115 3148 27160 3176
rect 27154 3136 27160 3148
rect 27212 3136 27218 3188
rect 28994 3176 29000 3188
rect 28955 3148 29000 3176
rect 28994 3136 29000 3148
rect 29052 3136 29058 3188
rect 29914 3136 29920 3188
rect 29972 3176 29978 3188
rect 30377 3179 30435 3185
rect 30377 3176 30389 3179
rect 29972 3148 30389 3176
rect 29972 3136 29978 3148
rect 30377 3145 30389 3148
rect 30423 3176 30435 3179
rect 30742 3176 30748 3188
rect 30423 3148 30748 3176
rect 30423 3145 30435 3148
rect 30377 3139 30435 3145
rect 30742 3136 30748 3148
rect 30800 3136 30806 3188
rect 32030 3176 32036 3188
rect 31991 3148 32036 3176
rect 32030 3136 32036 3148
rect 32088 3136 32094 3188
rect 32214 3136 32220 3188
rect 32272 3176 32278 3188
rect 33229 3179 33287 3185
rect 33229 3176 33241 3179
rect 32272 3148 33241 3176
rect 32272 3136 32278 3148
rect 33229 3145 33241 3148
rect 33275 3145 33287 3179
rect 33229 3139 33287 3145
rect 33870 3136 33876 3188
rect 33928 3176 33934 3188
rect 34241 3179 34299 3185
rect 34241 3176 34253 3179
rect 33928 3148 34253 3176
rect 33928 3136 33934 3148
rect 34241 3145 34253 3148
rect 34287 3145 34299 3179
rect 34241 3139 34299 3145
rect 37734 3136 37740 3188
rect 37792 3176 37798 3188
rect 38197 3179 38255 3185
rect 38197 3176 38209 3179
rect 37792 3148 38209 3176
rect 37792 3136 37798 3148
rect 38197 3145 38209 3148
rect 38243 3176 38255 3179
rect 39482 3176 39488 3188
rect 38243 3148 39488 3176
rect 38243 3145 38255 3148
rect 38197 3139 38255 3145
rect 39482 3136 39488 3148
rect 39540 3136 39546 3188
rect 16482 3108 16488 3120
rect 16443 3080 16488 3108
rect 16482 3068 16488 3080
rect 16540 3068 16546 3120
rect 18414 3068 18420 3120
rect 18472 3108 18478 3120
rect 20349 3111 20407 3117
rect 18472 3080 19288 3108
rect 18472 3068 18478 3080
rect 18966 3040 18972 3052
rect 18927 3012 18972 3040
rect 18966 3000 18972 3012
rect 19024 3000 19030 3052
rect 19260 3049 19288 3080
rect 20349 3077 20361 3111
rect 20395 3108 20407 3111
rect 21358 3108 21364 3120
rect 20395 3080 21364 3108
rect 20395 3077 20407 3080
rect 20349 3071 20407 3077
rect 21358 3068 21364 3080
rect 21416 3068 21422 3120
rect 22646 3108 22652 3120
rect 22607 3080 22652 3108
rect 22646 3068 22652 3080
rect 22704 3068 22710 3120
rect 19245 3043 19303 3049
rect 19245 3009 19257 3043
rect 19291 3009 19303 3043
rect 21174 3040 21180 3052
rect 21135 3012 21180 3040
rect 19245 3003 19303 3009
rect 21174 3000 21180 3012
rect 21232 3000 21238 3052
rect 25406 3040 25412 3052
rect 25367 3012 25412 3040
rect 25406 3000 25412 3012
rect 25464 3000 25470 3052
rect 27706 3040 27712 3052
rect 27667 3012 27712 3040
rect 27706 3000 27712 3012
rect 27764 3000 27770 3052
rect 28353 3043 28411 3049
rect 28353 3009 28365 3043
rect 28399 3040 28411 3043
rect 28810 3040 28816 3052
rect 28399 3012 28816 3040
rect 28399 3009 28411 3012
rect 28353 3003 28411 3009
rect 28810 3000 28816 3012
rect 28868 3000 28874 3052
rect 31202 3040 31208 3052
rect 31163 3012 31208 3040
rect 31202 3000 31208 3012
rect 31260 3000 31266 3052
rect 32048 3040 32076 3136
rect 32217 3043 32275 3049
rect 32217 3040 32229 3043
rect 32048 3012 32229 3040
rect 32217 3009 32229 3012
rect 32263 3009 32275 3043
rect 32217 3003 32275 3009
rect 36265 3043 36323 3049
rect 36265 3009 36277 3043
rect 36311 3040 36323 3043
rect 36354 3040 36360 3052
rect 36311 3012 36360 3040
rect 36311 3009 36323 3012
rect 36265 3003 36323 3009
rect 36354 3000 36360 3012
rect 36412 3040 36418 3052
rect 36909 3043 36967 3049
rect 36909 3040 36921 3043
rect 36412 3012 36921 3040
rect 36412 3000 36418 3012
rect 36909 3009 36921 3012
rect 36955 3009 36967 3043
rect 37182 3040 37188 3052
rect 37143 3012 37188 3040
rect 36909 3003 36967 3009
rect 15657 2975 15715 2981
rect 15657 2941 15669 2975
rect 15703 2941 15715 2975
rect 15657 2935 15715 2941
rect 16114 2932 16120 2984
rect 16172 2972 16178 2984
rect 16980 2975 17038 2981
rect 16980 2972 16992 2975
rect 16172 2944 16992 2972
rect 16172 2932 16178 2944
rect 16980 2941 16992 2944
rect 17026 2972 17038 2975
rect 17405 2975 17463 2981
rect 17405 2972 17417 2975
rect 17026 2944 17417 2972
rect 17026 2941 17038 2944
rect 16980 2935 17038 2941
rect 17405 2941 17417 2944
rect 17451 2941 17463 2975
rect 17405 2935 17463 2941
rect 23474 2932 23480 2984
rect 23532 2972 23538 2984
rect 23696 2975 23754 2981
rect 23696 2972 23708 2975
rect 23532 2944 23708 2972
rect 23532 2932 23538 2944
rect 23696 2941 23708 2944
rect 23742 2972 23754 2975
rect 24121 2975 24179 2981
rect 24121 2972 24133 2975
rect 23742 2944 24133 2972
rect 23742 2941 23754 2944
rect 23696 2935 23754 2941
rect 24121 2941 24133 2944
rect 24167 2941 24179 2975
rect 24121 2935 24179 2941
rect 26672 2975 26730 2981
rect 26672 2941 26684 2975
rect 26718 2972 26730 2975
rect 27154 2972 27160 2984
rect 26718 2944 27160 2972
rect 26718 2941 26730 2944
rect 26672 2935 26730 2941
rect 27154 2932 27160 2944
rect 27212 2932 27218 2984
rect 29508 2975 29566 2981
rect 29508 2941 29520 2975
rect 29554 2972 29566 2975
rect 30006 2972 30012 2984
rect 29554 2944 30012 2972
rect 29554 2941 29566 2944
rect 29508 2935 29566 2941
rect 30006 2932 30012 2944
rect 30064 2932 30070 2984
rect 31754 2972 31760 2984
rect 31667 2944 31760 2972
rect 31754 2932 31760 2944
rect 31812 2972 31818 2984
rect 32309 2975 32367 2981
rect 32309 2972 32321 2975
rect 31812 2944 32321 2972
rect 31812 2932 31818 2944
rect 32309 2941 32321 2944
rect 32355 2941 32367 2975
rect 33816 2975 33874 2981
rect 33816 2972 33828 2975
rect 32309 2935 32367 2941
rect 33612 2944 33828 2972
rect 9950 2864 9956 2916
rect 10008 2864 10014 2916
rect 11974 2864 11980 2916
rect 12032 2904 12038 2916
rect 13265 2907 13323 2913
rect 13265 2904 13277 2907
rect 12032 2876 13277 2904
rect 12032 2864 12038 2876
rect 13265 2873 13277 2876
rect 13311 2904 13323 2907
rect 13311 2876 13768 2904
rect 13311 2873 13323 2876
rect 13265 2867 13323 2873
rect 9030 2836 9036 2848
rect 8991 2808 9036 2836
rect 9030 2796 9036 2808
rect 9088 2836 9094 2848
rect 11882 2836 11888 2848
rect 9088 2808 11888 2836
rect 9088 2796 9094 2808
rect 11882 2796 11888 2808
rect 11940 2796 11946 2848
rect 13740 2836 13768 2876
rect 14550 2864 14556 2916
rect 14608 2864 14614 2916
rect 18785 2907 18843 2913
rect 18785 2873 18797 2907
rect 18831 2904 18843 2907
rect 19061 2907 19119 2913
rect 19061 2904 19073 2907
rect 18831 2876 19073 2904
rect 18831 2873 18843 2876
rect 18785 2867 18843 2873
rect 19061 2873 19073 2876
rect 19107 2904 19119 2907
rect 19426 2904 19432 2916
rect 19107 2876 19432 2904
rect 19107 2873 19119 2876
rect 19061 2867 19119 2873
rect 19426 2864 19432 2876
rect 19484 2864 19490 2916
rect 20714 2864 20720 2916
rect 20772 2904 20778 2916
rect 20990 2904 20996 2916
rect 20772 2876 20996 2904
rect 20772 2864 20778 2876
rect 20990 2864 20996 2876
rect 21048 2904 21054 2916
rect 21085 2907 21143 2913
rect 21085 2904 21097 2907
rect 21048 2876 21097 2904
rect 21048 2864 21054 2876
rect 21085 2873 21097 2876
rect 21131 2904 21143 2907
rect 21539 2907 21597 2913
rect 21539 2904 21551 2907
rect 21131 2876 21551 2904
rect 21131 2873 21143 2876
rect 21085 2867 21143 2873
rect 21539 2873 21551 2876
rect 21585 2904 21597 2907
rect 22646 2904 22652 2916
rect 21585 2876 22652 2904
rect 21585 2873 21597 2876
rect 21539 2867 21597 2873
rect 22646 2864 22652 2876
rect 22704 2864 22710 2916
rect 24762 2904 24768 2916
rect 24723 2876 24768 2904
rect 24762 2864 24768 2876
rect 24820 2864 24826 2916
rect 24857 2907 24915 2913
rect 24857 2873 24869 2907
rect 24903 2904 24915 2907
rect 27062 2904 27068 2916
rect 24903 2876 27068 2904
rect 24903 2873 24915 2876
rect 24857 2867 24915 2873
rect 14568 2836 14596 2864
rect 18230 2836 18236 2848
rect 13740 2808 14596 2836
rect 18191 2808 18236 2836
rect 18230 2796 18236 2808
rect 18288 2796 18294 2848
rect 22094 2836 22100 2848
rect 22055 2808 22100 2836
rect 22094 2796 22100 2808
rect 22152 2796 22158 2848
rect 24581 2839 24639 2845
rect 24581 2805 24593 2839
rect 24627 2836 24639 2839
rect 24872 2836 24900 2867
rect 27062 2864 27068 2876
rect 27120 2904 27126 2916
rect 27525 2907 27583 2913
rect 27525 2904 27537 2907
rect 27120 2876 27537 2904
rect 27120 2864 27126 2876
rect 27525 2873 27537 2876
rect 27571 2904 27583 2907
rect 27801 2907 27859 2913
rect 27801 2904 27813 2907
rect 27571 2876 27813 2904
rect 27571 2873 27583 2876
rect 27525 2867 27583 2873
rect 27801 2873 27813 2876
rect 27847 2904 27859 2907
rect 28350 2904 28356 2916
rect 27847 2876 28356 2904
rect 27847 2873 27859 2876
rect 27801 2867 27859 2873
rect 28350 2864 28356 2876
rect 28408 2864 28414 2916
rect 29595 2907 29653 2913
rect 29595 2873 29607 2907
rect 29641 2904 29653 2907
rect 30558 2904 30564 2916
rect 29641 2876 30564 2904
rect 29641 2873 29653 2876
rect 29595 2867 29653 2873
rect 30558 2864 30564 2876
rect 30616 2864 30622 2916
rect 30653 2907 30711 2913
rect 30653 2873 30665 2907
rect 30699 2904 30711 2907
rect 31938 2904 31944 2916
rect 30699 2876 31944 2904
rect 30699 2873 30711 2876
rect 30653 2867 30711 2873
rect 24627 2808 24900 2836
rect 24627 2805 24639 2808
rect 24581 2799 24639 2805
rect 25038 2796 25044 2848
rect 25096 2836 25102 2848
rect 25777 2839 25835 2845
rect 25777 2836 25789 2839
rect 25096 2808 25789 2836
rect 25096 2796 25102 2808
rect 25777 2805 25789 2808
rect 25823 2836 25835 2839
rect 28166 2836 28172 2848
rect 25823 2808 28172 2836
rect 25823 2805 25835 2808
rect 25777 2799 25835 2805
rect 28166 2796 28172 2808
rect 28224 2836 28230 2848
rect 28721 2839 28779 2845
rect 28721 2836 28733 2839
rect 28224 2808 28733 2836
rect 28224 2796 28230 2808
rect 28721 2805 28733 2808
rect 28767 2836 28779 2839
rect 30009 2839 30067 2845
rect 30009 2836 30021 2839
rect 28767 2808 30021 2836
rect 28767 2805 28779 2808
rect 28721 2799 28779 2805
rect 30009 2805 30021 2808
rect 30055 2836 30067 2839
rect 30668 2836 30696 2867
rect 31938 2864 31944 2876
rect 31996 2864 32002 2916
rect 33612 2848 33640 2944
rect 33816 2941 33828 2944
rect 33862 2941 33874 2975
rect 33816 2935 33874 2941
rect 34701 2975 34759 2981
rect 34701 2941 34713 2975
rect 34747 2972 34759 2975
rect 36170 2972 36176 2984
rect 34747 2944 36176 2972
rect 34747 2941 34759 2944
rect 34701 2935 34759 2941
rect 36170 2932 36176 2944
rect 36228 2932 36234 2984
rect 36924 2904 36952 3003
rect 37182 3000 37188 3012
rect 37240 3000 37246 3052
rect 37829 3043 37887 3049
rect 37829 3009 37841 3043
rect 37875 3040 37887 3043
rect 38102 3040 38108 3052
rect 37875 3012 38108 3040
rect 37875 3009 37887 3012
rect 37829 3003 37887 3009
rect 38102 3000 38108 3012
rect 38160 3000 38166 3052
rect 37277 2907 37335 2913
rect 37277 2904 37289 2907
rect 36924 2876 37289 2904
rect 37277 2873 37289 2876
rect 37323 2873 37335 2907
rect 37277 2867 37335 2873
rect 33594 2836 33600 2848
rect 30055 2808 30696 2836
rect 33555 2808 33600 2836
rect 30055 2805 30067 2808
rect 30009 2799 30067 2805
rect 33594 2796 33600 2808
rect 33652 2796 33658 2848
rect 33686 2796 33692 2848
rect 33744 2836 33750 2848
rect 33919 2839 33977 2845
rect 33919 2836 33931 2839
rect 33744 2808 33931 2836
rect 33744 2796 33750 2808
rect 33919 2805 33931 2808
rect 33965 2805 33977 2839
rect 35434 2836 35440 2848
rect 35395 2808 35440 2836
rect 33919 2799 33977 2805
rect 35434 2796 35440 2808
rect 35492 2796 35498 2848
rect 1104 2746 48852 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 48852 2746
rect 1104 2672 48852 2694
rect 9950 2592 9956 2644
rect 10008 2632 10014 2644
rect 11974 2632 11980 2644
rect 10008 2604 11980 2632
rect 10008 2592 10014 2604
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 12434 2632 12440 2644
rect 12395 2604 12440 2632
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 12894 2632 12900 2644
rect 12807 2604 12900 2632
rect 12894 2592 12900 2604
rect 12952 2632 12958 2644
rect 14182 2632 14188 2644
rect 12952 2604 14188 2632
rect 12952 2592 12958 2604
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 14274 2592 14280 2644
rect 14332 2632 14338 2644
rect 15654 2632 15660 2644
rect 14332 2604 14377 2632
rect 15615 2604 15660 2632
rect 14332 2592 14338 2604
rect 15654 2592 15660 2604
rect 15712 2592 15718 2644
rect 16117 2635 16175 2641
rect 16117 2601 16129 2635
rect 16163 2632 16175 2635
rect 16482 2632 16488 2644
rect 16163 2604 16488 2632
rect 16163 2601 16175 2604
rect 16117 2595 16175 2601
rect 16482 2592 16488 2604
rect 16540 2632 16546 2644
rect 16577 2635 16635 2641
rect 16577 2632 16589 2635
rect 16540 2604 16589 2632
rect 16540 2592 16546 2604
rect 16577 2601 16589 2604
rect 16623 2601 16635 2635
rect 16577 2595 16635 2601
rect 17129 2635 17187 2641
rect 17129 2601 17141 2635
rect 17175 2632 17187 2635
rect 18138 2632 18144 2644
rect 17175 2604 18144 2632
rect 17175 2601 17187 2604
rect 17129 2595 17187 2601
rect 10643 2567 10701 2573
rect 10643 2533 10655 2567
rect 10689 2564 10701 2567
rect 16390 2564 16396 2576
rect 10689 2536 16396 2564
rect 10689 2533 10701 2536
rect 10643 2527 10701 2533
rect 16390 2524 16396 2536
rect 16448 2524 16454 2576
rect 16592 2564 16620 2595
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 19426 2632 19432 2644
rect 19387 2604 19432 2632
rect 19426 2592 19432 2604
rect 19484 2592 19490 2644
rect 20990 2632 20996 2644
rect 20951 2604 20996 2632
rect 20990 2592 20996 2604
rect 21048 2632 21054 2644
rect 22281 2635 22339 2641
rect 21048 2604 21725 2632
rect 21048 2592 21054 2604
rect 21697 2573 21725 2604
rect 22281 2601 22293 2635
rect 22327 2632 22339 2635
rect 22830 2632 22836 2644
rect 22327 2604 22836 2632
rect 22327 2601 22339 2604
rect 22281 2595 22339 2601
rect 22830 2592 22836 2604
rect 22888 2592 22894 2644
rect 23290 2592 23296 2644
rect 23348 2632 23354 2644
rect 24397 2635 24455 2641
rect 24397 2632 24409 2635
rect 23348 2604 24409 2632
rect 23348 2592 23354 2604
rect 24397 2601 24409 2604
rect 24443 2632 24455 2635
rect 24443 2604 25084 2632
rect 24443 2601 24455 2604
rect 24397 2595 24455 2601
rect 25056 2573 25084 2604
rect 27706 2592 27712 2644
rect 27764 2632 27770 2644
rect 28583 2635 28641 2641
rect 28583 2632 28595 2635
rect 27764 2604 28595 2632
rect 27764 2592 27770 2604
rect 28583 2601 28595 2604
rect 28629 2601 28641 2635
rect 28583 2595 28641 2601
rect 30558 2592 30564 2644
rect 30616 2632 30622 2644
rect 31113 2635 31171 2641
rect 31113 2632 31125 2635
rect 30616 2604 31125 2632
rect 30616 2592 30622 2604
rect 31113 2601 31125 2604
rect 31159 2601 31171 2635
rect 31113 2595 31171 2601
rect 31619 2635 31677 2641
rect 31619 2601 31631 2635
rect 31665 2632 31677 2635
rect 31754 2632 31760 2644
rect 31665 2604 31760 2632
rect 31665 2601 31677 2604
rect 31619 2595 31677 2601
rect 31754 2592 31760 2604
rect 31812 2592 31818 2644
rect 34333 2635 34391 2641
rect 34333 2632 34345 2635
rect 33428 2604 34345 2632
rect 18049 2567 18107 2573
rect 18049 2564 18061 2567
rect 16592 2536 18061 2564
rect 18049 2533 18061 2536
rect 18095 2564 18107 2567
rect 18830 2567 18888 2573
rect 18830 2564 18842 2567
rect 18095 2536 18842 2564
rect 18095 2533 18107 2536
rect 18049 2527 18107 2533
rect 18830 2533 18842 2536
rect 18876 2533 18888 2567
rect 18830 2527 18888 2533
rect 21682 2567 21740 2573
rect 21682 2533 21694 2567
rect 21728 2533 21740 2567
rect 21682 2527 21740 2533
rect 25041 2567 25099 2573
rect 25041 2533 25053 2567
rect 25087 2533 25099 2567
rect 25041 2527 25099 2533
rect 25130 2524 25136 2576
rect 25188 2564 25194 2576
rect 26697 2567 26755 2573
rect 25188 2536 25233 2564
rect 25188 2524 25194 2536
rect 26697 2533 26709 2567
rect 26743 2564 26755 2567
rect 27062 2564 27068 2576
rect 26743 2536 27068 2564
rect 26743 2533 26755 2536
rect 26697 2527 26755 2533
rect 27062 2524 27068 2536
rect 27120 2524 27126 2576
rect 28258 2564 28264 2576
rect 28219 2536 28264 2564
rect 28258 2524 28264 2536
rect 28316 2524 28322 2576
rect 28350 2524 28356 2576
rect 28408 2564 28414 2576
rect 29549 2567 29607 2573
rect 29549 2564 29561 2567
rect 28408 2536 29561 2564
rect 28408 2524 28414 2536
rect 29549 2533 29561 2536
rect 29595 2564 29607 2567
rect 29914 2564 29920 2576
rect 29595 2536 29920 2564
rect 29595 2533 29607 2536
rect 29549 2527 29607 2533
rect 29914 2524 29920 2536
rect 29972 2524 29978 2576
rect 30650 2524 30656 2576
rect 30708 2564 30714 2576
rect 30745 2567 30803 2573
rect 30745 2564 30757 2567
rect 30708 2536 30757 2564
rect 30708 2524 30714 2536
rect 30745 2533 30757 2536
rect 30791 2533 30803 2567
rect 30745 2527 30803 2533
rect 10556 2499 10614 2505
rect 10556 2465 10568 2499
rect 10602 2496 10614 2499
rect 11054 2496 11060 2508
rect 10602 2468 11060 2496
rect 10602 2465 10614 2468
rect 10556 2459 10614 2465
rect 11054 2456 11060 2468
rect 11112 2456 11118 2508
rect 11422 2456 11428 2508
rect 11480 2496 11486 2508
rect 11552 2499 11610 2505
rect 11552 2496 11564 2499
rect 11480 2468 11564 2496
rect 11480 2456 11486 2468
rect 11552 2465 11564 2468
rect 11598 2465 11610 2499
rect 11552 2459 11610 2465
rect 12710 2456 12716 2508
rect 12768 2496 12774 2508
rect 13722 2496 13728 2508
rect 12768 2468 13728 2496
rect 12768 2456 12774 2468
rect 13722 2456 13728 2468
rect 13780 2496 13786 2508
rect 13817 2499 13875 2505
rect 13817 2496 13829 2499
rect 13780 2468 13829 2496
rect 13780 2456 13786 2468
rect 13817 2465 13829 2468
rect 13863 2465 13875 2499
rect 13817 2459 13875 2465
rect 14420 2499 14478 2505
rect 14420 2465 14432 2499
rect 14466 2496 14478 2499
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 14466 2468 14841 2496
rect 14466 2465 14478 2468
rect 14420 2459 14478 2465
rect 14829 2465 14841 2468
rect 14875 2496 14887 2499
rect 15562 2496 15568 2508
rect 14875 2468 15568 2496
rect 14875 2465 14887 2468
rect 14829 2459 14887 2465
rect 15562 2456 15568 2468
rect 15620 2456 15626 2508
rect 15654 2456 15660 2508
rect 15712 2496 15718 2508
rect 16209 2499 16267 2505
rect 16209 2496 16221 2499
rect 15712 2468 16221 2496
rect 15712 2456 15718 2468
rect 16209 2465 16221 2468
rect 16255 2465 16267 2499
rect 16209 2459 16267 2465
rect 17773 2499 17831 2505
rect 17773 2465 17785 2499
rect 17819 2496 17831 2499
rect 18506 2496 18512 2508
rect 17819 2468 18512 2496
rect 17819 2465 17831 2468
rect 17773 2459 17831 2465
rect 18506 2456 18512 2468
rect 18564 2456 18570 2508
rect 20625 2499 20683 2505
rect 20625 2465 20637 2499
rect 20671 2496 20683 2499
rect 21361 2499 21419 2505
rect 21361 2496 21373 2499
rect 20671 2468 21373 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 21361 2465 21373 2468
rect 21407 2496 21419 2499
rect 21450 2496 21456 2508
rect 21407 2468 21456 2496
rect 21407 2465 21419 2468
rect 21361 2459 21419 2465
rect 21450 2456 21456 2468
rect 21508 2456 21514 2508
rect 28276 2496 28304 2524
rect 31570 2505 31576 2508
rect 28480 2499 28538 2505
rect 28480 2496 28492 2499
rect 28276 2468 28492 2496
rect 28480 2465 28492 2468
rect 28526 2465 28538 2499
rect 31548 2499 31576 2505
rect 31548 2496 31560 2499
rect 31483 2468 31560 2496
rect 28480 2459 28538 2465
rect 31548 2465 31560 2468
rect 31628 2496 31634 2508
rect 31941 2499 31999 2505
rect 31941 2496 31953 2499
rect 31628 2468 31953 2496
rect 31548 2459 31576 2465
rect 31570 2456 31576 2459
rect 31628 2456 31634 2468
rect 31941 2465 31953 2468
rect 31987 2465 31999 2499
rect 31941 2459 31999 2465
rect 32401 2499 32459 2505
rect 32401 2465 32413 2499
rect 32447 2496 32459 2499
rect 33229 2499 33287 2505
rect 33229 2496 33241 2499
rect 32447 2468 33241 2496
rect 32447 2465 32459 2468
rect 32401 2459 32459 2465
rect 33229 2465 33241 2468
rect 33275 2496 33287 2499
rect 33428 2496 33456 2604
rect 34333 2601 34345 2604
rect 34379 2601 34391 2635
rect 35250 2632 35256 2644
rect 35211 2604 35256 2632
rect 34333 2595 34391 2601
rect 35250 2592 35256 2604
rect 35308 2592 35314 2644
rect 35434 2592 35440 2644
rect 35492 2632 35498 2644
rect 37139 2635 37197 2641
rect 37139 2632 37151 2635
rect 35492 2604 37151 2632
rect 35492 2592 35498 2604
rect 37139 2601 37151 2604
rect 37185 2601 37197 2635
rect 37139 2595 37197 2601
rect 37553 2635 37611 2641
rect 37553 2601 37565 2635
rect 37599 2632 37611 2635
rect 37734 2632 37740 2644
rect 37599 2604 37740 2632
rect 37599 2601 37611 2604
rect 37553 2595 37611 2601
rect 33778 2564 33784 2576
rect 33739 2536 33784 2564
rect 33778 2524 33784 2536
rect 33836 2524 33842 2576
rect 35268 2564 35296 2592
rect 35621 2567 35679 2573
rect 35621 2564 35633 2567
rect 35268 2536 35633 2564
rect 35621 2533 35633 2536
rect 35667 2533 35679 2567
rect 35621 2527 35679 2533
rect 36173 2567 36231 2573
rect 36173 2533 36185 2567
rect 36219 2564 36231 2567
rect 36814 2564 36820 2576
rect 36219 2536 36820 2564
rect 36219 2533 36231 2536
rect 36173 2527 36231 2533
rect 36814 2524 36820 2536
rect 36872 2524 36878 2576
rect 33275 2468 33456 2496
rect 34149 2499 34207 2505
rect 33275 2465 33287 2468
rect 33229 2459 33287 2465
rect 34149 2465 34161 2499
rect 34195 2496 34207 2499
rect 34609 2499 34667 2505
rect 34609 2496 34621 2499
rect 34195 2468 34621 2496
rect 34195 2465 34207 2468
rect 34149 2459 34207 2465
rect 34609 2465 34621 2468
rect 34655 2465 34667 2499
rect 34609 2459 34667 2465
rect 37068 2499 37126 2505
rect 37068 2465 37080 2499
rect 37114 2496 37126 2499
rect 37568 2496 37596 2595
rect 37734 2592 37740 2604
rect 37792 2592 37798 2644
rect 37114 2468 37596 2496
rect 37114 2465 37126 2468
rect 37068 2459 37126 2465
rect 13357 2431 13415 2437
rect 13357 2397 13369 2431
rect 13403 2428 13415 2431
rect 14507 2431 14565 2437
rect 13403 2400 13814 2428
rect 13403 2397 13415 2400
rect 13357 2391 13415 2397
rect 13786 2360 13814 2400
rect 14507 2397 14519 2431
rect 14553 2428 14565 2431
rect 16666 2428 16672 2440
rect 14553 2400 16672 2428
rect 14553 2397 14565 2400
rect 14507 2391 14565 2397
rect 16666 2388 16672 2400
rect 16724 2388 16730 2440
rect 24857 2431 24915 2437
rect 24857 2397 24869 2431
rect 24903 2428 24915 2431
rect 25130 2428 25136 2440
rect 24903 2400 25136 2428
rect 24903 2397 24915 2400
rect 24857 2391 24915 2397
rect 25130 2388 25136 2400
rect 25188 2388 25194 2440
rect 25406 2428 25412 2440
rect 25367 2400 25412 2428
rect 25406 2388 25412 2400
rect 25464 2388 25470 2440
rect 26234 2388 26240 2440
rect 26292 2428 26298 2440
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26292 2400 26985 2428
rect 26292 2388 26298 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 27249 2431 27307 2437
rect 27249 2428 27261 2431
rect 26973 2391 27031 2397
rect 27080 2400 27261 2428
rect 18230 2360 18236 2372
rect 13786 2332 18236 2360
rect 18230 2320 18236 2332
rect 18288 2320 18294 2372
rect 25590 2320 25596 2372
rect 25648 2360 25654 2372
rect 27080 2360 27108 2400
rect 27249 2397 27261 2400
rect 27295 2397 27307 2431
rect 27249 2391 27307 2397
rect 29825 2431 29883 2437
rect 29825 2397 29837 2431
rect 29871 2397 29883 2431
rect 30098 2428 30104 2440
rect 30059 2400 30104 2428
rect 29825 2391 29883 2397
rect 25648 2332 27108 2360
rect 25648 2320 25654 2332
rect 28442 2320 28448 2372
rect 28500 2360 28506 2372
rect 29089 2363 29147 2369
rect 29089 2360 29101 2363
rect 28500 2332 29101 2360
rect 28500 2320 28506 2332
rect 29089 2329 29101 2332
rect 29135 2360 29147 2363
rect 29840 2360 29868 2391
rect 30098 2388 30104 2400
rect 30156 2388 30162 2440
rect 31956 2428 31984 2459
rect 33318 2428 33324 2440
rect 31956 2400 33134 2428
rect 33279 2400 33324 2428
rect 29135 2332 29868 2360
rect 33106 2360 33134 2400
rect 33318 2388 33324 2400
rect 33376 2388 33382 2440
rect 34164 2360 34192 2459
rect 34330 2388 34336 2440
rect 34388 2428 34394 2440
rect 35529 2431 35587 2437
rect 35529 2428 35541 2431
rect 34388 2400 35541 2428
rect 34388 2388 34394 2400
rect 35529 2397 35541 2400
rect 35575 2428 35587 2431
rect 36449 2431 36507 2437
rect 36449 2428 36461 2431
rect 35575 2400 36461 2428
rect 35575 2397 35587 2400
rect 35529 2391 35587 2397
rect 36449 2397 36461 2400
rect 36495 2397 36507 2431
rect 36449 2391 36507 2397
rect 33106 2332 34192 2360
rect 29135 2329 29147 2332
rect 29089 2323 29147 2329
rect 5626 2252 5632 2304
rect 5684 2292 5690 2304
rect 9217 2295 9275 2301
rect 9217 2292 9229 2295
rect 5684 2264 9229 2292
rect 5684 2252 5690 2264
rect 9217 2261 9229 2264
rect 9263 2292 9275 2295
rect 10870 2292 10876 2304
rect 9263 2264 10876 2292
rect 9263 2261 9275 2264
rect 9217 2255 9275 2261
rect 10870 2252 10876 2264
rect 10928 2252 10934 2304
rect 11054 2292 11060 2304
rect 11015 2264 11060 2292
rect 11054 2252 11060 2264
rect 11112 2252 11118 2304
rect 11422 2292 11428 2304
rect 11383 2264 11428 2292
rect 11422 2252 11428 2264
rect 11480 2252 11486 2304
rect 11655 2295 11713 2301
rect 11655 2261 11667 2295
rect 11701 2292 11713 2295
rect 11882 2292 11888 2304
rect 11701 2264 11888 2292
rect 11701 2261 11713 2264
rect 11655 2255 11713 2261
rect 11882 2252 11888 2264
rect 11940 2252 11946 2304
rect 26234 2292 26240 2304
rect 26195 2264 26240 2292
rect 26234 2252 26240 2264
rect 26292 2252 26298 2304
rect 1104 2202 48852 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 48852 2202
rect 1104 2128 48852 2150
rect 33226 76 33232 128
rect 33284 116 33290 128
rect 33870 116 33876 128
rect 33284 88 33876 116
rect 33284 76 33290 88
rect 33870 76 33876 88
rect 33928 76 33934 128
rect 40034 76 40040 128
rect 40092 116 40098 128
rect 40954 116 40960 128
rect 40092 88 40960 116
rect 40092 76 40098 88
rect 40954 76 40960 88
rect 41012 76 41018 128
rect 41322 76 41328 128
rect 41380 116 41386 128
rect 48130 116 48136 128
rect 41380 88 48136 116
rect 41380 76 41386 88
rect 48130 76 48136 88
rect 48188 76 48194 128
<< via1 >>
rect 13820 49512 13872 49564
rect 16120 49512 16172 49564
rect 19432 49512 19484 49564
rect 20260 49512 20312 49564
rect 24216 49512 24268 49564
rect 24952 49512 25004 49564
rect 19606 47302 19658 47354
rect 19670 47302 19722 47354
rect 19734 47302 19786 47354
rect 19798 47302 19850 47354
rect 4246 46758 4298 46810
rect 4310 46758 4362 46810
rect 4374 46758 4426 46810
rect 4438 46758 4490 46810
rect 34966 46758 35018 46810
rect 35030 46758 35082 46810
rect 35094 46758 35146 46810
rect 35158 46758 35210 46810
rect 19606 46214 19658 46266
rect 19670 46214 19722 46266
rect 19734 46214 19786 46266
rect 19798 46214 19850 46266
rect 4246 45670 4298 45722
rect 4310 45670 4362 45722
rect 4374 45670 4426 45722
rect 4438 45670 4490 45722
rect 34966 45670 35018 45722
rect 35030 45670 35082 45722
rect 35094 45670 35146 45722
rect 35158 45670 35210 45722
rect 19606 45126 19658 45178
rect 19670 45126 19722 45178
rect 19734 45126 19786 45178
rect 19798 45126 19850 45178
rect 4246 44582 4298 44634
rect 4310 44582 4362 44634
rect 4374 44582 4426 44634
rect 4438 44582 4490 44634
rect 34966 44582 35018 44634
rect 35030 44582 35082 44634
rect 35094 44582 35146 44634
rect 35158 44582 35210 44634
rect 19606 44038 19658 44090
rect 19670 44038 19722 44090
rect 19734 44038 19786 44090
rect 19798 44038 19850 44090
rect 4246 43494 4298 43546
rect 4310 43494 4362 43546
rect 4374 43494 4426 43546
rect 4438 43494 4490 43546
rect 34966 43494 35018 43546
rect 35030 43494 35082 43546
rect 35094 43494 35146 43546
rect 35158 43494 35210 43546
rect 19606 42950 19658 43002
rect 19670 42950 19722 43002
rect 19734 42950 19786 43002
rect 19798 42950 19850 43002
rect 21824 42712 21876 42764
rect 21640 42508 21692 42560
rect 4246 42406 4298 42458
rect 4310 42406 4362 42458
rect 4374 42406 4426 42458
rect 4438 42406 4490 42458
rect 34966 42406 35018 42458
rect 35030 42406 35082 42458
rect 35094 42406 35146 42458
rect 35158 42406 35210 42458
rect 14188 42100 14240 42152
rect 24308 42100 24360 42152
rect 24860 42143 24912 42152
rect 24860 42109 24869 42143
rect 24869 42109 24903 42143
rect 24903 42109 24912 42143
rect 24860 42100 24912 42109
rect 21732 41964 21784 42016
rect 21824 42007 21876 42016
rect 21824 41973 21833 42007
rect 21833 41973 21867 42007
rect 21867 41973 21876 42007
rect 21824 41964 21876 41973
rect 24768 41964 24820 42016
rect 24860 41964 24912 42016
rect 30380 41964 30432 42016
rect 19606 41862 19658 41914
rect 19670 41862 19722 41914
rect 19734 41862 19786 41914
rect 19798 41862 19850 41914
rect 24768 41760 24820 41812
rect 21916 41692 21968 41744
rect 17500 41624 17552 41676
rect 19064 41624 19116 41676
rect 24216 41667 24268 41676
rect 24216 41633 24225 41667
rect 24225 41633 24259 41667
rect 24259 41633 24268 41667
rect 24216 41624 24268 41633
rect 25964 41624 26016 41676
rect 21640 41599 21692 41608
rect 21640 41565 21649 41599
rect 21649 41565 21683 41599
rect 21683 41565 21692 41599
rect 21640 41556 21692 41565
rect 22284 41599 22336 41608
rect 22284 41565 22293 41599
rect 22293 41565 22327 41599
rect 22327 41565 22336 41599
rect 22284 41556 22336 41565
rect 30196 41624 30248 41676
rect 32128 41624 32180 41676
rect 23204 41488 23256 41540
rect 27436 41556 27488 41608
rect 16488 41463 16540 41472
rect 16488 41429 16497 41463
rect 16497 41429 16531 41463
rect 16531 41429 16540 41463
rect 16488 41420 16540 41429
rect 16580 41420 16632 41472
rect 19156 41420 19208 41472
rect 19432 41463 19484 41472
rect 19432 41429 19441 41463
rect 19441 41429 19475 41463
rect 19475 41429 19484 41463
rect 19432 41420 19484 41429
rect 19708 41463 19760 41472
rect 19708 41429 19717 41463
rect 19717 41429 19751 41463
rect 19751 41429 19760 41463
rect 19708 41420 19760 41429
rect 24584 41420 24636 41472
rect 24952 41420 25004 41472
rect 26884 41420 26936 41472
rect 30104 41420 30156 41472
rect 32772 41420 32824 41472
rect 4246 41318 4298 41370
rect 4310 41318 4362 41370
rect 4374 41318 4426 41370
rect 4438 41318 4490 41370
rect 34966 41318 35018 41370
rect 35030 41318 35082 41370
rect 35094 41318 35146 41370
rect 35158 41318 35210 41370
rect 19064 41259 19116 41268
rect 19064 41225 19073 41259
rect 19073 41225 19107 41259
rect 19107 41225 19116 41259
rect 19064 41216 19116 41225
rect 21640 41216 21692 41268
rect 27436 41259 27488 41268
rect 27436 41225 27445 41259
rect 27445 41225 27479 41259
rect 27479 41225 27488 41259
rect 27436 41216 27488 41225
rect 19892 41191 19944 41200
rect 19892 41157 19901 41191
rect 19901 41157 19935 41191
rect 19935 41157 19944 41191
rect 19892 41148 19944 41157
rect 22284 41148 22336 41200
rect 24308 41148 24360 41200
rect 30932 41148 30984 41200
rect 32128 41148 32180 41200
rect 14556 41080 14608 41132
rect 16488 41080 16540 41132
rect 14280 41012 14332 41064
rect 19708 41080 19760 41132
rect 24768 41080 24820 41132
rect 27252 41080 27304 41132
rect 17500 41055 17552 41064
rect 17500 41021 17509 41055
rect 17509 41021 17543 41055
rect 17543 41021 17552 41055
rect 17500 41012 17552 41021
rect 18604 41012 18656 41064
rect 18788 41012 18840 41064
rect 18420 40944 18472 40996
rect 19432 40987 19484 40996
rect 19432 40953 19441 40987
rect 19441 40953 19475 40987
rect 19475 40953 19484 40987
rect 19432 40944 19484 40953
rect 21916 40944 21968 40996
rect 22100 40944 22152 40996
rect 14372 40876 14424 40928
rect 16488 40919 16540 40928
rect 16488 40885 16497 40919
rect 16497 40885 16531 40919
rect 16531 40885 16540 40919
rect 16488 40876 16540 40885
rect 18788 40919 18840 40928
rect 18788 40885 18797 40919
rect 18797 40885 18831 40919
rect 18831 40885 18840 40919
rect 18788 40876 18840 40885
rect 23020 40876 23072 40928
rect 30380 41012 30432 41064
rect 35532 41080 35584 41132
rect 25044 40987 25096 40996
rect 25044 40953 25053 40987
rect 25053 40953 25087 40987
rect 25087 40953 25096 40987
rect 25044 40944 25096 40953
rect 25964 40987 26016 40996
rect 25964 40953 25973 40987
rect 25973 40953 26007 40987
rect 26007 40953 26016 40987
rect 31668 40987 31720 40996
rect 25964 40944 26016 40953
rect 31668 40953 31677 40987
rect 31677 40953 31711 40987
rect 31711 40953 31720 40987
rect 31668 40944 31720 40953
rect 32864 41012 32916 41064
rect 33048 40987 33100 40996
rect 33048 40953 33057 40987
rect 33057 40953 33091 40987
rect 33091 40953 33100 40987
rect 33048 40944 33100 40953
rect 24308 40919 24360 40928
rect 24308 40885 24317 40919
rect 24317 40885 24351 40919
rect 24351 40885 24360 40919
rect 24308 40876 24360 40885
rect 26976 40876 27028 40928
rect 29920 40919 29972 40928
rect 29920 40885 29929 40919
rect 29929 40885 29963 40919
rect 29963 40885 29972 40919
rect 29920 40876 29972 40885
rect 30196 40919 30248 40928
rect 30196 40885 30205 40919
rect 30205 40885 30239 40919
rect 30239 40885 30248 40919
rect 30196 40876 30248 40885
rect 31484 40876 31536 40928
rect 32588 40876 32640 40928
rect 33784 40876 33836 40928
rect 19606 40774 19658 40826
rect 19670 40774 19722 40826
rect 19734 40774 19786 40826
rect 19798 40774 19850 40826
rect 24584 40715 24636 40724
rect 24584 40681 24593 40715
rect 24593 40681 24627 40715
rect 24627 40681 24636 40715
rect 24584 40672 24636 40681
rect 26884 40672 26936 40724
rect 16764 40604 16816 40656
rect 19432 40647 19484 40656
rect 19432 40613 19441 40647
rect 19441 40613 19475 40647
rect 19475 40613 19484 40647
rect 19432 40604 19484 40613
rect 21732 40647 21784 40656
rect 21732 40613 21741 40647
rect 21741 40613 21775 40647
rect 21775 40613 21784 40647
rect 21732 40604 21784 40613
rect 22008 40604 22060 40656
rect 25044 40647 25096 40656
rect 25044 40613 25053 40647
rect 25053 40613 25087 40647
rect 25087 40613 25096 40647
rect 25044 40604 25096 40613
rect 27068 40647 27120 40656
rect 27068 40613 27077 40647
rect 27077 40613 27111 40647
rect 27111 40613 27120 40647
rect 30196 40647 30248 40656
rect 27068 40604 27120 40613
rect 30196 40613 30205 40647
rect 30205 40613 30239 40647
rect 30239 40613 30248 40647
rect 30196 40604 30248 40613
rect 32680 40604 32732 40656
rect 17868 40536 17920 40588
rect 19064 40536 19116 40588
rect 23204 40579 23256 40588
rect 23204 40545 23213 40579
rect 23213 40545 23247 40579
rect 23247 40545 23256 40579
rect 23204 40536 23256 40545
rect 33968 40579 34020 40588
rect 33968 40545 33977 40579
rect 33977 40545 34011 40579
rect 34011 40545 34020 40579
rect 33968 40536 34020 40545
rect 35256 40536 35308 40588
rect 38292 40579 38344 40588
rect 38292 40545 38301 40579
rect 38301 40545 38335 40579
rect 38335 40545 38344 40579
rect 38292 40536 38344 40545
rect 14188 40468 14240 40520
rect 14648 40375 14700 40384
rect 14648 40341 14657 40375
rect 14657 40341 14691 40375
rect 14691 40341 14700 40375
rect 14648 40332 14700 40341
rect 16212 40332 16264 40384
rect 17224 40511 17276 40520
rect 17224 40477 17233 40511
rect 17233 40477 17267 40511
rect 17267 40477 17276 40511
rect 17224 40468 17276 40477
rect 19156 40468 19208 40520
rect 20536 40468 20588 40520
rect 22100 40468 22152 40520
rect 24952 40511 25004 40520
rect 24952 40477 24961 40511
rect 24961 40477 24995 40511
rect 24995 40477 25004 40511
rect 24952 40468 25004 40477
rect 26148 40468 26200 40520
rect 24308 40400 24360 40452
rect 29092 40468 29144 40520
rect 29920 40468 29972 40520
rect 31024 40468 31076 40520
rect 32496 40511 32548 40520
rect 32496 40477 32505 40511
rect 32505 40477 32539 40511
rect 32539 40477 32548 40511
rect 32496 40468 32548 40477
rect 32404 40400 32456 40452
rect 38752 40468 38804 40520
rect 33232 40400 33284 40452
rect 16672 40332 16724 40384
rect 22744 40332 22796 40384
rect 29920 40332 29972 40384
rect 32956 40332 33008 40384
rect 37464 40332 37516 40384
rect 38568 40332 38620 40384
rect 38844 40375 38896 40384
rect 38844 40341 38853 40375
rect 38853 40341 38887 40375
rect 38887 40341 38896 40375
rect 38844 40332 38896 40341
rect 4246 40230 4298 40282
rect 4310 40230 4362 40282
rect 4374 40230 4426 40282
rect 4438 40230 4490 40282
rect 34966 40230 35018 40282
rect 35030 40230 35082 40282
rect 35094 40230 35146 40282
rect 35158 40230 35210 40282
rect 14188 40171 14240 40180
rect 14188 40137 14197 40171
rect 14197 40137 14231 40171
rect 14231 40137 14240 40171
rect 14188 40128 14240 40137
rect 17868 40171 17920 40180
rect 17868 40137 17877 40171
rect 17877 40137 17911 40171
rect 17911 40137 17920 40171
rect 17868 40128 17920 40137
rect 19432 40128 19484 40180
rect 21732 40128 21784 40180
rect 22744 40171 22796 40180
rect 22744 40137 22753 40171
rect 22753 40137 22787 40171
rect 22787 40137 22796 40171
rect 22744 40128 22796 40137
rect 25044 40128 25096 40180
rect 26884 40128 26936 40180
rect 31024 40171 31076 40180
rect 31024 40137 31033 40171
rect 31033 40137 31067 40171
rect 31067 40137 31076 40171
rect 31024 40128 31076 40137
rect 33048 40128 33100 40180
rect 16028 40060 16080 40112
rect 22284 40103 22336 40112
rect 22284 40069 22293 40103
rect 22293 40069 22327 40103
rect 22327 40069 22336 40103
rect 22284 40060 22336 40069
rect 13360 40035 13412 40044
rect 13360 40001 13369 40035
rect 13369 40001 13403 40035
rect 13403 40001 13412 40035
rect 13360 39992 13412 40001
rect 14648 40035 14700 40044
rect 14648 40001 14657 40035
rect 14657 40001 14691 40035
rect 14691 40001 14700 40035
rect 14648 39992 14700 40001
rect 16580 39992 16632 40044
rect 24584 40060 24636 40112
rect 23204 40035 23256 40044
rect 23204 40001 23213 40035
rect 23213 40001 23247 40035
rect 23247 40001 23256 40035
rect 23204 39992 23256 40001
rect 27804 40060 27856 40112
rect 32220 40060 32272 40112
rect 33968 40103 34020 40112
rect 33968 40069 33977 40103
rect 33977 40069 34011 40103
rect 34011 40069 34020 40103
rect 33968 40060 34020 40069
rect 35256 40128 35308 40180
rect 39672 40128 39724 40180
rect 38292 40103 38344 40112
rect 38292 40069 38301 40103
rect 38301 40069 38335 40103
rect 38335 40069 38344 40103
rect 38292 40060 38344 40069
rect 39212 40060 39264 40112
rect 26976 40035 27028 40044
rect 26976 40001 26985 40035
rect 26985 40001 27019 40035
rect 27019 40001 27028 40035
rect 26976 39992 27028 40001
rect 27252 40035 27304 40044
rect 27252 40001 27261 40035
rect 27261 40001 27295 40035
rect 27295 40001 27304 40035
rect 27252 39992 27304 40001
rect 30104 40035 30156 40044
rect 30104 40001 30113 40035
rect 30113 40001 30147 40035
rect 30147 40001 30156 40035
rect 30104 39992 30156 40001
rect 32588 40035 32640 40044
rect 32588 40001 32597 40035
rect 32597 40001 32631 40035
rect 32631 40001 32640 40035
rect 32588 39992 32640 40001
rect 12992 39967 13044 39976
rect 12992 39933 13010 39967
rect 13010 39933 13044 39967
rect 12992 39924 13044 39933
rect 14740 39899 14792 39908
rect 14740 39865 14749 39899
rect 14749 39865 14783 39899
rect 14783 39865 14792 39899
rect 14740 39856 14792 39865
rect 15292 39899 15344 39908
rect 15292 39865 15301 39899
rect 15301 39865 15335 39899
rect 15335 39865 15344 39899
rect 15292 39856 15344 39865
rect 16764 39856 16816 39908
rect 13176 39788 13228 39840
rect 16396 39788 16448 39840
rect 17500 39856 17552 39908
rect 35532 39924 35584 39976
rect 37464 39967 37516 39976
rect 19432 39899 19484 39908
rect 19432 39865 19441 39899
rect 19441 39865 19475 39899
rect 19475 39865 19484 39899
rect 19432 39856 19484 39865
rect 19984 39899 20036 39908
rect 19984 39865 19993 39899
rect 19993 39865 20027 39899
rect 20027 39865 20036 39899
rect 19984 39856 20036 39865
rect 18788 39831 18840 39840
rect 18788 39797 18797 39831
rect 18797 39797 18831 39831
rect 18831 39797 18840 39831
rect 18788 39788 18840 39797
rect 25044 39856 25096 39908
rect 27068 39899 27120 39908
rect 27068 39865 27088 39899
rect 27088 39865 27120 39899
rect 27068 39856 27120 39865
rect 30196 39899 30248 39908
rect 30196 39865 30205 39899
rect 30205 39865 30239 39899
rect 30239 39865 30248 39899
rect 30196 39856 30248 39865
rect 22008 39788 22060 39840
rect 24952 39788 25004 39840
rect 29092 39831 29144 39840
rect 29092 39797 29101 39831
rect 29101 39797 29135 39831
rect 29135 39797 29144 39831
rect 29092 39788 29144 39797
rect 30012 39788 30064 39840
rect 31760 39788 31812 39840
rect 32588 39856 32640 39908
rect 35716 39856 35768 39908
rect 37464 39933 37473 39967
rect 37473 39933 37507 39967
rect 37507 39933 37516 39967
rect 37464 39924 37516 39933
rect 37740 39899 37792 39908
rect 37740 39865 37749 39899
rect 37749 39865 37783 39899
rect 37783 39865 37792 39899
rect 37740 39856 37792 39865
rect 38752 39899 38804 39908
rect 38752 39865 38761 39899
rect 38761 39865 38795 39899
rect 38795 39865 38804 39899
rect 38752 39856 38804 39865
rect 38844 39899 38896 39908
rect 38844 39865 38853 39899
rect 38853 39865 38887 39899
rect 38887 39865 38896 39899
rect 38844 39856 38896 39865
rect 42156 39856 42208 39908
rect 33140 39788 33192 39840
rect 36084 39788 36136 39840
rect 19606 39686 19658 39738
rect 19670 39686 19722 39738
rect 19734 39686 19786 39738
rect 19798 39686 19850 39738
rect 13176 39516 13228 39568
rect 14740 39584 14792 39636
rect 16212 39584 16264 39636
rect 16488 39584 16540 39636
rect 19432 39627 19484 39636
rect 19432 39593 19441 39627
rect 19441 39593 19475 39627
rect 19475 39593 19484 39627
rect 19432 39584 19484 39593
rect 24308 39627 24360 39636
rect 24308 39593 24317 39627
rect 24317 39593 24351 39627
rect 24351 39593 24360 39627
rect 24308 39584 24360 39593
rect 25044 39584 25096 39636
rect 30104 39584 30156 39636
rect 32496 39627 32548 39636
rect 32496 39593 32505 39627
rect 32505 39593 32539 39627
rect 32539 39593 32548 39627
rect 32496 39584 32548 39593
rect 36084 39584 36136 39636
rect 14004 39559 14056 39568
rect 14004 39525 14013 39559
rect 14013 39525 14047 39559
rect 14047 39525 14056 39559
rect 14004 39516 14056 39525
rect 16028 39516 16080 39568
rect 16396 39516 16448 39568
rect 16672 39559 16724 39568
rect 16672 39525 16681 39559
rect 16681 39525 16715 39559
rect 16715 39525 16724 39559
rect 16672 39516 16724 39525
rect 16764 39559 16816 39568
rect 16764 39525 16773 39559
rect 16773 39525 16807 39559
rect 16807 39525 16816 39559
rect 16764 39516 16816 39525
rect 18696 39516 18748 39568
rect 19156 39516 19208 39568
rect 22008 39516 22060 39568
rect 27068 39559 27120 39568
rect 27068 39525 27077 39559
rect 27077 39525 27111 39559
rect 27111 39525 27120 39559
rect 27068 39516 27120 39525
rect 29000 39516 29052 39568
rect 32680 39516 32732 39568
rect 36452 39516 36504 39568
rect 38568 39516 38620 39568
rect 38844 39559 38896 39568
rect 38844 39525 38853 39559
rect 38853 39525 38887 39559
rect 38887 39525 38896 39559
rect 38844 39516 38896 39525
rect 11888 39448 11940 39500
rect 15660 39491 15712 39500
rect 15660 39457 15678 39491
rect 15678 39457 15712 39491
rect 15660 39448 15712 39457
rect 30932 39448 30984 39500
rect 34428 39448 34480 39500
rect 40776 39448 40828 39500
rect 15292 39380 15344 39432
rect 15936 39380 15988 39432
rect 18512 39423 18564 39432
rect 18512 39389 18521 39423
rect 18521 39389 18555 39423
rect 18555 39389 18564 39423
rect 18512 39380 18564 39389
rect 21824 39423 21876 39432
rect 21824 39389 21833 39423
rect 21833 39389 21867 39423
rect 21867 39389 21876 39423
rect 21824 39380 21876 39389
rect 23940 39423 23992 39432
rect 19432 39312 19484 39364
rect 19984 39312 20036 39364
rect 23940 39389 23949 39423
rect 23949 39389 23983 39423
rect 23983 39389 23992 39423
rect 23940 39380 23992 39389
rect 26976 39423 27028 39432
rect 26976 39389 26985 39423
rect 26985 39389 27019 39423
rect 27019 39389 27028 39423
rect 26976 39380 27028 39389
rect 27804 39380 27856 39432
rect 29184 39423 29236 39432
rect 29184 39389 29193 39423
rect 29193 39389 29227 39423
rect 29227 39389 29236 39423
rect 29184 39380 29236 39389
rect 32864 39423 32916 39432
rect 32864 39389 32873 39423
rect 32873 39389 32907 39423
rect 32907 39389 32916 39423
rect 32864 39380 32916 39389
rect 36820 39423 36872 39432
rect 22284 39312 22336 39364
rect 32404 39312 32456 39364
rect 36820 39389 36829 39423
rect 36829 39389 36863 39423
rect 36863 39389 36872 39423
rect 36820 39380 36872 39389
rect 41420 39380 41472 39432
rect 13268 39244 13320 39296
rect 23756 39287 23808 39296
rect 23756 39253 23765 39287
rect 23765 39253 23799 39287
rect 23799 39253 23808 39287
rect 23756 39244 23808 39253
rect 25228 39287 25280 39296
rect 25228 39253 25237 39287
rect 25237 39253 25271 39287
rect 25271 39253 25280 39287
rect 25228 39244 25280 39253
rect 30104 39287 30156 39296
rect 30104 39253 30113 39287
rect 30113 39253 30147 39287
rect 30147 39253 30156 39287
rect 30104 39244 30156 39253
rect 30748 39244 30800 39296
rect 33048 39244 33100 39296
rect 40960 39244 41012 39296
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 34966 39142 35018 39194
rect 35030 39142 35082 39194
rect 35094 39142 35146 39194
rect 35158 39142 35210 39194
rect 13176 39040 13228 39092
rect 14740 39040 14792 39092
rect 15660 39083 15712 39092
rect 15660 39049 15669 39083
rect 15669 39049 15703 39083
rect 15703 39049 15712 39083
rect 15660 39040 15712 39049
rect 16764 39040 16816 39092
rect 18696 39040 18748 39092
rect 10508 38836 10560 38888
rect 13728 38904 13780 38956
rect 14372 38904 14424 38956
rect 16488 38904 16540 38956
rect 11336 38879 11388 38888
rect 11336 38845 11345 38879
rect 11345 38845 11379 38879
rect 11379 38845 11388 38879
rect 11336 38836 11388 38845
rect 12624 38836 12676 38888
rect 15384 38836 15436 38888
rect 17224 38836 17276 38888
rect 21824 39040 21876 39092
rect 26976 39040 27028 39092
rect 29000 39040 29052 39092
rect 30656 39083 30708 39092
rect 30656 39049 30665 39083
rect 30665 39049 30699 39083
rect 30699 39049 30708 39083
rect 30656 39040 30708 39049
rect 32864 39040 32916 39092
rect 35624 39083 35676 39092
rect 35624 39049 35633 39083
rect 35633 39049 35667 39083
rect 35667 39049 35676 39083
rect 35624 39040 35676 39049
rect 38568 39040 38620 39092
rect 41512 39040 41564 39092
rect 11704 38768 11756 38820
rect 11888 38743 11940 38752
rect 11888 38709 11897 38743
rect 11897 38709 11931 38743
rect 11931 38709 11940 38743
rect 11888 38700 11940 38709
rect 13452 38700 13504 38752
rect 14740 38811 14792 38820
rect 14740 38777 14749 38811
rect 14749 38777 14783 38811
rect 14783 38777 14792 38811
rect 14740 38768 14792 38777
rect 18696 38768 18748 38820
rect 17868 38743 17920 38752
rect 17868 38709 17877 38743
rect 17877 38709 17911 38743
rect 17911 38709 17920 38743
rect 17868 38700 17920 38709
rect 19248 38836 19300 38888
rect 20444 38879 20496 38888
rect 20444 38845 20453 38879
rect 20453 38845 20487 38879
rect 20487 38845 20496 38879
rect 20444 38836 20496 38845
rect 24308 38904 24360 38956
rect 24768 38904 24820 38956
rect 25228 38947 25280 38956
rect 25228 38913 25237 38947
rect 25237 38913 25271 38947
rect 25271 38913 25280 38947
rect 25228 38904 25280 38913
rect 20628 38768 20680 38820
rect 22652 38879 22704 38888
rect 22652 38845 22661 38879
rect 22661 38845 22695 38879
rect 22695 38845 22704 38879
rect 22652 38836 22704 38845
rect 23480 38879 23532 38888
rect 23480 38845 23489 38879
rect 23489 38845 23523 38879
rect 23523 38845 23532 38879
rect 23480 38836 23532 38845
rect 22008 38768 22060 38820
rect 23204 38768 23256 38820
rect 23756 38836 23808 38888
rect 25320 38836 25372 38888
rect 31668 38972 31720 39024
rect 32404 38972 32456 39024
rect 33140 38972 33192 39024
rect 36820 38972 36872 39024
rect 37832 38972 37884 39024
rect 29276 38879 29328 38888
rect 25504 38811 25556 38820
rect 19984 38743 20036 38752
rect 19984 38709 19993 38743
rect 19993 38709 20027 38743
rect 20027 38709 20036 38743
rect 19984 38700 20036 38709
rect 23388 38700 23440 38752
rect 23940 38743 23992 38752
rect 23940 38709 23949 38743
rect 23949 38709 23983 38743
rect 23983 38709 23992 38743
rect 23940 38700 23992 38709
rect 25504 38777 25513 38811
rect 25513 38777 25547 38811
rect 25547 38777 25556 38811
rect 25504 38768 25556 38777
rect 29276 38845 29285 38879
rect 29285 38845 29319 38879
rect 29319 38845 29328 38879
rect 29276 38836 29328 38845
rect 33048 38904 33100 38956
rect 30012 38836 30064 38888
rect 30748 38836 30800 38888
rect 34428 38879 34480 38888
rect 34428 38845 34437 38879
rect 34437 38845 34471 38879
rect 34471 38845 34480 38879
rect 34428 38836 34480 38845
rect 35624 38836 35676 38888
rect 39304 38836 39356 38888
rect 39948 38836 40000 38888
rect 41328 38836 41380 38888
rect 46940 38836 46992 38888
rect 30656 38768 30708 38820
rect 27068 38700 27120 38752
rect 29000 38743 29052 38752
rect 29000 38709 29009 38743
rect 29009 38709 29043 38743
rect 29043 38709 29052 38743
rect 29000 38700 29052 38709
rect 29184 38700 29236 38752
rect 31760 38743 31812 38752
rect 31760 38709 31769 38743
rect 31769 38709 31803 38743
rect 31803 38709 31812 38743
rect 31760 38700 31812 38709
rect 32680 38743 32732 38752
rect 32680 38709 32689 38743
rect 32689 38709 32723 38743
rect 32723 38709 32732 38743
rect 36452 38768 36504 38820
rect 37004 38768 37056 38820
rect 38844 38768 38896 38820
rect 32680 38700 32732 38709
rect 35900 38700 35952 38752
rect 38568 38700 38620 38752
rect 40776 38768 40828 38820
rect 40868 38700 40920 38752
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 11336 38496 11388 38548
rect 11704 38496 11756 38548
rect 12624 38539 12676 38548
rect 12624 38505 12633 38539
rect 12633 38505 12667 38539
rect 12667 38505 12676 38539
rect 12624 38496 12676 38505
rect 13728 38496 13780 38548
rect 16672 38539 16724 38548
rect 16672 38505 16681 38539
rect 16681 38505 16715 38539
rect 16715 38505 16724 38539
rect 16672 38496 16724 38505
rect 17868 38496 17920 38548
rect 18512 38539 18564 38548
rect 18512 38505 18521 38539
rect 18521 38505 18555 38539
rect 18555 38505 18564 38539
rect 18512 38496 18564 38505
rect 20444 38539 20496 38548
rect 20444 38505 20453 38539
rect 20453 38505 20487 38539
rect 20487 38505 20496 38539
rect 20444 38496 20496 38505
rect 23388 38496 23440 38548
rect 25228 38496 25280 38548
rect 25504 38496 25556 38548
rect 29000 38496 29052 38548
rect 30288 38496 30340 38548
rect 30932 38496 30984 38548
rect 33048 38496 33100 38548
rect 38108 38539 38160 38548
rect 38108 38505 38117 38539
rect 38117 38505 38151 38539
rect 38151 38505 38160 38539
rect 38108 38496 38160 38505
rect 38752 38496 38804 38548
rect 13268 38471 13320 38480
rect 13268 38437 13277 38471
rect 13277 38437 13311 38471
rect 13311 38437 13320 38471
rect 13268 38428 13320 38437
rect 13452 38428 13504 38480
rect 15476 38471 15528 38480
rect 15476 38437 15485 38471
rect 15485 38437 15519 38471
rect 15519 38437 15528 38471
rect 15476 38428 15528 38437
rect 21824 38428 21876 38480
rect 23204 38428 23256 38480
rect 27068 38471 27120 38480
rect 27068 38437 27077 38471
rect 27077 38437 27111 38471
rect 27111 38437 27120 38471
rect 27068 38428 27120 38437
rect 27712 38428 27764 38480
rect 29552 38428 29604 38480
rect 30104 38428 30156 38480
rect 31576 38428 31628 38480
rect 32588 38471 32640 38480
rect 32588 38437 32597 38471
rect 32597 38437 32631 38471
rect 32631 38437 32640 38471
rect 32588 38428 32640 38437
rect 32864 38428 32916 38480
rect 35808 38428 35860 38480
rect 41052 38428 41104 38480
rect 18420 38403 18472 38412
rect 18420 38369 18429 38403
rect 18429 38369 18463 38403
rect 18463 38369 18472 38403
rect 18420 38360 18472 38369
rect 19156 38360 19208 38412
rect 25136 38403 25188 38412
rect 25136 38369 25145 38403
rect 25145 38369 25179 38403
rect 25179 38369 25188 38403
rect 25136 38360 25188 38369
rect 25320 38403 25372 38412
rect 25320 38369 25329 38403
rect 25329 38369 25363 38403
rect 25363 38369 25372 38403
rect 25320 38360 25372 38369
rect 28448 38403 28500 38412
rect 28448 38369 28457 38403
rect 28457 38369 28491 38403
rect 28491 38369 28500 38403
rect 28448 38360 28500 38369
rect 33968 38360 34020 38412
rect 35900 38360 35952 38412
rect 37740 38403 37792 38412
rect 37740 38369 37749 38403
rect 37749 38369 37783 38403
rect 37783 38369 37792 38403
rect 37740 38360 37792 38369
rect 38844 38360 38896 38412
rect 39580 38360 39632 38412
rect 11520 38292 11572 38344
rect 12624 38292 12676 38344
rect 15844 38292 15896 38344
rect 16028 38335 16080 38344
rect 16028 38301 16037 38335
rect 16037 38301 16071 38335
rect 16071 38301 16080 38335
rect 16028 38292 16080 38301
rect 16948 38335 17000 38344
rect 16948 38301 16957 38335
rect 16957 38301 16991 38335
rect 16991 38301 17000 38335
rect 16948 38292 17000 38301
rect 17224 38335 17276 38344
rect 17224 38301 17233 38335
rect 17233 38301 17267 38335
rect 17267 38301 17276 38335
rect 17224 38292 17276 38301
rect 22192 38292 22244 38344
rect 22284 38335 22336 38344
rect 22284 38301 22293 38335
rect 22293 38301 22327 38335
rect 22327 38301 22336 38335
rect 22284 38292 22336 38301
rect 23204 38292 23256 38344
rect 23664 38335 23716 38344
rect 23664 38301 23673 38335
rect 23673 38301 23707 38335
rect 23707 38301 23716 38335
rect 23664 38292 23716 38301
rect 28080 38292 28132 38344
rect 29920 38292 29972 38344
rect 31852 38292 31904 38344
rect 32036 38292 32088 38344
rect 32864 38335 32916 38344
rect 32864 38301 32873 38335
rect 32873 38301 32907 38335
rect 32907 38301 32916 38335
rect 32864 38292 32916 38301
rect 34244 38292 34296 38344
rect 35256 38335 35308 38344
rect 35256 38301 35265 38335
rect 35265 38301 35299 38335
rect 35299 38301 35308 38335
rect 35256 38292 35308 38301
rect 40868 38335 40920 38344
rect 40868 38301 40877 38335
rect 40877 38301 40911 38335
rect 40911 38301 40920 38335
rect 40868 38292 40920 38301
rect 27528 38267 27580 38276
rect 27528 38233 27537 38267
rect 27537 38233 27571 38267
rect 27571 38233 27580 38267
rect 27528 38224 27580 38233
rect 41420 38267 41472 38276
rect 41420 38233 41429 38267
rect 41429 38233 41463 38267
rect 41463 38233 41472 38267
rect 41420 38224 41472 38233
rect 12348 38199 12400 38208
rect 12348 38165 12357 38199
rect 12357 38165 12391 38199
rect 12391 38165 12400 38199
rect 12348 38156 12400 38165
rect 12532 38156 12584 38208
rect 19156 38156 19208 38208
rect 19984 38156 20036 38208
rect 25136 38156 25188 38208
rect 29276 38199 29328 38208
rect 29276 38165 29285 38199
rect 29285 38165 29319 38199
rect 29319 38165 29328 38199
rect 29276 38156 29328 38165
rect 31944 38156 31996 38208
rect 35716 38156 35768 38208
rect 36452 38199 36504 38208
rect 36452 38165 36461 38199
rect 36461 38165 36495 38199
rect 36495 38165 36504 38199
rect 36452 38156 36504 38165
rect 36544 38156 36596 38208
rect 38936 38199 38988 38208
rect 38936 38165 38945 38199
rect 38945 38165 38979 38199
rect 38979 38165 38988 38199
rect 38936 38156 38988 38165
rect 42524 38199 42576 38208
rect 42524 38165 42533 38199
rect 42533 38165 42567 38199
rect 42567 38165 42576 38199
rect 42524 38156 42576 38165
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 13452 37995 13504 38004
rect 13452 37961 13461 37995
rect 13461 37961 13495 37995
rect 13495 37961 13504 37995
rect 13452 37952 13504 37961
rect 17684 37952 17736 38004
rect 18420 37995 18472 38004
rect 18420 37961 18429 37995
rect 18429 37961 18463 37995
rect 18463 37961 18472 37995
rect 18420 37952 18472 37961
rect 20628 37952 20680 38004
rect 22192 37995 22244 38004
rect 22192 37961 22201 37995
rect 22201 37961 22235 37995
rect 22235 37961 22244 37995
rect 22192 37952 22244 37961
rect 23296 37995 23348 38004
rect 23296 37961 23305 37995
rect 23305 37961 23339 37995
rect 23339 37961 23348 37995
rect 23296 37952 23348 37961
rect 24768 37995 24820 38004
rect 24768 37961 24777 37995
rect 24777 37961 24811 37995
rect 24811 37961 24820 37995
rect 24768 37952 24820 37961
rect 27712 37995 27764 38004
rect 27712 37961 27721 37995
rect 27721 37961 27755 37995
rect 27755 37961 27764 37995
rect 27712 37952 27764 37961
rect 28080 37995 28132 38004
rect 28080 37961 28089 37995
rect 28089 37961 28123 37995
rect 28123 37961 28132 37995
rect 28080 37952 28132 37961
rect 29552 37995 29604 38004
rect 29552 37961 29561 37995
rect 29561 37961 29595 37995
rect 29595 37961 29604 37995
rect 29552 37952 29604 37961
rect 29920 37952 29972 38004
rect 31760 37952 31812 38004
rect 32588 37952 32640 38004
rect 32864 37952 32916 38004
rect 33968 37995 34020 38004
rect 33968 37961 33977 37995
rect 33977 37961 34011 37995
rect 34011 37961 34020 37995
rect 33968 37952 34020 37961
rect 37740 37952 37792 38004
rect 38844 37952 38896 38004
rect 40868 37952 40920 38004
rect 12532 37859 12584 37868
rect 12532 37825 12541 37859
rect 12541 37825 12575 37859
rect 12575 37825 12584 37859
rect 12532 37816 12584 37825
rect 12624 37816 12676 37868
rect 13268 37884 13320 37936
rect 15844 37884 15896 37936
rect 17224 37884 17276 37936
rect 10232 37612 10284 37664
rect 11336 37791 11388 37800
rect 11336 37757 11345 37791
rect 11345 37757 11379 37791
rect 11379 37757 11388 37791
rect 11336 37748 11388 37757
rect 14740 37748 14792 37800
rect 15936 37791 15988 37800
rect 15936 37757 15945 37791
rect 15945 37757 15979 37791
rect 15979 37757 15988 37791
rect 15936 37748 15988 37757
rect 17224 37791 17276 37800
rect 17224 37757 17233 37791
rect 17233 37757 17267 37791
rect 17267 37757 17276 37791
rect 17224 37748 17276 37757
rect 19340 37791 19392 37800
rect 19340 37757 19349 37791
rect 19349 37757 19383 37791
rect 19383 37757 19392 37791
rect 19340 37748 19392 37757
rect 20628 37791 20680 37800
rect 11520 37723 11572 37732
rect 11520 37689 11529 37723
rect 11529 37689 11563 37723
rect 11563 37689 11572 37723
rect 11520 37680 11572 37689
rect 11704 37612 11756 37664
rect 11980 37612 12032 37664
rect 12348 37612 12400 37664
rect 15292 37723 15344 37732
rect 14740 37655 14792 37664
rect 14740 37621 14749 37655
rect 14749 37621 14783 37655
rect 14783 37621 14792 37655
rect 14740 37612 14792 37621
rect 15292 37689 15301 37723
rect 15301 37689 15335 37723
rect 15335 37689 15344 37723
rect 15292 37680 15344 37689
rect 15476 37680 15528 37732
rect 16948 37680 17000 37732
rect 17592 37680 17644 37732
rect 19156 37680 19208 37732
rect 20628 37757 20637 37791
rect 20637 37757 20671 37791
rect 20671 37757 20680 37791
rect 20628 37748 20680 37757
rect 25136 37884 25188 37936
rect 22560 37748 22612 37800
rect 20720 37680 20772 37732
rect 21824 37655 21876 37664
rect 21824 37621 21833 37655
rect 21833 37621 21867 37655
rect 21867 37621 21876 37655
rect 21824 37612 21876 37621
rect 23388 37612 23440 37664
rect 26516 37816 26568 37868
rect 28448 37859 28500 37868
rect 28448 37825 28457 37859
rect 28457 37825 28491 37859
rect 28491 37825 28500 37859
rect 28448 37816 28500 37825
rect 24768 37748 24820 37800
rect 30748 37859 30800 37868
rect 30748 37825 30757 37859
rect 30757 37825 30791 37859
rect 30791 37825 30800 37859
rect 30748 37816 30800 37825
rect 31668 37884 31720 37936
rect 31944 37816 31996 37868
rect 32772 37859 32824 37868
rect 32772 37825 32781 37859
rect 32781 37825 32815 37859
rect 32815 37825 32824 37859
rect 32772 37816 32824 37825
rect 33232 37816 33284 37868
rect 30104 37748 30156 37800
rect 24676 37680 24728 37732
rect 25504 37680 25556 37732
rect 24308 37612 24360 37664
rect 26608 37612 26660 37664
rect 26700 37612 26752 37664
rect 26884 37723 26936 37732
rect 26884 37689 26893 37723
rect 26893 37689 26927 37723
rect 26927 37689 26936 37723
rect 26884 37680 26936 37689
rect 27804 37680 27856 37732
rect 29736 37680 29788 37732
rect 32864 37723 32916 37732
rect 32864 37689 32873 37723
rect 32873 37689 32907 37723
rect 32907 37689 32916 37723
rect 33416 37723 33468 37732
rect 32864 37680 32916 37689
rect 33416 37689 33425 37723
rect 33425 37689 33459 37723
rect 33459 37689 33468 37723
rect 33416 37680 33468 37689
rect 32036 37612 32088 37664
rect 35808 37884 35860 37936
rect 38108 37884 38160 37936
rect 40040 37884 40092 37936
rect 42156 37884 42208 37936
rect 36544 37816 36596 37868
rect 38936 37816 38988 37868
rect 40960 37859 41012 37868
rect 40960 37825 40969 37859
rect 40969 37825 41003 37859
rect 41003 37825 41012 37859
rect 40960 37816 41012 37825
rect 41236 37859 41288 37868
rect 41236 37825 41245 37859
rect 41245 37825 41279 37859
rect 41279 37825 41288 37859
rect 41236 37816 41288 37825
rect 35992 37791 36044 37800
rect 35992 37757 36001 37791
rect 36001 37757 36035 37791
rect 36035 37757 36044 37791
rect 35992 37748 36044 37757
rect 39580 37748 39632 37800
rect 40684 37748 40736 37800
rect 36452 37680 36504 37732
rect 37188 37680 37240 37732
rect 38844 37680 38896 37732
rect 39304 37723 39356 37732
rect 39304 37689 39313 37723
rect 39313 37689 39347 37723
rect 39347 37689 39356 37723
rect 39304 37680 39356 37689
rect 41052 37723 41104 37732
rect 41052 37689 41061 37723
rect 41061 37689 41095 37723
rect 41095 37689 41104 37723
rect 41052 37680 41104 37689
rect 42524 37723 42576 37732
rect 42524 37689 42533 37723
rect 42533 37689 42567 37723
rect 42567 37689 42576 37723
rect 42524 37680 42576 37689
rect 40868 37612 40920 37664
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 10876 37451 10928 37460
rect 10876 37417 10885 37451
rect 10885 37417 10919 37451
rect 10919 37417 10928 37451
rect 10876 37408 10928 37417
rect 11336 37408 11388 37460
rect 11520 37451 11572 37460
rect 11520 37417 11529 37451
rect 11529 37417 11563 37451
rect 11563 37417 11572 37451
rect 11520 37408 11572 37417
rect 12532 37408 12584 37460
rect 15292 37408 15344 37460
rect 15844 37408 15896 37460
rect 17592 37451 17644 37460
rect 17592 37417 17601 37451
rect 17601 37417 17635 37451
rect 17635 37417 17644 37451
rect 17592 37408 17644 37417
rect 20628 37451 20680 37460
rect 20628 37417 20637 37451
rect 20637 37417 20671 37451
rect 20671 37417 20680 37451
rect 20628 37408 20680 37417
rect 25136 37451 25188 37460
rect 25136 37417 25145 37451
rect 25145 37417 25179 37451
rect 25179 37417 25188 37451
rect 25136 37408 25188 37417
rect 25320 37408 25372 37460
rect 29000 37408 29052 37460
rect 29644 37408 29696 37460
rect 30012 37451 30064 37460
rect 30012 37417 30021 37451
rect 30021 37417 30055 37451
rect 30055 37417 30064 37451
rect 30012 37408 30064 37417
rect 31576 37408 31628 37460
rect 32496 37451 32548 37460
rect 32496 37417 32505 37451
rect 32505 37417 32539 37451
rect 32539 37417 32548 37451
rect 32496 37408 32548 37417
rect 33232 37408 33284 37460
rect 35256 37451 35308 37460
rect 35256 37417 35265 37451
rect 35265 37417 35299 37451
rect 35299 37417 35308 37451
rect 35256 37408 35308 37417
rect 36452 37451 36504 37460
rect 36452 37417 36461 37451
rect 36461 37417 36495 37451
rect 36495 37417 36504 37451
rect 36452 37408 36504 37417
rect 40868 37451 40920 37460
rect 40868 37417 40877 37451
rect 40877 37417 40911 37451
rect 40911 37417 40920 37451
rect 40868 37408 40920 37417
rect 40960 37408 41012 37460
rect 12164 37340 12216 37392
rect 14280 37340 14332 37392
rect 17224 37340 17276 37392
rect 21824 37340 21876 37392
rect 23664 37340 23716 37392
rect 24768 37383 24820 37392
rect 24768 37349 24777 37383
rect 24777 37349 24811 37383
rect 24811 37349 24820 37383
rect 24768 37340 24820 37349
rect 13452 37272 13504 37324
rect 16028 37272 16080 37324
rect 16488 37272 16540 37324
rect 17040 37272 17092 37324
rect 11244 37204 11296 37256
rect 12164 37247 12216 37256
rect 12164 37213 12173 37247
rect 12173 37213 12207 37247
rect 12207 37213 12216 37247
rect 12164 37204 12216 37213
rect 12624 37247 12676 37256
rect 12624 37213 12633 37247
rect 12633 37213 12667 37247
rect 12667 37213 12676 37247
rect 12624 37204 12676 37213
rect 17316 37247 17368 37256
rect 17316 37213 17325 37247
rect 17325 37213 17359 37247
rect 17359 37213 17368 37247
rect 17316 37204 17368 37213
rect 18144 37315 18196 37324
rect 18144 37281 18153 37315
rect 18153 37281 18187 37315
rect 18187 37281 18196 37315
rect 18144 37272 18196 37281
rect 24032 37315 24084 37324
rect 24032 37281 24041 37315
rect 24041 37281 24075 37315
rect 24075 37281 24084 37315
rect 24032 37272 24084 37281
rect 24584 37315 24636 37324
rect 24584 37281 24593 37315
rect 24593 37281 24627 37315
rect 24627 37281 24636 37315
rect 26792 37340 26844 37392
rect 28632 37383 28684 37392
rect 28632 37349 28641 37383
rect 28641 37349 28675 37383
rect 28675 37349 28684 37383
rect 28632 37340 28684 37349
rect 31392 37340 31444 37392
rect 32312 37340 32364 37392
rect 24584 37272 24636 37281
rect 30748 37272 30800 37324
rect 30840 37315 30892 37324
rect 30840 37281 30849 37315
rect 30849 37281 30883 37315
rect 30883 37281 30892 37315
rect 30840 37272 30892 37281
rect 32680 37272 32732 37324
rect 40040 37340 40092 37392
rect 41604 37340 41656 37392
rect 35716 37315 35768 37324
rect 35716 37281 35725 37315
rect 35725 37281 35759 37315
rect 35759 37281 35768 37315
rect 35716 37272 35768 37281
rect 35900 37315 35952 37324
rect 35900 37281 35909 37315
rect 35909 37281 35943 37315
rect 35943 37281 35952 37315
rect 35900 37272 35952 37281
rect 38844 37315 38896 37324
rect 18696 37247 18748 37256
rect 14372 37068 14424 37120
rect 18420 37068 18472 37120
rect 18696 37213 18705 37247
rect 18705 37213 18739 37247
rect 18739 37213 18748 37247
rect 18696 37204 18748 37213
rect 19708 37204 19760 37256
rect 23388 37204 23440 37256
rect 26976 37247 27028 37256
rect 26976 37213 26985 37247
rect 26985 37213 27019 37247
rect 27019 37213 27028 37247
rect 26976 37204 27028 37213
rect 27252 37247 27304 37256
rect 27252 37213 27261 37247
rect 27261 37213 27295 37247
rect 27295 37213 27304 37247
rect 27252 37204 27304 37213
rect 28540 37247 28592 37256
rect 28540 37213 28549 37247
rect 28549 37213 28583 37247
rect 28583 37213 28592 37247
rect 28540 37204 28592 37213
rect 28816 37247 28868 37256
rect 28816 37213 28825 37247
rect 28825 37213 28859 37247
rect 28859 37213 28868 37247
rect 28816 37204 28868 37213
rect 32312 37204 32364 37256
rect 33784 37204 33836 37256
rect 34244 37247 34296 37256
rect 34244 37213 34253 37247
rect 34253 37213 34287 37247
rect 34287 37213 34296 37247
rect 34244 37204 34296 37213
rect 23204 37136 23256 37188
rect 31576 37136 31628 37188
rect 38844 37281 38853 37315
rect 38853 37281 38887 37315
rect 38887 37281 38896 37315
rect 38844 37272 38896 37281
rect 40132 37204 40184 37256
rect 41788 37247 41840 37256
rect 41788 37213 41797 37247
rect 41797 37213 41831 37247
rect 41831 37213 41840 37247
rect 41788 37204 41840 37213
rect 42616 37204 42668 37256
rect 39028 37136 39080 37188
rect 19156 37111 19208 37120
rect 19156 37077 19165 37111
rect 19165 37077 19199 37111
rect 19199 37077 19208 37111
rect 19156 37068 19208 37077
rect 19248 37068 19300 37120
rect 21732 37068 21784 37120
rect 24768 37068 24820 37120
rect 26700 37111 26752 37120
rect 26700 37077 26709 37111
rect 26709 37077 26743 37111
rect 26743 37077 26752 37111
rect 26700 37068 26752 37077
rect 33692 37111 33744 37120
rect 33692 37077 33701 37111
rect 33701 37077 33735 37111
rect 33735 37077 33744 37111
rect 33692 37068 33744 37077
rect 36820 37111 36872 37120
rect 36820 37077 36829 37111
rect 36829 37077 36863 37111
rect 36863 37077 36872 37111
rect 36820 37068 36872 37077
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 12164 36907 12216 36916
rect 12164 36873 12173 36907
rect 12173 36873 12207 36907
rect 12207 36873 12216 36907
rect 12164 36864 12216 36873
rect 13452 36907 13504 36916
rect 13452 36873 13461 36907
rect 13461 36873 13495 36907
rect 13495 36873 13504 36907
rect 13452 36864 13504 36873
rect 16028 36864 16080 36916
rect 17040 36907 17092 36916
rect 17040 36873 17049 36907
rect 17049 36873 17083 36907
rect 17083 36873 17092 36907
rect 17040 36864 17092 36873
rect 18788 36864 18840 36916
rect 19708 36864 19760 36916
rect 21824 36907 21876 36916
rect 13268 36796 13320 36848
rect 13820 36728 13872 36780
rect 15936 36796 15988 36848
rect 21824 36873 21833 36907
rect 21833 36873 21867 36907
rect 21867 36873 21876 36907
rect 21824 36864 21876 36873
rect 23388 36864 23440 36916
rect 24032 36864 24084 36916
rect 26700 36864 26752 36916
rect 30840 36864 30892 36916
rect 32680 36907 32732 36916
rect 32680 36873 32689 36907
rect 32689 36873 32723 36907
rect 32723 36873 32732 36907
rect 32680 36864 32732 36873
rect 33784 36864 33836 36916
rect 26516 36796 26568 36848
rect 26792 36796 26844 36848
rect 27068 36796 27120 36848
rect 28632 36796 28684 36848
rect 16764 36728 16816 36780
rect 18696 36771 18748 36780
rect 18696 36737 18705 36771
rect 18705 36737 18739 36771
rect 18739 36737 18748 36771
rect 18696 36728 18748 36737
rect 20536 36771 20588 36780
rect 20536 36737 20545 36771
rect 20545 36737 20579 36771
rect 20579 36737 20588 36771
rect 20536 36728 20588 36737
rect 22560 36728 22612 36780
rect 32220 36796 32272 36848
rect 33416 36796 33468 36848
rect 31392 36771 31444 36780
rect 13728 36635 13780 36644
rect 13728 36601 13737 36635
rect 13737 36601 13771 36635
rect 13771 36601 13780 36635
rect 13728 36592 13780 36601
rect 15200 36635 15252 36644
rect 15200 36601 15209 36635
rect 15209 36601 15243 36635
rect 15243 36601 15252 36635
rect 15200 36592 15252 36601
rect 11244 36524 11296 36576
rect 11612 36524 11664 36576
rect 14464 36524 14516 36576
rect 18788 36592 18840 36644
rect 16488 36524 16540 36576
rect 17408 36524 17460 36576
rect 18144 36524 18196 36576
rect 21732 36660 21784 36712
rect 23296 36660 23348 36712
rect 24308 36660 24360 36712
rect 31392 36737 31401 36771
rect 31401 36737 31435 36771
rect 31435 36737 31444 36771
rect 31392 36728 31444 36737
rect 31668 36771 31720 36780
rect 31668 36737 31677 36771
rect 31677 36737 31711 36771
rect 31711 36737 31720 36771
rect 31668 36728 31720 36737
rect 32956 36771 33008 36780
rect 32956 36737 32965 36771
rect 32965 36737 32999 36771
rect 32999 36737 33008 36771
rect 32956 36728 33008 36737
rect 33692 36728 33744 36780
rect 35900 36728 35952 36780
rect 37464 36864 37516 36916
rect 37004 36796 37056 36848
rect 38936 36864 38988 36916
rect 39028 36907 39080 36916
rect 39028 36873 39037 36907
rect 39037 36873 39071 36907
rect 39071 36873 39080 36907
rect 41604 36907 41656 36916
rect 39028 36864 39080 36873
rect 41604 36873 41613 36907
rect 41613 36873 41647 36907
rect 41647 36873 41656 36907
rect 41604 36864 41656 36873
rect 42524 36864 42576 36916
rect 38844 36796 38896 36848
rect 41788 36796 41840 36848
rect 36912 36771 36964 36780
rect 36912 36737 36921 36771
rect 36921 36737 36955 36771
rect 36955 36737 36964 36771
rect 36912 36728 36964 36737
rect 37280 36728 37332 36780
rect 27528 36703 27580 36712
rect 27528 36669 27537 36703
rect 27537 36669 27571 36703
rect 27571 36669 27580 36703
rect 27528 36660 27580 36669
rect 34704 36703 34756 36712
rect 21180 36635 21232 36644
rect 21180 36601 21189 36635
rect 21189 36601 21223 36635
rect 21223 36601 21232 36635
rect 21180 36592 21232 36601
rect 23112 36592 23164 36644
rect 24216 36592 24268 36644
rect 24584 36592 24636 36644
rect 21916 36524 21968 36576
rect 23572 36524 23624 36576
rect 26792 36524 26844 36576
rect 27068 36592 27120 36644
rect 29000 36567 29052 36576
rect 29000 36533 29009 36567
rect 29009 36533 29043 36567
rect 29043 36533 29052 36567
rect 34704 36669 34713 36703
rect 34713 36669 34747 36703
rect 34747 36669 34756 36703
rect 34704 36660 34756 36669
rect 35440 36703 35492 36712
rect 35440 36669 35449 36703
rect 35449 36669 35483 36703
rect 35483 36669 35492 36703
rect 35440 36660 35492 36669
rect 35716 36660 35768 36712
rect 36268 36660 36320 36712
rect 38016 36660 38068 36712
rect 29644 36592 29696 36644
rect 30748 36592 30800 36644
rect 30472 36567 30524 36576
rect 29000 36524 29052 36533
rect 30472 36533 30481 36567
rect 30481 36533 30515 36567
rect 30515 36533 30524 36567
rect 30472 36524 30524 36533
rect 31484 36635 31536 36644
rect 31484 36601 31493 36635
rect 31493 36601 31527 36635
rect 31527 36601 31536 36635
rect 31484 36592 31536 36601
rect 32680 36592 32732 36644
rect 35624 36635 35676 36644
rect 35624 36601 35633 36635
rect 35633 36601 35667 36635
rect 35667 36601 35676 36635
rect 35624 36592 35676 36601
rect 36820 36592 36872 36644
rect 41144 36660 41196 36712
rect 41696 36660 41748 36712
rect 31576 36524 31628 36576
rect 31852 36524 31904 36576
rect 32496 36524 32548 36576
rect 33232 36524 33284 36576
rect 42340 36592 42392 36644
rect 38016 36524 38068 36576
rect 40040 36567 40092 36576
rect 40040 36533 40049 36567
rect 40049 36533 40083 36567
rect 40083 36533 40092 36567
rect 40040 36524 40092 36533
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 13728 36320 13780 36372
rect 14004 36363 14056 36372
rect 14004 36329 14013 36363
rect 14013 36329 14047 36363
rect 14047 36329 14056 36363
rect 14004 36320 14056 36329
rect 15200 36320 15252 36372
rect 16304 36320 16356 36372
rect 20536 36363 20588 36372
rect 20536 36329 20545 36363
rect 20545 36329 20579 36363
rect 20579 36329 20588 36363
rect 20536 36320 20588 36329
rect 12716 36295 12768 36304
rect 12716 36261 12725 36295
rect 12725 36261 12759 36295
rect 12759 36261 12768 36295
rect 12716 36252 12768 36261
rect 13268 36295 13320 36304
rect 13268 36261 13277 36295
rect 13277 36261 13311 36295
rect 13311 36261 13320 36295
rect 13268 36252 13320 36261
rect 18788 36252 18840 36304
rect 19892 36295 19944 36304
rect 19892 36261 19901 36295
rect 19901 36261 19935 36295
rect 19935 36261 19944 36295
rect 19892 36252 19944 36261
rect 22100 36252 22152 36304
rect 26976 36320 27028 36372
rect 27068 36320 27120 36372
rect 30472 36320 30524 36372
rect 30748 36363 30800 36372
rect 30748 36329 30757 36363
rect 30757 36329 30791 36363
rect 30791 36329 30800 36363
rect 30748 36320 30800 36329
rect 32312 36363 32364 36372
rect 32312 36329 32321 36363
rect 32321 36329 32355 36363
rect 32355 36329 32364 36363
rect 32312 36320 32364 36329
rect 35624 36363 35676 36372
rect 35624 36329 35633 36363
rect 35633 36329 35667 36363
rect 35667 36329 35676 36363
rect 35624 36320 35676 36329
rect 36176 36363 36228 36372
rect 36176 36329 36185 36363
rect 36185 36329 36219 36363
rect 36219 36329 36228 36363
rect 36176 36320 36228 36329
rect 37740 36320 37792 36372
rect 40132 36363 40184 36372
rect 22744 36252 22796 36304
rect 23020 36252 23072 36304
rect 10416 36227 10468 36236
rect 10416 36193 10425 36227
rect 10425 36193 10459 36227
rect 10459 36193 10468 36227
rect 10416 36184 10468 36193
rect 10876 36227 10928 36236
rect 10876 36193 10885 36227
rect 10885 36193 10919 36227
rect 10919 36193 10928 36227
rect 10876 36184 10928 36193
rect 14096 36227 14148 36236
rect 14096 36193 14105 36227
rect 14105 36193 14139 36227
rect 14139 36193 14148 36227
rect 14096 36184 14148 36193
rect 15292 36184 15344 36236
rect 10968 36159 11020 36168
rect 10968 36125 10977 36159
rect 10977 36125 11011 36159
rect 11011 36125 11020 36159
rect 10968 36116 11020 36125
rect 12164 36116 12216 36168
rect 12624 36159 12676 36168
rect 12624 36125 12633 36159
rect 12633 36125 12667 36159
rect 12667 36125 12676 36159
rect 12624 36116 12676 36125
rect 16396 36159 16448 36168
rect 16396 36125 16405 36159
rect 16405 36125 16439 36159
rect 16439 36125 16448 36159
rect 16396 36116 16448 36125
rect 17316 36184 17368 36236
rect 18328 36184 18380 36236
rect 21732 36184 21784 36236
rect 24216 36227 24268 36236
rect 20996 36116 21048 36168
rect 21916 36159 21968 36168
rect 21916 36125 21925 36159
rect 21925 36125 21959 36159
rect 21959 36125 21968 36159
rect 21916 36116 21968 36125
rect 16488 36048 16540 36100
rect 23388 36048 23440 36100
rect 24216 36193 24225 36227
rect 24225 36193 24259 36227
rect 24259 36193 24268 36227
rect 24216 36184 24268 36193
rect 24768 36184 24820 36236
rect 25412 36227 25464 36236
rect 29000 36252 29052 36304
rect 29644 36252 29696 36304
rect 31852 36252 31904 36304
rect 32036 36252 32088 36304
rect 32864 36295 32916 36304
rect 32864 36261 32873 36295
rect 32873 36261 32907 36295
rect 32907 36261 32916 36295
rect 32864 36252 32916 36261
rect 33140 36252 33192 36304
rect 37832 36295 37884 36304
rect 37832 36261 37841 36295
rect 37841 36261 37875 36295
rect 37875 36261 37884 36295
rect 37832 36252 37884 36261
rect 40132 36329 40141 36363
rect 40141 36329 40175 36363
rect 40175 36329 40184 36363
rect 40132 36320 40184 36329
rect 38016 36252 38068 36304
rect 41236 36320 41288 36372
rect 41788 36363 41840 36372
rect 40868 36295 40920 36304
rect 40868 36261 40877 36295
rect 40877 36261 40911 36295
rect 40911 36261 40920 36295
rect 40868 36252 40920 36261
rect 41788 36329 41797 36363
rect 41797 36329 41831 36363
rect 41831 36329 41840 36363
rect 41788 36320 41840 36329
rect 25412 36193 25456 36227
rect 25456 36193 25464 36227
rect 25412 36184 25464 36193
rect 27068 36184 27120 36236
rect 28356 36184 28408 36236
rect 28448 36227 28500 36236
rect 28448 36193 28457 36227
rect 28457 36193 28491 36227
rect 28491 36193 28500 36227
rect 28448 36184 28500 36193
rect 29460 36184 29512 36236
rect 30012 36184 30064 36236
rect 31484 36184 31536 36236
rect 34336 36227 34388 36236
rect 34336 36193 34345 36227
rect 34345 36193 34379 36227
rect 34379 36193 34388 36227
rect 34336 36184 34388 36193
rect 39672 36227 39724 36236
rect 39672 36193 39681 36227
rect 39681 36193 39715 36227
rect 39715 36193 39724 36227
rect 39672 36184 39724 36193
rect 24308 36159 24360 36168
rect 24308 36125 24317 36159
rect 24317 36125 24351 36159
rect 24351 36125 24360 36159
rect 24308 36116 24360 36125
rect 28540 36116 28592 36168
rect 29552 36159 29604 36168
rect 29552 36125 29561 36159
rect 29561 36125 29595 36159
rect 29595 36125 29604 36159
rect 29552 36116 29604 36125
rect 35808 36159 35860 36168
rect 28356 36048 28408 36100
rect 31392 36048 31444 36100
rect 35808 36125 35817 36159
rect 35817 36125 35851 36159
rect 35851 36125 35860 36159
rect 35808 36116 35860 36125
rect 36912 36048 36964 36100
rect 41696 36116 41748 36168
rect 38476 36048 38528 36100
rect 12072 36023 12124 36032
rect 12072 35989 12081 36023
rect 12081 35989 12115 36023
rect 12115 35989 12124 36023
rect 12072 35980 12124 35989
rect 14648 35980 14700 36032
rect 16580 35980 16632 36032
rect 18420 35980 18472 36032
rect 19524 36023 19576 36032
rect 19524 35989 19533 36023
rect 19533 35989 19567 36023
rect 19567 35989 19576 36023
rect 19524 35980 19576 35989
rect 24768 36023 24820 36032
rect 24768 35989 24777 36023
rect 24777 35989 24811 36023
rect 24811 35989 24820 36023
rect 24768 35980 24820 35989
rect 27712 36023 27764 36032
rect 27712 35989 27721 36023
rect 27721 35989 27755 36023
rect 27755 35989 27764 36023
rect 27712 35980 27764 35989
rect 34796 35980 34848 36032
rect 35440 35980 35492 36032
rect 37004 35980 37056 36032
rect 40776 35980 40828 36032
rect 41420 35980 41472 36032
rect 42432 35980 42484 36032
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 9680 35776 9732 35828
rect 10416 35819 10468 35828
rect 10416 35785 10425 35819
rect 10425 35785 10459 35819
rect 10459 35785 10468 35819
rect 10416 35776 10468 35785
rect 10876 35776 10928 35828
rect 11336 35776 11388 35828
rect 13728 35776 13780 35828
rect 16304 35819 16356 35828
rect 16304 35785 16313 35819
rect 16313 35785 16347 35819
rect 16347 35785 16356 35819
rect 16304 35776 16356 35785
rect 18328 35819 18380 35828
rect 18328 35785 18337 35819
rect 18337 35785 18371 35819
rect 18371 35785 18380 35819
rect 18328 35776 18380 35785
rect 18788 35776 18840 35828
rect 19524 35776 19576 35828
rect 19892 35776 19944 35828
rect 20996 35819 21048 35828
rect 12532 35708 12584 35760
rect 14004 35708 14056 35760
rect 14096 35683 14148 35692
rect 14096 35649 14105 35683
rect 14105 35649 14139 35683
rect 14139 35649 14148 35683
rect 14096 35640 14148 35649
rect 14372 35683 14424 35692
rect 14372 35649 14381 35683
rect 14381 35649 14415 35683
rect 14415 35649 14424 35683
rect 14372 35640 14424 35649
rect 20996 35785 21005 35819
rect 21005 35785 21039 35819
rect 21039 35785 21048 35819
rect 20996 35776 21048 35785
rect 23112 35819 23164 35828
rect 23112 35785 23121 35819
rect 23121 35785 23155 35819
rect 23155 35785 23164 35819
rect 23112 35776 23164 35785
rect 23388 35819 23440 35828
rect 23388 35785 23397 35819
rect 23397 35785 23431 35819
rect 23431 35785 23440 35819
rect 23388 35776 23440 35785
rect 24676 35776 24728 35828
rect 25412 35776 25464 35828
rect 27068 35819 27120 35828
rect 27068 35785 27077 35819
rect 27077 35785 27111 35819
rect 27111 35785 27120 35819
rect 27068 35776 27120 35785
rect 28448 35776 28500 35828
rect 29552 35776 29604 35828
rect 29644 35776 29696 35828
rect 32496 35776 32548 35828
rect 34336 35776 34388 35828
rect 16580 35640 16632 35692
rect 16764 35683 16816 35692
rect 16764 35649 16773 35683
rect 16773 35649 16807 35683
rect 16807 35649 16816 35683
rect 16764 35640 16816 35649
rect 28816 35708 28868 35760
rect 19892 35683 19944 35692
rect 19892 35649 19901 35683
rect 19901 35649 19935 35683
rect 19935 35649 19944 35683
rect 19892 35640 19944 35649
rect 22008 35640 22060 35692
rect 23572 35640 23624 35692
rect 24768 35640 24820 35692
rect 26148 35683 26200 35692
rect 26148 35649 26157 35683
rect 26157 35649 26191 35683
rect 26191 35649 26200 35683
rect 26148 35640 26200 35649
rect 26424 35683 26476 35692
rect 26424 35649 26433 35683
rect 26433 35649 26467 35683
rect 26467 35649 26476 35683
rect 26424 35640 26476 35649
rect 28172 35640 28224 35692
rect 28356 35640 28408 35692
rect 28724 35683 28776 35692
rect 28724 35649 28733 35683
rect 28733 35649 28767 35683
rect 28767 35649 28776 35683
rect 28724 35640 28776 35649
rect 32404 35708 32456 35760
rect 36820 35776 36872 35828
rect 37740 35819 37792 35828
rect 37740 35785 37749 35819
rect 37749 35785 37783 35819
rect 37783 35785 37792 35819
rect 37740 35776 37792 35785
rect 38384 35776 38436 35828
rect 39672 35819 39724 35828
rect 39672 35785 39681 35819
rect 39681 35785 39715 35819
rect 39715 35785 39724 35819
rect 39672 35776 39724 35785
rect 41696 35819 41748 35828
rect 41696 35785 41705 35819
rect 41705 35785 41739 35819
rect 41739 35785 41748 35819
rect 41696 35776 41748 35785
rect 31300 35683 31352 35692
rect 31300 35649 31309 35683
rect 31309 35649 31343 35683
rect 31343 35649 31352 35683
rect 31300 35640 31352 35649
rect 31668 35640 31720 35692
rect 33048 35640 33100 35692
rect 37280 35708 37332 35760
rect 35624 35640 35676 35692
rect 35808 35640 35860 35692
rect 39304 35708 39356 35760
rect 38476 35683 38528 35692
rect 38476 35649 38485 35683
rect 38485 35649 38519 35683
rect 38519 35649 38528 35683
rect 38476 35640 38528 35649
rect 40776 35683 40828 35692
rect 40776 35649 40785 35683
rect 40785 35649 40819 35683
rect 40819 35649 40828 35683
rect 40776 35640 40828 35649
rect 41420 35683 41472 35692
rect 41420 35649 41429 35683
rect 41429 35649 41463 35683
rect 41463 35649 41472 35683
rect 41420 35640 41472 35649
rect 42616 35683 42668 35692
rect 42616 35649 42625 35683
rect 42625 35649 42659 35683
rect 42659 35649 42668 35683
rect 42616 35640 42668 35649
rect 11336 35615 11388 35624
rect 11336 35581 11345 35615
rect 11345 35581 11379 35615
rect 11379 35581 11388 35615
rect 11336 35572 11388 35581
rect 11980 35504 12032 35556
rect 13360 35504 13412 35556
rect 14464 35547 14516 35556
rect 14464 35513 14473 35547
rect 14473 35513 14507 35547
rect 14507 35513 14516 35547
rect 14464 35504 14516 35513
rect 15936 35504 15988 35556
rect 15292 35479 15344 35488
rect 15292 35445 15301 35479
rect 15301 35445 15335 35479
rect 15335 35445 15344 35479
rect 15292 35436 15344 35445
rect 16580 35547 16632 35556
rect 16580 35513 16589 35547
rect 16589 35513 16623 35547
rect 16623 35513 16632 35547
rect 16580 35504 16632 35513
rect 19708 35547 19760 35556
rect 19708 35513 19717 35547
rect 19717 35513 19751 35547
rect 19751 35513 19760 35547
rect 19708 35504 19760 35513
rect 22100 35504 22152 35556
rect 22376 35436 22428 35488
rect 24676 35479 24728 35488
rect 24676 35445 24685 35479
rect 24685 35445 24719 35479
rect 24719 35445 24728 35479
rect 24676 35436 24728 35445
rect 25228 35479 25280 35488
rect 25228 35445 25237 35479
rect 25237 35445 25271 35479
rect 25271 35445 25280 35479
rect 25228 35436 25280 35445
rect 25872 35479 25924 35488
rect 25872 35445 25881 35479
rect 25881 35445 25915 35479
rect 25915 35445 25924 35479
rect 27712 35504 27764 35556
rect 25872 35436 25924 35445
rect 26516 35436 26568 35488
rect 29736 35615 29788 35624
rect 29736 35581 29745 35615
rect 29745 35581 29779 35615
rect 29779 35581 29788 35615
rect 29736 35572 29788 35581
rect 30748 35547 30800 35556
rect 30748 35513 30757 35547
rect 30757 35513 30791 35547
rect 30791 35513 30800 35547
rect 30748 35504 30800 35513
rect 33140 35504 33192 35556
rect 36176 35504 36228 35556
rect 40868 35547 40920 35556
rect 28724 35436 28776 35488
rect 40868 35513 40877 35547
rect 40877 35513 40911 35547
rect 40911 35513 40920 35547
rect 40868 35504 40920 35513
rect 38660 35436 38712 35488
rect 42064 35479 42116 35488
rect 42064 35445 42073 35479
rect 42073 35445 42107 35479
rect 42107 35445 42116 35479
rect 42432 35547 42484 35556
rect 42432 35513 42441 35547
rect 42441 35513 42475 35547
rect 42475 35513 42484 35547
rect 42432 35504 42484 35513
rect 42064 35436 42116 35445
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 10876 35232 10928 35284
rect 12164 35275 12216 35284
rect 12164 35241 12173 35275
rect 12173 35241 12207 35275
rect 12207 35241 12216 35275
rect 12164 35232 12216 35241
rect 12716 35232 12768 35284
rect 14372 35232 14424 35284
rect 16396 35232 16448 35284
rect 22008 35275 22060 35284
rect 22008 35241 22017 35275
rect 22017 35241 22051 35275
rect 22051 35241 22060 35275
rect 22008 35232 22060 35241
rect 23112 35232 23164 35284
rect 23848 35232 23900 35284
rect 24676 35275 24728 35284
rect 24676 35241 24685 35275
rect 24685 35241 24719 35275
rect 24719 35241 24728 35275
rect 24676 35232 24728 35241
rect 25872 35232 25924 35284
rect 26148 35275 26200 35284
rect 26148 35241 26157 35275
rect 26157 35241 26191 35275
rect 26191 35241 26200 35275
rect 26148 35232 26200 35241
rect 11980 35164 12032 35216
rect 13360 35164 13412 35216
rect 15660 35164 15712 35216
rect 16304 35164 16356 35216
rect 19340 35164 19392 35216
rect 21088 35207 21140 35216
rect 21088 35173 21097 35207
rect 21097 35173 21131 35207
rect 21131 35173 21140 35207
rect 21088 35164 21140 35173
rect 22100 35164 22152 35216
rect 25412 35164 25464 35216
rect 27160 35164 27212 35216
rect 27344 35232 27396 35284
rect 27712 35232 27764 35284
rect 32864 35275 32916 35284
rect 32864 35241 32873 35275
rect 32873 35241 32907 35275
rect 32907 35241 32916 35275
rect 32864 35232 32916 35241
rect 37832 35232 37884 35284
rect 38660 35275 38712 35284
rect 38660 35241 38669 35275
rect 38669 35241 38703 35275
rect 38703 35241 38712 35275
rect 38660 35232 38712 35241
rect 29552 35164 29604 35216
rect 33140 35207 33192 35216
rect 33140 35173 33149 35207
rect 33149 35173 33183 35207
rect 33183 35173 33192 35207
rect 33140 35164 33192 35173
rect 35808 35164 35860 35216
rect 36176 35164 36228 35216
rect 37924 35164 37976 35216
rect 40776 35232 40828 35284
rect 40868 35207 40920 35216
rect 40868 35173 40877 35207
rect 40877 35173 40911 35207
rect 40911 35173 40920 35207
rect 41512 35207 41564 35216
rect 40868 35164 40920 35173
rect 41512 35173 41521 35207
rect 41521 35173 41555 35207
rect 41555 35173 41564 35207
rect 41512 35164 41564 35173
rect 42432 35164 42484 35216
rect 10968 35096 11020 35148
rect 12072 35096 12124 35148
rect 14464 35096 14516 35148
rect 17316 35139 17368 35148
rect 17316 35105 17325 35139
rect 17325 35105 17359 35139
rect 17359 35105 17368 35139
rect 17316 35096 17368 35105
rect 17776 35139 17828 35148
rect 17776 35105 17785 35139
rect 17785 35105 17819 35139
rect 17819 35105 17828 35139
rect 17776 35096 17828 35105
rect 24308 35139 24360 35148
rect 24308 35105 24317 35139
rect 24317 35105 24351 35139
rect 24351 35105 24360 35139
rect 24308 35096 24360 35105
rect 29000 35139 29052 35148
rect 29000 35105 29009 35139
rect 29009 35105 29043 35139
rect 29043 35105 29052 35139
rect 29000 35096 29052 35105
rect 29460 35139 29512 35148
rect 29460 35105 29469 35139
rect 29469 35105 29503 35139
rect 29503 35105 29512 35139
rect 29460 35096 29512 35105
rect 30472 35139 30524 35148
rect 30472 35105 30481 35139
rect 30481 35105 30515 35139
rect 30515 35105 30524 35139
rect 30472 35096 30524 35105
rect 34520 35139 34572 35148
rect 12440 35028 12492 35080
rect 15568 35071 15620 35080
rect 15568 35037 15577 35071
rect 15577 35037 15611 35071
rect 15611 35037 15620 35071
rect 15568 35028 15620 35037
rect 19432 35028 19484 35080
rect 20996 35071 21048 35080
rect 18052 34960 18104 35012
rect 20996 35037 21005 35071
rect 21005 35037 21039 35071
rect 21039 35037 21048 35071
rect 20996 35028 21048 35037
rect 19892 34960 19944 35012
rect 21180 34960 21232 35012
rect 22376 35028 22428 35080
rect 23664 35028 23716 35080
rect 27160 35071 27212 35080
rect 27160 35037 27169 35071
rect 27169 35037 27203 35071
rect 27203 35037 27212 35071
rect 27160 35028 27212 35037
rect 28724 35028 28776 35080
rect 30564 35028 30616 35080
rect 34520 35105 34529 35139
rect 34529 35105 34563 35139
rect 34563 35105 34572 35139
rect 34520 35096 34572 35105
rect 35440 35096 35492 35148
rect 35992 35096 36044 35148
rect 31208 35071 31260 35080
rect 31208 35037 31217 35071
rect 31217 35037 31251 35071
rect 31251 35037 31260 35071
rect 31208 35028 31260 35037
rect 33048 35071 33100 35080
rect 33048 35037 33057 35071
rect 33057 35037 33091 35071
rect 33091 35037 33100 35071
rect 33048 35028 33100 35037
rect 33416 35071 33468 35080
rect 33416 35037 33425 35071
rect 33425 35037 33459 35071
rect 33459 35037 33468 35071
rect 33416 35028 33468 35037
rect 38108 35028 38160 35080
rect 39580 35071 39632 35080
rect 39580 35037 39589 35071
rect 39589 35037 39623 35071
rect 39623 35037 39632 35071
rect 39580 35028 39632 35037
rect 41420 35071 41472 35080
rect 41420 35037 41429 35071
rect 41429 35037 41463 35071
rect 41463 35037 41472 35071
rect 41420 35028 41472 35037
rect 27252 34960 27304 35012
rect 32404 35003 32456 35012
rect 32404 34969 32413 35003
rect 32413 34969 32447 35003
rect 32447 34969 32456 35003
rect 37188 35003 37240 35012
rect 32404 34960 32456 34969
rect 37188 34969 37197 35003
rect 37197 34969 37231 35003
rect 37231 34969 37240 35003
rect 42156 35096 42208 35148
rect 37188 34960 37240 34969
rect 16488 34935 16540 34944
rect 16488 34901 16497 34935
rect 16497 34901 16531 34935
rect 16531 34901 16540 34935
rect 16488 34892 16540 34901
rect 23848 34935 23900 34944
rect 23848 34901 23857 34935
rect 23857 34901 23891 34935
rect 23891 34901 23900 34935
rect 23848 34892 23900 34901
rect 28172 34935 28224 34944
rect 28172 34901 28181 34935
rect 28181 34901 28215 34935
rect 28215 34901 28224 34935
rect 28172 34892 28224 34901
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 11980 34688 12032 34740
rect 12440 34552 12492 34604
rect 13452 34688 13504 34740
rect 14096 34731 14148 34740
rect 14096 34697 14105 34731
rect 14105 34697 14139 34731
rect 14139 34697 14148 34731
rect 14096 34688 14148 34697
rect 14464 34731 14516 34740
rect 14464 34697 14473 34731
rect 14473 34697 14507 34731
rect 14507 34697 14516 34731
rect 14464 34688 14516 34697
rect 14556 34688 14608 34740
rect 17776 34688 17828 34740
rect 18604 34731 18656 34740
rect 18604 34697 18613 34731
rect 18613 34697 18647 34731
rect 18647 34697 18656 34731
rect 18604 34688 18656 34697
rect 18788 34688 18840 34740
rect 21088 34688 21140 34740
rect 22376 34688 22428 34740
rect 24676 34688 24728 34740
rect 25228 34731 25280 34740
rect 25228 34697 25237 34731
rect 25237 34697 25271 34731
rect 25271 34697 25280 34731
rect 25228 34688 25280 34697
rect 13360 34663 13412 34672
rect 13360 34629 13369 34663
rect 13369 34629 13403 34663
rect 13403 34629 13412 34663
rect 15660 34663 15712 34672
rect 13360 34620 13412 34629
rect 15660 34629 15669 34663
rect 15669 34629 15703 34663
rect 15703 34629 15712 34663
rect 15660 34620 15712 34629
rect 16764 34663 16816 34672
rect 16764 34629 16773 34663
rect 16773 34629 16807 34663
rect 16807 34629 16816 34663
rect 16764 34620 16816 34629
rect 17316 34620 17368 34672
rect 28172 34688 28224 34740
rect 14648 34595 14700 34604
rect 14648 34561 14657 34595
rect 14657 34561 14691 34595
rect 14691 34561 14700 34595
rect 14648 34552 14700 34561
rect 15384 34552 15436 34604
rect 16672 34552 16724 34604
rect 17776 34595 17828 34604
rect 17776 34561 17785 34595
rect 17785 34561 17819 34595
rect 17819 34561 17828 34595
rect 17776 34552 17828 34561
rect 19156 34552 19208 34604
rect 19432 34552 19484 34604
rect 10876 34484 10928 34536
rect 13084 34484 13136 34536
rect 14096 34484 14148 34536
rect 18604 34484 18656 34536
rect 20076 34484 20128 34536
rect 28356 34620 28408 34672
rect 29000 34663 29052 34672
rect 29000 34629 29009 34663
rect 29009 34629 29043 34663
rect 29043 34629 29052 34663
rect 32588 34688 32640 34740
rect 33048 34688 33100 34740
rect 38108 34731 38160 34740
rect 29000 34620 29052 34629
rect 24768 34552 24820 34604
rect 25412 34595 25464 34604
rect 25412 34561 25421 34595
rect 25421 34561 25455 34595
rect 25455 34561 25464 34595
rect 25412 34552 25464 34561
rect 26424 34552 26476 34604
rect 27344 34552 27396 34604
rect 27528 34552 27580 34604
rect 28540 34552 28592 34604
rect 29460 34552 29512 34604
rect 31300 34595 31352 34604
rect 31300 34561 31309 34595
rect 31309 34561 31343 34595
rect 31343 34561 31352 34595
rect 31300 34552 31352 34561
rect 23848 34484 23900 34536
rect 24952 34484 25004 34536
rect 14464 34416 14516 34468
rect 10600 34348 10652 34400
rect 12900 34348 12952 34400
rect 13912 34348 13964 34400
rect 16488 34416 16540 34468
rect 19248 34459 19300 34468
rect 19248 34425 19257 34459
rect 19257 34425 19291 34459
rect 19291 34425 19300 34459
rect 19248 34416 19300 34425
rect 19432 34416 19484 34468
rect 22008 34459 22060 34468
rect 22008 34425 22017 34459
rect 22017 34425 22051 34459
rect 22051 34425 22060 34459
rect 22008 34416 22060 34425
rect 22100 34459 22152 34468
rect 22100 34425 22109 34459
rect 22109 34425 22143 34459
rect 22143 34425 22152 34459
rect 22100 34416 22152 34425
rect 16580 34348 16632 34400
rect 17316 34391 17368 34400
rect 17316 34357 17325 34391
rect 17325 34357 17359 34391
rect 17359 34357 17368 34391
rect 17316 34348 17368 34357
rect 17776 34348 17828 34400
rect 19340 34348 19392 34400
rect 25228 34348 25280 34400
rect 26976 34391 27028 34400
rect 26976 34357 26985 34391
rect 26985 34357 27019 34391
rect 27019 34357 27028 34391
rect 27344 34459 27396 34468
rect 27344 34425 27353 34459
rect 27353 34425 27387 34459
rect 27387 34425 27396 34459
rect 27344 34416 27396 34425
rect 27712 34416 27764 34468
rect 30472 34459 30524 34468
rect 30472 34425 30481 34459
rect 30481 34425 30515 34459
rect 30515 34425 30524 34459
rect 30472 34416 30524 34425
rect 26976 34348 27028 34357
rect 29828 34391 29880 34400
rect 29828 34357 29837 34391
rect 29837 34357 29871 34391
rect 29871 34357 29880 34391
rect 29828 34348 29880 34357
rect 30748 34459 30800 34468
rect 30748 34425 30757 34459
rect 30757 34425 30791 34459
rect 30791 34425 30800 34459
rect 30748 34416 30800 34425
rect 31760 34552 31812 34604
rect 32404 34595 32456 34604
rect 32404 34561 32413 34595
rect 32413 34561 32447 34595
rect 32447 34561 32456 34595
rect 32404 34552 32456 34561
rect 36636 34620 36688 34672
rect 38108 34697 38117 34731
rect 38117 34697 38151 34731
rect 38151 34697 38160 34731
rect 38108 34688 38160 34697
rect 41512 34688 41564 34740
rect 41696 34688 41748 34740
rect 41972 34620 42024 34672
rect 35532 34595 35584 34604
rect 35532 34561 35541 34595
rect 35541 34561 35575 34595
rect 35575 34561 35584 34595
rect 35532 34552 35584 34561
rect 36452 34552 36504 34604
rect 36912 34595 36964 34604
rect 36912 34561 36921 34595
rect 36921 34561 36955 34595
rect 36955 34561 36964 34595
rect 36912 34552 36964 34561
rect 37924 34552 37976 34604
rect 39580 34595 39632 34604
rect 39580 34561 39589 34595
rect 39589 34561 39623 34595
rect 39623 34561 39632 34595
rect 39580 34552 39632 34561
rect 42064 34552 42116 34604
rect 35440 34527 35492 34536
rect 35440 34493 35449 34527
rect 35449 34493 35483 34527
rect 35483 34493 35492 34527
rect 35440 34484 35492 34493
rect 39304 34527 39356 34536
rect 32128 34391 32180 34400
rect 32128 34357 32137 34391
rect 32137 34357 32171 34391
rect 32171 34357 32180 34391
rect 32588 34416 32640 34468
rect 34520 34416 34572 34468
rect 35900 34416 35952 34468
rect 32128 34348 32180 34357
rect 33140 34348 33192 34400
rect 35992 34348 36044 34400
rect 36728 34459 36780 34468
rect 36728 34425 36737 34459
rect 36737 34425 36771 34459
rect 36771 34425 36780 34459
rect 38660 34459 38712 34468
rect 36728 34416 36780 34425
rect 38660 34425 38669 34459
rect 38669 34425 38703 34459
rect 38703 34425 38712 34459
rect 39304 34493 39313 34527
rect 39313 34493 39347 34527
rect 39347 34493 39356 34527
rect 39304 34484 39356 34493
rect 38660 34416 38712 34425
rect 42432 34484 42484 34536
rect 37188 34348 37240 34400
rect 40132 34348 40184 34400
rect 42248 34391 42300 34400
rect 42248 34357 42257 34391
rect 42257 34357 42291 34391
rect 42291 34357 42300 34391
rect 42248 34348 42300 34357
rect 42340 34348 42392 34400
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 10968 34187 11020 34196
rect 10968 34153 10977 34187
rect 10977 34153 11011 34187
rect 11011 34153 11020 34187
rect 10968 34144 11020 34153
rect 14648 34187 14700 34196
rect 14648 34153 14657 34187
rect 14657 34153 14691 34187
rect 14691 34153 14700 34187
rect 14648 34144 14700 34153
rect 10876 34076 10928 34128
rect 15568 34144 15620 34196
rect 16672 34187 16724 34196
rect 16672 34153 16681 34187
rect 16681 34153 16715 34187
rect 16715 34153 16724 34187
rect 16672 34144 16724 34153
rect 19248 34187 19300 34196
rect 19248 34153 19257 34187
rect 19257 34153 19291 34187
rect 19291 34153 19300 34187
rect 19248 34144 19300 34153
rect 19340 34144 19392 34196
rect 20076 34187 20128 34196
rect 20076 34153 20085 34187
rect 20085 34153 20119 34187
rect 20119 34153 20128 34187
rect 20076 34144 20128 34153
rect 20996 34144 21048 34196
rect 21824 34187 21876 34196
rect 21824 34153 21833 34187
rect 21833 34153 21867 34187
rect 21867 34153 21876 34187
rect 21824 34144 21876 34153
rect 22100 34144 22152 34196
rect 24308 34187 24360 34196
rect 24308 34153 24317 34187
rect 24317 34153 24351 34187
rect 24351 34153 24360 34187
rect 24308 34144 24360 34153
rect 27160 34144 27212 34196
rect 30748 34144 30800 34196
rect 33048 34144 33100 34196
rect 36728 34144 36780 34196
rect 41420 34187 41472 34196
rect 41420 34153 41429 34187
rect 41429 34153 41463 34187
rect 41463 34153 41472 34187
rect 41420 34144 41472 34153
rect 42340 34144 42392 34196
rect 15476 34119 15528 34128
rect 15476 34085 15485 34119
rect 15485 34085 15519 34119
rect 15519 34085 15528 34119
rect 15476 34076 15528 34085
rect 26976 34076 27028 34128
rect 27344 34119 27396 34128
rect 27344 34085 27353 34119
rect 27353 34085 27387 34119
rect 27387 34085 27396 34119
rect 27344 34076 27396 34085
rect 29644 34076 29696 34128
rect 30564 34076 30616 34128
rect 32312 34076 32364 34128
rect 36544 34076 36596 34128
rect 37924 34076 37976 34128
rect 11888 34051 11940 34060
rect 11888 34017 11897 34051
rect 11897 34017 11931 34051
rect 11931 34017 11940 34051
rect 11888 34008 11940 34017
rect 13728 34051 13780 34060
rect 13728 34017 13737 34051
rect 13737 34017 13771 34051
rect 13771 34017 13780 34051
rect 13728 34008 13780 34017
rect 14096 34008 14148 34060
rect 14556 34008 14608 34060
rect 17500 34008 17552 34060
rect 18052 34008 18104 34060
rect 15384 33983 15436 33992
rect 15384 33949 15393 33983
rect 15393 33949 15427 33983
rect 15427 33949 15436 33983
rect 15384 33940 15436 33949
rect 18880 33983 18932 33992
rect 18880 33949 18889 33983
rect 18889 33949 18923 33983
rect 18923 33949 18932 33983
rect 18880 33940 18932 33949
rect 21456 33983 21508 33992
rect 21456 33949 21465 33983
rect 21465 33949 21499 33983
rect 21499 33949 21508 33983
rect 21456 33940 21508 33949
rect 24952 34008 25004 34060
rect 25688 34008 25740 34060
rect 31208 34008 31260 34060
rect 33876 34008 33928 34060
rect 35624 34008 35676 34060
rect 38200 34076 38252 34128
rect 38660 34076 38712 34128
rect 39028 34051 39080 34060
rect 39028 34017 39037 34051
rect 39037 34017 39071 34051
rect 39071 34017 39080 34051
rect 39028 34008 39080 34017
rect 39396 34008 39448 34060
rect 40316 34008 40368 34060
rect 41696 34051 41748 34060
rect 41696 34017 41705 34051
rect 41705 34017 41739 34051
rect 41739 34017 41748 34051
rect 41696 34008 41748 34017
rect 42156 34051 42208 34060
rect 42156 34017 42165 34051
rect 42165 34017 42199 34051
rect 42199 34017 42208 34051
rect 42156 34008 42208 34017
rect 25596 33983 25648 33992
rect 25596 33949 25605 33983
rect 25605 33949 25639 33983
rect 25639 33949 25648 33983
rect 25596 33940 25648 33949
rect 27620 33940 27672 33992
rect 29460 33983 29512 33992
rect 29460 33949 29469 33983
rect 29469 33949 29503 33983
rect 29503 33949 29512 33983
rect 29460 33940 29512 33949
rect 35532 33983 35584 33992
rect 35532 33949 35541 33983
rect 35541 33949 35575 33983
rect 35575 33949 35584 33983
rect 35532 33940 35584 33949
rect 38476 33940 38528 33992
rect 39764 33983 39816 33992
rect 39764 33949 39773 33983
rect 39773 33949 39807 33983
rect 39807 33949 39816 33983
rect 39764 33940 39816 33949
rect 42616 33940 42668 33992
rect 15936 33915 15988 33924
rect 15936 33881 15945 33915
rect 15945 33881 15979 33915
rect 15979 33881 15988 33915
rect 15936 33872 15988 33881
rect 16764 33872 16816 33924
rect 22192 33872 22244 33924
rect 23296 33872 23348 33924
rect 27712 33872 27764 33924
rect 27804 33915 27856 33924
rect 27804 33881 27813 33915
rect 27813 33881 27847 33915
rect 27847 33881 27856 33915
rect 27804 33872 27856 33881
rect 31760 33872 31812 33924
rect 33324 33872 33376 33924
rect 34520 33915 34572 33924
rect 34520 33881 34529 33915
rect 34529 33881 34563 33915
rect 34563 33881 34572 33915
rect 34520 33872 34572 33881
rect 35440 33872 35492 33924
rect 39304 33872 39356 33924
rect 12532 33804 12584 33856
rect 17868 33804 17920 33856
rect 18420 33847 18472 33856
rect 18420 33813 18429 33847
rect 18429 33813 18463 33847
rect 18463 33813 18472 33847
rect 18420 33804 18472 33813
rect 22928 33804 22980 33856
rect 27528 33804 27580 33856
rect 33048 33847 33100 33856
rect 33048 33813 33057 33847
rect 33057 33813 33091 33847
rect 33091 33813 33100 33847
rect 33048 33804 33100 33813
rect 37924 33804 37976 33856
rect 40776 33804 40828 33856
rect 43628 33847 43680 33856
rect 43628 33813 43637 33847
rect 43637 33813 43671 33847
rect 43671 33813 43680 33847
rect 43628 33804 43680 33813
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 10508 33643 10560 33652
rect 10508 33609 10517 33643
rect 10517 33609 10551 33643
rect 10551 33609 10560 33643
rect 10508 33600 10560 33609
rect 11888 33643 11940 33652
rect 11888 33609 11897 33643
rect 11897 33609 11931 33643
rect 11931 33609 11940 33643
rect 11888 33600 11940 33609
rect 13728 33643 13780 33652
rect 13728 33609 13737 33643
rect 13737 33609 13771 33643
rect 13771 33609 13780 33643
rect 14096 33643 14148 33652
rect 13728 33600 13780 33609
rect 14096 33609 14105 33643
rect 14105 33609 14139 33643
rect 14139 33609 14148 33643
rect 14096 33600 14148 33609
rect 15384 33600 15436 33652
rect 16028 33643 16080 33652
rect 16028 33609 16037 33643
rect 16037 33609 16071 33643
rect 16071 33609 16080 33643
rect 16028 33600 16080 33609
rect 17500 33643 17552 33652
rect 17500 33609 17509 33643
rect 17509 33609 17543 33643
rect 17543 33609 17552 33643
rect 17500 33600 17552 33609
rect 17960 33600 18012 33652
rect 19432 33643 19484 33652
rect 19432 33609 19441 33643
rect 19441 33609 19475 33643
rect 19475 33609 19484 33643
rect 19432 33600 19484 33609
rect 20352 33600 20404 33652
rect 21824 33600 21876 33652
rect 22008 33600 22060 33652
rect 25688 33600 25740 33652
rect 27344 33643 27396 33652
rect 27344 33609 27353 33643
rect 27353 33609 27387 33643
rect 27387 33609 27396 33643
rect 27344 33600 27396 33609
rect 27620 33643 27672 33652
rect 27620 33609 27629 33643
rect 27629 33609 27663 33643
rect 27663 33609 27672 33643
rect 27620 33600 27672 33609
rect 29644 33600 29696 33652
rect 30380 33600 30432 33652
rect 32128 33600 32180 33652
rect 12532 33507 12584 33516
rect 12532 33473 12541 33507
rect 12541 33473 12575 33507
rect 12575 33473 12584 33507
rect 12532 33464 12584 33473
rect 13912 33464 13964 33516
rect 14740 33507 14792 33516
rect 14740 33473 14749 33507
rect 14749 33473 14783 33507
rect 14783 33473 14792 33507
rect 14740 33464 14792 33473
rect 18880 33464 18932 33516
rect 21456 33464 21508 33516
rect 27804 33532 27856 33584
rect 24676 33464 24728 33516
rect 10508 33396 10560 33448
rect 10968 33396 11020 33448
rect 17960 33396 18012 33448
rect 18328 33439 18380 33448
rect 18328 33405 18337 33439
rect 18337 33405 18371 33439
rect 18371 33405 18380 33439
rect 18328 33396 18380 33405
rect 18420 33396 18472 33448
rect 21180 33439 21232 33448
rect 21180 33405 21189 33439
rect 21189 33405 21223 33439
rect 21223 33405 21232 33439
rect 21180 33396 21232 33405
rect 11428 33328 11480 33380
rect 12716 33328 12768 33380
rect 13176 33371 13228 33380
rect 13176 33337 13185 33371
rect 13185 33337 13219 33371
rect 13219 33337 13228 33371
rect 13176 33328 13228 33337
rect 15384 33371 15436 33380
rect 14556 33303 14608 33312
rect 14556 33269 14565 33303
rect 14565 33269 14599 33303
rect 14599 33269 14608 33303
rect 15384 33337 15393 33371
rect 15393 33337 15427 33371
rect 15427 33337 15436 33371
rect 15384 33328 15436 33337
rect 19248 33328 19300 33380
rect 21732 33396 21784 33448
rect 22928 33439 22980 33448
rect 22928 33405 22937 33439
rect 22937 33405 22971 33439
rect 22971 33405 22980 33439
rect 22928 33396 22980 33405
rect 25596 33464 25648 33516
rect 26056 33507 26108 33516
rect 26056 33473 26065 33507
rect 26065 33473 26099 33507
rect 26099 33473 26108 33507
rect 26056 33464 26108 33473
rect 25228 33371 25280 33380
rect 14556 33260 14608 33269
rect 14924 33260 14976 33312
rect 15476 33260 15528 33312
rect 16948 33260 17000 33312
rect 24400 33303 24452 33312
rect 24400 33269 24409 33303
rect 24409 33269 24443 33303
rect 24443 33269 24452 33303
rect 25228 33337 25237 33371
rect 25237 33337 25271 33371
rect 25271 33337 25280 33371
rect 25228 33328 25280 33337
rect 27528 33396 27580 33448
rect 28264 33439 28316 33448
rect 28264 33405 28273 33439
rect 28273 33405 28307 33439
rect 28307 33405 28316 33439
rect 28264 33396 28316 33405
rect 28632 33396 28684 33448
rect 30564 33396 30616 33448
rect 31116 33439 31168 33448
rect 31116 33405 31125 33439
rect 31125 33405 31159 33439
rect 31159 33405 31168 33439
rect 31116 33396 31168 33405
rect 33048 33600 33100 33652
rect 33876 33643 33928 33652
rect 33876 33609 33885 33643
rect 33885 33609 33919 33643
rect 33919 33609 33928 33643
rect 33876 33600 33928 33609
rect 35532 33600 35584 33652
rect 38200 33600 38252 33652
rect 39028 33600 39080 33652
rect 40040 33600 40092 33652
rect 40316 33643 40368 33652
rect 40316 33609 40325 33643
rect 40325 33609 40359 33643
rect 40359 33609 40368 33643
rect 40316 33600 40368 33609
rect 41512 33600 41564 33652
rect 41696 33643 41748 33652
rect 41696 33609 41705 33643
rect 41705 33609 41739 33643
rect 41739 33609 41748 33643
rect 41696 33600 41748 33609
rect 42156 33643 42208 33652
rect 42156 33609 42165 33643
rect 42165 33609 42199 33643
rect 42199 33609 42208 33643
rect 42156 33600 42208 33609
rect 37464 33532 37516 33584
rect 33324 33507 33376 33516
rect 33324 33473 33333 33507
rect 33333 33473 33367 33507
rect 33367 33473 33376 33507
rect 33324 33464 33376 33473
rect 36084 33464 36136 33516
rect 32312 33371 32364 33380
rect 32312 33337 32321 33371
rect 32321 33337 32355 33371
rect 32355 33337 32364 33371
rect 32312 33328 32364 33337
rect 24400 33260 24452 33269
rect 29460 33260 29512 33312
rect 36452 33396 36504 33448
rect 37924 33507 37976 33516
rect 37924 33473 37933 33507
rect 37933 33473 37967 33507
rect 37967 33473 37976 33507
rect 37924 33464 37976 33473
rect 38292 33464 38344 33516
rect 44180 33532 44232 33584
rect 40776 33507 40828 33516
rect 40776 33473 40785 33507
rect 40785 33473 40819 33507
rect 40819 33473 40828 33507
rect 40776 33464 40828 33473
rect 43628 33507 43680 33516
rect 43628 33473 43637 33507
rect 43637 33473 43671 33507
rect 43671 33473 43680 33507
rect 43628 33464 43680 33473
rect 37648 33396 37700 33448
rect 39212 33396 39264 33448
rect 41972 33396 42024 33448
rect 32772 33328 32824 33380
rect 34612 33328 34664 33380
rect 36544 33260 36596 33312
rect 40868 33371 40920 33380
rect 40868 33337 40877 33371
rect 40877 33337 40911 33371
rect 40911 33337 40920 33371
rect 40868 33328 40920 33337
rect 38108 33260 38160 33312
rect 40500 33260 40552 33312
rect 44088 33328 44140 33380
rect 44272 33371 44324 33380
rect 44272 33337 44281 33371
rect 44281 33337 44315 33371
rect 44315 33337 44324 33371
rect 44272 33328 44324 33337
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 14740 33099 14792 33108
rect 14740 33065 14749 33099
rect 14749 33065 14783 33099
rect 14783 33065 14792 33099
rect 14740 33056 14792 33065
rect 16028 33056 16080 33108
rect 18052 33099 18104 33108
rect 18052 33065 18061 33099
rect 18061 33065 18095 33099
rect 18095 33065 18104 33099
rect 18052 33056 18104 33065
rect 24400 33099 24452 33108
rect 24400 33065 24409 33099
rect 24409 33065 24443 33099
rect 24443 33065 24452 33099
rect 24400 33056 24452 33065
rect 24952 33099 25004 33108
rect 24952 33065 24961 33099
rect 24961 33065 24995 33099
rect 24995 33065 25004 33099
rect 24952 33056 25004 33065
rect 26056 33099 26108 33108
rect 26056 33065 26065 33099
rect 26065 33065 26099 33099
rect 26099 33065 26108 33099
rect 26056 33056 26108 33065
rect 32220 33099 32272 33108
rect 32220 33065 32229 33099
rect 32229 33065 32263 33099
rect 32263 33065 32272 33099
rect 32220 33056 32272 33065
rect 33232 33099 33284 33108
rect 33232 33065 33241 33099
rect 33241 33065 33275 33099
rect 33275 33065 33284 33099
rect 33232 33056 33284 33065
rect 34796 33056 34848 33108
rect 36544 33056 36596 33108
rect 37832 33056 37884 33108
rect 11980 32988 12032 33040
rect 12900 32988 12952 33040
rect 13452 33031 13504 33040
rect 13452 32997 13461 33031
rect 13461 32997 13495 33031
rect 13495 32997 13504 33031
rect 13452 32988 13504 32997
rect 13544 33031 13596 33040
rect 13544 32997 13553 33031
rect 13553 32997 13587 33031
rect 13587 32997 13596 33031
rect 13544 32988 13596 32997
rect 14556 32988 14608 33040
rect 17500 32988 17552 33040
rect 19248 32988 19300 33040
rect 15752 32920 15804 32972
rect 19064 32963 19116 32972
rect 19064 32929 19073 32963
rect 19073 32929 19107 32963
rect 19107 32929 19116 32963
rect 19064 32920 19116 32929
rect 20076 32988 20128 33040
rect 20352 32988 20404 33040
rect 23112 32988 23164 33040
rect 24768 32988 24820 33040
rect 26424 32988 26476 33040
rect 28816 33031 28868 33040
rect 28816 32997 28825 33031
rect 28825 32997 28859 33031
rect 28859 32997 28868 33031
rect 28816 32988 28868 32997
rect 29828 32988 29880 33040
rect 34336 32988 34388 33040
rect 39396 33056 39448 33108
rect 42064 33056 42116 33108
rect 43628 33056 43680 33108
rect 44088 33056 44140 33108
rect 38568 32988 38620 33040
rect 38936 32988 38988 33040
rect 39856 32988 39908 33040
rect 40132 32988 40184 33040
rect 40868 32988 40920 33040
rect 22284 32920 22336 32972
rect 22468 32963 22520 32972
rect 22468 32929 22477 32963
rect 22477 32929 22511 32963
rect 22511 32929 22520 32963
rect 22468 32920 22520 32929
rect 25228 32920 25280 32972
rect 28080 32963 28132 32972
rect 28080 32929 28089 32963
rect 28089 32929 28123 32963
rect 28123 32929 28132 32963
rect 28080 32920 28132 32929
rect 28264 32920 28316 32972
rect 30472 32963 30524 32972
rect 10140 32895 10192 32904
rect 10140 32861 10149 32895
rect 10149 32861 10183 32895
rect 10183 32861 10192 32895
rect 10140 32852 10192 32861
rect 11428 32852 11480 32904
rect 13728 32895 13780 32904
rect 13728 32861 13737 32895
rect 13737 32861 13771 32895
rect 13771 32861 13780 32895
rect 13728 32852 13780 32861
rect 17040 32852 17092 32904
rect 23296 32852 23348 32904
rect 26884 32895 26936 32904
rect 26332 32784 26384 32836
rect 26884 32861 26893 32895
rect 26893 32861 26927 32895
rect 26927 32861 26936 32895
rect 26884 32852 26936 32861
rect 28632 32852 28684 32904
rect 27436 32784 27488 32836
rect 30472 32929 30481 32963
rect 30481 32929 30515 32963
rect 30515 32929 30524 32963
rect 30472 32920 30524 32929
rect 30748 32963 30800 32972
rect 30748 32929 30757 32963
rect 30757 32929 30791 32963
rect 30791 32929 30800 32963
rect 30748 32920 30800 32929
rect 31116 32920 31168 32972
rect 32128 32920 32180 32972
rect 32496 32920 32548 32972
rect 32680 32963 32732 32972
rect 32680 32929 32689 32963
rect 32689 32929 32723 32963
rect 32723 32929 32732 32963
rect 32680 32920 32732 32929
rect 36268 32963 36320 32972
rect 36268 32929 36277 32963
rect 36277 32929 36311 32963
rect 36311 32929 36320 32963
rect 36268 32920 36320 32929
rect 36544 32963 36596 32972
rect 36544 32929 36553 32963
rect 36553 32929 36587 32963
rect 36587 32929 36596 32963
rect 36544 32920 36596 32929
rect 39396 32920 39448 32972
rect 42616 32920 42668 32972
rect 32312 32852 32364 32904
rect 35992 32852 36044 32904
rect 36728 32852 36780 32904
rect 37188 32852 37240 32904
rect 39764 32895 39816 32904
rect 39764 32861 39773 32895
rect 39773 32861 39807 32895
rect 39807 32861 39816 32895
rect 39764 32852 39816 32861
rect 41604 32895 41656 32904
rect 41604 32861 41613 32895
rect 41613 32861 41647 32895
rect 41647 32861 41656 32895
rect 41604 32852 41656 32861
rect 42984 32852 43036 32904
rect 45100 32895 45152 32904
rect 45100 32861 45109 32895
rect 45109 32861 45143 32895
rect 45143 32861 45152 32895
rect 45100 32852 45152 32861
rect 32404 32784 32456 32836
rect 38108 32784 38160 32836
rect 38568 32784 38620 32836
rect 10692 32759 10744 32768
rect 10692 32725 10701 32759
rect 10701 32725 10735 32759
rect 10735 32725 10744 32759
rect 10692 32716 10744 32725
rect 10968 32716 11020 32768
rect 12532 32759 12584 32768
rect 12532 32725 12541 32759
rect 12541 32725 12575 32759
rect 12575 32725 12584 32759
rect 12532 32716 12584 32725
rect 17684 32759 17736 32768
rect 17684 32725 17693 32759
rect 17693 32725 17727 32759
rect 17727 32725 17736 32759
rect 17684 32716 17736 32725
rect 18328 32759 18380 32768
rect 18328 32725 18337 32759
rect 18337 32725 18371 32759
rect 18371 32725 18380 32759
rect 18328 32716 18380 32725
rect 21548 32716 21600 32768
rect 23572 32716 23624 32768
rect 25688 32759 25740 32768
rect 25688 32725 25697 32759
rect 25697 32725 25731 32759
rect 25731 32725 25740 32759
rect 25688 32716 25740 32725
rect 27988 32716 28040 32768
rect 28264 32759 28316 32768
rect 28264 32725 28288 32759
rect 28288 32725 28316 32759
rect 28264 32716 28316 32725
rect 28448 32716 28500 32768
rect 30012 32716 30064 32768
rect 31576 32759 31628 32768
rect 31576 32725 31585 32759
rect 31585 32725 31619 32759
rect 31619 32725 31628 32759
rect 31576 32716 31628 32725
rect 36084 32716 36136 32768
rect 37556 32716 37608 32768
rect 42156 32784 42208 32836
rect 40868 32716 40920 32768
rect 41052 32716 41104 32768
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 10140 32512 10192 32564
rect 10508 32308 10560 32360
rect 11980 32444 12032 32496
rect 13452 32512 13504 32564
rect 17500 32555 17552 32564
rect 17500 32521 17509 32555
rect 17509 32521 17543 32555
rect 17543 32521 17552 32555
rect 17500 32512 17552 32521
rect 20352 32512 20404 32564
rect 21732 32555 21784 32564
rect 21732 32521 21741 32555
rect 21741 32521 21775 32555
rect 21775 32521 21784 32555
rect 21732 32512 21784 32521
rect 22468 32512 22520 32564
rect 13544 32487 13596 32496
rect 13544 32453 13553 32487
rect 13553 32453 13587 32487
rect 13587 32453 13596 32487
rect 13544 32444 13596 32453
rect 21548 32487 21600 32496
rect 13176 32419 13228 32428
rect 13176 32385 13185 32419
rect 13185 32385 13219 32419
rect 13219 32385 13228 32419
rect 13176 32376 13228 32385
rect 15384 32419 15436 32428
rect 15384 32385 15393 32419
rect 15393 32385 15427 32419
rect 15427 32385 15436 32419
rect 15384 32376 15436 32385
rect 15844 32376 15896 32428
rect 16488 32419 16540 32428
rect 16488 32385 16497 32419
rect 16497 32385 16531 32419
rect 16531 32385 16540 32419
rect 16488 32376 16540 32385
rect 17776 32376 17828 32428
rect 18788 32376 18840 32428
rect 19892 32376 19944 32428
rect 21548 32453 21557 32487
rect 21557 32453 21591 32487
rect 21591 32453 21600 32487
rect 21548 32444 21600 32453
rect 20996 32376 21048 32428
rect 18880 32308 18932 32360
rect 20260 32351 20312 32360
rect 20260 32317 20269 32351
rect 20269 32317 20303 32351
rect 20303 32317 20312 32351
rect 20260 32308 20312 32317
rect 21732 32308 21784 32360
rect 24032 32512 24084 32564
rect 23112 32487 23164 32496
rect 23112 32453 23121 32487
rect 23121 32453 23155 32487
rect 23155 32453 23164 32487
rect 23112 32444 23164 32453
rect 23940 32487 23992 32496
rect 23940 32453 23949 32487
rect 23949 32453 23983 32487
rect 23983 32453 23992 32487
rect 23940 32444 23992 32453
rect 22744 32376 22796 32428
rect 24952 32512 25004 32564
rect 27988 32512 28040 32564
rect 32680 32512 32732 32564
rect 34060 32512 34112 32564
rect 34336 32512 34388 32564
rect 37188 32555 37240 32564
rect 37188 32521 37197 32555
rect 37197 32521 37231 32555
rect 37231 32521 37240 32555
rect 37188 32512 37240 32521
rect 37832 32555 37884 32564
rect 37832 32521 37841 32555
rect 37841 32521 37875 32555
rect 37875 32521 37884 32555
rect 37832 32512 37884 32521
rect 39764 32512 39816 32564
rect 42616 32555 42668 32564
rect 42616 32521 42625 32555
rect 42625 32521 42659 32555
rect 42659 32521 42668 32555
rect 42616 32512 42668 32521
rect 43628 32555 43680 32564
rect 25136 32376 25188 32428
rect 25688 32376 25740 32428
rect 27436 32376 27488 32428
rect 12624 32283 12676 32292
rect 12624 32249 12633 32283
rect 12633 32249 12667 32283
rect 12667 32249 12676 32283
rect 12624 32240 12676 32249
rect 13544 32240 13596 32292
rect 14740 32283 14792 32292
rect 14740 32249 14749 32283
rect 14749 32249 14783 32283
rect 14783 32249 14792 32283
rect 14740 32240 14792 32249
rect 14832 32283 14884 32292
rect 14832 32249 14841 32283
rect 14841 32249 14875 32283
rect 14875 32249 14884 32283
rect 14832 32240 14884 32249
rect 17132 32283 17184 32292
rect 15752 32215 15804 32224
rect 15752 32181 15761 32215
rect 15761 32181 15795 32215
rect 15795 32181 15804 32215
rect 15752 32172 15804 32181
rect 17132 32249 17141 32283
rect 17141 32249 17175 32283
rect 17175 32249 17184 32283
rect 17132 32240 17184 32249
rect 17684 32240 17736 32292
rect 17224 32172 17276 32224
rect 17868 32240 17920 32292
rect 18144 32283 18196 32292
rect 18144 32249 18153 32283
rect 18153 32249 18187 32283
rect 18187 32249 18196 32283
rect 18144 32240 18196 32249
rect 19064 32172 19116 32224
rect 19984 32172 20036 32224
rect 20996 32172 21048 32224
rect 23112 32240 23164 32292
rect 26608 32240 26660 32292
rect 28264 32308 28316 32360
rect 39856 32487 39908 32496
rect 39856 32453 39865 32487
rect 39865 32453 39899 32487
rect 39899 32453 39908 32487
rect 43628 32521 43637 32555
rect 43637 32521 43671 32555
rect 43671 32521 43680 32555
rect 43628 32512 43680 32521
rect 44364 32487 44416 32496
rect 39856 32444 39908 32453
rect 44364 32453 44373 32487
rect 44373 32453 44407 32487
rect 44407 32453 44416 32487
rect 44364 32444 44416 32453
rect 31576 32376 31628 32428
rect 31300 32351 31352 32360
rect 31300 32317 31309 32351
rect 31309 32317 31343 32351
rect 31343 32317 31352 32351
rect 32772 32376 32824 32428
rect 34796 32376 34848 32428
rect 35440 32419 35492 32428
rect 35440 32385 35449 32419
rect 35449 32385 35483 32419
rect 35483 32385 35492 32419
rect 35440 32376 35492 32385
rect 38476 32419 38528 32428
rect 38476 32385 38485 32419
rect 38485 32385 38519 32419
rect 38519 32385 38528 32419
rect 38476 32376 38528 32385
rect 41144 32376 41196 32428
rect 45100 32512 45152 32564
rect 31300 32308 31352 32317
rect 31944 32351 31996 32360
rect 31944 32317 31953 32351
rect 31953 32317 31987 32351
rect 31987 32317 31996 32351
rect 31944 32308 31996 32317
rect 32680 32308 32732 32360
rect 27528 32240 27580 32292
rect 29920 32240 29972 32292
rect 30012 32283 30064 32292
rect 30012 32249 30021 32283
rect 30021 32249 30055 32283
rect 30055 32249 30064 32283
rect 30564 32283 30616 32292
rect 30012 32240 30064 32249
rect 30564 32249 30573 32283
rect 30573 32249 30607 32283
rect 30607 32249 30616 32283
rect 30564 32240 30616 32249
rect 32128 32283 32180 32292
rect 32128 32249 32137 32283
rect 32137 32249 32171 32283
rect 32171 32249 32180 32283
rect 32128 32240 32180 32249
rect 21364 32172 21416 32224
rect 22284 32215 22336 32224
rect 22284 32181 22293 32215
rect 22293 32181 22327 32215
rect 22327 32181 22336 32215
rect 22284 32172 22336 32181
rect 24768 32172 24820 32224
rect 26424 32172 26476 32224
rect 26700 32215 26752 32224
rect 26700 32181 26709 32215
rect 26709 32181 26743 32215
rect 26743 32181 26752 32215
rect 26700 32172 26752 32181
rect 27436 32215 27488 32224
rect 27436 32181 27445 32215
rect 27445 32181 27479 32215
rect 27479 32181 27488 32215
rect 27436 32172 27488 32181
rect 27804 32172 27856 32224
rect 28632 32215 28684 32224
rect 28632 32181 28641 32215
rect 28641 32181 28675 32215
rect 28675 32181 28684 32215
rect 28632 32172 28684 32181
rect 30472 32172 30524 32224
rect 32312 32172 32364 32224
rect 32588 32172 32640 32224
rect 33048 32172 33100 32224
rect 34520 32172 34572 32224
rect 42156 32308 42208 32360
rect 38568 32283 38620 32292
rect 38568 32249 38577 32283
rect 38577 32249 38611 32283
rect 38611 32249 38620 32283
rect 38568 32240 38620 32249
rect 41052 32283 41104 32292
rect 41052 32249 41061 32283
rect 41061 32249 41095 32283
rect 41095 32249 41104 32283
rect 41052 32240 41104 32249
rect 41696 32283 41748 32292
rect 36268 32172 36320 32224
rect 36544 32215 36596 32224
rect 36544 32181 36553 32215
rect 36553 32181 36587 32215
rect 36587 32181 36596 32215
rect 36544 32172 36596 32181
rect 36820 32172 36872 32224
rect 37740 32172 37792 32224
rect 38016 32172 38068 32224
rect 40868 32215 40920 32224
rect 40868 32181 40877 32215
rect 40877 32181 40911 32215
rect 40911 32181 40920 32215
rect 41696 32249 41705 32283
rect 41705 32249 41739 32283
rect 41739 32249 41748 32283
rect 41696 32240 41748 32249
rect 44088 32240 44140 32292
rect 40868 32172 40920 32181
rect 43628 32172 43680 32224
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 10508 32011 10560 32020
rect 10508 31977 10517 32011
rect 10517 31977 10551 32011
rect 10551 31977 10560 32011
rect 10508 31968 10560 31977
rect 11428 32011 11480 32020
rect 11428 31977 11437 32011
rect 11437 31977 11471 32011
rect 11471 31977 11480 32011
rect 11428 31968 11480 31977
rect 12624 32011 12676 32020
rect 12624 31977 12633 32011
rect 12633 31977 12667 32011
rect 12667 31977 12676 32011
rect 12624 31968 12676 31977
rect 13176 31968 13228 32020
rect 16488 32011 16540 32020
rect 16488 31977 16497 32011
rect 16497 31977 16531 32011
rect 16531 31977 16540 32011
rect 16488 31968 16540 31977
rect 18236 32011 18288 32020
rect 18236 31977 18245 32011
rect 18245 31977 18279 32011
rect 18279 31977 18288 32011
rect 18236 31968 18288 31977
rect 18880 31968 18932 32020
rect 12532 31900 12584 31952
rect 13452 31900 13504 31952
rect 14832 31900 14884 31952
rect 15476 31943 15528 31952
rect 15476 31909 15485 31943
rect 15485 31909 15519 31943
rect 15519 31909 15528 31943
rect 15476 31900 15528 31909
rect 16948 31900 17000 31952
rect 17224 31943 17276 31952
rect 17224 31909 17233 31943
rect 17233 31909 17267 31943
rect 17267 31909 17276 31943
rect 20076 31968 20128 32020
rect 23112 31968 23164 32020
rect 23296 32011 23348 32020
rect 23296 31977 23305 32011
rect 23305 31977 23339 32011
rect 23339 31977 23348 32011
rect 23296 31968 23348 31977
rect 23940 31968 23992 32020
rect 24032 32011 24084 32020
rect 24032 31977 24041 32011
rect 24041 31977 24075 32011
rect 24075 31977 24084 32011
rect 24032 31968 24084 31977
rect 25228 31968 25280 32020
rect 26332 32011 26384 32020
rect 26332 31977 26341 32011
rect 26341 31977 26375 32011
rect 26375 31977 26384 32011
rect 26332 31968 26384 31977
rect 26424 31968 26476 32020
rect 30748 32011 30800 32020
rect 30748 31977 30757 32011
rect 30757 31977 30791 32011
rect 30791 31977 30800 32011
rect 30748 31968 30800 31977
rect 31944 31968 31996 32020
rect 32496 32011 32548 32020
rect 32496 31977 32505 32011
rect 32505 31977 32539 32011
rect 32539 31977 32548 32011
rect 32496 31968 32548 31977
rect 38476 31968 38528 32020
rect 41604 31968 41656 32020
rect 43720 31968 43772 32020
rect 17224 31900 17276 31909
rect 21548 31900 21600 31952
rect 9680 31832 9732 31884
rect 10416 31875 10468 31884
rect 10416 31841 10425 31875
rect 10425 31841 10459 31875
rect 10459 31841 10468 31875
rect 10416 31832 10468 31841
rect 10692 31832 10744 31884
rect 12348 31832 12400 31884
rect 12992 31832 13044 31884
rect 19340 31832 19392 31884
rect 20812 31832 20864 31884
rect 22192 31832 22244 31884
rect 23480 31900 23532 31952
rect 22652 31875 22704 31884
rect 22652 31841 22661 31875
rect 22661 31841 22695 31875
rect 22695 31841 22704 31875
rect 22652 31832 22704 31841
rect 24860 31900 24912 31952
rect 25136 31943 25188 31952
rect 25136 31909 25145 31943
rect 25145 31909 25179 31943
rect 25179 31909 25188 31943
rect 25136 31900 25188 31909
rect 26608 31900 26660 31952
rect 28080 31900 28132 31952
rect 28448 31943 28500 31952
rect 24492 31832 24544 31884
rect 24952 31875 25004 31884
rect 24952 31841 24961 31875
rect 24961 31841 24995 31875
rect 24995 31841 25004 31875
rect 24952 31832 25004 31841
rect 26424 31875 26476 31884
rect 26424 31841 26433 31875
rect 26433 31841 26467 31875
rect 26467 31841 26476 31875
rect 26424 31832 26476 31841
rect 27528 31832 27580 31884
rect 28448 31909 28457 31943
rect 28457 31909 28491 31943
rect 28491 31909 28500 31943
rect 28448 31900 28500 31909
rect 30012 31900 30064 31952
rect 34520 31900 34572 31952
rect 36084 31943 36136 31952
rect 36084 31909 36093 31943
rect 36093 31909 36127 31943
rect 36127 31909 36136 31943
rect 36084 31900 36136 31909
rect 36176 31943 36228 31952
rect 36176 31909 36185 31943
rect 36185 31909 36219 31943
rect 36219 31909 36228 31943
rect 36176 31900 36228 31909
rect 37740 31900 37792 31952
rect 38108 31943 38160 31952
rect 38108 31909 38117 31943
rect 38117 31909 38151 31943
rect 38151 31909 38160 31943
rect 38108 31900 38160 31909
rect 40316 31900 40368 31952
rect 40868 31943 40920 31952
rect 40868 31909 40877 31943
rect 40877 31909 40911 31943
rect 40911 31909 40920 31943
rect 40868 31900 40920 31909
rect 43996 31900 44048 31952
rect 38936 31832 38988 31884
rect 39856 31832 39908 31884
rect 42248 31875 42300 31884
rect 42248 31841 42257 31875
rect 42257 31841 42291 31875
rect 42291 31841 42300 31875
rect 42248 31832 42300 31841
rect 45100 31832 45152 31884
rect 13820 31764 13872 31816
rect 15384 31807 15436 31816
rect 15384 31773 15393 31807
rect 15393 31773 15427 31807
rect 15427 31773 15436 31807
rect 15384 31764 15436 31773
rect 19616 31807 19668 31816
rect 13728 31739 13780 31748
rect 13728 31705 13737 31739
rect 13737 31705 13771 31739
rect 13771 31705 13780 31739
rect 13728 31696 13780 31705
rect 15936 31739 15988 31748
rect 15936 31705 15945 31739
rect 15945 31705 15979 31739
rect 15979 31705 15988 31739
rect 19616 31773 19625 31807
rect 19625 31773 19659 31807
rect 19659 31773 19668 31807
rect 19616 31764 19668 31773
rect 20996 31764 21048 31816
rect 26700 31764 26752 31816
rect 27160 31764 27212 31816
rect 15936 31696 15988 31705
rect 17500 31696 17552 31748
rect 19892 31696 19944 31748
rect 26332 31696 26384 31748
rect 12992 31628 13044 31680
rect 14740 31628 14792 31680
rect 17040 31628 17092 31680
rect 19432 31671 19484 31680
rect 19432 31637 19456 31671
rect 19456 31637 19484 31671
rect 19432 31628 19484 31637
rect 20352 31671 20404 31680
rect 20352 31637 20361 31671
rect 20361 31637 20395 31671
rect 20395 31637 20404 31671
rect 20352 31628 20404 31637
rect 21364 31628 21416 31680
rect 25412 31671 25464 31680
rect 25412 31637 25421 31671
rect 25421 31637 25455 31671
rect 25455 31637 25464 31671
rect 25412 31628 25464 31637
rect 25872 31628 25924 31680
rect 27804 31764 27856 31816
rect 29552 31764 29604 31816
rect 32128 31807 32180 31816
rect 32128 31773 32137 31807
rect 32137 31773 32171 31807
rect 32171 31773 32180 31807
rect 32128 31764 32180 31773
rect 32680 31764 32732 31816
rect 33968 31764 34020 31816
rect 28172 31696 28224 31748
rect 30288 31696 30340 31748
rect 35256 31764 35308 31816
rect 38384 31807 38436 31816
rect 38384 31773 38393 31807
rect 38393 31773 38427 31807
rect 38427 31773 38436 31807
rect 38384 31764 38436 31773
rect 40776 31807 40828 31816
rect 40776 31773 40785 31807
rect 40785 31773 40819 31807
rect 40819 31773 40828 31807
rect 40776 31764 40828 31773
rect 41144 31807 41196 31816
rect 41144 31773 41153 31807
rect 41153 31773 41187 31807
rect 41187 31773 41196 31807
rect 41144 31764 41196 31773
rect 42616 31764 42668 31816
rect 44180 31807 44232 31816
rect 44180 31773 44189 31807
rect 44189 31773 44223 31807
rect 44223 31773 44232 31807
rect 44180 31764 44232 31773
rect 45284 31764 45336 31816
rect 35348 31696 35400 31748
rect 44088 31696 44140 31748
rect 27988 31671 28040 31680
rect 27988 31637 27997 31671
rect 27997 31637 28031 31671
rect 28031 31637 28040 31671
rect 27988 31628 28040 31637
rect 29276 31671 29328 31680
rect 29276 31637 29285 31671
rect 29285 31637 29319 31671
rect 29319 31637 29328 31671
rect 29276 31628 29328 31637
rect 32864 31628 32916 31680
rect 34796 31628 34848 31680
rect 41144 31628 41196 31680
rect 44272 31628 44324 31680
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 12992 31424 13044 31476
rect 13452 31467 13504 31476
rect 13452 31433 13461 31467
rect 13461 31433 13495 31467
rect 13495 31433 13504 31467
rect 13452 31424 13504 31433
rect 13820 31467 13872 31476
rect 13820 31433 13829 31467
rect 13829 31433 13863 31467
rect 13863 31433 13872 31467
rect 13820 31424 13872 31433
rect 15476 31424 15528 31476
rect 17224 31424 17276 31476
rect 19156 31424 19208 31476
rect 21732 31424 21784 31476
rect 23480 31424 23532 31476
rect 26424 31424 26476 31476
rect 30012 31424 30064 31476
rect 31576 31424 31628 31476
rect 32864 31424 32916 31476
rect 34520 31424 34572 31476
rect 35900 31424 35952 31476
rect 13636 31356 13688 31408
rect 16120 31356 16172 31408
rect 12532 31331 12584 31340
rect 12532 31297 12541 31331
rect 12541 31297 12575 31331
rect 12575 31297 12584 31331
rect 12532 31288 12584 31297
rect 13176 31288 13228 31340
rect 15384 31288 15436 31340
rect 17040 31331 17092 31340
rect 17040 31297 17049 31331
rect 17049 31297 17083 31331
rect 17083 31297 17092 31331
rect 17040 31288 17092 31297
rect 19616 31356 19668 31408
rect 19800 31399 19852 31408
rect 19800 31365 19809 31399
rect 19809 31365 19843 31399
rect 19843 31365 19852 31399
rect 19800 31356 19852 31365
rect 20812 31399 20864 31408
rect 20812 31365 20821 31399
rect 20821 31365 20855 31399
rect 20855 31365 20864 31399
rect 20812 31356 20864 31365
rect 20996 31356 21048 31408
rect 22652 31356 22704 31408
rect 12808 31152 12860 31204
rect 12900 31152 12952 31204
rect 15292 31220 15344 31272
rect 16488 31220 16540 31272
rect 18236 31220 18288 31272
rect 19432 31220 19484 31272
rect 20444 31220 20496 31272
rect 20904 31220 20956 31272
rect 27436 31356 27488 31408
rect 36176 31356 36228 31408
rect 25780 31288 25832 31340
rect 24952 31263 25004 31272
rect 24952 31229 24961 31263
rect 24961 31229 24995 31263
rect 24995 31229 25004 31263
rect 24952 31220 25004 31229
rect 27988 31288 28040 31340
rect 29276 31331 29328 31340
rect 29276 31297 29285 31331
rect 29285 31297 29319 31331
rect 29319 31297 29328 31331
rect 29276 31288 29328 31297
rect 32220 31288 32272 31340
rect 34244 31288 34296 31340
rect 35164 31288 35216 31340
rect 35440 31331 35492 31340
rect 35440 31297 35449 31331
rect 35449 31297 35483 31331
rect 35483 31297 35492 31331
rect 35440 31288 35492 31297
rect 28172 31263 28224 31272
rect 17408 31152 17460 31204
rect 17868 31152 17920 31204
rect 19156 31152 19208 31204
rect 20352 31152 20404 31204
rect 25412 31195 25464 31204
rect 10416 31127 10468 31136
rect 10416 31093 10425 31127
rect 10425 31093 10459 31127
rect 10459 31093 10468 31127
rect 10416 31084 10468 31093
rect 10692 31084 10744 31136
rect 11704 31084 11756 31136
rect 12348 31084 12400 31136
rect 13084 31084 13136 31136
rect 14924 31127 14976 31136
rect 14924 31093 14933 31127
rect 14933 31093 14967 31127
rect 14967 31093 14976 31127
rect 14924 31084 14976 31093
rect 18972 31084 19024 31136
rect 22284 31084 22336 31136
rect 23940 31127 23992 31136
rect 23940 31093 23949 31127
rect 23949 31093 23983 31127
rect 23983 31093 23992 31127
rect 23940 31084 23992 31093
rect 25412 31161 25421 31195
rect 25421 31161 25455 31195
rect 25455 31161 25464 31195
rect 25412 31152 25464 31161
rect 25964 31195 26016 31204
rect 25964 31161 25973 31195
rect 25973 31161 26007 31195
rect 26007 31161 26016 31195
rect 25964 31152 26016 31161
rect 27620 31152 27672 31204
rect 28172 31229 28181 31263
rect 28181 31229 28215 31263
rect 28215 31229 28224 31263
rect 28172 31220 28224 31229
rect 28632 31220 28684 31272
rect 30932 31263 30984 31272
rect 30932 31229 30941 31263
rect 30941 31229 30975 31263
rect 30975 31229 30984 31263
rect 30932 31220 30984 31229
rect 38108 31424 38160 31476
rect 40316 31467 40368 31476
rect 40316 31433 40325 31467
rect 40325 31433 40359 31467
rect 40359 31433 40368 31467
rect 40316 31424 40368 31433
rect 41052 31424 41104 31476
rect 42616 31467 42668 31476
rect 42616 31433 42625 31467
rect 42625 31433 42659 31467
rect 42659 31433 42668 31467
rect 42616 31424 42668 31433
rect 43720 31424 43772 31476
rect 44088 31424 44140 31476
rect 40592 31356 40644 31408
rect 40868 31356 40920 31408
rect 42984 31356 43036 31408
rect 37372 31331 37424 31340
rect 37372 31297 37381 31331
rect 37381 31297 37415 31331
rect 37415 31297 37424 31331
rect 37372 31288 37424 31297
rect 43628 31331 43680 31340
rect 36912 31220 36964 31272
rect 43628 31297 43637 31331
rect 43637 31297 43671 31331
rect 43671 31297 43680 31331
rect 43628 31288 43680 31297
rect 26240 31084 26292 31136
rect 27712 31084 27764 31136
rect 28724 31127 28776 31136
rect 28724 31093 28733 31127
rect 28733 31093 28767 31127
rect 28767 31093 28776 31127
rect 28724 31084 28776 31093
rect 29000 31127 29052 31136
rect 29000 31093 29009 31127
rect 29009 31093 29043 31127
rect 29043 31093 29052 31127
rect 29000 31084 29052 31093
rect 30380 31084 30432 31136
rect 32496 31152 32548 31204
rect 34704 31152 34756 31204
rect 34796 31152 34848 31204
rect 33416 31084 33468 31136
rect 33968 31127 34020 31136
rect 33968 31093 33977 31127
rect 33977 31093 34011 31127
rect 34011 31093 34020 31127
rect 33968 31084 34020 31093
rect 35164 31152 35216 31204
rect 35532 31084 35584 31136
rect 39948 31220 40000 31272
rect 40316 31220 40368 31272
rect 39580 31195 39632 31204
rect 39580 31161 39589 31195
rect 39589 31161 39623 31195
rect 39623 31161 39632 31195
rect 39580 31152 39632 31161
rect 40776 31152 40828 31204
rect 41236 31152 41288 31204
rect 39856 31127 39908 31136
rect 39856 31093 39865 31127
rect 39865 31093 39899 31127
rect 39899 31093 39908 31127
rect 39856 31084 39908 31093
rect 40868 31084 40920 31136
rect 44732 31220 44784 31272
rect 45100 31263 45152 31272
rect 45100 31229 45109 31263
rect 45109 31229 45143 31263
rect 45143 31229 45152 31263
rect 45100 31220 45152 31229
rect 43720 31195 43772 31204
rect 43720 31161 43729 31195
rect 43729 31161 43763 31195
rect 43763 31161 43772 31195
rect 43720 31152 43772 31161
rect 42340 31127 42392 31136
rect 42340 31093 42349 31127
rect 42349 31093 42383 31127
rect 42383 31093 42392 31127
rect 42340 31084 42392 31093
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 13728 30923 13780 30932
rect 13728 30889 13737 30923
rect 13737 30889 13771 30923
rect 13771 30889 13780 30923
rect 13728 30880 13780 30889
rect 11980 30855 12032 30864
rect 11980 30821 11989 30855
rect 11989 30821 12023 30855
rect 12023 30821 12032 30855
rect 11980 30812 12032 30821
rect 12532 30855 12584 30864
rect 12532 30821 12541 30855
rect 12541 30821 12575 30855
rect 12575 30821 12584 30855
rect 12532 30812 12584 30821
rect 15476 30855 15528 30864
rect 15476 30821 15485 30855
rect 15485 30821 15519 30855
rect 15519 30821 15528 30855
rect 15476 30812 15528 30821
rect 16948 30880 17000 30932
rect 18144 30880 18196 30932
rect 19064 30923 19116 30932
rect 19064 30889 19073 30923
rect 19073 30889 19107 30923
rect 19107 30889 19116 30923
rect 19064 30880 19116 30889
rect 20444 30923 20496 30932
rect 20444 30889 20453 30923
rect 20453 30889 20487 30923
rect 20487 30889 20496 30923
rect 20444 30880 20496 30889
rect 23940 30880 23992 30932
rect 24492 30923 24544 30932
rect 24492 30889 24501 30923
rect 24501 30889 24535 30923
rect 24535 30889 24544 30923
rect 24492 30880 24544 30889
rect 28264 30880 28316 30932
rect 30012 30880 30064 30932
rect 17132 30812 17184 30864
rect 17592 30855 17644 30864
rect 17592 30821 17601 30855
rect 17601 30821 17635 30855
rect 17635 30821 17644 30855
rect 17592 30812 17644 30821
rect 22928 30855 22980 30864
rect 22928 30821 22937 30855
rect 22937 30821 22971 30855
rect 22971 30821 22980 30855
rect 22928 30812 22980 30821
rect 24952 30812 25004 30864
rect 25964 30812 26016 30864
rect 32220 30880 32272 30932
rect 32680 30923 32732 30932
rect 32680 30889 32689 30923
rect 32689 30889 32723 30923
rect 32723 30889 32732 30923
rect 32680 30880 32732 30889
rect 32864 30880 32916 30932
rect 30472 30812 30524 30864
rect 33048 30855 33100 30864
rect 33048 30821 33057 30855
rect 33057 30821 33091 30855
rect 33091 30821 33100 30855
rect 33048 30812 33100 30821
rect 33324 30880 33376 30932
rect 37740 30880 37792 30932
rect 41236 30923 41288 30932
rect 41236 30889 41245 30923
rect 41245 30889 41279 30923
rect 41279 30889 41288 30923
rect 41236 30880 41288 30889
rect 41696 30923 41748 30932
rect 41696 30889 41705 30923
rect 41705 30889 41739 30923
rect 41739 30889 41748 30923
rect 41696 30880 41748 30889
rect 34704 30855 34756 30864
rect 34704 30821 34713 30855
rect 34713 30821 34747 30855
rect 34747 30821 34756 30855
rect 34704 30812 34756 30821
rect 35256 30855 35308 30864
rect 35256 30821 35265 30855
rect 35265 30821 35299 30855
rect 35299 30821 35308 30855
rect 35256 30812 35308 30821
rect 35992 30855 36044 30864
rect 35992 30821 36001 30855
rect 36001 30821 36035 30855
rect 36035 30821 36044 30855
rect 35992 30812 36044 30821
rect 36820 30855 36872 30864
rect 36820 30821 36829 30855
rect 36829 30821 36863 30855
rect 36863 30821 36872 30855
rect 36820 30812 36872 30821
rect 38476 30855 38528 30864
rect 38476 30821 38485 30855
rect 38485 30821 38519 30855
rect 38519 30821 38528 30855
rect 38476 30812 38528 30821
rect 40408 30855 40460 30864
rect 40408 30821 40417 30855
rect 40417 30821 40451 30855
rect 40451 30821 40460 30855
rect 40408 30812 40460 30821
rect 40684 30812 40736 30864
rect 43904 30812 43956 30864
rect 44272 30812 44324 30864
rect 45008 30855 45060 30864
rect 45008 30821 45017 30855
rect 45017 30821 45051 30855
rect 45051 30821 45060 30855
rect 45008 30812 45060 30821
rect 45100 30855 45152 30864
rect 45100 30821 45109 30855
rect 45109 30821 45143 30855
rect 45143 30821 45152 30855
rect 45100 30812 45152 30821
rect 10508 30787 10560 30796
rect 10508 30753 10517 30787
rect 10517 30753 10551 30787
rect 10551 30753 10560 30787
rect 10508 30744 10560 30753
rect 10692 30787 10744 30796
rect 10692 30753 10701 30787
rect 10701 30753 10735 30787
rect 10735 30753 10744 30787
rect 10692 30744 10744 30753
rect 13636 30744 13688 30796
rect 14648 30744 14700 30796
rect 18328 30744 18380 30796
rect 18972 30787 19024 30796
rect 18972 30753 18981 30787
rect 18981 30753 19015 30787
rect 19015 30753 19024 30787
rect 18972 30744 19024 30753
rect 19432 30787 19484 30796
rect 10784 30719 10836 30728
rect 10784 30685 10793 30719
rect 10793 30685 10827 30719
rect 10827 30685 10836 30719
rect 10784 30676 10836 30685
rect 11888 30719 11940 30728
rect 11888 30685 11897 30719
rect 11897 30685 11931 30719
rect 11931 30685 11940 30719
rect 11888 30676 11940 30685
rect 15016 30676 15068 30728
rect 17500 30719 17552 30728
rect 17500 30685 17509 30719
rect 17509 30685 17543 30719
rect 17543 30685 17552 30719
rect 17500 30676 17552 30685
rect 12808 30583 12860 30592
rect 12808 30549 12817 30583
rect 12817 30549 12851 30583
rect 12851 30549 12860 30583
rect 12808 30540 12860 30549
rect 14372 30540 14424 30592
rect 18972 30608 19024 30660
rect 16396 30583 16448 30592
rect 16396 30549 16405 30583
rect 16405 30549 16439 30583
rect 16439 30549 16448 30583
rect 19432 30753 19441 30787
rect 19441 30753 19475 30787
rect 19475 30753 19484 30787
rect 19432 30744 19484 30753
rect 19892 30744 19944 30796
rect 20628 30744 20680 30796
rect 21180 30787 21232 30796
rect 21180 30753 21189 30787
rect 21189 30753 21223 30787
rect 21223 30753 21232 30787
rect 21180 30744 21232 30753
rect 21640 30787 21692 30796
rect 21640 30753 21649 30787
rect 21649 30753 21683 30787
rect 21683 30753 21692 30787
rect 21640 30744 21692 30753
rect 22192 30676 22244 30728
rect 22652 30676 22704 30728
rect 23480 30719 23532 30728
rect 23480 30685 23489 30719
rect 23489 30685 23523 30719
rect 23523 30685 23532 30719
rect 24124 30719 24176 30728
rect 23480 30676 23532 30685
rect 24124 30685 24133 30719
rect 24133 30685 24167 30719
rect 24167 30685 24176 30719
rect 24124 30676 24176 30685
rect 20352 30608 20404 30660
rect 27528 30744 27580 30796
rect 29092 30744 29144 30796
rect 36360 30744 36412 30796
rect 42248 30787 42300 30796
rect 42248 30753 42292 30787
rect 42292 30753 42300 30787
rect 42248 30744 42300 30753
rect 27436 30719 27488 30728
rect 27436 30685 27445 30719
rect 27445 30685 27479 30719
rect 27479 30685 27488 30719
rect 27436 30676 27488 30685
rect 28632 30676 28684 30728
rect 30104 30719 30156 30728
rect 30104 30685 30113 30719
rect 30113 30685 30147 30719
rect 30147 30685 30156 30719
rect 30104 30676 30156 30685
rect 30840 30676 30892 30728
rect 29552 30608 29604 30660
rect 30564 30608 30616 30660
rect 33232 30676 33284 30728
rect 33508 30676 33560 30728
rect 33692 30719 33744 30728
rect 33692 30685 33701 30719
rect 33701 30685 33735 30719
rect 33735 30685 33744 30719
rect 33692 30676 33744 30685
rect 37464 30676 37516 30728
rect 38384 30719 38436 30728
rect 38384 30685 38393 30719
rect 38393 30685 38427 30719
rect 38427 30685 38436 30719
rect 38384 30676 38436 30685
rect 38568 30676 38620 30728
rect 32956 30608 33008 30660
rect 40776 30676 40828 30728
rect 41144 30676 41196 30728
rect 43444 30719 43496 30728
rect 43444 30685 43453 30719
rect 43453 30685 43487 30719
rect 43487 30685 43496 30719
rect 43444 30676 43496 30685
rect 45284 30719 45336 30728
rect 45284 30685 45293 30719
rect 45293 30685 45327 30719
rect 45327 30685 45336 30719
rect 45284 30676 45336 30685
rect 41880 30608 41932 30660
rect 16396 30540 16448 30549
rect 21824 30540 21876 30592
rect 25780 30583 25832 30592
rect 25780 30549 25789 30583
rect 25789 30549 25823 30583
rect 25823 30549 25832 30583
rect 25780 30540 25832 30549
rect 27068 30540 27120 30592
rect 27620 30540 27672 30592
rect 29644 30540 29696 30592
rect 30932 30540 30984 30592
rect 35256 30540 35308 30592
rect 41696 30540 41748 30592
rect 44272 30540 44324 30592
rect 44456 30583 44508 30592
rect 44456 30549 44465 30583
rect 44465 30549 44499 30583
rect 44499 30549 44508 30583
rect 44456 30540 44508 30549
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 12808 30336 12860 30388
rect 13360 30336 13412 30388
rect 14280 30336 14332 30388
rect 14648 30379 14700 30388
rect 14648 30345 14657 30379
rect 14657 30345 14691 30379
rect 14691 30345 14700 30379
rect 14648 30336 14700 30345
rect 17316 30379 17368 30388
rect 17316 30345 17325 30379
rect 17325 30345 17359 30379
rect 17359 30345 17368 30379
rect 17316 30336 17368 30345
rect 17592 30379 17644 30388
rect 17592 30345 17601 30379
rect 17601 30345 17635 30379
rect 17635 30345 17644 30379
rect 17592 30336 17644 30345
rect 19432 30336 19484 30388
rect 20628 30379 20680 30388
rect 20628 30345 20637 30379
rect 20637 30345 20671 30379
rect 20671 30345 20680 30379
rect 20628 30336 20680 30345
rect 22652 30336 22704 30388
rect 22928 30336 22980 30388
rect 24124 30336 24176 30388
rect 11888 30268 11940 30320
rect 10784 30200 10836 30252
rect 11796 30243 11848 30252
rect 11796 30209 11805 30243
rect 11805 30209 11839 30243
rect 11839 30209 11848 30243
rect 11796 30200 11848 30209
rect 11980 30200 12032 30252
rect 15844 30311 15896 30320
rect 15844 30277 15853 30311
rect 15853 30277 15887 30311
rect 15887 30277 15896 30311
rect 15844 30268 15896 30277
rect 19064 30200 19116 30252
rect 11244 30132 11296 30184
rect 13360 30132 13412 30184
rect 14372 30175 14424 30184
rect 14372 30141 14381 30175
rect 14381 30141 14415 30175
rect 14415 30141 14424 30175
rect 14372 30132 14424 30141
rect 17316 30132 17368 30184
rect 17684 30132 17736 30184
rect 19892 30132 19944 30184
rect 21364 30175 21416 30184
rect 21364 30141 21373 30175
rect 21373 30141 21407 30175
rect 21407 30141 21416 30175
rect 21364 30132 21416 30141
rect 11336 30064 11388 30116
rect 13728 30107 13780 30116
rect 13728 30073 13737 30107
rect 13737 30073 13771 30107
rect 13771 30073 13780 30107
rect 13728 30064 13780 30073
rect 13820 30107 13872 30116
rect 13820 30073 13829 30107
rect 13829 30073 13863 30107
rect 13863 30073 13872 30107
rect 13820 30064 13872 30073
rect 15476 30064 15528 30116
rect 18512 30064 18564 30116
rect 25872 30336 25924 30388
rect 21824 30175 21876 30184
rect 21824 30141 21833 30175
rect 21833 30141 21867 30175
rect 21867 30141 21876 30175
rect 21824 30132 21876 30141
rect 23756 30132 23808 30184
rect 25596 30132 25648 30184
rect 26332 30243 26384 30252
rect 26332 30209 26341 30243
rect 26341 30209 26375 30243
rect 26375 30209 26384 30243
rect 26332 30200 26384 30209
rect 29552 30336 29604 30388
rect 30104 30336 30156 30388
rect 30472 30379 30524 30388
rect 30472 30345 30481 30379
rect 30481 30345 30515 30379
rect 30515 30345 30524 30379
rect 30472 30336 30524 30345
rect 32864 30336 32916 30388
rect 33048 30379 33100 30388
rect 33048 30345 33057 30379
rect 33057 30345 33091 30379
rect 33091 30345 33100 30379
rect 33048 30336 33100 30345
rect 36360 30336 36412 30388
rect 37832 30336 37884 30388
rect 38476 30336 38528 30388
rect 40408 30336 40460 30388
rect 29644 30268 29696 30320
rect 29092 30243 29144 30252
rect 29092 30209 29101 30243
rect 29101 30209 29135 30243
rect 29135 30209 29144 30243
rect 29092 30200 29144 30209
rect 30196 30200 30248 30252
rect 30840 30243 30892 30252
rect 30840 30209 30849 30243
rect 30849 30209 30883 30243
rect 30883 30209 30892 30243
rect 30840 30200 30892 30209
rect 31300 30200 31352 30252
rect 33968 30268 34020 30320
rect 35256 30200 35308 30252
rect 35348 30243 35400 30252
rect 35348 30209 35357 30243
rect 35357 30209 35391 30243
rect 35391 30209 35400 30243
rect 37372 30243 37424 30252
rect 35348 30200 35400 30209
rect 37372 30209 37381 30243
rect 37381 30209 37415 30243
rect 37415 30209 37424 30243
rect 37372 30200 37424 30209
rect 38384 30268 38436 30320
rect 41512 30268 41564 30320
rect 42248 30311 42300 30320
rect 41696 30200 41748 30252
rect 22468 30064 22520 30116
rect 22928 30064 22980 30116
rect 24952 30064 25004 30116
rect 9496 30039 9548 30048
rect 9496 30005 9505 30039
rect 9505 30005 9539 30039
rect 9539 30005 9548 30039
rect 9496 29996 9548 30005
rect 10048 30039 10100 30048
rect 10048 30005 10057 30039
rect 10057 30005 10091 30039
rect 10091 30005 10100 30039
rect 10048 29996 10100 30005
rect 16304 29996 16356 30048
rect 18328 30039 18380 30048
rect 18328 30005 18337 30039
rect 18337 30005 18371 30039
rect 18371 30005 18380 30039
rect 18328 29996 18380 30005
rect 18880 29996 18932 30048
rect 23756 29996 23808 30048
rect 25412 29996 25464 30048
rect 27436 29996 27488 30048
rect 27620 30039 27672 30048
rect 27620 30005 27629 30039
rect 27629 30005 27663 30039
rect 27663 30005 27672 30039
rect 27620 29996 27672 30005
rect 29552 30132 29604 30184
rect 30012 30132 30064 30184
rect 39028 30132 39080 30184
rect 42248 30277 42257 30311
rect 42257 30277 42291 30311
rect 42291 30277 42300 30311
rect 42248 30268 42300 30277
rect 43444 30336 43496 30388
rect 44456 30336 44508 30388
rect 46572 30379 46624 30388
rect 46572 30345 46581 30379
rect 46581 30345 46615 30379
rect 46615 30345 46624 30379
rect 46572 30336 46624 30345
rect 42984 30268 43036 30320
rect 44364 30311 44416 30320
rect 44364 30277 44373 30311
rect 44373 30277 44407 30311
rect 44407 30277 44416 30311
rect 44364 30268 44416 30277
rect 43628 30200 43680 30252
rect 45008 30268 45060 30320
rect 45100 30243 45152 30252
rect 45100 30209 45109 30243
rect 45109 30209 45143 30243
rect 45143 30209 45152 30243
rect 45100 30200 45152 30209
rect 42800 30175 42852 30184
rect 42800 30141 42818 30175
rect 42818 30141 42852 30175
rect 42800 30132 42852 30141
rect 44456 30132 44508 30184
rect 46572 30132 46624 30184
rect 30932 30107 30984 30116
rect 30932 30073 30941 30107
rect 30941 30073 30975 30107
rect 30975 30073 30984 30107
rect 30932 30064 30984 30073
rect 33324 30107 33376 30116
rect 28816 29996 28868 30048
rect 31392 29996 31444 30048
rect 33324 30073 33333 30107
rect 33333 30073 33367 30107
rect 33367 30073 33376 30107
rect 33324 30064 33376 30073
rect 33416 30107 33468 30116
rect 33416 30073 33425 30107
rect 33425 30073 33459 30107
rect 33459 30073 33468 30107
rect 33416 30064 33468 30073
rect 33692 30064 33744 30116
rect 34336 30064 34388 30116
rect 34980 29996 35032 30048
rect 37832 30064 37884 30116
rect 41328 30107 41380 30116
rect 41328 30073 41337 30107
rect 41337 30073 41371 30107
rect 41371 30073 41380 30107
rect 41880 30107 41932 30116
rect 41328 30064 41380 30073
rect 41880 30073 41889 30107
rect 41889 30073 41923 30107
rect 41923 30073 41932 30107
rect 41880 30064 41932 30073
rect 43904 30107 43956 30116
rect 43904 30073 43913 30107
rect 43913 30073 43947 30107
rect 43947 30073 43956 30107
rect 43904 30064 43956 30073
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 10508 29792 10560 29844
rect 10784 29835 10836 29844
rect 10784 29801 10793 29835
rect 10793 29801 10827 29835
rect 10827 29801 10836 29835
rect 10784 29792 10836 29801
rect 11796 29835 11848 29844
rect 11796 29801 11805 29835
rect 11805 29801 11839 29835
rect 11839 29801 11848 29835
rect 11796 29792 11848 29801
rect 13820 29792 13872 29844
rect 15016 29835 15068 29844
rect 15016 29801 15025 29835
rect 15025 29801 15059 29835
rect 15059 29801 15068 29835
rect 15016 29792 15068 29801
rect 17316 29835 17368 29844
rect 11336 29724 11388 29776
rect 13452 29724 13504 29776
rect 17316 29801 17325 29835
rect 17325 29801 17359 29835
rect 17359 29801 17368 29835
rect 17316 29792 17368 29801
rect 17592 29792 17644 29844
rect 19064 29792 19116 29844
rect 22468 29792 22520 29844
rect 24952 29835 25004 29844
rect 24952 29801 24961 29835
rect 24961 29801 24995 29835
rect 24995 29801 25004 29835
rect 24952 29792 25004 29801
rect 25412 29792 25464 29844
rect 25780 29792 25832 29844
rect 27528 29835 27580 29844
rect 27528 29801 27537 29835
rect 27537 29801 27571 29835
rect 27571 29801 27580 29835
rect 27528 29792 27580 29801
rect 30104 29835 30156 29844
rect 30104 29801 30113 29835
rect 30113 29801 30147 29835
rect 30147 29801 30156 29835
rect 30104 29792 30156 29801
rect 33324 29792 33376 29844
rect 34980 29835 35032 29844
rect 34980 29801 34989 29835
rect 34989 29801 35023 29835
rect 35023 29801 35032 29835
rect 34980 29792 35032 29801
rect 36636 29792 36688 29844
rect 37372 29835 37424 29844
rect 37372 29801 37381 29835
rect 37381 29801 37415 29835
rect 37415 29801 37424 29835
rect 37372 29792 37424 29801
rect 40408 29835 40460 29844
rect 40408 29801 40417 29835
rect 40417 29801 40451 29835
rect 40451 29801 40460 29835
rect 40408 29792 40460 29801
rect 40776 29835 40828 29844
rect 40776 29801 40785 29835
rect 40785 29801 40819 29835
rect 40819 29801 40828 29835
rect 40776 29792 40828 29801
rect 41328 29792 41380 29844
rect 15476 29767 15528 29776
rect 15476 29733 15485 29767
rect 15485 29733 15519 29767
rect 15519 29733 15528 29767
rect 15476 29724 15528 29733
rect 17500 29724 17552 29776
rect 18880 29767 18932 29776
rect 18880 29733 18889 29767
rect 18889 29733 18923 29767
rect 18923 29733 18932 29767
rect 18880 29724 18932 29733
rect 24124 29767 24176 29776
rect 24124 29733 24133 29767
rect 24133 29733 24167 29767
rect 24167 29733 24176 29767
rect 26332 29767 26384 29776
rect 24124 29724 24176 29733
rect 26332 29733 26341 29767
rect 26341 29733 26375 29767
rect 26375 29733 26384 29767
rect 26332 29724 26384 29733
rect 30380 29767 30432 29776
rect 30380 29733 30389 29767
rect 30389 29733 30423 29767
rect 30423 29733 30432 29767
rect 30380 29724 30432 29733
rect 31944 29724 31996 29776
rect 12900 29656 12952 29708
rect 14372 29656 14424 29708
rect 21088 29656 21140 29708
rect 9864 29588 9916 29640
rect 10876 29631 10928 29640
rect 10876 29597 10885 29631
rect 10885 29597 10919 29631
rect 10919 29597 10928 29631
rect 10876 29588 10928 29597
rect 12992 29631 13044 29640
rect 12992 29597 13001 29631
rect 13001 29597 13035 29631
rect 13035 29597 13044 29631
rect 12992 29588 13044 29597
rect 14648 29588 14700 29640
rect 16304 29588 16356 29640
rect 16948 29631 17000 29640
rect 16948 29597 16957 29631
rect 16957 29597 16991 29631
rect 16991 29597 17000 29631
rect 16948 29588 17000 29597
rect 18788 29631 18840 29640
rect 18788 29597 18797 29631
rect 18797 29597 18831 29631
rect 18831 29597 18840 29631
rect 18788 29588 18840 29597
rect 18972 29588 19024 29640
rect 22192 29631 22244 29640
rect 22192 29597 22201 29631
rect 22201 29597 22235 29631
rect 22235 29597 22244 29631
rect 22192 29588 22244 29597
rect 26608 29656 26660 29708
rect 28356 29699 28408 29708
rect 28356 29665 28365 29699
rect 28365 29665 28399 29699
rect 28399 29665 28408 29699
rect 28356 29656 28408 29665
rect 28724 29699 28776 29708
rect 28724 29665 28733 29699
rect 28733 29665 28767 29699
rect 28767 29665 28776 29699
rect 28724 29656 28776 29665
rect 31484 29656 31536 29708
rect 32128 29699 32180 29708
rect 32128 29665 32137 29699
rect 32137 29665 32171 29699
rect 32171 29665 32180 29699
rect 32128 29656 32180 29665
rect 32496 29724 32548 29776
rect 34152 29767 34204 29776
rect 34152 29733 34161 29767
rect 34161 29733 34195 29767
rect 34195 29733 34204 29767
rect 34152 29724 34204 29733
rect 37832 29724 37884 29776
rect 39396 29724 39448 29776
rect 41144 29724 41196 29776
rect 43904 29792 43956 29844
rect 45100 29792 45152 29844
rect 43444 29724 43496 29776
rect 32588 29699 32640 29708
rect 32588 29665 32597 29699
rect 32597 29665 32631 29699
rect 32631 29665 32640 29699
rect 32588 29656 32640 29665
rect 33416 29656 33468 29708
rect 35532 29699 35584 29708
rect 35532 29665 35541 29699
rect 35541 29665 35575 29699
rect 35575 29665 35584 29699
rect 35532 29656 35584 29665
rect 36452 29656 36504 29708
rect 24032 29631 24084 29640
rect 24032 29597 24041 29631
rect 24041 29597 24075 29631
rect 24075 29597 24084 29631
rect 24032 29588 24084 29597
rect 15936 29563 15988 29572
rect 15936 29529 15945 29563
rect 15945 29529 15979 29563
rect 15979 29529 15988 29563
rect 15936 29520 15988 29529
rect 23296 29520 23348 29572
rect 23480 29520 23532 29572
rect 29184 29588 29236 29640
rect 30288 29631 30340 29640
rect 30288 29597 30297 29631
rect 30297 29597 30331 29631
rect 30331 29597 30340 29631
rect 30288 29588 30340 29597
rect 25228 29520 25280 29572
rect 27068 29563 27120 29572
rect 27068 29529 27077 29563
rect 27077 29529 27111 29563
rect 27111 29529 27120 29563
rect 27068 29520 27120 29529
rect 28448 29520 28500 29572
rect 31392 29588 31444 29640
rect 33048 29588 33100 29640
rect 34336 29631 34388 29640
rect 34336 29597 34345 29631
rect 34345 29597 34379 29631
rect 34379 29597 34388 29631
rect 34336 29588 34388 29597
rect 37740 29631 37792 29640
rect 37740 29597 37749 29631
rect 37749 29597 37783 29631
rect 37783 29597 37792 29631
rect 37740 29588 37792 29597
rect 39580 29656 39632 29708
rect 45100 29699 45152 29708
rect 45100 29665 45109 29699
rect 45109 29665 45143 29699
rect 45143 29665 45152 29699
rect 45100 29656 45152 29665
rect 39856 29588 39908 29640
rect 41236 29631 41288 29640
rect 41236 29597 41245 29631
rect 41245 29597 41279 29631
rect 41279 29597 41288 29631
rect 41236 29588 41288 29597
rect 43352 29631 43404 29640
rect 43352 29597 43361 29631
rect 43361 29597 43395 29631
rect 43395 29597 43404 29631
rect 43352 29588 43404 29597
rect 31300 29563 31352 29572
rect 31300 29529 31309 29563
rect 31309 29529 31343 29563
rect 31343 29529 31352 29563
rect 31300 29520 31352 29529
rect 35440 29520 35492 29572
rect 10140 29452 10192 29504
rect 12532 29495 12584 29504
rect 12532 29461 12541 29495
rect 12541 29461 12575 29495
rect 12575 29461 12584 29495
rect 12532 29452 12584 29461
rect 20444 29452 20496 29504
rect 21640 29495 21692 29504
rect 21640 29461 21649 29495
rect 21649 29461 21683 29495
rect 21683 29461 21692 29495
rect 21640 29452 21692 29461
rect 29276 29495 29328 29504
rect 29276 29461 29285 29495
rect 29285 29461 29319 29495
rect 29319 29461 29328 29495
rect 29276 29452 29328 29461
rect 35348 29495 35400 29504
rect 35348 29461 35357 29495
rect 35357 29461 35391 29495
rect 35391 29461 35400 29495
rect 35348 29452 35400 29461
rect 35900 29452 35952 29504
rect 35992 29452 36044 29504
rect 38660 29495 38712 29504
rect 38660 29461 38669 29495
rect 38669 29461 38703 29495
rect 38703 29461 38712 29495
rect 38660 29452 38712 29461
rect 44824 29452 44876 29504
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 10232 29248 10284 29300
rect 12440 29248 12492 29300
rect 13452 29291 13504 29300
rect 13452 29257 13461 29291
rect 13461 29257 13495 29291
rect 13495 29257 13504 29291
rect 13452 29248 13504 29257
rect 14648 29291 14700 29300
rect 14648 29257 14657 29291
rect 14657 29257 14691 29291
rect 14691 29257 14700 29291
rect 14648 29248 14700 29257
rect 15476 29248 15528 29300
rect 18420 29248 18472 29300
rect 18880 29291 18932 29300
rect 18880 29257 18889 29291
rect 18889 29257 18923 29291
rect 18923 29257 18932 29291
rect 18880 29248 18932 29257
rect 19156 29248 19208 29300
rect 24032 29248 24084 29300
rect 28356 29248 28408 29300
rect 28724 29248 28776 29300
rect 32588 29291 32640 29300
rect 32588 29257 32597 29291
rect 32597 29257 32631 29291
rect 32631 29257 32640 29291
rect 32588 29248 32640 29257
rect 34152 29248 34204 29300
rect 36728 29248 36780 29300
rect 44824 29291 44876 29300
rect 11336 29223 11388 29232
rect 11336 29189 11345 29223
rect 11345 29189 11379 29223
rect 11379 29189 11388 29223
rect 11336 29180 11388 29189
rect 18788 29180 18840 29232
rect 20444 29223 20496 29232
rect 20444 29189 20453 29223
rect 20453 29189 20487 29223
rect 20487 29189 20496 29223
rect 20444 29180 20496 29189
rect 10876 29112 10928 29164
rect 12992 29155 13044 29164
rect 12992 29121 13001 29155
rect 13001 29121 13035 29155
rect 13035 29121 13044 29155
rect 12992 29112 13044 29121
rect 16948 29112 17000 29164
rect 18696 29112 18748 29164
rect 19984 29155 20036 29164
rect 19984 29121 19993 29155
rect 19993 29121 20027 29155
rect 20027 29121 20036 29155
rect 19984 29112 20036 29121
rect 20904 29112 20956 29164
rect 21088 29112 21140 29164
rect 22468 29112 22520 29164
rect 24124 29112 24176 29164
rect 26056 29155 26108 29164
rect 26056 29121 26065 29155
rect 26065 29121 26099 29155
rect 26099 29121 26108 29155
rect 26056 29112 26108 29121
rect 32772 29180 32824 29232
rect 33508 29180 33560 29232
rect 27620 29112 27672 29164
rect 30564 29112 30616 29164
rect 31300 29112 31352 29164
rect 31392 29155 31444 29164
rect 31392 29121 31401 29155
rect 31401 29121 31435 29155
rect 31435 29121 31444 29155
rect 31392 29112 31444 29121
rect 10232 29087 10284 29096
rect 10232 29053 10241 29087
rect 10241 29053 10275 29087
rect 10275 29053 10284 29087
rect 10232 29044 10284 29053
rect 12440 29087 12492 29096
rect 9496 28976 9548 29028
rect 10692 28976 10744 29028
rect 12440 29053 12449 29087
rect 12449 29053 12483 29087
rect 12483 29053 12492 29087
rect 12440 29044 12492 29053
rect 12532 29044 12584 29096
rect 14464 29044 14516 29096
rect 14924 29044 14976 29096
rect 16212 29087 16264 29096
rect 16212 29053 16221 29087
rect 16221 29053 16255 29087
rect 16255 29053 16264 29087
rect 16212 29044 16264 29053
rect 16580 29044 16632 29096
rect 16304 28976 16356 29028
rect 18420 29044 18472 29096
rect 21548 29044 21600 29096
rect 17316 28976 17368 29028
rect 18512 28976 18564 29028
rect 20352 28976 20404 29028
rect 20904 29019 20956 29028
rect 20904 28985 20913 29019
rect 20913 28985 20947 29019
rect 20947 28985 20956 29019
rect 20904 28976 20956 28985
rect 21640 28976 21692 29028
rect 26240 29044 26292 29096
rect 27804 29044 27856 29096
rect 28908 29044 28960 29096
rect 29276 29087 29328 29096
rect 29276 29053 29285 29087
rect 29285 29053 29319 29087
rect 29319 29053 29328 29087
rect 29276 29044 29328 29053
rect 25228 28976 25280 29028
rect 15016 28908 15068 28960
rect 17500 28908 17552 28960
rect 21548 28951 21600 28960
rect 21548 28917 21557 28951
rect 21557 28917 21591 28951
rect 21591 28917 21600 28951
rect 21548 28908 21600 28917
rect 21824 28951 21876 28960
rect 21824 28917 21833 28951
rect 21833 28917 21867 28951
rect 21867 28917 21876 28951
rect 21824 28908 21876 28917
rect 26608 29019 26660 29028
rect 25412 28908 25464 28960
rect 26608 28985 26617 29019
rect 26617 28985 26651 29019
rect 26651 28985 26660 29019
rect 26608 28976 26660 28985
rect 29000 28951 29052 28960
rect 29000 28917 29009 28951
rect 29009 28917 29043 28951
rect 29043 28917 29052 28951
rect 29000 28908 29052 28917
rect 30196 28908 30248 28960
rect 30380 28908 30432 28960
rect 31944 29112 31996 29164
rect 32956 29112 33008 29164
rect 35348 29112 35400 29164
rect 35440 29155 35492 29164
rect 35440 29121 35449 29155
rect 35449 29121 35483 29155
rect 35483 29121 35492 29155
rect 35440 29112 35492 29121
rect 36636 29087 36688 29096
rect 36636 29053 36645 29087
rect 36645 29053 36679 29087
rect 36679 29053 36688 29087
rect 36636 29044 36688 29053
rect 36820 29044 36872 29096
rect 37740 29112 37792 29164
rect 37832 29155 37884 29164
rect 37832 29121 37841 29155
rect 37841 29121 37875 29155
rect 37875 29121 37884 29155
rect 38568 29155 38620 29164
rect 37832 29112 37884 29121
rect 38568 29121 38577 29155
rect 38577 29121 38611 29155
rect 38611 29121 38620 29155
rect 38568 29112 38620 29121
rect 39396 29112 39448 29164
rect 32128 28951 32180 28960
rect 32128 28917 32137 28951
rect 32137 28917 32171 28951
rect 32171 28917 32180 28951
rect 32128 28908 32180 28917
rect 32956 29019 33008 29028
rect 32956 28985 32965 29019
rect 32965 28985 32999 29019
rect 32999 28985 33008 29019
rect 32956 28976 33008 28985
rect 35072 29019 35124 29028
rect 35072 28985 35081 29019
rect 35081 28985 35115 29019
rect 35115 28985 35124 29019
rect 35072 28976 35124 28985
rect 35440 28976 35492 29028
rect 36452 29019 36504 29028
rect 36452 28985 36461 29019
rect 36461 28985 36495 29019
rect 36495 28985 36504 29019
rect 36452 28976 36504 28985
rect 38292 29019 38344 29028
rect 38292 28985 38301 29019
rect 38301 28985 38335 29019
rect 38335 28985 38344 29019
rect 38292 28976 38344 28985
rect 38660 28976 38712 29028
rect 35532 28908 35584 28960
rect 44824 29257 44833 29291
rect 44833 29257 44867 29291
rect 44867 29257 44876 29291
rect 44824 29248 44876 29257
rect 42984 29180 43036 29232
rect 42432 29112 42484 29164
rect 42708 29155 42760 29164
rect 41052 29044 41104 29096
rect 42708 29121 42717 29155
rect 42717 29121 42751 29155
rect 42751 29121 42760 29155
rect 42708 29112 42760 29121
rect 43352 29112 43404 29164
rect 41236 29019 41288 29028
rect 41236 28985 41245 29019
rect 41245 28985 41279 29019
rect 41279 28985 41288 29019
rect 41236 28976 41288 28985
rect 43904 29019 43956 29028
rect 43904 28985 43913 29019
rect 43913 28985 43947 29019
rect 43947 28985 43956 29019
rect 43904 28976 43956 28985
rect 41144 28908 41196 28960
rect 43352 28951 43404 28960
rect 43352 28917 43361 28951
rect 43361 28917 43395 28951
rect 43395 28917 43404 28951
rect 43352 28908 43404 28917
rect 44364 28908 44416 28960
rect 45100 28951 45152 28960
rect 45100 28917 45109 28951
rect 45109 28917 45143 28951
rect 45143 28917 45152 28951
rect 45100 28908 45152 28917
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 9864 28747 9916 28756
rect 9864 28713 9873 28747
rect 9873 28713 9907 28747
rect 9907 28713 9916 28747
rect 9864 28704 9916 28713
rect 15016 28747 15068 28756
rect 15016 28713 15025 28747
rect 15025 28713 15059 28747
rect 15059 28713 15068 28747
rect 15016 28704 15068 28713
rect 12164 28679 12216 28688
rect 12164 28645 12173 28679
rect 12173 28645 12207 28679
rect 12207 28645 12216 28679
rect 12164 28636 12216 28645
rect 16304 28704 16356 28756
rect 21456 28704 21508 28756
rect 15476 28679 15528 28688
rect 15476 28645 15485 28679
rect 15485 28645 15519 28679
rect 15519 28645 15528 28679
rect 15476 28636 15528 28645
rect 17224 28636 17276 28688
rect 22192 28704 22244 28756
rect 29184 28704 29236 28756
rect 30104 28747 30156 28756
rect 30104 28713 30113 28747
rect 30113 28713 30147 28747
rect 30147 28713 30156 28747
rect 30104 28704 30156 28713
rect 30932 28704 30984 28756
rect 31300 28747 31352 28756
rect 31300 28713 31309 28747
rect 31309 28713 31343 28747
rect 31343 28713 31352 28747
rect 31300 28704 31352 28713
rect 31944 28747 31996 28756
rect 31944 28713 31953 28747
rect 31953 28713 31987 28747
rect 31987 28713 31996 28747
rect 31944 28704 31996 28713
rect 33416 28747 33468 28756
rect 33416 28713 33425 28747
rect 33425 28713 33459 28747
rect 33459 28713 33468 28747
rect 33416 28704 33468 28713
rect 34152 28704 34204 28756
rect 22468 28636 22520 28688
rect 23112 28679 23164 28688
rect 10324 28611 10376 28620
rect 10324 28577 10333 28611
rect 10333 28577 10367 28611
rect 10367 28577 10376 28611
rect 10324 28568 10376 28577
rect 10600 28568 10652 28620
rect 14280 28568 14332 28620
rect 17960 28568 18012 28620
rect 18604 28568 18656 28620
rect 23112 28645 23121 28679
rect 23121 28645 23155 28679
rect 23155 28645 23164 28679
rect 23112 28636 23164 28645
rect 25044 28679 25096 28688
rect 25044 28645 25053 28679
rect 25053 28645 25087 28679
rect 25087 28645 25096 28679
rect 25044 28636 25096 28645
rect 25596 28679 25648 28688
rect 25596 28645 25605 28679
rect 25605 28645 25639 28679
rect 25639 28645 25648 28679
rect 25596 28636 25648 28645
rect 26700 28679 26752 28688
rect 26700 28645 26709 28679
rect 26709 28645 26743 28679
rect 26743 28645 26752 28679
rect 26700 28636 26752 28645
rect 28908 28679 28960 28688
rect 28908 28645 28917 28679
rect 28917 28645 28951 28679
rect 28951 28645 28960 28679
rect 28908 28636 28960 28645
rect 32496 28636 32548 28688
rect 35072 28704 35124 28756
rect 36820 28704 36872 28756
rect 37740 28704 37792 28756
rect 38660 28704 38712 28756
rect 39580 28747 39632 28756
rect 39580 28713 39589 28747
rect 39589 28713 39623 28747
rect 39623 28713 39632 28747
rect 39580 28704 39632 28713
rect 41236 28704 41288 28756
rect 42432 28747 42484 28756
rect 42432 28713 42441 28747
rect 42441 28713 42475 28747
rect 42475 28713 42484 28747
rect 42432 28704 42484 28713
rect 43904 28747 43956 28756
rect 43904 28713 43913 28747
rect 43913 28713 43947 28747
rect 43947 28713 43956 28747
rect 43904 28704 43956 28713
rect 35256 28636 35308 28688
rect 38292 28636 38344 28688
rect 27896 28568 27948 28620
rect 28724 28611 28776 28620
rect 28724 28577 28733 28611
rect 28733 28577 28767 28611
rect 28767 28577 28776 28611
rect 28724 28568 28776 28577
rect 29368 28568 29420 28620
rect 30288 28568 30340 28620
rect 33048 28611 33100 28620
rect 33048 28577 33057 28611
rect 33057 28577 33091 28611
rect 33091 28577 33100 28611
rect 33048 28568 33100 28577
rect 33692 28568 33744 28620
rect 35624 28568 35676 28620
rect 36820 28568 36872 28620
rect 37188 28568 37240 28620
rect 38568 28568 38620 28620
rect 40684 28636 40736 28688
rect 41052 28636 41104 28688
rect 42708 28636 42760 28688
rect 10876 28543 10928 28552
rect 10876 28509 10885 28543
rect 10885 28509 10919 28543
rect 10919 28509 10928 28543
rect 10876 28500 10928 28509
rect 12072 28543 12124 28552
rect 12072 28509 12081 28543
rect 12081 28509 12115 28543
rect 12115 28509 12124 28543
rect 12072 28500 12124 28509
rect 12808 28500 12860 28552
rect 15660 28543 15712 28552
rect 15660 28509 15669 28543
rect 15669 28509 15703 28543
rect 15703 28509 15712 28543
rect 15660 28500 15712 28509
rect 17500 28500 17552 28552
rect 17592 28543 17644 28552
rect 17592 28509 17601 28543
rect 17601 28509 17635 28543
rect 17635 28509 17644 28543
rect 21180 28543 21232 28552
rect 17592 28500 17644 28509
rect 21180 28509 21189 28543
rect 21189 28509 21223 28543
rect 21223 28509 21232 28543
rect 21180 28500 21232 28509
rect 23296 28543 23348 28552
rect 23296 28509 23305 28543
rect 23305 28509 23339 28543
rect 23339 28509 23348 28543
rect 23296 28500 23348 28509
rect 24768 28543 24820 28552
rect 24768 28509 24777 28543
rect 24777 28509 24811 28543
rect 24811 28509 24820 28543
rect 24768 28500 24820 28509
rect 26608 28543 26660 28552
rect 26608 28509 26617 28543
rect 26617 28509 26651 28543
rect 26651 28509 26660 28543
rect 26608 28500 26660 28509
rect 29736 28543 29788 28552
rect 23664 28432 23716 28484
rect 25964 28432 26016 28484
rect 29736 28509 29745 28543
rect 29745 28509 29779 28543
rect 29779 28509 29788 28543
rect 29736 28500 29788 28509
rect 35256 28500 35308 28552
rect 35992 28500 36044 28552
rect 37648 28500 37700 28552
rect 39304 28500 39356 28552
rect 40224 28500 40276 28552
rect 41052 28543 41104 28552
rect 41052 28509 41061 28543
rect 41061 28509 41095 28543
rect 41095 28509 41104 28543
rect 41052 28500 41104 28509
rect 42340 28568 42392 28620
rect 43260 28611 43312 28620
rect 43260 28577 43269 28611
rect 43269 28577 43303 28611
rect 43303 28577 43312 28611
rect 43260 28568 43312 28577
rect 43628 28568 43680 28620
rect 44640 28568 44692 28620
rect 42524 28500 42576 28552
rect 42800 28500 42852 28552
rect 39580 28432 39632 28484
rect 41144 28432 41196 28484
rect 43352 28432 43404 28484
rect 10508 28364 10560 28416
rect 15016 28364 15068 28416
rect 18144 28407 18196 28416
rect 18144 28373 18153 28407
rect 18153 28373 18187 28407
rect 18187 28373 18196 28407
rect 18144 28364 18196 28373
rect 18696 28364 18748 28416
rect 19708 28407 19760 28416
rect 19708 28373 19717 28407
rect 19717 28373 19751 28407
rect 19751 28373 19760 28407
rect 19708 28364 19760 28373
rect 20352 28407 20404 28416
rect 20352 28373 20361 28407
rect 20361 28373 20395 28407
rect 20395 28373 20404 28407
rect 20352 28364 20404 28373
rect 23020 28364 23072 28416
rect 27712 28364 27764 28416
rect 32220 28364 32272 28416
rect 32864 28407 32916 28416
rect 32864 28373 32873 28407
rect 32873 28373 32907 28407
rect 32907 28373 32916 28407
rect 32864 28364 32916 28373
rect 37832 28364 37884 28416
rect 38936 28364 38988 28416
rect 41328 28364 41380 28416
rect 42248 28364 42300 28416
rect 43720 28364 43772 28416
rect 45468 28364 45520 28416
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 12532 28160 12584 28212
rect 17500 28160 17552 28212
rect 22560 28160 22612 28212
rect 23112 28203 23164 28212
rect 23112 28169 23121 28203
rect 23121 28169 23155 28203
rect 23155 28169 23164 28203
rect 23112 28160 23164 28169
rect 19708 28092 19760 28144
rect 24768 28160 24820 28212
rect 26608 28160 26660 28212
rect 27344 28160 27396 28212
rect 28632 28160 28684 28212
rect 29092 28160 29144 28212
rect 30196 28203 30248 28212
rect 30196 28169 30205 28203
rect 30205 28169 30239 28203
rect 30239 28169 30248 28203
rect 30196 28160 30248 28169
rect 32496 28160 32548 28212
rect 33692 28203 33744 28212
rect 33692 28169 33701 28203
rect 33701 28169 33735 28203
rect 33735 28169 33744 28203
rect 33692 28160 33744 28169
rect 34152 28160 34204 28212
rect 35900 28203 35952 28212
rect 25044 28092 25096 28144
rect 10508 28067 10560 28076
rect 10508 28033 10517 28067
rect 10517 28033 10551 28067
rect 10551 28033 10560 28067
rect 10508 28024 10560 28033
rect 11796 28024 11848 28076
rect 12164 28024 12216 28076
rect 13268 28024 13320 28076
rect 14188 28024 14240 28076
rect 15292 28024 15344 28076
rect 17592 28024 17644 28076
rect 21180 28067 21232 28076
rect 21180 28033 21189 28067
rect 21189 28033 21223 28067
rect 21223 28033 21232 28067
rect 21180 28024 21232 28033
rect 9864 27820 9916 27872
rect 11336 27956 11388 28008
rect 14280 27999 14332 28008
rect 14280 27965 14289 27999
rect 14289 27965 14323 27999
rect 14323 27965 14332 27999
rect 14280 27956 14332 27965
rect 17684 27956 17736 28008
rect 18144 27999 18196 28008
rect 18144 27965 18153 27999
rect 18153 27965 18187 27999
rect 18187 27965 18196 27999
rect 18144 27956 18196 27965
rect 11704 27888 11756 27940
rect 12532 27888 12584 27940
rect 11428 27863 11480 27872
rect 11428 27829 11437 27863
rect 11437 27829 11471 27863
rect 11471 27829 11480 27863
rect 11428 27820 11480 27829
rect 13084 27820 13136 27872
rect 13268 27931 13320 27940
rect 13268 27897 13277 27931
rect 13277 27897 13311 27931
rect 13311 27897 13320 27931
rect 15108 27931 15160 27940
rect 13268 27888 13320 27897
rect 15108 27897 15117 27931
rect 15117 27897 15151 27931
rect 15151 27897 15160 27931
rect 15108 27888 15160 27897
rect 13728 27820 13780 27872
rect 15476 27888 15528 27940
rect 15752 27931 15804 27940
rect 15752 27897 15761 27931
rect 15761 27897 15795 27931
rect 15795 27897 15804 27931
rect 15752 27888 15804 27897
rect 17224 27888 17276 27940
rect 18604 27888 18656 27940
rect 20904 27956 20956 28008
rect 21640 27956 21692 28008
rect 21732 27956 21784 28008
rect 22560 27956 22612 28008
rect 16948 27820 17000 27872
rect 18512 27863 18564 27872
rect 18512 27829 18521 27863
rect 18521 27829 18555 27863
rect 18555 27829 18564 27863
rect 18512 27820 18564 27829
rect 18788 27820 18840 27872
rect 20260 27863 20312 27872
rect 20260 27829 20269 27863
rect 20269 27829 20303 27863
rect 20303 27829 20312 27863
rect 20260 27820 20312 27829
rect 21456 27863 21508 27872
rect 21456 27829 21465 27863
rect 21465 27829 21499 27863
rect 21499 27829 21508 27863
rect 21456 27820 21508 27829
rect 22560 27820 22612 27872
rect 26700 28092 26752 28144
rect 32864 28092 32916 28144
rect 33416 28135 33468 28144
rect 33416 28101 33425 28135
rect 33425 28101 33459 28135
rect 33459 28101 33468 28135
rect 33416 28092 33468 28101
rect 25596 28024 25648 28076
rect 29184 28024 29236 28076
rect 26056 27999 26108 28008
rect 26056 27965 26065 27999
rect 26065 27965 26099 27999
rect 26099 27965 26108 27999
rect 27344 27999 27396 28008
rect 26056 27956 26108 27965
rect 27344 27965 27353 27999
rect 27353 27965 27387 27999
rect 27387 27965 27396 27999
rect 27344 27956 27396 27965
rect 25320 27820 25372 27872
rect 27896 27820 27948 27872
rect 28264 27820 28316 27872
rect 29000 27863 29052 27872
rect 29000 27829 29009 27863
rect 29009 27829 29043 27863
rect 29043 27829 29052 27863
rect 29736 27888 29788 27940
rect 29000 27820 29052 27829
rect 30104 27820 30156 27872
rect 32220 27956 32272 28008
rect 33416 27888 33468 27940
rect 35900 28169 35909 28203
rect 35909 28169 35943 28203
rect 35943 28169 35952 28203
rect 35900 28160 35952 28169
rect 37188 28203 37240 28212
rect 37188 28169 37197 28203
rect 37197 28169 37231 28203
rect 37231 28169 37240 28203
rect 37188 28160 37240 28169
rect 39304 28203 39356 28212
rect 39304 28169 39313 28203
rect 39313 28169 39347 28203
rect 39347 28169 39356 28203
rect 39304 28160 39356 28169
rect 40684 28203 40736 28212
rect 40684 28169 40693 28203
rect 40693 28169 40727 28203
rect 40727 28169 40736 28203
rect 40684 28160 40736 28169
rect 41144 28203 41196 28212
rect 41144 28169 41153 28203
rect 41153 28169 41187 28203
rect 41187 28169 41196 28203
rect 41144 28160 41196 28169
rect 43260 28160 43312 28212
rect 44640 28203 44692 28212
rect 44640 28169 44649 28203
rect 44649 28169 44683 28203
rect 44683 28169 44692 28203
rect 44640 28160 44692 28169
rect 38568 28092 38620 28144
rect 41328 28067 41380 28076
rect 41328 28033 41337 28067
rect 41337 28033 41371 28067
rect 41371 28033 41380 28067
rect 41328 28024 41380 28033
rect 43720 28067 43772 28076
rect 43720 28033 43729 28067
rect 43729 28033 43763 28067
rect 43763 28033 43772 28067
rect 43720 28024 43772 28033
rect 43812 28024 43864 28076
rect 31668 27863 31720 27872
rect 31668 27829 31677 27863
rect 31677 27829 31711 27863
rect 31711 27829 31720 27863
rect 31668 27820 31720 27829
rect 33232 27820 33284 27872
rect 36820 27820 36872 27872
rect 41880 27956 41932 28008
rect 38660 27888 38712 27940
rect 38844 27888 38896 27940
rect 41144 27888 41196 27940
rect 41512 27888 41564 27940
rect 38016 27820 38068 27872
rect 38752 27820 38804 27872
rect 40224 27863 40276 27872
rect 40224 27829 40233 27863
rect 40233 27829 40267 27863
rect 40267 27829 40276 27863
rect 40224 27820 40276 27829
rect 42524 27863 42576 27872
rect 42524 27829 42533 27863
rect 42533 27829 42567 27863
rect 42567 27829 42576 27863
rect 42524 27820 42576 27829
rect 43628 27820 43680 27872
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 11428 27616 11480 27668
rect 12624 27616 12676 27668
rect 10324 27548 10376 27600
rect 10876 27523 10928 27532
rect 10876 27489 10885 27523
rect 10885 27489 10919 27523
rect 10919 27489 10928 27523
rect 10876 27480 10928 27489
rect 11336 27548 11388 27600
rect 13728 27616 13780 27668
rect 14188 27591 14240 27600
rect 14188 27557 14197 27591
rect 14197 27557 14231 27591
rect 14231 27557 14240 27591
rect 14188 27548 14240 27557
rect 11796 27523 11848 27532
rect 11796 27489 11805 27523
rect 11805 27489 11839 27523
rect 11839 27489 11848 27523
rect 11796 27480 11848 27489
rect 13820 27412 13872 27464
rect 12164 27344 12216 27396
rect 12256 27387 12308 27396
rect 12256 27353 12265 27387
rect 12265 27353 12299 27387
rect 12299 27353 12308 27387
rect 20260 27616 20312 27668
rect 23664 27659 23716 27668
rect 23664 27625 23673 27659
rect 23673 27625 23707 27659
rect 23707 27625 23716 27659
rect 23664 27616 23716 27625
rect 25596 27659 25648 27668
rect 25596 27625 25605 27659
rect 25605 27625 25639 27659
rect 25639 27625 25648 27659
rect 25596 27616 25648 27625
rect 26608 27616 26660 27668
rect 32220 27659 32272 27668
rect 32220 27625 32229 27659
rect 32229 27625 32263 27659
rect 32263 27625 32272 27659
rect 32220 27616 32272 27625
rect 35256 27616 35308 27668
rect 38108 27659 38160 27668
rect 38108 27625 38117 27659
rect 38117 27625 38151 27659
rect 38151 27625 38160 27659
rect 38108 27616 38160 27625
rect 38660 27659 38712 27668
rect 38660 27625 38669 27659
rect 38669 27625 38703 27659
rect 38703 27625 38712 27659
rect 38660 27616 38712 27625
rect 39488 27616 39540 27668
rect 41512 27659 41564 27668
rect 15476 27591 15528 27600
rect 15476 27557 15485 27591
rect 15485 27557 15519 27591
rect 15519 27557 15528 27591
rect 15476 27548 15528 27557
rect 16948 27548 17000 27600
rect 17224 27591 17276 27600
rect 17224 27557 17233 27591
rect 17233 27557 17267 27591
rect 17267 27557 17276 27591
rect 17224 27548 17276 27557
rect 18696 27591 18748 27600
rect 18696 27557 18705 27591
rect 18705 27557 18739 27591
rect 18739 27557 18748 27591
rect 18696 27548 18748 27557
rect 18788 27591 18840 27600
rect 18788 27557 18797 27591
rect 18797 27557 18831 27591
rect 18831 27557 18840 27591
rect 18788 27548 18840 27557
rect 20444 27548 20496 27600
rect 22560 27548 22612 27600
rect 23020 27548 23072 27600
rect 25136 27591 25188 27600
rect 25136 27557 25145 27591
rect 25145 27557 25179 27591
rect 25179 27557 25188 27591
rect 25136 27548 25188 27557
rect 30380 27548 30432 27600
rect 34796 27548 34848 27600
rect 39580 27591 39632 27600
rect 39580 27557 39589 27591
rect 39589 27557 39623 27591
rect 39623 27557 39632 27591
rect 39580 27548 39632 27557
rect 41512 27625 41521 27659
rect 41521 27625 41555 27659
rect 41555 27625 41564 27659
rect 41512 27616 41564 27625
rect 42248 27616 42300 27668
rect 43628 27548 43680 27600
rect 45468 27591 45520 27600
rect 45468 27557 45477 27591
rect 45477 27557 45511 27591
rect 45511 27557 45520 27591
rect 45468 27548 45520 27557
rect 45560 27591 45612 27600
rect 45560 27557 45569 27591
rect 45569 27557 45603 27591
rect 45603 27557 45612 27591
rect 45560 27548 45612 27557
rect 21088 27523 21140 27532
rect 21088 27489 21097 27523
rect 21097 27489 21131 27523
rect 21131 27489 21140 27523
rect 21088 27480 21140 27489
rect 21640 27523 21692 27532
rect 21640 27489 21649 27523
rect 21649 27489 21683 27523
rect 21683 27489 21692 27523
rect 21640 27480 21692 27489
rect 24860 27480 24912 27532
rect 27252 27523 27304 27532
rect 27252 27489 27261 27523
rect 27261 27489 27295 27523
rect 27295 27489 27304 27523
rect 27252 27480 27304 27489
rect 28724 27480 28776 27532
rect 29368 27523 29420 27532
rect 29368 27489 29377 27523
rect 29377 27489 29411 27523
rect 29411 27489 29420 27523
rect 29368 27480 29420 27489
rect 29736 27480 29788 27532
rect 15384 27455 15436 27464
rect 15384 27421 15393 27455
rect 15393 27421 15427 27455
rect 15427 27421 15436 27455
rect 15384 27412 15436 27421
rect 15752 27455 15804 27464
rect 15752 27421 15761 27455
rect 15761 27421 15795 27455
rect 15795 27421 15804 27455
rect 15752 27412 15804 27421
rect 17132 27412 17184 27464
rect 18880 27412 18932 27464
rect 21824 27455 21876 27464
rect 21824 27421 21833 27455
rect 21833 27421 21867 27455
rect 21867 27421 21876 27455
rect 21824 27412 21876 27421
rect 27528 27412 27580 27464
rect 32312 27480 32364 27532
rect 32588 27523 32640 27532
rect 31208 27412 31260 27464
rect 32588 27489 32597 27523
rect 32597 27489 32631 27523
rect 32631 27489 32640 27523
rect 32588 27480 32640 27489
rect 34060 27480 34112 27532
rect 34704 27480 34756 27532
rect 36176 27523 36228 27532
rect 36176 27489 36185 27523
rect 36185 27489 36219 27523
rect 36219 27489 36228 27523
rect 36176 27480 36228 27489
rect 32864 27412 32916 27464
rect 35716 27412 35768 27464
rect 37096 27480 37148 27532
rect 38936 27480 38988 27532
rect 41052 27480 41104 27532
rect 37464 27412 37516 27464
rect 43904 27455 43956 27464
rect 23296 27387 23348 27396
rect 12256 27344 12308 27353
rect 23296 27353 23305 27387
rect 23305 27353 23339 27387
rect 23339 27353 23348 27387
rect 23296 27344 23348 27353
rect 28724 27344 28776 27396
rect 36636 27344 36688 27396
rect 39212 27344 39264 27396
rect 43904 27421 43913 27455
rect 43913 27421 43947 27455
rect 43947 27421 43956 27455
rect 43904 27412 43956 27421
rect 44824 27412 44876 27464
rect 43812 27344 43864 27396
rect 9956 27276 10008 27328
rect 10600 27276 10652 27328
rect 12072 27319 12124 27328
rect 12072 27285 12081 27319
rect 12081 27285 12115 27319
rect 12115 27285 12124 27319
rect 12072 27276 12124 27285
rect 13084 27319 13136 27328
rect 13084 27285 13093 27319
rect 13093 27285 13127 27319
rect 13127 27285 13136 27319
rect 13084 27276 13136 27285
rect 15108 27319 15160 27328
rect 15108 27285 15117 27319
rect 15117 27285 15151 27319
rect 15151 27285 15160 27319
rect 15108 27276 15160 27285
rect 18236 27276 18288 27328
rect 24952 27276 25004 27328
rect 27160 27276 27212 27328
rect 27620 27276 27672 27328
rect 30196 27319 30248 27328
rect 30196 27285 30205 27319
rect 30205 27285 30239 27319
rect 30239 27285 30248 27319
rect 30196 27276 30248 27285
rect 36728 27276 36780 27328
rect 40224 27276 40276 27328
rect 42064 27319 42116 27328
rect 42064 27285 42073 27319
rect 42073 27285 42107 27319
rect 42107 27285 42116 27319
rect 42064 27276 42116 27285
rect 43628 27319 43680 27328
rect 43628 27285 43637 27319
rect 43637 27285 43671 27319
rect 43671 27285 43680 27319
rect 43628 27276 43680 27285
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 10876 27072 10928 27124
rect 12164 27115 12216 27124
rect 12164 27081 12173 27115
rect 12173 27081 12207 27115
rect 12207 27081 12216 27115
rect 12164 27072 12216 27081
rect 10508 27004 10560 27056
rect 11152 27047 11204 27056
rect 11152 27013 11161 27047
rect 11161 27013 11195 27047
rect 11195 27013 11204 27047
rect 11152 27004 11204 27013
rect 11336 27004 11388 27056
rect 13820 27115 13872 27124
rect 13820 27081 13829 27115
rect 13829 27081 13863 27115
rect 13863 27081 13872 27115
rect 13820 27072 13872 27081
rect 15108 27072 15160 27124
rect 17224 27072 17276 27124
rect 18788 27072 18840 27124
rect 19156 27072 19208 27124
rect 20444 27072 20496 27124
rect 23020 27115 23072 27124
rect 23020 27081 23029 27115
rect 23029 27081 23063 27115
rect 23063 27081 23072 27115
rect 23020 27072 23072 27081
rect 24492 27072 24544 27124
rect 24860 27115 24912 27124
rect 24860 27081 24869 27115
rect 24869 27081 24903 27115
rect 24903 27081 24912 27115
rect 24860 27072 24912 27081
rect 27620 27072 27672 27124
rect 28724 27072 28776 27124
rect 29368 27072 29420 27124
rect 32588 27072 32640 27124
rect 34704 27115 34756 27124
rect 34704 27081 34713 27115
rect 34713 27081 34747 27115
rect 34747 27081 34756 27115
rect 34704 27072 34756 27081
rect 35716 27115 35768 27124
rect 35716 27081 35725 27115
rect 35725 27081 35759 27115
rect 35759 27081 35768 27115
rect 35716 27072 35768 27081
rect 38108 27072 38160 27124
rect 39488 27115 39540 27124
rect 39488 27081 39497 27115
rect 39497 27081 39531 27115
rect 39531 27081 39540 27115
rect 39488 27072 39540 27081
rect 39580 27072 39632 27124
rect 41512 27115 41564 27124
rect 41512 27081 41521 27115
rect 41521 27081 41555 27115
rect 41555 27081 41564 27115
rect 41512 27072 41564 27081
rect 42064 27072 42116 27124
rect 45468 27072 45520 27124
rect 12716 27004 12768 27056
rect 12808 26979 12860 26988
rect 12808 26945 12817 26979
rect 12817 26945 12851 26979
rect 12851 26945 12860 26979
rect 12808 26936 12860 26945
rect 15016 26979 15068 26988
rect 15016 26945 15025 26979
rect 15025 26945 15059 26979
rect 15059 26945 15068 26979
rect 15016 26936 15068 26945
rect 15660 26979 15712 26988
rect 15660 26945 15669 26979
rect 15669 26945 15703 26979
rect 15703 26945 15712 26979
rect 15660 26936 15712 26945
rect 9864 26868 9916 26920
rect 10416 26868 10468 26920
rect 20996 27004 21048 27056
rect 22560 27004 22612 27056
rect 25228 27004 25280 27056
rect 25964 27004 26016 27056
rect 26056 27004 26108 27056
rect 26792 27004 26844 27056
rect 20904 26936 20956 26988
rect 21824 26979 21876 26988
rect 21824 26945 21833 26979
rect 21833 26945 21867 26979
rect 21867 26945 21876 26979
rect 21824 26936 21876 26945
rect 26700 26936 26752 26988
rect 10600 26800 10652 26852
rect 12624 26843 12676 26852
rect 12624 26809 12633 26843
rect 12633 26809 12667 26843
rect 12667 26809 12676 26843
rect 12624 26800 12676 26809
rect 13268 26800 13320 26852
rect 9956 26775 10008 26784
rect 9956 26741 9965 26775
rect 9965 26741 9999 26775
rect 9999 26741 10008 26775
rect 9956 26732 10008 26741
rect 18236 26868 18288 26920
rect 20076 26868 20128 26920
rect 24400 26911 24452 26920
rect 24400 26877 24409 26911
rect 24409 26877 24443 26911
rect 24443 26877 24452 26911
rect 24400 26868 24452 26877
rect 28356 26868 28408 26920
rect 29092 26868 29144 26920
rect 32128 27004 32180 27056
rect 32404 26979 32456 26988
rect 32404 26945 32413 26979
rect 32413 26945 32447 26979
rect 32447 26945 32456 26979
rect 32404 26936 32456 26945
rect 39764 27004 39816 27056
rect 30196 26868 30248 26920
rect 15476 26732 15528 26784
rect 17868 26775 17920 26784
rect 17868 26741 17877 26775
rect 17877 26741 17911 26775
rect 17911 26741 17920 26775
rect 17868 26732 17920 26741
rect 18144 26775 18196 26784
rect 18144 26741 18153 26775
rect 18153 26741 18187 26775
rect 18187 26741 18196 26775
rect 18144 26732 18196 26741
rect 20536 26775 20588 26784
rect 20536 26741 20545 26775
rect 20545 26741 20579 26775
rect 20579 26741 20588 26775
rect 20536 26732 20588 26741
rect 21088 26775 21140 26784
rect 21088 26741 21097 26775
rect 21097 26741 21131 26775
rect 21131 26741 21140 26775
rect 21088 26732 21140 26741
rect 21456 26732 21508 26784
rect 24860 26800 24912 26852
rect 25136 26843 25188 26852
rect 25136 26809 25145 26843
rect 25145 26809 25179 26843
rect 25179 26809 25188 26843
rect 25136 26800 25188 26809
rect 22744 26732 22796 26784
rect 26976 26800 27028 26852
rect 30840 26843 30892 26852
rect 30840 26809 30849 26843
rect 30849 26809 30883 26843
rect 30883 26809 30892 26843
rect 30840 26800 30892 26809
rect 31668 26868 31720 26920
rect 33508 26936 33560 26988
rect 33876 26936 33928 26988
rect 33324 26868 33376 26920
rect 37096 26911 37148 26920
rect 33968 26843 34020 26852
rect 33968 26809 33977 26843
rect 33977 26809 34011 26843
rect 34011 26809 34020 26843
rect 33968 26800 34020 26809
rect 36452 26843 36504 26852
rect 36452 26809 36461 26843
rect 36461 26809 36495 26843
rect 36495 26809 36504 26843
rect 37096 26877 37105 26911
rect 37105 26877 37139 26911
rect 37139 26877 37148 26911
rect 37096 26868 37148 26877
rect 37372 26843 37424 26852
rect 36452 26800 36504 26809
rect 37372 26809 37381 26843
rect 37381 26809 37415 26843
rect 37415 26809 37424 26843
rect 37372 26800 37424 26809
rect 27252 26732 27304 26784
rect 27528 26775 27580 26784
rect 27528 26741 27537 26775
rect 27537 26741 27571 26775
rect 27571 26741 27580 26775
rect 27528 26732 27580 26741
rect 31208 26775 31260 26784
rect 31208 26741 31217 26775
rect 31217 26741 31251 26775
rect 31251 26741 31260 26775
rect 31208 26732 31260 26741
rect 32220 26732 32272 26784
rect 32864 26732 32916 26784
rect 34888 26775 34940 26784
rect 34888 26741 34897 26775
rect 34897 26741 34931 26775
rect 34931 26741 34940 26775
rect 34888 26732 34940 26741
rect 36176 26775 36228 26784
rect 36176 26741 36185 26775
rect 36185 26741 36219 26775
rect 36219 26741 36228 26775
rect 36176 26732 36228 26741
rect 38936 26936 38988 26988
rect 40224 26936 40276 26988
rect 41328 26936 41380 26988
rect 42248 26936 42300 26988
rect 42432 26979 42484 26988
rect 42432 26945 42441 26979
rect 42441 26945 42475 26979
rect 42475 26945 42484 26979
rect 42432 26936 42484 26945
rect 38660 26800 38712 26852
rect 39120 26800 39172 26852
rect 44272 26936 44324 26988
rect 45560 26936 45612 26988
rect 44180 26843 44232 26852
rect 42064 26732 42116 26784
rect 44180 26809 44189 26843
rect 44189 26809 44223 26843
rect 44223 26809 44232 26843
rect 44180 26800 44232 26809
rect 44272 26843 44324 26852
rect 44272 26809 44281 26843
rect 44281 26809 44315 26843
rect 44315 26809 44324 26843
rect 44824 26843 44876 26852
rect 44272 26800 44324 26809
rect 44824 26809 44833 26843
rect 44833 26809 44867 26843
rect 44867 26809 44876 26843
rect 44824 26800 44876 26809
rect 43628 26775 43680 26784
rect 43628 26741 43637 26775
rect 43637 26741 43671 26775
rect 43671 26741 43680 26775
rect 43628 26732 43680 26741
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 13084 26528 13136 26580
rect 15016 26571 15068 26580
rect 15016 26537 15025 26571
rect 15025 26537 15059 26571
rect 15059 26537 15068 26571
rect 15016 26528 15068 26537
rect 15384 26528 15436 26580
rect 16948 26528 17000 26580
rect 18788 26528 18840 26580
rect 20076 26528 20128 26580
rect 21824 26571 21876 26580
rect 21824 26537 21833 26571
rect 21833 26537 21867 26571
rect 21867 26537 21876 26571
rect 21824 26528 21876 26537
rect 24860 26528 24912 26580
rect 26700 26571 26752 26580
rect 26700 26537 26709 26571
rect 26709 26537 26743 26571
rect 26743 26537 26752 26571
rect 26700 26528 26752 26537
rect 28356 26571 28408 26580
rect 28356 26537 28365 26571
rect 28365 26537 28399 26571
rect 28399 26537 28408 26571
rect 28356 26528 28408 26537
rect 11336 26460 11388 26512
rect 12072 26460 12124 26512
rect 16028 26503 16080 26512
rect 16028 26469 16037 26503
rect 16037 26469 16071 26503
rect 16071 26469 16080 26503
rect 16028 26460 16080 26469
rect 16212 26460 16264 26512
rect 10048 26392 10100 26444
rect 10508 26435 10560 26444
rect 10508 26401 10517 26435
rect 10517 26401 10551 26435
rect 10551 26401 10560 26435
rect 10508 26392 10560 26401
rect 12808 26392 12860 26444
rect 13176 26392 13228 26444
rect 14372 26392 14424 26444
rect 17500 26435 17552 26444
rect 17500 26401 17509 26435
rect 17509 26401 17543 26435
rect 17543 26401 17552 26435
rect 17500 26392 17552 26401
rect 18236 26392 18288 26444
rect 19524 26392 19576 26444
rect 22744 26460 22796 26512
rect 24952 26503 25004 26512
rect 24952 26469 24961 26503
rect 24961 26469 24995 26503
rect 24995 26469 25004 26503
rect 24952 26460 25004 26469
rect 25136 26460 25188 26512
rect 25688 26460 25740 26512
rect 27988 26503 28040 26512
rect 27988 26469 27997 26503
rect 27997 26469 28031 26503
rect 28031 26469 28040 26503
rect 30196 26528 30248 26580
rect 30840 26571 30892 26580
rect 30840 26537 30849 26571
rect 30849 26537 30883 26571
rect 30883 26537 30892 26571
rect 30840 26528 30892 26537
rect 33968 26528 34020 26580
rect 34796 26571 34848 26580
rect 34796 26537 34805 26571
rect 34805 26537 34839 26571
rect 34839 26537 34848 26571
rect 34796 26528 34848 26537
rect 35348 26528 35400 26580
rect 37096 26571 37148 26580
rect 37096 26537 37105 26571
rect 37105 26537 37139 26571
rect 37139 26537 37148 26571
rect 37096 26528 37148 26537
rect 37464 26571 37516 26580
rect 37464 26537 37473 26571
rect 37473 26537 37507 26571
rect 37507 26537 37516 26571
rect 37464 26528 37516 26537
rect 41052 26528 41104 26580
rect 43904 26528 43956 26580
rect 44180 26528 44232 26580
rect 27988 26460 28040 26469
rect 28908 26460 28960 26512
rect 32312 26503 32364 26512
rect 32312 26469 32321 26503
rect 32321 26469 32355 26503
rect 32355 26469 32364 26503
rect 32312 26460 32364 26469
rect 32496 26460 32548 26512
rect 35808 26460 35860 26512
rect 38108 26460 38160 26512
rect 41880 26503 41932 26512
rect 41880 26469 41889 26503
rect 41889 26469 41923 26503
rect 41923 26469 41932 26503
rect 41880 26460 41932 26469
rect 42156 26460 42208 26512
rect 21088 26392 21140 26444
rect 11888 26324 11940 26376
rect 15200 26324 15252 26376
rect 18052 26367 18104 26376
rect 15660 26256 15712 26308
rect 18052 26333 18061 26367
rect 18061 26333 18095 26367
rect 18095 26333 18104 26367
rect 18052 26324 18104 26333
rect 19156 26324 19208 26376
rect 19616 26367 19668 26376
rect 19616 26333 19625 26367
rect 19625 26333 19659 26367
rect 19659 26333 19668 26367
rect 19616 26324 19668 26333
rect 19984 26324 20036 26376
rect 22192 26324 22244 26376
rect 23940 26392 23992 26444
rect 27252 26435 27304 26444
rect 27252 26401 27261 26435
rect 27261 26401 27295 26435
rect 27295 26401 27304 26435
rect 27252 26392 27304 26401
rect 29092 26392 29144 26444
rect 30932 26435 30984 26444
rect 30932 26401 30941 26435
rect 30941 26401 30975 26435
rect 30975 26401 30984 26435
rect 30932 26392 30984 26401
rect 33968 26435 34020 26444
rect 33968 26401 33977 26435
rect 33977 26401 34011 26435
rect 34011 26401 34020 26435
rect 33968 26392 34020 26401
rect 36544 26435 36596 26444
rect 36544 26401 36553 26435
rect 36553 26401 36587 26435
rect 36587 26401 36596 26435
rect 36544 26392 36596 26401
rect 37372 26392 37424 26444
rect 39764 26435 39816 26444
rect 39764 26401 39773 26435
rect 39773 26401 39807 26435
rect 39807 26401 39816 26435
rect 39764 26392 39816 26401
rect 40224 26435 40276 26444
rect 40224 26401 40233 26435
rect 40233 26401 40267 26435
rect 40267 26401 40276 26435
rect 40224 26392 40276 26401
rect 44272 26460 44324 26512
rect 43720 26392 43772 26444
rect 44364 26435 44416 26444
rect 44364 26401 44373 26435
rect 44373 26401 44407 26435
rect 44407 26401 44416 26435
rect 44364 26392 44416 26401
rect 27620 26367 27672 26376
rect 27620 26333 27629 26367
rect 27629 26333 27663 26367
rect 27663 26333 27672 26367
rect 27620 26324 27672 26333
rect 29276 26367 29328 26376
rect 29276 26333 29285 26367
rect 29285 26333 29319 26367
rect 29319 26333 29328 26367
rect 29276 26324 29328 26333
rect 30012 26324 30064 26376
rect 31852 26324 31904 26376
rect 17776 26256 17828 26308
rect 20444 26256 20496 26308
rect 34888 26324 34940 26376
rect 36084 26324 36136 26376
rect 40500 26367 40552 26376
rect 40500 26333 40509 26367
rect 40509 26333 40543 26367
rect 40543 26333 40552 26367
rect 40500 26324 40552 26333
rect 41788 26367 41840 26376
rect 41788 26333 41797 26367
rect 41797 26333 41831 26367
rect 41831 26333 41840 26367
rect 41788 26324 41840 26333
rect 42064 26367 42116 26376
rect 42064 26333 42073 26367
rect 42073 26333 42107 26367
rect 42107 26333 42116 26367
rect 42064 26324 42116 26333
rect 42432 26324 42484 26376
rect 35256 26256 35308 26308
rect 35624 26299 35676 26308
rect 35624 26265 35633 26299
rect 35633 26265 35667 26299
rect 35667 26265 35676 26299
rect 35624 26256 35676 26265
rect 9864 26188 9916 26240
rect 18972 26231 19024 26240
rect 18972 26197 18981 26231
rect 18981 26197 19015 26231
rect 19015 26197 19024 26231
rect 18972 26188 19024 26197
rect 21640 26188 21692 26240
rect 22100 26188 22152 26240
rect 23020 26231 23072 26240
rect 23020 26197 23029 26231
rect 23029 26197 23063 26231
rect 23063 26197 23072 26231
rect 23020 26188 23072 26197
rect 26516 26188 26568 26240
rect 27160 26231 27212 26240
rect 27160 26197 27169 26231
rect 27169 26197 27203 26231
rect 27203 26197 27212 26231
rect 27160 26188 27212 26197
rect 27804 26188 27856 26240
rect 33324 26231 33376 26240
rect 33324 26197 33333 26231
rect 33333 26197 33367 26231
rect 33367 26197 33376 26231
rect 33324 26188 33376 26197
rect 34704 26188 34756 26240
rect 38936 26231 38988 26240
rect 38936 26197 38945 26231
rect 38945 26197 38979 26231
rect 38979 26197 38988 26231
rect 38936 26188 38988 26197
rect 39212 26231 39264 26240
rect 39212 26197 39221 26231
rect 39221 26197 39255 26231
rect 39255 26197 39264 26231
rect 39212 26188 39264 26197
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 10232 25984 10284 26036
rect 11888 26027 11940 26036
rect 11888 25993 11897 26027
rect 11897 25993 11931 26027
rect 11931 25993 11940 26027
rect 11888 25984 11940 25993
rect 14372 25984 14424 26036
rect 17684 25984 17736 26036
rect 19616 26027 19668 26036
rect 19616 25993 19625 26027
rect 19625 25993 19659 26027
rect 19659 25993 19668 26027
rect 19616 25984 19668 25993
rect 20444 25984 20496 26036
rect 25136 25984 25188 26036
rect 11336 25916 11388 25968
rect 14924 25916 14976 25968
rect 16028 25916 16080 25968
rect 17500 25959 17552 25968
rect 17500 25925 17509 25959
rect 17509 25925 17543 25959
rect 17543 25925 17552 25959
rect 17500 25916 17552 25925
rect 19248 25916 19300 25968
rect 23940 25959 23992 25968
rect 13268 25891 13320 25900
rect 13268 25857 13277 25891
rect 13277 25857 13311 25891
rect 13311 25857 13320 25891
rect 15292 25891 15344 25900
rect 13268 25848 13320 25857
rect 15292 25857 15301 25891
rect 15301 25857 15335 25891
rect 15335 25857 15344 25891
rect 15292 25848 15344 25857
rect 16856 25848 16908 25900
rect 17132 25848 17184 25900
rect 17776 25848 17828 25900
rect 18880 25848 18932 25900
rect 23940 25925 23949 25959
rect 23949 25925 23983 25959
rect 23983 25925 23992 25959
rect 28540 25984 28592 26036
rect 29276 25984 29328 26036
rect 36084 26027 36136 26036
rect 36084 25993 36093 26027
rect 36093 25993 36127 26027
rect 36127 25993 36136 26027
rect 36084 25984 36136 25993
rect 37372 25984 37424 26036
rect 38936 25984 38988 26036
rect 39764 25984 39816 26036
rect 41788 25984 41840 26036
rect 43720 26027 43772 26036
rect 43720 25993 43729 26027
rect 43729 25993 43763 26027
rect 43763 25993 43772 26027
rect 43720 25984 43772 25993
rect 23940 25916 23992 25925
rect 22192 25891 22244 25900
rect 22192 25857 22201 25891
rect 22201 25857 22235 25891
rect 22235 25857 22244 25891
rect 22192 25848 22244 25857
rect 25228 25848 25280 25900
rect 25412 25891 25464 25900
rect 25412 25857 25421 25891
rect 25421 25857 25455 25891
rect 25455 25857 25464 25891
rect 25412 25848 25464 25857
rect 26516 25891 26568 25900
rect 26516 25857 26525 25891
rect 26525 25857 26559 25891
rect 26559 25857 26568 25891
rect 26516 25848 26568 25857
rect 26792 25848 26844 25900
rect 30932 25916 30984 25968
rect 31208 25916 31260 25968
rect 36452 25916 36504 25968
rect 36544 25959 36596 25968
rect 36544 25925 36553 25959
rect 36553 25925 36587 25959
rect 36587 25925 36596 25959
rect 36544 25916 36596 25925
rect 40040 25916 40092 25968
rect 41880 25916 41932 25968
rect 44732 25984 44784 26036
rect 28356 25848 28408 25900
rect 29000 25848 29052 25900
rect 30656 25848 30708 25900
rect 30840 25848 30892 25900
rect 32220 25848 32272 25900
rect 34796 25848 34848 25900
rect 35348 25848 35400 25900
rect 36728 25891 36780 25900
rect 36728 25857 36737 25891
rect 36737 25857 36771 25891
rect 36771 25857 36780 25891
rect 36728 25848 36780 25857
rect 36912 25848 36964 25900
rect 39212 25848 39264 25900
rect 42064 25848 42116 25900
rect 10232 25823 10284 25832
rect 10232 25789 10241 25823
rect 10241 25789 10275 25823
rect 10275 25789 10284 25823
rect 10232 25780 10284 25789
rect 10600 25823 10652 25832
rect 10600 25789 10609 25823
rect 10609 25789 10643 25823
rect 10643 25789 10652 25823
rect 10600 25780 10652 25789
rect 20076 25823 20128 25832
rect 20076 25789 20085 25823
rect 20085 25789 20119 25823
rect 20119 25789 20128 25823
rect 20076 25780 20128 25789
rect 20536 25823 20588 25832
rect 20536 25789 20545 25823
rect 20545 25789 20579 25823
rect 20579 25789 20588 25823
rect 20536 25780 20588 25789
rect 21640 25823 21692 25832
rect 21640 25789 21649 25823
rect 21649 25789 21683 25823
rect 21683 25789 21692 25823
rect 21640 25780 21692 25789
rect 22100 25823 22152 25832
rect 22100 25789 22109 25823
rect 22109 25789 22143 25823
rect 22143 25789 22152 25823
rect 22100 25780 22152 25789
rect 28540 25780 28592 25832
rect 28816 25780 28868 25832
rect 31484 25780 31536 25832
rect 33232 25823 33284 25832
rect 33232 25789 33241 25823
rect 33241 25789 33275 25823
rect 33275 25789 33284 25823
rect 33232 25780 33284 25789
rect 35624 25780 35676 25832
rect 43352 25780 43404 25832
rect 43996 25891 44048 25900
rect 43996 25857 44005 25891
rect 44005 25857 44039 25891
rect 44039 25857 44048 25891
rect 43996 25848 44048 25857
rect 44088 25848 44140 25900
rect 10784 25755 10836 25764
rect 10784 25721 10793 25755
rect 10793 25721 10827 25755
rect 10827 25721 10836 25755
rect 10784 25712 10836 25721
rect 13544 25712 13596 25764
rect 13912 25755 13964 25764
rect 13912 25721 13921 25755
rect 13921 25721 13955 25755
rect 13955 25721 13964 25755
rect 13912 25712 13964 25721
rect 14832 25755 14884 25764
rect 14832 25721 14841 25755
rect 14841 25721 14875 25755
rect 14875 25721 14884 25755
rect 14832 25712 14884 25721
rect 14924 25755 14976 25764
rect 14924 25721 14933 25755
rect 14933 25721 14967 25755
rect 14967 25721 14976 25755
rect 14924 25712 14976 25721
rect 16028 25712 16080 25764
rect 16488 25755 16540 25764
rect 16488 25721 16497 25755
rect 16497 25721 16531 25755
rect 16531 25721 16540 25755
rect 16488 25712 16540 25721
rect 18972 25712 19024 25764
rect 19064 25712 19116 25764
rect 22284 25712 22336 25764
rect 24768 25712 24820 25764
rect 9404 25644 9456 25696
rect 10508 25644 10560 25696
rect 11060 25687 11112 25696
rect 11060 25653 11069 25687
rect 11069 25653 11103 25687
rect 11103 25653 11112 25687
rect 11060 25644 11112 25653
rect 11336 25644 11388 25696
rect 13176 25644 13228 25696
rect 18236 25687 18288 25696
rect 18236 25653 18245 25687
rect 18245 25653 18279 25687
rect 18279 25653 18288 25687
rect 18236 25644 18288 25653
rect 20168 25687 20220 25696
rect 20168 25653 20177 25687
rect 20177 25653 20211 25687
rect 20211 25653 20220 25687
rect 20168 25644 20220 25653
rect 20628 25644 20680 25696
rect 21640 25644 21692 25696
rect 22744 25687 22796 25696
rect 22744 25653 22753 25687
rect 22753 25653 22787 25687
rect 22787 25653 22796 25687
rect 22744 25644 22796 25653
rect 26516 25712 26568 25764
rect 26700 25712 26752 25764
rect 30656 25712 30708 25764
rect 26884 25644 26936 25696
rect 27620 25687 27672 25696
rect 27620 25653 27629 25687
rect 27629 25653 27663 25687
rect 27663 25653 27672 25687
rect 27620 25644 27672 25653
rect 27804 25644 27856 25696
rect 28540 25644 28592 25696
rect 28908 25644 28960 25696
rect 31668 25687 31720 25696
rect 31668 25653 31677 25687
rect 31677 25653 31711 25687
rect 31711 25653 31720 25687
rect 31668 25644 31720 25653
rect 32312 25687 32364 25696
rect 32312 25653 32321 25687
rect 32321 25653 32355 25687
rect 32355 25653 32364 25687
rect 32312 25644 32364 25653
rect 33416 25644 33468 25696
rect 33968 25687 34020 25696
rect 33968 25653 33977 25687
rect 33977 25653 34011 25687
rect 34011 25653 34020 25687
rect 33968 25644 34020 25653
rect 34428 25644 34480 25696
rect 37004 25712 37056 25764
rect 39028 25755 39080 25764
rect 39028 25721 39037 25755
rect 39037 25721 39071 25755
rect 39071 25721 39080 25755
rect 39580 25755 39632 25764
rect 39028 25712 39080 25721
rect 39580 25721 39589 25755
rect 39589 25721 39623 25755
rect 39623 25721 39632 25755
rect 39580 25712 39632 25721
rect 39764 25712 39816 25764
rect 40224 25755 40276 25764
rect 40224 25721 40233 25755
rect 40233 25721 40267 25755
rect 40267 25721 40276 25755
rect 40224 25712 40276 25721
rect 41420 25755 41472 25764
rect 41420 25721 41429 25755
rect 41429 25721 41463 25755
rect 41463 25721 41472 25755
rect 41420 25712 41472 25721
rect 35808 25687 35860 25696
rect 35808 25653 35817 25687
rect 35817 25653 35851 25687
rect 35851 25653 35860 25687
rect 35808 25644 35860 25653
rect 38108 25687 38160 25696
rect 38108 25653 38117 25687
rect 38117 25653 38151 25687
rect 38151 25653 38160 25687
rect 38108 25644 38160 25653
rect 44272 25712 44324 25764
rect 41696 25644 41748 25696
rect 43812 25644 43864 25696
rect 44364 25644 44416 25696
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 11336 25483 11388 25492
rect 11336 25449 11345 25483
rect 11345 25449 11379 25483
rect 11379 25449 11388 25483
rect 11336 25440 11388 25449
rect 14832 25440 14884 25492
rect 16488 25483 16540 25492
rect 16488 25449 16497 25483
rect 16497 25449 16531 25483
rect 16531 25449 16540 25483
rect 16488 25440 16540 25449
rect 17776 25483 17828 25492
rect 17776 25449 17785 25483
rect 17785 25449 17819 25483
rect 17819 25449 17828 25483
rect 17776 25440 17828 25449
rect 18972 25440 19024 25492
rect 19156 25440 19208 25492
rect 20076 25483 20128 25492
rect 10324 25372 10376 25424
rect 11152 25372 11204 25424
rect 10232 25304 10284 25356
rect 11888 25304 11940 25356
rect 10784 25236 10836 25288
rect 10048 25143 10100 25152
rect 10048 25109 10057 25143
rect 10057 25109 10091 25143
rect 10091 25109 10100 25143
rect 10048 25100 10100 25109
rect 12072 25100 12124 25152
rect 13268 25372 13320 25424
rect 15292 25372 15344 25424
rect 15476 25372 15528 25424
rect 18512 25372 18564 25424
rect 13636 25304 13688 25356
rect 14188 25347 14240 25356
rect 14188 25313 14232 25347
rect 14232 25313 14240 25347
rect 14188 25304 14240 25313
rect 18052 25304 18104 25356
rect 20076 25449 20085 25483
rect 20085 25449 20119 25483
rect 20119 25449 20128 25483
rect 20076 25440 20128 25449
rect 22192 25483 22244 25492
rect 22192 25449 22201 25483
rect 22201 25449 22235 25483
rect 22235 25449 22244 25483
rect 22192 25440 22244 25449
rect 24952 25440 25004 25492
rect 25228 25440 25280 25492
rect 26792 25483 26844 25492
rect 26792 25449 26801 25483
rect 26801 25449 26835 25483
rect 26835 25449 26844 25483
rect 26792 25440 26844 25449
rect 28356 25483 28408 25492
rect 28356 25449 28365 25483
rect 28365 25449 28399 25483
rect 28399 25449 28408 25483
rect 28356 25440 28408 25449
rect 31852 25483 31904 25492
rect 31852 25449 31861 25483
rect 31861 25449 31895 25483
rect 31895 25449 31904 25483
rect 31852 25440 31904 25449
rect 34520 25440 34572 25492
rect 19432 25372 19484 25424
rect 23020 25372 23072 25424
rect 25044 25415 25096 25424
rect 25044 25381 25053 25415
rect 25053 25381 25087 25415
rect 25087 25381 25096 25415
rect 25044 25372 25096 25381
rect 25136 25372 25188 25424
rect 25688 25372 25740 25424
rect 29920 25415 29972 25424
rect 29920 25381 29929 25415
rect 29929 25381 29963 25415
rect 29963 25381 29972 25415
rect 29920 25372 29972 25381
rect 32312 25415 32364 25424
rect 32312 25381 32321 25415
rect 32321 25381 32355 25415
rect 32355 25381 32364 25415
rect 32312 25372 32364 25381
rect 34704 25372 34756 25424
rect 36728 25440 36780 25492
rect 41420 25483 41472 25492
rect 41420 25449 41429 25483
rect 41429 25449 41463 25483
rect 41463 25449 41472 25483
rect 41420 25440 41472 25449
rect 35808 25372 35860 25424
rect 37004 25415 37056 25424
rect 37004 25381 37013 25415
rect 37013 25381 37047 25415
rect 37047 25381 37056 25415
rect 37004 25372 37056 25381
rect 38936 25415 38988 25424
rect 38936 25381 38945 25415
rect 38945 25381 38979 25415
rect 38979 25381 38988 25415
rect 38936 25372 38988 25381
rect 41696 25415 41748 25424
rect 41696 25381 41705 25415
rect 41705 25381 41739 25415
rect 41739 25381 41748 25415
rect 41696 25372 41748 25381
rect 43628 25372 43680 25424
rect 12808 25236 12860 25288
rect 15108 25236 15160 25288
rect 20352 25304 20404 25356
rect 26424 25304 26476 25356
rect 27068 25304 27120 25356
rect 33600 25304 33652 25356
rect 36452 25304 36504 25356
rect 37648 25304 37700 25356
rect 40316 25304 40368 25356
rect 20076 25236 20128 25288
rect 23296 25279 23348 25288
rect 23296 25245 23305 25279
rect 23305 25245 23339 25279
rect 23339 25245 23348 25279
rect 23296 25236 23348 25245
rect 25136 25236 25188 25288
rect 13912 25168 13964 25220
rect 16304 25168 16356 25220
rect 25412 25236 25464 25288
rect 28172 25236 28224 25288
rect 28540 25236 28592 25288
rect 30104 25236 30156 25288
rect 32588 25236 32640 25288
rect 29368 25168 29420 25220
rect 30380 25211 30432 25220
rect 30380 25177 30389 25211
rect 30389 25177 30423 25211
rect 30423 25177 30432 25211
rect 35808 25236 35860 25288
rect 38844 25279 38896 25288
rect 38844 25245 38853 25279
rect 38853 25245 38887 25279
rect 38887 25245 38896 25279
rect 38844 25236 38896 25245
rect 39028 25236 39080 25288
rect 39580 25236 39632 25288
rect 41604 25279 41656 25288
rect 41604 25245 41613 25279
rect 41613 25245 41647 25279
rect 41647 25245 41656 25279
rect 41604 25236 41656 25245
rect 30380 25168 30432 25177
rect 15200 25100 15252 25152
rect 16212 25143 16264 25152
rect 16212 25109 16221 25143
rect 16221 25109 16255 25143
rect 16255 25109 16264 25143
rect 16212 25100 16264 25109
rect 16856 25143 16908 25152
rect 16856 25109 16865 25143
rect 16865 25109 16899 25143
rect 16899 25109 16908 25143
rect 16856 25100 16908 25109
rect 19340 25100 19392 25152
rect 20536 25100 20588 25152
rect 22100 25100 22152 25152
rect 22652 25100 22704 25152
rect 23940 25100 23992 25152
rect 26516 25100 26568 25152
rect 27252 25100 27304 25152
rect 28908 25143 28960 25152
rect 28908 25109 28917 25143
rect 28917 25109 28951 25143
rect 28951 25109 28960 25143
rect 28908 25100 28960 25109
rect 30932 25100 30984 25152
rect 35440 25168 35492 25220
rect 35992 25168 36044 25220
rect 39212 25168 39264 25220
rect 43720 25236 43772 25288
rect 44640 25236 44692 25288
rect 44088 25168 44140 25220
rect 34704 25100 34756 25152
rect 36544 25100 36596 25152
rect 38200 25143 38252 25152
rect 38200 25109 38209 25143
rect 38209 25109 38243 25143
rect 38243 25109 38252 25143
rect 38200 25100 38252 25109
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 10324 24939 10376 24948
rect 10324 24905 10333 24939
rect 10333 24905 10367 24939
rect 10367 24905 10376 24939
rect 10324 24896 10376 24905
rect 12808 24896 12860 24948
rect 13544 24939 13596 24948
rect 13544 24905 13553 24939
rect 13553 24905 13587 24939
rect 13587 24905 13596 24939
rect 13544 24896 13596 24905
rect 14556 24896 14608 24948
rect 15476 24939 15528 24948
rect 15476 24905 15485 24939
rect 15485 24905 15519 24939
rect 15519 24905 15528 24939
rect 15476 24896 15528 24905
rect 18052 24896 18104 24948
rect 23020 24939 23072 24948
rect 23020 24905 23029 24939
rect 23029 24905 23063 24939
rect 23063 24905 23072 24939
rect 23020 24896 23072 24905
rect 25044 24896 25096 24948
rect 26608 24939 26660 24948
rect 26608 24905 26617 24939
rect 26617 24905 26651 24939
rect 26651 24905 26660 24939
rect 26608 24896 26660 24905
rect 27068 24939 27120 24948
rect 27068 24905 27077 24939
rect 27077 24905 27111 24939
rect 27111 24905 27120 24939
rect 27068 24896 27120 24905
rect 34520 24896 34572 24948
rect 34796 24896 34848 24948
rect 36452 24896 36504 24948
rect 37004 24896 37056 24948
rect 37648 24896 37700 24948
rect 38936 24939 38988 24948
rect 38936 24905 38945 24939
rect 38945 24905 38979 24939
rect 38979 24905 38988 24939
rect 38936 24896 38988 24905
rect 39488 24896 39540 24948
rect 40316 24896 40368 24948
rect 41696 24939 41748 24948
rect 41696 24905 41705 24939
rect 41705 24905 41739 24939
rect 41739 24905 41748 24939
rect 41696 24896 41748 24905
rect 43628 24939 43680 24948
rect 43628 24905 43637 24939
rect 43637 24905 43671 24939
rect 43671 24905 43680 24939
rect 43628 24896 43680 24905
rect 43996 24896 44048 24948
rect 44456 24896 44508 24948
rect 44640 24939 44692 24948
rect 44640 24905 44649 24939
rect 44649 24905 44683 24939
rect 44683 24905 44692 24939
rect 44640 24896 44692 24905
rect 11244 24828 11296 24880
rect 10048 24760 10100 24812
rect 10600 24760 10652 24812
rect 10416 24735 10468 24744
rect 10416 24701 10425 24735
rect 10425 24701 10459 24735
rect 10459 24701 10468 24735
rect 10416 24692 10468 24701
rect 12624 24735 12676 24744
rect 12624 24701 12633 24735
rect 12633 24701 12667 24735
rect 12667 24701 12676 24735
rect 12624 24692 12676 24701
rect 14372 24735 14424 24744
rect 14372 24701 14381 24735
rect 14381 24701 14415 24735
rect 14415 24701 14424 24735
rect 14372 24692 14424 24701
rect 18236 24828 18288 24880
rect 16120 24760 16172 24812
rect 17132 24760 17184 24812
rect 18512 24760 18564 24812
rect 20168 24803 20220 24812
rect 11152 24667 11204 24676
rect 11152 24633 11161 24667
rect 11161 24633 11195 24667
rect 11195 24633 11204 24667
rect 11152 24624 11204 24633
rect 13452 24624 13504 24676
rect 17868 24692 17920 24744
rect 18052 24735 18104 24744
rect 18052 24701 18061 24735
rect 18061 24701 18095 24735
rect 18095 24701 18104 24735
rect 18052 24692 18104 24701
rect 20168 24769 20177 24803
rect 20177 24769 20211 24803
rect 20211 24769 20220 24803
rect 20168 24760 20220 24769
rect 15108 24667 15160 24676
rect 15108 24633 15117 24667
rect 15117 24633 15151 24667
rect 15151 24633 15160 24667
rect 15108 24624 15160 24633
rect 14188 24599 14240 24608
rect 14188 24565 14197 24599
rect 14197 24565 14231 24599
rect 14231 24565 14240 24599
rect 14188 24556 14240 24565
rect 16212 24624 16264 24676
rect 16304 24624 16356 24676
rect 19064 24624 19116 24676
rect 18144 24599 18196 24608
rect 18144 24565 18153 24599
rect 18153 24565 18187 24599
rect 18187 24565 18196 24599
rect 18144 24556 18196 24565
rect 19340 24556 19392 24608
rect 21272 24692 21324 24744
rect 27896 24828 27948 24880
rect 23940 24803 23992 24812
rect 23940 24769 23949 24803
rect 23949 24769 23983 24803
rect 23983 24769 23992 24803
rect 23940 24760 23992 24769
rect 29368 24803 29420 24812
rect 29368 24769 29377 24803
rect 29377 24769 29411 24803
rect 29411 24769 29420 24803
rect 29368 24760 29420 24769
rect 29828 24760 29880 24812
rect 22652 24692 22704 24744
rect 25688 24735 25740 24744
rect 25688 24701 25697 24735
rect 25697 24701 25731 24735
rect 25731 24701 25740 24735
rect 25688 24692 25740 24701
rect 27436 24735 27488 24744
rect 27436 24701 27445 24735
rect 27445 24701 27479 24735
rect 27479 24701 27488 24735
rect 27436 24692 27488 24701
rect 27988 24735 28040 24744
rect 27988 24701 27997 24735
rect 27997 24701 28031 24735
rect 28031 24701 28040 24735
rect 27988 24692 28040 24701
rect 35348 24828 35400 24880
rect 38844 24828 38896 24880
rect 44824 24828 44876 24880
rect 34704 24760 34756 24812
rect 35256 24803 35308 24812
rect 35256 24769 35265 24803
rect 35265 24769 35299 24803
rect 35299 24769 35308 24803
rect 35256 24760 35308 24769
rect 37740 24803 37792 24812
rect 37740 24769 37749 24803
rect 37749 24769 37783 24803
rect 37783 24769 37792 24803
rect 37740 24760 37792 24769
rect 38200 24760 38252 24812
rect 36360 24692 36412 24744
rect 39856 24692 39908 24744
rect 40868 24735 40920 24744
rect 40868 24701 40912 24735
rect 40912 24701 40920 24735
rect 40868 24692 40920 24701
rect 22744 24624 22796 24676
rect 24216 24624 24268 24676
rect 28172 24667 28224 24676
rect 20720 24556 20772 24608
rect 20996 24556 21048 24608
rect 28172 24633 28181 24667
rect 28181 24633 28215 24667
rect 28215 24633 28224 24667
rect 28172 24624 28224 24633
rect 28908 24624 28960 24676
rect 31760 24667 31812 24676
rect 28264 24556 28316 24608
rect 31760 24633 31769 24667
rect 31769 24633 31803 24667
rect 31803 24633 31812 24667
rect 31760 24624 31812 24633
rect 32404 24667 32456 24676
rect 29920 24556 29972 24608
rect 31668 24556 31720 24608
rect 32404 24633 32413 24667
rect 32413 24633 32447 24667
rect 32447 24633 32456 24667
rect 32404 24624 32456 24633
rect 32588 24624 32640 24676
rect 34520 24624 34572 24676
rect 35072 24667 35124 24676
rect 35072 24633 35081 24667
rect 35081 24633 35115 24667
rect 35115 24633 35124 24667
rect 35072 24624 35124 24633
rect 38016 24667 38068 24676
rect 38016 24633 38025 24667
rect 38025 24633 38059 24667
rect 38059 24633 38068 24667
rect 38016 24624 38068 24633
rect 44272 24692 44324 24744
rect 33600 24556 33652 24608
rect 36360 24556 36412 24608
rect 38660 24599 38712 24608
rect 38660 24565 38669 24599
rect 38669 24565 38703 24599
rect 38703 24565 38712 24599
rect 38660 24556 38712 24565
rect 41696 24556 41748 24608
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 10416 24395 10468 24404
rect 10416 24361 10425 24395
rect 10425 24361 10459 24395
rect 10459 24361 10468 24395
rect 10416 24352 10468 24361
rect 10784 24395 10836 24404
rect 10784 24361 10793 24395
rect 10793 24361 10827 24395
rect 10827 24361 10836 24395
rect 10784 24352 10836 24361
rect 12072 24395 12124 24404
rect 12072 24361 12081 24395
rect 12081 24361 12115 24395
rect 12115 24361 12124 24395
rect 12072 24352 12124 24361
rect 12624 24352 12676 24404
rect 13360 24352 13412 24404
rect 14372 24395 14424 24404
rect 11244 24284 11296 24336
rect 12440 24216 12492 24268
rect 13268 24216 13320 24268
rect 13452 24259 13504 24268
rect 13452 24225 13461 24259
rect 13461 24225 13495 24259
rect 13495 24225 13504 24259
rect 13452 24216 13504 24225
rect 14372 24361 14381 24395
rect 14381 24361 14415 24395
rect 14415 24361 14424 24395
rect 14372 24352 14424 24361
rect 15108 24352 15160 24404
rect 16856 24352 16908 24404
rect 20168 24395 20220 24404
rect 20168 24361 20177 24395
rect 20177 24361 20211 24395
rect 20211 24361 20220 24395
rect 20168 24352 20220 24361
rect 21180 24395 21232 24404
rect 21180 24361 21189 24395
rect 21189 24361 21223 24395
rect 21223 24361 21232 24395
rect 21180 24352 21232 24361
rect 23296 24395 23348 24404
rect 23296 24361 23305 24395
rect 23305 24361 23339 24395
rect 23339 24361 23348 24395
rect 23296 24352 23348 24361
rect 24216 24395 24268 24404
rect 24216 24361 24225 24395
rect 24225 24361 24259 24395
rect 24259 24361 24268 24395
rect 24216 24352 24268 24361
rect 24768 24395 24820 24404
rect 24768 24361 24777 24395
rect 24777 24361 24811 24395
rect 24811 24361 24820 24395
rect 24768 24352 24820 24361
rect 25136 24395 25188 24404
rect 25136 24361 25145 24395
rect 25145 24361 25179 24395
rect 25179 24361 25188 24395
rect 25136 24352 25188 24361
rect 27988 24352 28040 24404
rect 28172 24395 28224 24404
rect 28172 24361 28181 24395
rect 28181 24361 28215 24395
rect 28215 24361 28224 24395
rect 28172 24352 28224 24361
rect 28816 24395 28868 24404
rect 28816 24361 28825 24395
rect 28825 24361 28859 24395
rect 28859 24361 28868 24395
rect 28816 24352 28868 24361
rect 30104 24395 30156 24404
rect 30104 24361 30113 24395
rect 30113 24361 30147 24395
rect 30147 24361 30156 24395
rect 30104 24352 30156 24361
rect 31760 24395 31812 24404
rect 31760 24361 31769 24395
rect 31769 24361 31803 24395
rect 31803 24361 31812 24395
rect 31760 24352 31812 24361
rect 32588 24395 32640 24404
rect 32588 24361 32597 24395
rect 32597 24361 32631 24395
rect 32631 24361 32640 24395
rect 32588 24352 32640 24361
rect 35072 24395 35124 24404
rect 35072 24361 35081 24395
rect 35081 24361 35115 24395
rect 35115 24361 35124 24395
rect 35072 24352 35124 24361
rect 36452 24395 36504 24404
rect 36452 24361 36461 24395
rect 36461 24361 36495 24395
rect 36495 24361 36504 24395
rect 36452 24352 36504 24361
rect 37372 24352 37424 24404
rect 38936 24352 38988 24404
rect 16120 24327 16172 24336
rect 16120 24293 16129 24327
rect 16129 24293 16163 24327
rect 16163 24293 16172 24327
rect 16120 24284 16172 24293
rect 18512 24284 18564 24336
rect 20536 24284 20588 24336
rect 16028 24216 16080 24268
rect 17408 24216 17460 24268
rect 18144 24216 18196 24268
rect 19892 24216 19944 24268
rect 21272 24216 21324 24268
rect 22652 24284 22704 24336
rect 30472 24327 30524 24336
rect 22192 24216 22244 24268
rect 22284 24216 22336 24268
rect 22928 24216 22980 24268
rect 11152 24191 11204 24200
rect 11152 24157 11161 24191
rect 11161 24157 11195 24191
rect 11195 24157 11204 24191
rect 11152 24148 11204 24157
rect 15200 24148 15252 24200
rect 14372 24080 14424 24132
rect 18420 24080 18472 24132
rect 18788 24080 18840 24132
rect 12348 24012 12400 24064
rect 18880 24055 18932 24064
rect 18880 24021 18889 24055
rect 18889 24021 18923 24055
rect 18923 24021 18932 24055
rect 18880 24012 18932 24021
rect 19156 24055 19208 24064
rect 19156 24021 19165 24055
rect 19165 24021 19199 24055
rect 19199 24021 19208 24055
rect 19156 24012 19208 24021
rect 21640 24012 21692 24064
rect 25412 24216 25464 24268
rect 26424 24216 26476 24268
rect 28724 24259 28776 24268
rect 28724 24225 28733 24259
rect 28733 24225 28767 24259
rect 28767 24225 28776 24259
rect 28724 24216 28776 24225
rect 30472 24293 30481 24327
rect 30481 24293 30515 24327
rect 30515 24293 30524 24327
rect 30472 24284 30524 24293
rect 35348 24327 35400 24336
rect 35348 24293 35357 24327
rect 35357 24293 35391 24327
rect 35391 24293 35400 24327
rect 35348 24284 35400 24293
rect 35624 24284 35676 24336
rect 38108 24284 38160 24336
rect 41236 24284 41288 24336
rect 41604 24352 41656 24404
rect 41696 24327 41748 24336
rect 41696 24293 41705 24327
rect 41705 24293 41739 24327
rect 41739 24293 41748 24327
rect 41696 24284 41748 24293
rect 43260 24284 43312 24336
rect 29460 24216 29512 24268
rect 31760 24216 31812 24268
rect 33784 24259 33836 24268
rect 23848 24191 23900 24200
rect 23848 24157 23857 24191
rect 23857 24157 23891 24191
rect 23891 24157 23900 24191
rect 23848 24148 23900 24157
rect 27436 24191 27488 24200
rect 27436 24157 27445 24191
rect 27445 24157 27479 24191
rect 27479 24157 27488 24191
rect 27436 24148 27488 24157
rect 30380 24191 30432 24200
rect 30380 24157 30389 24191
rect 30389 24157 30423 24191
rect 30423 24157 30432 24191
rect 30380 24148 30432 24157
rect 31024 24191 31076 24200
rect 31024 24157 31033 24191
rect 31033 24157 31067 24191
rect 31067 24157 31076 24191
rect 31024 24148 31076 24157
rect 32680 24148 32732 24200
rect 33784 24225 33793 24259
rect 33793 24225 33827 24259
rect 33827 24225 33836 24259
rect 33784 24216 33836 24225
rect 34060 24259 34112 24268
rect 34060 24225 34069 24259
rect 34069 24225 34103 24259
rect 34103 24225 34112 24259
rect 34060 24216 34112 24225
rect 40500 24259 40552 24268
rect 40500 24225 40509 24259
rect 40509 24225 40543 24259
rect 40543 24225 40552 24259
rect 40500 24216 40552 24225
rect 42800 24216 42852 24268
rect 34336 24191 34388 24200
rect 34336 24157 34345 24191
rect 34345 24157 34379 24191
rect 34379 24157 34388 24191
rect 34336 24148 34388 24157
rect 36360 24148 36412 24200
rect 37924 24191 37976 24200
rect 37924 24157 37933 24191
rect 37933 24157 37967 24191
rect 37967 24157 37976 24191
rect 37924 24148 37976 24157
rect 43444 24191 43496 24200
rect 43444 24157 43453 24191
rect 43453 24157 43487 24191
rect 43487 24157 43496 24191
rect 43444 24148 43496 24157
rect 44088 24191 44140 24200
rect 44088 24157 44097 24191
rect 44097 24157 44131 24191
rect 44131 24157 44140 24191
rect 44088 24148 44140 24157
rect 24032 24012 24084 24064
rect 25688 24055 25740 24064
rect 25688 24021 25697 24055
rect 25697 24021 25731 24055
rect 25731 24021 25740 24055
rect 25688 24012 25740 24021
rect 27344 24012 27396 24064
rect 29736 24055 29788 24064
rect 29736 24021 29745 24055
rect 29745 24021 29779 24055
rect 29779 24021 29788 24055
rect 29736 24012 29788 24021
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 11152 23808 11204 23860
rect 12256 23851 12308 23860
rect 12256 23817 12265 23851
rect 12265 23817 12299 23851
rect 12299 23817 12308 23851
rect 12256 23808 12308 23817
rect 13268 23808 13320 23860
rect 17408 23851 17460 23860
rect 11244 23783 11296 23792
rect 11244 23749 11253 23783
rect 11253 23749 11287 23783
rect 11287 23749 11296 23783
rect 11244 23740 11296 23749
rect 15568 23740 15620 23792
rect 12348 23672 12400 23724
rect 12992 23715 13044 23724
rect 10416 23604 10468 23656
rect 12256 23604 12308 23656
rect 12992 23681 13001 23715
rect 13001 23681 13035 23715
rect 13035 23681 13044 23715
rect 12992 23672 13044 23681
rect 9956 23536 10008 23588
rect 14372 23672 14424 23724
rect 17408 23817 17417 23851
rect 17417 23817 17451 23851
rect 17451 23817 17460 23851
rect 17408 23808 17460 23817
rect 18144 23808 18196 23860
rect 18512 23808 18564 23860
rect 18880 23808 18932 23860
rect 19892 23851 19944 23860
rect 19892 23817 19901 23851
rect 19901 23817 19935 23851
rect 19935 23817 19944 23851
rect 19892 23808 19944 23817
rect 20536 23851 20588 23860
rect 20536 23817 20545 23851
rect 20545 23817 20579 23851
rect 20579 23817 20588 23851
rect 20536 23808 20588 23817
rect 21272 23808 21324 23860
rect 22192 23851 22244 23860
rect 22192 23817 22201 23851
rect 22201 23817 22235 23851
rect 22235 23817 22244 23851
rect 22192 23808 22244 23817
rect 22928 23851 22980 23860
rect 22928 23817 22937 23851
rect 22937 23817 22971 23851
rect 22971 23817 22980 23851
rect 22928 23808 22980 23817
rect 24216 23808 24268 23860
rect 26424 23851 26476 23860
rect 26424 23817 26433 23851
rect 26433 23817 26467 23851
rect 26467 23817 26476 23851
rect 26424 23808 26476 23817
rect 27620 23808 27672 23860
rect 27896 23808 27948 23860
rect 28724 23851 28776 23860
rect 28724 23817 28733 23851
rect 28733 23817 28767 23851
rect 28767 23817 28776 23851
rect 28724 23808 28776 23817
rect 29460 23851 29512 23860
rect 29460 23817 29469 23851
rect 29469 23817 29503 23851
rect 29503 23817 29512 23851
rect 29460 23808 29512 23817
rect 30472 23808 30524 23860
rect 33784 23808 33836 23860
rect 34244 23808 34296 23860
rect 36544 23851 36596 23860
rect 36544 23817 36553 23851
rect 36553 23817 36587 23851
rect 36587 23817 36596 23851
rect 36544 23808 36596 23817
rect 36636 23808 36688 23860
rect 19432 23783 19484 23792
rect 19432 23749 19441 23783
rect 19441 23749 19475 23783
rect 19475 23749 19484 23783
rect 19432 23740 19484 23749
rect 20076 23740 20128 23792
rect 21732 23740 21784 23792
rect 31024 23740 31076 23792
rect 35808 23783 35860 23792
rect 35808 23749 35817 23783
rect 35817 23749 35851 23783
rect 35851 23749 35860 23783
rect 35808 23740 35860 23749
rect 14464 23647 14516 23656
rect 14464 23613 14473 23647
rect 14473 23613 14507 23647
rect 14507 23613 14516 23647
rect 14464 23604 14516 23613
rect 18144 23672 18196 23724
rect 19156 23672 19208 23724
rect 21180 23672 21232 23724
rect 25688 23672 25740 23724
rect 29828 23715 29880 23724
rect 23940 23647 23992 23656
rect 23940 23613 23949 23647
rect 23949 23613 23983 23647
rect 23983 23613 23992 23647
rect 23940 23604 23992 23613
rect 24032 23604 24084 23656
rect 27620 23647 27672 23656
rect 27620 23613 27629 23647
rect 27629 23613 27663 23647
rect 27663 23613 27672 23647
rect 27620 23604 27672 23613
rect 29828 23681 29837 23715
rect 29837 23681 29871 23715
rect 29871 23681 29880 23715
rect 29828 23672 29880 23681
rect 30104 23672 30156 23724
rect 33232 23672 33284 23724
rect 27988 23604 28040 23656
rect 36360 23604 36412 23656
rect 38660 23808 38712 23860
rect 40500 23808 40552 23860
rect 41236 23851 41288 23860
rect 41236 23817 41245 23851
rect 41245 23817 41279 23851
rect 41279 23817 41288 23851
rect 41236 23808 41288 23817
rect 43444 23808 43496 23860
rect 43260 23740 43312 23792
rect 37740 23715 37792 23724
rect 37740 23681 37749 23715
rect 37749 23681 37783 23715
rect 37783 23681 37792 23715
rect 37740 23672 37792 23681
rect 39120 23672 39172 23724
rect 42156 23672 42208 23724
rect 37188 23604 37240 23656
rect 38200 23604 38252 23656
rect 40776 23647 40828 23656
rect 40776 23613 40820 23647
rect 40820 23613 40828 23647
rect 40776 23604 40828 23613
rect 14740 23536 14792 23588
rect 15108 23579 15160 23588
rect 15108 23545 15117 23579
rect 15117 23545 15151 23579
rect 15151 23545 15160 23579
rect 15108 23536 15160 23545
rect 15568 23536 15620 23588
rect 15844 23536 15896 23588
rect 16028 23579 16080 23588
rect 16028 23545 16037 23579
rect 16037 23545 16071 23579
rect 16071 23545 16080 23579
rect 16028 23536 16080 23545
rect 18880 23536 18932 23588
rect 16120 23468 16172 23520
rect 20720 23468 20772 23520
rect 28080 23579 28132 23588
rect 28080 23545 28089 23579
rect 28089 23545 28123 23579
rect 28123 23545 28132 23579
rect 28080 23536 28132 23545
rect 29000 23536 29052 23588
rect 21456 23468 21508 23520
rect 29736 23468 29788 23520
rect 31760 23468 31812 23520
rect 33324 23536 33376 23588
rect 34060 23536 34112 23588
rect 35348 23579 35400 23588
rect 35348 23545 35350 23579
rect 35350 23545 35384 23579
rect 35384 23545 35400 23579
rect 35348 23536 35400 23545
rect 38844 23579 38896 23588
rect 38844 23545 38853 23579
rect 38853 23545 38887 23579
rect 38887 23545 38896 23579
rect 38844 23536 38896 23545
rect 39028 23536 39080 23588
rect 32956 23468 33008 23520
rect 38108 23511 38160 23520
rect 38108 23477 38117 23511
rect 38117 23477 38151 23511
rect 38151 23477 38160 23511
rect 38108 23468 38160 23477
rect 41972 23579 42024 23588
rect 41972 23545 41981 23579
rect 41981 23545 42015 23579
rect 42015 23545 42024 23579
rect 41972 23536 42024 23545
rect 42800 23511 42852 23520
rect 42800 23477 42809 23511
rect 42809 23477 42843 23511
rect 42843 23477 42852 23511
rect 42800 23468 42852 23477
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 13452 23264 13504 23316
rect 15108 23307 15160 23316
rect 15108 23273 15117 23307
rect 15117 23273 15151 23307
rect 15151 23273 15160 23307
rect 15108 23264 15160 23273
rect 15568 23264 15620 23316
rect 15936 23264 15988 23316
rect 18788 23307 18840 23316
rect 18788 23273 18797 23307
rect 18797 23273 18831 23307
rect 18831 23273 18840 23307
rect 18788 23264 18840 23273
rect 19248 23264 19300 23316
rect 19984 23264 20036 23316
rect 20352 23264 20404 23316
rect 20812 23264 20864 23316
rect 17224 23196 17276 23248
rect 19064 23239 19116 23248
rect 19064 23205 19073 23239
rect 19073 23205 19107 23239
rect 19107 23205 19116 23239
rect 19064 23196 19116 23205
rect 20996 23196 21048 23248
rect 11888 23171 11940 23180
rect 11888 23137 11897 23171
rect 11897 23137 11931 23171
rect 11931 23137 11940 23171
rect 11888 23128 11940 23137
rect 12348 23171 12400 23180
rect 12348 23137 12357 23171
rect 12357 23137 12391 23171
rect 12391 23137 12400 23171
rect 12348 23128 12400 23137
rect 14280 23128 14332 23180
rect 12440 23103 12492 23112
rect 12440 23069 12449 23103
rect 12449 23069 12483 23103
rect 12483 23069 12492 23103
rect 12440 23060 12492 23069
rect 15384 23103 15436 23112
rect 15384 23069 15393 23103
rect 15393 23069 15427 23103
rect 15427 23069 15436 23103
rect 15384 23060 15436 23069
rect 15844 23060 15896 23112
rect 17040 23103 17092 23112
rect 17040 23069 17049 23103
rect 17049 23069 17083 23103
rect 17083 23069 17092 23103
rect 17040 23060 17092 23069
rect 18972 23103 19024 23112
rect 18972 23069 18981 23103
rect 18981 23069 19015 23103
rect 19015 23069 19024 23103
rect 18972 23060 19024 23069
rect 19616 23103 19668 23112
rect 19616 23069 19625 23103
rect 19625 23069 19659 23103
rect 19659 23069 19668 23103
rect 19616 23060 19668 23069
rect 23848 23264 23900 23316
rect 27896 23264 27948 23316
rect 30104 23264 30156 23316
rect 30472 23264 30524 23316
rect 32956 23264 33008 23316
rect 37096 23307 37148 23316
rect 37096 23273 37105 23307
rect 37105 23273 37139 23307
rect 37139 23273 37148 23307
rect 37096 23264 37148 23273
rect 37924 23264 37976 23316
rect 39212 23307 39264 23316
rect 39212 23273 39221 23307
rect 39221 23273 39255 23307
rect 39255 23273 39264 23307
rect 39212 23264 39264 23273
rect 41236 23307 41288 23316
rect 41236 23273 41245 23307
rect 41245 23273 41279 23307
rect 41279 23273 41288 23307
rect 41236 23264 41288 23273
rect 41972 23264 42024 23316
rect 42156 23264 42208 23316
rect 44088 23264 44140 23316
rect 28264 23196 28316 23248
rect 32588 23196 32640 23248
rect 34428 23196 34480 23248
rect 34704 23196 34756 23248
rect 22928 23171 22980 23180
rect 22928 23137 22937 23171
rect 22937 23137 22971 23171
rect 22971 23137 22980 23171
rect 22928 23128 22980 23137
rect 23388 23128 23440 23180
rect 24032 23128 24084 23180
rect 24492 23171 24544 23180
rect 24492 23137 24501 23171
rect 24501 23137 24535 23171
rect 24535 23137 24544 23171
rect 24492 23128 24544 23137
rect 25228 23171 25280 23180
rect 25228 23137 25237 23171
rect 25237 23137 25271 23171
rect 25271 23137 25280 23171
rect 25228 23128 25280 23137
rect 26332 23128 26384 23180
rect 26976 23128 27028 23180
rect 30380 23128 30432 23180
rect 36268 23171 36320 23180
rect 36268 23137 36277 23171
rect 36277 23137 36311 23171
rect 36311 23137 36320 23171
rect 36268 23128 36320 23137
rect 37924 23171 37976 23180
rect 37924 23137 37933 23171
rect 37933 23137 37967 23171
rect 37967 23137 37976 23171
rect 37924 23128 37976 23137
rect 38292 23171 38344 23180
rect 38292 23137 38301 23171
rect 38301 23137 38335 23171
rect 38335 23137 38344 23171
rect 38292 23128 38344 23137
rect 39304 23171 39356 23180
rect 39304 23137 39313 23171
rect 39313 23137 39347 23171
rect 39347 23137 39356 23171
rect 39304 23128 39356 23137
rect 39764 23171 39816 23180
rect 39764 23137 39773 23171
rect 39773 23137 39807 23171
rect 39807 23137 39816 23171
rect 39764 23128 39816 23137
rect 40224 23128 40276 23180
rect 42800 23128 42852 23180
rect 15660 22924 15712 22976
rect 19432 22992 19484 23044
rect 26424 23060 26476 23112
rect 27712 23103 27764 23112
rect 27712 23069 27721 23103
rect 27721 23069 27755 23103
rect 27755 23069 27764 23103
rect 27712 23060 27764 23069
rect 28816 23060 28868 23112
rect 32128 23103 32180 23112
rect 32128 23069 32137 23103
rect 32137 23069 32171 23103
rect 32171 23069 32180 23103
rect 32128 23060 32180 23069
rect 34520 23103 34572 23112
rect 34520 23069 34529 23103
rect 34529 23069 34563 23103
rect 34563 23069 34572 23103
rect 34520 23060 34572 23069
rect 41696 23060 41748 23112
rect 21548 23035 21600 23044
rect 21548 23001 21557 23035
rect 21557 23001 21591 23035
rect 21591 23001 21600 23035
rect 21548 22992 21600 23001
rect 25320 22992 25372 23044
rect 31024 22992 31076 23044
rect 17776 22924 17828 22976
rect 26700 22967 26752 22976
rect 26700 22933 26709 22967
rect 26709 22933 26743 22967
rect 26743 22933 26752 22967
rect 26700 22924 26752 22933
rect 28632 22967 28684 22976
rect 28632 22933 28641 22967
rect 28641 22933 28675 22967
rect 28675 22933 28684 22967
rect 28632 22924 28684 22933
rect 35348 22924 35400 22976
rect 35808 22924 35860 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 14280 22763 14332 22772
rect 14280 22729 14289 22763
rect 14289 22729 14323 22763
rect 14323 22729 14332 22763
rect 14280 22720 14332 22729
rect 17040 22720 17092 22772
rect 15476 22652 15528 22704
rect 15660 22695 15712 22704
rect 15660 22661 15669 22695
rect 15669 22661 15703 22695
rect 15703 22661 15712 22695
rect 15660 22652 15712 22661
rect 12440 22627 12492 22636
rect 12440 22593 12449 22627
rect 12449 22593 12483 22627
rect 12483 22593 12492 22627
rect 12440 22584 12492 22593
rect 15108 22627 15160 22636
rect 15108 22593 15117 22627
rect 15117 22593 15151 22627
rect 15151 22593 15160 22627
rect 15108 22584 15160 22593
rect 16120 22584 16172 22636
rect 17316 22720 17368 22772
rect 19432 22720 19484 22772
rect 20996 22763 21048 22772
rect 20996 22729 21005 22763
rect 21005 22729 21039 22763
rect 21039 22729 21048 22763
rect 20996 22720 21048 22729
rect 22928 22763 22980 22772
rect 22928 22729 22937 22763
rect 22937 22729 22971 22763
rect 22971 22729 22980 22763
rect 22928 22720 22980 22729
rect 23388 22763 23440 22772
rect 23388 22729 23397 22763
rect 23397 22729 23431 22763
rect 23431 22729 23440 22763
rect 23388 22720 23440 22729
rect 24492 22763 24544 22772
rect 24492 22729 24501 22763
rect 24501 22729 24535 22763
rect 24535 22729 24544 22763
rect 24492 22720 24544 22729
rect 28264 22720 28316 22772
rect 28816 22720 28868 22772
rect 31024 22720 31076 22772
rect 32680 22720 32732 22772
rect 36268 22763 36320 22772
rect 36268 22729 36277 22763
rect 36277 22729 36311 22763
rect 36311 22729 36320 22763
rect 36268 22720 36320 22729
rect 38292 22720 38344 22772
rect 39764 22763 39816 22772
rect 39764 22729 39773 22763
rect 39773 22729 39807 22763
rect 39807 22729 39816 22763
rect 39764 22720 39816 22729
rect 41236 22720 41288 22772
rect 41696 22763 41748 22772
rect 41696 22729 41705 22763
rect 41705 22729 41739 22763
rect 41739 22729 41748 22763
rect 41696 22720 41748 22729
rect 17776 22652 17828 22704
rect 19616 22652 19668 22704
rect 18788 22627 18840 22636
rect 18788 22593 18797 22627
rect 18797 22593 18831 22627
rect 18831 22593 18840 22627
rect 18788 22584 18840 22593
rect 19064 22627 19116 22636
rect 19064 22593 19073 22627
rect 19073 22593 19107 22627
rect 19107 22593 19116 22627
rect 19064 22584 19116 22593
rect 19984 22584 20036 22636
rect 21548 22627 21600 22636
rect 21548 22593 21557 22627
rect 21557 22593 21591 22627
rect 21591 22593 21600 22627
rect 21548 22584 21600 22593
rect 23940 22652 23992 22704
rect 23572 22559 23624 22568
rect 23572 22525 23581 22559
rect 23581 22525 23615 22559
rect 23615 22525 23624 22559
rect 23572 22516 23624 22525
rect 25228 22516 25280 22568
rect 26148 22559 26200 22568
rect 10508 22448 10560 22500
rect 11888 22448 11940 22500
rect 12808 22448 12860 22500
rect 11244 22380 11296 22432
rect 15476 22448 15528 22500
rect 17224 22448 17276 22500
rect 18880 22491 18932 22500
rect 18880 22457 18889 22491
rect 18889 22457 18923 22491
rect 18923 22457 18932 22491
rect 18880 22448 18932 22457
rect 15752 22380 15804 22432
rect 15936 22380 15988 22432
rect 21456 22448 21508 22500
rect 24676 22491 24728 22500
rect 24676 22457 24685 22491
rect 24685 22457 24719 22491
rect 24719 22457 24728 22491
rect 24676 22448 24728 22457
rect 26148 22525 26157 22559
rect 26157 22525 26191 22559
rect 26191 22525 26200 22559
rect 27620 22584 27672 22636
rect 27712 22584 27764 22636
rect 28724 22652 28776 22704
rect 30104 22652 30156 22704
rect 30012 22584 30064 22636
rect 30932 22584 30984 22636
rect 26148 22516 26200 22525
rect 27988 22516 28040 22568
rect 32772 22652 32824 22704
rect 33600 22652 33652 22704
rect 33968 22652 34020 22704
rect 32128 22584 32180 22636
rect 35256 22584 35308 22636
rect 38568 22652 38620 22704
rect 38752 22652 38804 22704
rect 39304 22695 39356 22704
rect 39304 22661 39313 22695
rect 39313 22661 39347 22695
rect 39347 22661 39356 22695
rect 39304 22652 39356 22661
rect 43444 22652 43496 22704
rect 31668 22516 31720 22568
rect 33324 22516 33376 22568
rect 33784 22559 33836 22568
rect 26332 22448 26384 22500
rect 28632 22448 28684 22500
rect 29828 22448 29880 22500
rect 30104 22448 30156 22500
rect 33784 22525 33828 22559
rect 33828 22525 33836 22559
rect 33784 22516 33836 22525
rect 34888 22448 34940 22500
rect 35348 22491 35400 22500
rect 35348 22457 35357 22491
rect 35357 22457 35391 22491
rect 35391 22457 35400 22491
rect 35348 22448 35400 22457
rect 23664 22380 23716 22432
rect 25780 22423 25832 22432
rect 25780 22389 25789 22423
rect 25789 22389 25823 22423
rect 25823 22389 25832 22423
rect 25780 22380 25832 22389
rect 26424 22423 26476 22432
rect 26424 22389 26433 22423
rect 26433 22389 26467 22423
rect 26467 22389 26476 22423
rect 26424 22380 26476 22389
rect 28264 22380 28316 22432
rect 29644 22423 29696 22432
rect 29644 22389 29653 22423
rect 29653 22389 29687 22423
rect 29687 22389 29696 22423
rect 29644 22380 29696 22389
rect 32588 22423 32640 22432
rect 32588 22389 32597 22423
rect 32597 22389 32631 22423
rect 32631 22389 32640 22423
rect 32588 22380 32640 22389
rect 34704 22380 34756 22432
rect 35716 22380 35768 22432
rect 36176 22380 36228 22432
rect 37096 22516 37148 22568
rect 39028 22516 39080 22568
rect 42524 22516 42576 22568
rect 43812 22559 43864 22568
rect 43812 22525 43821 22559
rect 43821 22525 43855 22559
rect 43855 22525 43864 22559
rect 43812 22516 43864 22525
rect 37648 22491 37700 22500
rect 37648 22457 37657 22491
rect 37657 22457 37691 22491
rect 37691 22457 37700 22491
rect 37648 22448 37700 22457
rect 38384 22448 38436 22500
rect 37924 22423 37976 22432
rect 37924 22389 37933 22423
rect 37933 22389 37967 22423
rect 37967 22389 37976 22423
rect 37924 22380 37976 22389
rect 38016 22380 38068 22432
rect 38752 22380 38804 22432
rect 43720 22380 43772 22432
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 12440 22219 12492 22228
rect 12440 22185 12449 22219
rect 12449 22185 12483 22219
rect 12483 22185 12492 22219
rect 12440 22176 12492 22185
rect 14832 22176 14884 22228
rect 15384 22176 15436 22228
rect 18972 22176 19024 22228
rect 20260 22176 20312 22228
rect 23572 22176 23624 22228
rect 29000 22219 29052 22228
rect 29000 22185 29009 22219
rect 29009 22185 29043 22219
rect 29043 22185 29052 22219
rect 29000 22176 29052 22185
rect 29828 22219 29880 22228
rect 29828 22185 29837 22219
rect 29837 22185 29871 22219
rect 29871 22185 29880 22219
rect 29828 22176 29880 22185
rect 30012 22176 30064 22228
rect 31668 22219 31720 22228
rect 31668 22185 31677 22219
rect 31677 22185 31711 22219
rect 31711 22185 31720 22219
rect 31668 22176 31720 22185
rect 34520 22219 34572 22228
rect 34520 22185 34529 22219
rect 34529 22185 34563 22219
rect 34563 22185 34572 22219
rect 34520 22176 34572 22185
rect 34888 22219 34940 22228
rect 34888 22185 34897 22219
rect 34897 22185 34931 22219
rect 34931 22185 34940 22219
rect 34888 22176 34940 22185
rect 12808 22108 12860 22160
rect 14464 22108 14516 22160
rect 15108 22151 15160 22160
rect 15108 22117 15117 22151
rect 15117 22117 15151 22151
rect 15151 22117 15160 22151
rect 15108 22108 15160 22117
rect 15752 22108 15804 22160
rect 15844 22108 15896 22160
rect 17224 22151 17276 22160
rect 17224 22117 17233 22151
rect 17233 22117 17267 22151
rect 17267 22117 17276 22151
rect 17224 22108 17276 22117
rect 17776 22151 17828 22160
rect 17776 22117 17785 22151
rect 17785 22117 17819 22151
rect 17819 22117 17828 22151
rect 17776 22108 17828 22117
rect 19156 22108 19208 22160
rect 21272 22151 21324 22160
rect 21272 22117 21281 22151
rect 21281 22117 21315 22151
rect 21315 22117 21324 22151
rect 21272 22108 21324 22117
rect 10048 22040 10100 22092
rect 11796 22040 11848 22092
rect 12992 22083 13044 22092
rect 11244 21904 11296 21956
rect 12992 22049 13001 22083
rect 13001 22049 13035 22083
rect 13035 22049 13044 22083
rect 12992 22040 13044 22049
rect 18604 22083 18656 22092
rect 18604 22049 18613 22083
rect 18613 22049 18647 22083
rect 18647 22049 18656 22083
rect 18604 22040 18656 22049
rect 19616 22083 19668 22092
rect 19616 22049 19625 22083
rect 19625 22049 19659 22083
rect 19659 22049 19668 22083
rect 19616 22040 19668 22049
rect 22744 22040 22796 22092
rect 26424 22108 26476 22160
rect 28264 22108 28316 22160
rect 33416 22151 33468 22160
rect 24492 22083 24544 22092
rect 24492 22049 24501 22083
rect 24501 22049 24535 22083
rect 24535 22049 24544 22083
rect 24492 22040 24544 22049
rect 24676 22083 24728 22092
rect 24676 22049 24685 22083
rect 24685 22049 24719 22083
rect 24719 22049 24728 22083
rect 24676 22040 24728 22049
rect 26976 22083 27028 22092
rect 26976 22049 26985 22083
rect 26985 22049 27019 22083
rect 27019 22049 27028 22083
rect 26976 22040 27028 22049
rect 30932 22040 30984 22092
rect 33416 22117 33425 22151
rect 33425 22117 33459 22151
rect 33459 22117 33468 22151
rect 33416 22108 33468 22117
rect 35808 22176 35860 22228
rect 38292 22219 38344 22228
rect 38292 22185 38301 22219
rect 38301 22185 38335 22219
rect 38335 22185 38344 22219
rect 38292 22176 38344 22185
rect 38660 22176 38712 22228
rect 35348 22108 35400 22160
rect 35900 22108 35952 22160
rect 40040 22151 40092 22160
rect 40040 22117 40049 22151
rect 40049 22117 40083 22151
rect 40083 22117 40092 22151
rect 40040 22108 40092 22117
rect 43628 22108 43680 22160
rect 32404 22040 32456 22092
rect 36636 22083 36688 22092
rect 36636 22049 36645 22083
rect 36645 22049 36679 22083
rect 36679 22049 36688 22083
rect 36636 22040 36688 22049
rect 37004 22040 37056 22092
rect 37648 22040 37700 22092
rect 41420 22083 41472 22092
rect 41420 22049 41429 22083
rect 41429 22049 41463 22083
rect 41463 22049 41472 22083
rect 41420 22040 41472 22049
rect 12900 21972 12952 22024
rect 14740 21972 14792 22024
rect 16580 21972 16632 22024
rect 17132 22015 17184 22024
rect 17132 21981 17141 22015
rect 17141 21981 17175 22015
rect 17175 21981 17184 22015
rect 17132 21972 17184 21981
rect 19064 21972 19116 22024
rect 21180 22015 21232 22024
rect 21180 21981 21189 22015
rect 21189 21981 21223 22015
rect 21223 21981 21232 22015
rect 21180 21972 21232 21981
rect 21548 22015 21600 22024
rect 21548 21981 21557 22015
rect 21557 21981 21591 22015
rect 21591 21981 21600 22015
rect 21548 21972 21600 21981
rect 24124 21972 24176 22024
rect 27068 21972 27120 22024
rect 27528 21972 27580 22024
rect 27712 21972 27764 22024
rect 28080 22015 28132 22024
rect 28080 21981 28089 22015
rect 28089 21981 28123 22015
rect 28123 21981 28132 22015
rect 28080 21972 28132 21981
rect 28816 21972 28868 22024
rect 31576 21972 31628 22024
rect 33324 22015 33376 22024
rect 33324 21981 33333 22015
rect 33333 21981 33367 22015
rect 33367 21981 33376 22015
rect 33324 21972 33376 21981
rect 33692 22015 33744 22024
rect 33692 21981 33701 22015
rect 33701 21981 33735 22015
rect 33735 21981 33744 22015
rect 33692 21972 33744 21981
rect 36912 21972 36964 22024
rect 39948 22015 40000 22024
rect 39948 21981 39957 22015
rect 39957 21981 39991 22015
rect 39991 21981 40000 22015
rect 39948 21972 40000 21981
rect 41512 21972 41564 22024
rect 12348 21904 12400 21956
rect 21456 21904 21508 21956
rect 23572 21904 23624 21956
rect 27620 21947 27672 21956
rect 15936 21836 15988 21888
rect 18972 21836 19024 21888
rect 19432 21836 19484 21888
rect 23112 21879 23164 21888
rect 23112 21845 23121 21879
rect 23121 21845 23155 21879
rect 23155 21845 23164 21879
rect 23112 21836 23164 21845
rect 27620 21913 27629 21947
rect 27629 21913 27663 21947
rect 27663 21913 27672 21947
rect 27620 21904 27672 21913
rect 29552 21904 29604 21956
rect 34244 21904 34296 21956
rect 34428 21904 34480 21956
rect 42156 22015 42208 22024
rect 42156 21981 42165 22015
rect 42165 21981 42199 22015
rect 42199 21981 42208 22015
rect 42156 21972 42208 21981
rect 43444 22015 43496 22024
rect 43444 21981 43453 22015
rect 43453 21981 43487 22015
rect 43487 21981 43496 22015
rect 43444 21972 43496 21981
rect 42248 21904 42300 21956
rect 43260 21904 43312 21956
rect 32772 21836 32824 21888
rect 33048 21879 33100 21888
rect 33048 21845 33057 21879
rect 33057 21845 33091 21879
rect 33091 21845 33100 21879
rect 33048 21836 33100 21845
rect 37004 21836 37056 21888
rect 37096 21879 37148 21888
rect 37096 21845 37105 21879
rect 37105 21845 37139 21879
rect 37139 21845 37148 21879
rect 37096 21836 37148 21845
rect 39028 21836 39080 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 11244 21675 11296 21684
rect 11244 21641 11253 21675
rect 11253 21641 11287 21675
rect 11287 21641 11296 21675
rect 11244 21632 11296 21641
rect 12716 21632 12768 21684
rect 12808 21675 12860 21684
rect 12808 21641 12817 21675
rect 12817 21641 12851 21675
rect 12851 21641 12860 21675
rect 12808 21632 12860 21641
rect 12992 21632 13044 21684
rect 16580 21675 16632 21684
rect 16580 21641 16589 21675
rect 16589 21641 16623 21675
rect 16623 21641 16632 21675
rect 16580 21632 16632 21641
rect 17132 21632 17184 21684
rect 17224 21632 17276 21684
rect 17592 21675 17644 21684
rect 17592 21641 17601 21675
rect 17601 21641 17635 21675
rect 17635 21641 17644 21675
rect 17592 21632 17644 21641
rect 18604 21675 18656 21684
rect 18604 21641 18613 21675
rect 18613 21641 18647 21675
rect 18647 21641 18656 21675
rect 18604 21632 18656 21641
rect 21272 21632 21324 21684
rect 22744 21675 22796 21684
rect 22744 21641 22753 21675
rect 22753 21641 22787 21675
rect 22787 21641 22796 21675
rect 22744 21632 22796 21641
rect 24492 21675 24544 21684
rect 24492 21641 24501 21675
rect 24501 21641 24535 21675
rect 24535 21641 24544 21675
rect 24492 21632 24544 21641
rect 24676 21632 24728 21684
rect 27160 21675 27212 21684
rect 27160 21641 27169 21675
rect 27169 21641 27203 21675
rect 27203 21641 27212 21675
rect 27160 21632 27212 21641
rect 28264 21632 28316 21684
rect 30932 21632 30984 21684
rect 31208 21632 31260 21684
rect 32496 21632 32548 21684
rect 33324 21632 33376 21684
rect 33416 21632 33468 21684
rect 34060 21632 34112 21684
rect 35900 21675 35952 21684
rect 35900 21641 35909 21675
rect 35909 21641 35943 21675
rect 35943 21641 35952 21675
rect 35900 21632 35952 21641
rect 37648 21632 37700 21684
rect 39948 21632 40000 21684
rect 41420 21675 41472 21684
rect 41420 21641 41429 21675
rect 41429 21641 41463 21675
rect 41463 21641 41472 21675
rect 41420 21632 41472 21641
rect 43444 21632 43496 21684
rect 17316 21607 17368 21616
rect 17316 21573 17325 21607
rect 17325 21573 17359 21607
rect 17359 21573 17368 21607
rect 17316 21564 17368 21573
rect 12900 21471 12952 21480
rect 12900 21437 12909 21471
rect 12909 21437 12943 21471
rect 12943 21437 12952 21471
rect 12900 21428 12952 21437
rect 19432 21496 19484 21548
rect 19984 21496 20036 21548
rect 18788 21471 18840 21480
rect 18788 21437 18797 21471
rect 18797 21437 18831 21471
rect 18831 21437 18840 21471
rect 18788 21428 18840 21437
rect 18972 21428 19024 21480
rect 20536 21428 20588 21480
rect 12808 21360 12860 21412
rect 11796 21292 11848 21344
rect 15752 21360 15804 21412
rect 16028 21360 16080 21412
rect 18236 21360 18288 21412
rect 19616 21360 19668 21412
rect 24124 21496 24176 21548
rect 21364 21428 21416 21480
rect 22376 21428 22428 21480
rect 26148 21564 26200 21616
rect 27528 21564 27580 21616
rect 27896 21607 27948 21616
rect 27896 21573 27905 21607
rect 27905 21573 27939 21607
rect 27939 21573 27948 21607
rect 27896 21564 27948 21573
rect 40500 21564 40552 21616
rect 41236 21564 41288 21616
rect 27712 21496 27764 21548
rect 30656 21496 30708 21548
rect 32404 21539 32456 21548
rect 32404 21505 32413 21539
rect 32413 21505 32447 21539
rect 32447 21505 32456 21539
rect 32404 21496 32456 21505
rect 32772 21496 32824 21548
rect 33692 21539 33744 21548
rect 33692 21505 33701 21539
rect 33701 21505 33735 21539
rect 33735 21505 33744 21539
rect 33692 21496 33744 21505
rect 34980 21539 35032 21548
rect 34980 21505 34989 21539
rect 34989 21505 35023 21539
rect 35023 21505 35032 21539
rect 34980 21496 35032 21505
rect 35256 21539 35308 21548
rect 35256 21505 35265 21539
rect 35265 21505 35299 21539
rect 35299 21505 35308 21539
rect 35256 21496 35308 21505
rect 37188 21496 37240 21548
rect 37280 21539 37332 21548
rect 37280 21505 37289 21539
rect 37289 21505 37323 21539
rect 37323 21505 37332 21539
rect 37280 21496 37332 21505
rect 40040 21496 40092 21548
rect 26148 21471 26200 21480
rect 26148 21437 26157 21471
rect 26157 21437 26191 21471
rect 26191 21437 26200 21471
rect 26148 21428 26200 21437
rect 27620 21471 27672 21480
rect 27620 21437 27629 21471
rect 27629 21437 27663 21471
rect 27663 21437 27672 21471
rect 27620 21428 27672 21437
rect 29552 21471 29604 21480
rect 29552 21437 29561 21471
rect 29561 21437 29595 21471
rect 29595 21437 29604 21471
rect 29552 21428 29604 21437
rect 29736 21471 29788 21480
rect 29736 21437 29745 21471
rect 29745 21437 29779 21471
rect 29779 21437 29788 21471
rect 29736 21428 29788 21437
rect 31208 21428 31260 21480
rect 31484 21428 31536 21480
rect 32864 21471 32916 21480
rect 32864 21437 32873 21471
rect 32873 21437 32907 21471
rect 32907 21437 32916 21471
rect 32864 21428 32916 21437
rect 40316 21428 40368 21480
rect 26240 21403 26292 21412
rect 18144 21292 18196 21344
rect 18512 21292 18564 21344
rect 18972 21335 19024 21344
rect 18972 21301 18981 21335
rect 18981 21301 19015 21335
rect 19015 21301 19024 21335
rect 18972 21292 19024 21301
rect 20720 21335 20772 21344
rect 20720 21301 20729 21335
rect 20729 21301 20763 21335
rect 20763 21301 20772 21335
rect 26240 21369 26249 21403
rect 26249 21369 26283 21403
rect 26283 21369 26292 21403
rect 26240 21360 26292 21369
rect 30012 21403 30064 21412
rect 30012 21369 30021 21403
rect 30021 21369 30055 21403
rect 30055 21369 30064 21403
rect 30012 21360 30064 21369
rect 20720 21292 20772 21301
rect 23572 21292 23624 21344
rect 26976 21292 27028 21344
rect 27528 21335 27580 21344
rect 27528 21301 27537 21335
rect 27537 21301 27571 21335
rect 27571 21301 27580 21335
rect 27528 21292 27580 21301
rect 29828 21292 29880 21344
rect 32128 21292 32180 21344
rect 32956 21292 33008 21344
rect 36912 21360 36964 21412
rect 38936 21403 38988 21412
rect 38936 21369 38945 21403
rect 38945 21369 38979 21403
rect 38979 21369 38988 21403
rect 38936 21360 38988 21369
rect 39028 21403 39080 21412
rect 39028 21369 39037 21403
rect 39037 21369 39071 21403
rect 39071 21369 39080 21403
rect 39580 21403 39632 21412
rect 39028 21360 39080 21369
rect 39580 21369 39589 21403
rect 39589 21369 39623 21403
rect 39623 21369 39632 21403
rect 39580 21360 39632 21369
rect 36452 21292 36504 21344
rect 36636 21335 36688 21344
rect 36636 21301 36645 21335
rect 36645 21301 36679 21335
rect 36679 21301 36688 21335
rect 36636 21292 36688 21301
rect 36820 21292 36872 21344
rect 38292 21292 38344 21344
rect 42156 21539 42208 21548
rect 42156 21505 42165 21539
rect 42165 21505 42199 21539
rect 42199 21505 42208 21539
rect 42156 21496 42208 21505
rect 43720 21496 43772 21548
rect 44180 21496 44232 21548
rect 42984 21292 43036 21344
rect 43628 21292 43680 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 12900 21088 12952 21140
rect 17132 21131 17184 21140
rect 17132 21097 17141 21131
rect 17141 21097 17175 21131
rect 17175 21097 17184 21131
rect 17132 21088 17184 21097
rect 21180 21088 21232 21140
rect 26148 21088 26200 21140
rect 27160 21088 27212 21140
rect 28816 21131 28868 21140
rect 11612 21020 11664 21072
rect 12164 21020 12216 21072
rect 10600 20995 10652 21004
rect 10600 20961 10609 20995
rect 10609 20961 10643 20995
rect 10643 20961 10652 20995
rect 10600 20952 10652 20961
rect 12532 20952 12584 21004
rect 12808 21020 12860 21072
rect 15844 21020 15896 21072
rect 17592 21063 17644 21072
rect 17592 21029 17601 21063
rect 17601 21029 17635 21063
rect 17635 21029 17644 21063
rect 17592 21020 17644 21029
rect 19156 21020 19208 21072
rect 20720 21020 20772 21072
rect 21088 21063 21140 21072
rect 21088 21029 21097 21063
rect 21097 21029 21131 21063
rect 21131 21029 21140 21063
rect 21088 21020 21140 21029
rect 24768 21063 24820 21072
rect 24768 21029 24777 21063
rect 24777 21029 24811 21063
rect 24811 21029 24820 21063
rect 24768 21020 24820 21029
rect 28816 21097 28825 21131
rect 28825 21097 28859 21131
rect 28859 21097 28868 21131
rect 28816 21088 28868 21097
rect 32404 21088 32456 21140
rect 32588 21088 32640 21140
rect 32772 21088 32824 21140
rect 34980 21131 35032 21140
rect 34980 21097 34989 21131
rect 34989 21097 35023 21131
rect 35023 21097 35032 21131
rect 34980 21088 35032 21097
rect 35808 21088 35860 21140
rect 38936 21131 38988 21140
rect 38936 21097 38945 21131
rect 38945 21097 38979 21131
rect 38979 21097 38988 21131
rect 38936 21088 38988 21097
rect 42248 21131 42300 21140
rect 42248 21097 42257 21131
rect 42257 21097 42291 21131
rect 42291 21097 42300 21131
rect 42248 21088 42300 21097
rect 43720 21088 43772 21140
rect 14004 20952 14056 21004
rect 18972 20952 19024 21004
rect 23572 20995 23624 21004
rect 23572 20961 23581 20995
rect 23581 20961 23615 20995
rect 23615 20961 23624 20995
rect 23572 20952 23624 20961
rect 26332 20952 26384 21004
rect 27620 20952 27672 21004
rect 29736 21020 29788 21072
rect 34060 21063 34112 21072
rect 34060 21029 34069 21063
rect 34069 21029 34103 21063
rect 34103 21029 34112 21063
rect 34060 21020 34112 21029
rect 34244 21020 34296 21072
rect 35256 21020 35308 21072
rect 36452 21063 36504 21072
rect 36452 21029 36461 21063
rect 36461 21029 36495 21063
rect 36495 21029 36504 21063
rect 36452 21020 36504 21029
rect 39028 21020 39080 21072
rect 40040 21020 40092 21072
rect 41604 21020 41656 21072
rect 43628 21020 43680 21072
rect 28264 20952 28316 21004
rect 29092 20952 29144 21004
rect 30104 20952 30156 21004
rect 30932 20995 30984 21004
rect 15200 20884 15252 20936
rect 16948 20884 17000 20936
rect 17500 20927 17552 20936
rect 17500 20893 17509 20927
rect 17509 20893 17543 20927
rect 17543 20893 17552 20927
rect 17500 20884 17552 20893
rect 12808 20816 12860 20868
rect 16212 20816 16264 20868
rect 21916 20884 21968 20936
rect 24400 20884 24452 20936
rect 21548 20859 21600 20868
rect 21548 20825 21557 20859
rect 21557 20825 21591 20859
rect 21591 20825 21600 20859
rect 21548 20816 21600 20825
rect 23296 20816 23348 20868
rect 26884 20884 26936 20936
rect 26976 20884 27028 20936
rect 28632 20884 28684 20936
rect 27436 20816 27488 20868
rect 30932 20961 30941 20995
rect 30941 20961 30975 20995
rect 30975 20961 30984 20995
rect 30932 20952 30984 20961
rect 33048 20995 33100 21004
rect 33048 20961 33057 20995
rect 33057 20961 33091 20995
rect 33091 20961 33100 20995
rect 33048 20952 33100 20961
rect 35716 20995 35768 21004
rect 35716 20961 35725 20995
rect 35725 20961 35759 20995
rect 35759 20961 35768 20995
rect 35716 20952 35768 20961
rect 36176 20995 36228 21004
rect 36176 20961 36185 20995
rect 36185 20961 36219 20995
rect 36219 20961 36228 20995
rect 36176 20952 36228 20961
rect 38844 20952 38896 21004
rect 32036 20884 32088 20936
rect 34612 20884 34664 20936
rect 37004 20884 37056 20936
rect 39672 20884 39724 20936
rect 40040 20927 40092 20936
rect 40040 20893 40049 20927
rect 40049 20893 40083 20927
rect 40083 20893 40092 20927
rect 40040 20884 40092 20893
rect 41144 20884 41196 20936
rect 41512 20884 41564 20936
rect 43260 20884 43312 20936
rect 43444 20927 43496 20936
rect 43444 20893 43453 20927
rect 43453 20893 43487 20927
rect 43487 20893 43496 20927
rect 43444 20884 43496 20893
rect 31116 20816 31168 20868
rect 41236 20816 41288 20868
rect 41972 20816 42024 20868
rect 10968 20791 11020 20800
rect 10968 20757 10977 20791
rect 10977 20757 11011 20791
rect 11011 20757 11020 20791
rect 10968 20748 11020 20757
rect 16396 20748 16448 20800
rect 18788 20748 18840 20800
rect 23388 20791 23440 20800
rect 23388 20757 23397 20791
rect 23397 20757 23431 20791
rect 23431 20757 23440 20791
rect 23388 20748 23440 20757
rect 23756 20748 23808 20800
rect 27712 20791 27764 20800
rect 27712 20757 27721 20791
rect 27721 20757 27755 20791
rect 27755 20757 27764 20791
rect 27712 20748 27764 20757
rect 28080 20791 28132 20800
rect 28080 20757 28089 20791
rect 28089 20757 28123 20791
rect 28123 20757 28132 20791
rect 28080 20748 28132 20757
rect 31484 20748 31536 20800
rect 33692 20791 33744 20800
rect 33692 20757 33701 20791
rect 33701 20757 33735 20791
rect 33735 20757 33744 20791
rect 33692 20748 33744 20757
rect 36912 20791 36964 20800
rect 36912 20757 36921 20791
rect 36921 20757 36955 20791
rect 36955 20757 36964 20791
rect 36912 20748 36964 20757
rect 37188 20791 37240 20800
rect 37188 20757 37197 20791
rect 37197 20757 37231 20791
rect 37231 20757 37240 20791
rect 37188 20748 37240 20757
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 10140 20587 10192 20596
rect 10140 20553 10149 20587
rect 10149 20553 10183 20587
rect 10183 20553 10192 20587
rect 10140 20544 10192 20553
rect 12532 20544 12584 20596
rect 14004 20587 14056 20596
rect 14004 20553 14013 20587
rect 14013 20553 14047 20587
rect 14047 20553 14056 20587
rect 14004 20544 14056 20553
rect 14832 20587 14884 20596
rect 14832 20553 14841 20587
rect 14841 20553 14875 20587
rect 14875 20553 14884 20587
rect 14832 20544 14884 20553
rect 16948 20587 17000 20596
rect 16948 20553 16957 20587
rect 16957 20553 16991 20587
rect 16991 20553 17000 20587
rect 16948 20544 17000 20553
rect 17592 20544 17644 20596
rect 16212 20519 16264 20528
rect 16212 20485 16221 20519
rect 16221 20485 16255 20519
rect 16255 20485 16264 20519
rect 16212 20476 16264 20485
rect 15844 20408 15896 20460
rect 12624 20340 12676 20392
rect 13176 20340 13228 20392
rect 10692 20315 10744 20324
rect 10692 20281 10701 20315
rect 10701 20281 10735 20315
rect 10735 20281 10744 20315
rect 10692 20272 10744 20281
rect 13728 20315 13780 20324
rect 13728 20281 13737 20315
rect 13737 20281 13771 20315
rect 13771 20281 13780 20315
rect 13728 20272 13780 20281
rect 15384 20247 15436 20256
rect 15384 20213 15393 20247
rect 15393 20213 15427 20247
rect 15427 20213 15436 20247
rect 15752 20315 15804 20324
rect 15752 20281 15761 20315
rect 15761 20281 15795 20315
rect 15795 20281 15804 20315
rect 15752 20272 15804 20281
rect 16304 20272 16356 20324
rect 18972 20544 19024 20596
rect 21088 20544 21140 20596
rect 21916 20587 21968 20596
rect 21916 20553 21925 20587
rect 21925 20553 21959 20587
rect 21959 20553 21968 20587
rect 21916 20544 21968 20553
rect 22376 20544 22428 20596
rect 23388 20587 23440 20596
rect 23388 20553 23397 20587
rect 23397 20553 23431 20587
rect 23431 20553 23440 20587
rect 23388 20544 23440 20553
rect 24768 20587 24820 20596
rect 24768 20553 24777 20587
rect 24777 20553 24811 20587
rect 24811 20553 24820 20587
rect 24768 20544 24820 20553
rect 25504 20544 25556 20596
rect 28264 20544 28316 20596
rect 28632 20587 28684 20596
rect 28632 20553 28641 20587
rect 28641 20553 28675 20587
rect 28675 20553 28684 20587
rect 28632 20544 28684 20553
rect 29092 20587 29144 20596
rect 29092 20553 29101 20587
rect 29101 20553 29135 20587
rect 29135 20553 29144 20587
rect 29092 20544 29144 20553
rect 30932 20544 30984 20596
rect 32036 20587 32088 20596
rect 32036 20553 32045 20587
rect 32045 20553 32079 20587
rect 32079 20553 32088 20587
rect 32036 20544 32088 20553
rect 32496 20587 32548 20596
rect 32496 20553 32505 20587
rect 32505 20553 32539 20587
rect 32539 20553 32548 20587
rect 32496 20544 32548 20553
rect 32680 20544 32732 20596
rect 34060 20544 34112 20596
rect 34612 20587 34664 20596
rect 34612 20553 34621 20587
rect 34621 20553 34655 20587
rect 34655 20553 34664 20587
rect 34612 20544 34664 20553
rect 35440 20587 35492 20596
rect 35440 20553 35449 20587
rect 35449 20553 35483 20587
rect 35483 20553 35492 20587
rect 35440 20544 35492 20553
rect 36176 20544 36228 20596
rect 38844 20544 38896 20596
rect 39028 20544 39080 20596
rect 39672 20587 39724 20596
rect 39672 20553 39681 20587
rect 39681 20553 39715 20587
rect 39715 20553 39724 20587
rect 39672 20544 39724 20553
rect 43444 20544 43496 20596
rect 44272 20587 44324 20596
rect 44272 20553 44281 20587
rect 44281 20553 44315 20587
rect 44315 20553 44324 20587
rect 44272 20544 44324 20553
rect 19156 20519 19208 20528
rect 19156 20485 19165 20519
rect 19165 20485 19199 20519
rect 19199 20485 19208 20519
rect 19156 20476 19208 20485
rect 23572 20476 23624 20528
rect 27436 20476 27488 20528
rect 28080 20476 28132 20528
rect 31116 20519 31168 20528
rect 31116 20485 31125 20519
rect 31125 20485 31159 20519
rect 31159 20485 31168 20519
rect 31116 20476 31168 20485
rect 32772 20476 32824 20528
rect 36636 20476 36688 20528
rect 15384 20204 15436 20213
rect 16028 20204 16080 20256
rect 19064 20272 19116 20324
rect 21364 20408 21416 20460
rect 23204 20408 23256 20460
rect 26516 20408 26568 20460
rect 19984 20204 20036 20256
rect 20352 20247 20404 20256
rect 20352 20213 20361 20247
rect 20361 20213 20395 20247
rect 20395 20213 20404 20247
rect 20628 20340 20680 20392
rect 21548 20340 21600 20392
rect 26700 20340 26752 20392
rect 23756 20315 23808 20324
rect 23756 20281 23765 20315
rect 23765 20281 23799 20315
rect 23799 20281 23808 20315
rect 23756 20272 23808 20281
rect 20352 20204 20404 20213
rect 23388 20204 23440 20256
rect 26148 20204 26200 20256
rect 27712 20272 27764 20324
rect 30012 20408 30064 20460
rect 33692 20408 33744 20460
rect 33784 20451 33836 20460
rect 33784 20417 33793 20451
rect 33793 20417 33827 20451
rect 33827 20417 33836 20451
rect 33784 20408 33836 20417
rect 34704 20408 34756 20460
rect 29828 20340 29880 20392
rect 30104 20272 30156 20324
rect 32680 20340 32732 20392
rect 35440 20340 35492 20392
rect 27436 20247 27488 20256
rect 27436 20213 27445 20247
rect 27445 20213 27479 20247
rect 27479 20213 27488 20247
rect 27436 20204 27488 20213
rect 29920 20204 29972 20256
rect 30656 20204 30708 20256
rect 31116 20272 31168 20324
rect 33324 20272 33376 20324
rect 36452 20408 36504 20460
rect 38108 20408 38160 20460
rect 40040 20408 40092 20460
rect 41972 20408 42024 20460
rect 42892 20383 42944 20392
rect 42892 20349 42910 20383
rect 42910 20349 42944 20383
rect 43904 20476 43956 20528
rect 42892 20340 42944 20349
rect 43812 20340 43864 20392
rect 44272 20340 44324 20392
rect 32404 20204 32456 20256
rect 33140 20204 33192 20256
rect 36820 20272 36872 20324
rect 36268 20204 36320 20256
rect 36912 20204 36964 20256
rect 39212 20272 39264 20324
rect 41328 20315 41380 20324
rect 41328 20281 41337 20315
rect 41337 20281 41371 20315
rect 41371 20281 41380 20315
rect 41328 20272 41380 20281
rect 41604 20272 41656 20324
rect 43444 20272 43496 20324
rect 41052 20247 41104 20256
rect 41052 20213 41061 20247
rect 41061 20213 41095 20247
rect 41095 20213 41104 20247
rect 41052 20204 41104 20213
rect 41144 20204 41196 20256
rect 43628 20247 43680 20256
rect 43628 20213 43637 20247
rect 43637 20213 43671 20247
rect 43671 20213 43680 20247
rect 43628 20204 43680 20213
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 10600 20043 10652 20052
rect 10600 20009 10609 20043
rect 10609 20009 10643 20043
rect 10643 20009 10652 20043
rect 10600 20000 10652 20009
rect 16304 20043 16356 20052
rect 16304 20009 16313 20043
rect 16313 20009 16347 20043
rect 16347 20009 16356 20043
rect 16304 20000 16356 20009
rect 16948 20000 17000 20052
rect 17500 20043 17552 20052
rect 10968 19932 11020 19984
rect 13268 19975 13320 19984
rect 13268 19941 13277 19975
rect 13277 19941 13311 19975
rect 13311 19941 13320 19975
rect 13268 19932 13320 19941
rect 15200 19932 15252 19984
rect 15844 19932 15896 19984
rect 16028 19975 16080 19984
rect 16028 19941 16037 19975
rect 16037 19941 16071 19975
rect 16071 19941 16080 19975
rect 16028 19932 16080 19941
rect 17500 20009 17509 20043
rect 17509 20009 17543 20043
rect 17543 20009 17552 20043
rect 17500 20000 17552 20009
rect 18420 20000 18472 20052
rect 20352 20000 20404 20052
rect 20536 20043 20588 20052
rect 20536 20009 20545 20043
rect 20545 20009 20579 20043
rect 20579 20009 20588 20043
rect 20536 20000 20588 20009
rect 19340 19932 19392 19984
rect 20168 19932 20220 19984
rect 20812 19932 20864 19984
rect 10140 19864 10192 19916
rect 16764 19864 16816 19916
rect 17960 19907 18012 19916
rect 17960 19873 17969 19907
rect 17969 19873 18003 19907
rect 18003 19873 18012 19907
rect 17960 19864 18012 19873
rect 19248 19907 19300 19916
rect 19248 19873 19257 19907
rect 19257 19873 19291 19907
rect 19291 19873 19300 19907
rect 19248 19864 19300 19873
rect 11244 19796 11296 19848
rect 13176 19839 13228 19848
rect 11520 19771 11572 19780
rect 11520 19737 11529 19771
rect 11529 19737 11563 19771
rect 11563 19737 11572 19771
rect 11520 19728 11572 19737
rect 13176 19805 13185 19839
rect 13185 19805 13219 19839
rect 13219 19805 13228 19839
rect 13176 19796 13228 19805
rect 13360 19728 13412 19780
rect 19064 19796 19116 19848
rect 20996 19796 21048 19848
rect 26148 20000 26200 20052
rect 26332 20043 26384 20052
rect 26332 20009 26341 20043
rect 26341 20009 26375 20043
rect 26375 20009 26384 20043
rect 26332 20000 26384 20009
rect 27620 20000 27672 20052
rect 30012 20043 30064 20052
rect 30012 20009 30021 20043
rect 30021 20009 30055 20043
rect 30055 20009 30064 20043
rect 30012 20000 30064 20009
rect 33692 20000 33744 20052
rect 40500 20043 40552 20052
rect 40500 20009 40509 20043
rect 40509 20009 40543 20043
rect 40543 20009 40552 20043
rect 40500 20000 40552 20009
rect 42984 20000 43036 20052
rect 23112 19932 23164 19984
rect 26240 19932 26292 19984
rect 30656 19975 30708 19984
rect 30656 19941 30665 19975
rect 30665 19941 30699 19975
rect 30699 19941 30708 19975
rect 30656 19932 30708 19941
rect 33140 19932 33192 19984
rect 27344 19864 27396 19916
rect 28632 19864 28684 19916
rect 29460 19907 29512 19916
rect 29460 19873 29469 19907
rect 29469 19873 29503 19907
rect 29503 19873 29512 19907
rect 29460 19864 29512 19873
rect 32772 19864 32824 19916
rect 32864 19864 32916 19916
rect 34060 19932 34112 19984
rect 35992 19932 36044 19984
rect 36268 19975 36320 19984
rect 36268 19941 36277 19975
rect 36277 19941 36311 19975
rect 36311 19941 36320 19975
rect 36268 19932 36320 19941
rect 37924 19932 37976 19984
rect 38660 19932 38712 19984
rect 40868 19932 40920 19984
rect 43444 19975 43496 19984
rect 41052 19907 41104 19916
rect 41052 19873 41061 19907
rect 41061 19873 41095 19907
rect 41095 19873 41104 19907
rect 41052 19864 41104 19873
rect 41604 19864 41656 19916
rect 43444 19941 43453 19975
rect 43453 19941 43487 19975
rect 43487 19941 43496 19975
rect 43444 19932 43496 19941
rect 43628 19932 43680 19984
rect 44088 19932 44140 19984
rect 42708 19864 42760 19916
rect 44916 19907 44968 19916
rect 44916 19873 44960 19907
rect 44960 19873 44968 19907
rect 44916 19864 44968 19873
rect 23296 19839 23348 19848
rect 23296 19805 23305 19839
rect 23305 19805 23339 19839
rect 23339 19805 23348 19839
rect 23296 19796 23348 19805
rect 19156 19728 19208 19780
rect 20352 19728 20404 19780
rect 23204 19728 23256 19780
rect 25044 19796 25096 19848
rect 25596 19839 25648 19848
rect 25596 19805 25605 19839
rect 25605 19805 25639 19839
rect 25639 19805 25648 19839
rect 25596 19796 25648 19805
rect 26700 19796 26752 19848
rect 26884 19839 26936 19848
rect 26884 19805 26893 19839
rect 26893 19805 26927 19839
rect 26927 19805 26936 19839
rect 26884 19796 26936 19805
rect 31392 19796 31444 19848
rect 32128 19796 32180 19848
rect 33692 19839 33744 19848
rect 33692 19805 33701 19839
rect 33701 19805 33735 19839
rect 33735 19805 33744 19839
rect 33692 19796 33744 19805
rect 33784 19796 33836 19848
rect 36820 19839 36872 19848
rect 36820 19805 36829 19839
rect 36829 19805 36863 19839
rect 36863 19805 36872 19839
rect 36820 19796 36872 19805
rect 38752 19796 38804 19848
rect 39212 19796 39264 19848
rect 40132 19839 40184 19848
rect 40132 19805 40141 19839
rect 40141 19805 40175 19839
rect 40175 19805 40184 19839
rect 40132 19796 40184 19805
rect 40776 19796 40828 19848
rect 42524 19796 42576 19848
rect 43720 19839 43772 19848
rect 43720 19805 43729 19839
rect 43729 19805 43763 19839
rect 43763 19805 43772 19839
rect 43720 19796 43772 19805
rect 23756 19728 23808 19780
rect 31208 19728 31260 19780
rect 33324 19728 33376 19780
rect 35716 19771 35768 19780
rect 35716 19737 35725 19771
rect 35725 19737 35759 19771
rect 35759 19737 35768 19771
rect 35716 19728 35768 19737
rect 41512 19728 41564 19780
rect 42248 19728 42300 19780
rect 43812 19728 43864 19780
rect 14096 19703 14148 19712
rect 14096 19669 14105 19703
rect 14105 19669 14139 19703
rect 14139 19669 14148 19703
rect 14096 19660 14148 19669
rect 16948 19660 17000 19712
rect 19340 19660 19392 19712
rect 19524 19703 19576 19712
rect 19524 19669 19533 19703
rect 19533 19669 19567 19703
rect 19567 19669 19576 19703
rect 19524 19660 19576 19669
rect 20168 19660 20220 19712
rect 21088 19660 21140 19712
rect 21180 19703 21232 19712
rect 21180 19669 21189 19703
rect 21189 19669 21223 19703
rect 21223 19669 21232 19703
rect 24216 19703 24268 19712
rect 21180 19660 21232 19669
rect 24216 19669 24225 19703
rect 24225 19669 24259 19703
rect 24259 19669 24268 19703
rect 24216 19660 24268 19669
rect 24400 19660 24452 19712
rect 26884 19660 26936 19712
rect 27436 19660 27488 19712
rect 27896 19660 27948 19712
rect 29460 19660 29512 19712
rect 37372 19660 37424 19712
rect 38108 19660 38160 19712
rect 41328 19703 41380 19712
rect 41328 19669 41337 19703
rect 41337 19669 41371 19703
rect 41371 19669 41380 19703
rect 41328 19660 41380 19669
rect 41788 19703 41840 19712
rect 41788 19669 41797 19703
rect 41797 19669 41831 19703
rect 41831 19669 41840 19703
rect 41788 19660 41840 19669
rect 43260 19660 43312 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 10140 19456 10192 19508
rect 10692 19499 10744 19508
rect 10692 19465 10701 19499
rect 10701 19465 10735 19499
rect 10735 19465 10744 19499
rect 10692 19456 10744 19465
rect 12164 19499 12216 19508
rect 12164 19465 12173 19499
rect 12173 19465 12207 19499
rect 12207 19465 12216 19499
rect 12164 19456 12216 19465
rect 12624 19499 12676 19508
rect 12624 19465 12633 19499
rect 12633 19465 12667 19499
rect 12667 19465 12676 19499
rect 12624 19456 12676 19465
rect 15200 19499 15252 19508
rect 15200 19465 15209 19499
rect 15209 19465 15243 19499
rect 15243 19465 15252 19499
rect 15200 19456 15252 19465
rect 15844 19499 15896 19508
rect 15844 19465 15853 19499
rect 15853 19465 15887 19499
rect 15887 19465 15896 19499
rect 15844 19456 15896 19465
rect 16764 19456 16816 19508
rect 17408 19499 17460 19508
rect 17408 19465 17417 19499
rect 17417 19465 17451 19499
rect 17451 19465 17460 19499
rect 17408 19456 17460 19465
rect 17500 19456 17552 19508
rect 18880 19456 18932 19508
rect 19984 19456 20036 19508
rect 21088 19456 21140 19508
rect 23112 19499 23164 19508
rect 23112 19465 23121 19499
rect 23121 19465 23155 19499
rect 23155 19465 23164 19499
rect 23112 19456 23164 19465
rect 26240 19456 26292 19508
rect 28264 19499 28316 19508
rect 28264 19465 28273 19499
rect 28273 19465 28307 19499
rect 28307 19465 28316 19499
rect 28264 19456 28316 19465
rect 28632 19499 28684 19508
rect 28632 19465 28641 19499
rect 28641 19465 28675 19499
rect 28675 19465 28684 19499
rect 28632 19456 28684 19465
rect 29460 19456 29512 19508
rect 31392 19499 31444 19508
rect 31392 19465 31401 19499
rect 31401 19465 31435 19499
rect 31435 19465 31444 19499
rect 31392 19456 31444 19465
rect 32772 19499 32824 19508
rect 32772 19465 32781 19499
rect 32781 19465 32815 19499
rect 32815 19465 32824 19499
rect 32772 19456 32824 19465
rect 33692 19456 33744 19508
rect 35992 19456 36044 19508
rect 36268 19456 36320 19508
rect 14280 19431 14332 19440
rect 14280 19397 14289 19431
rect 14289 19397 14323 19431
rect 14323 19397 14332 19431
rect 14280 19388 14332 19397
rect 19340 19388 19392 19440
rect 20812 19388 20864 19440
rect 30656 19388 30708 19440
rect 32864 19388 32916 19440
rect 33140 19431 33192 19440
rect 33140 19397 33149 19431
rect 33149 19397 33183 19431
rect 33183 19397 33192 19431
rect 33140 19388 33192 19397
rect 11060 19320 11112 19372
rect 11520 19363 11572 19372
rect 11520 19329 11529 19363
rect 11529 19329 11563 19363
rect 11563 19329 11572 19363
rect 11520 19320 11572 19329
rect 15384 19363 15436 19372
rect 15384 19329 15393 19363
rect 15393 19329 15427 19363
rect 15427 19329 15436 19363
rect 15384 19320 15436 19329
rect 19892 19320 19944 19372
rect 12164 19252 12216 19304
rect 16948 19295 17000 19304
rect 16948 19261 16957 19295
rect 16957 19261 16991 19295
rect 16991 19261 17000 19295
rect 16948 19252 17000 19261
rect 10692 19116 10744 19168
rect 13820 19227 13872 19236
rect 13820 19193 13829 19227
rect 13829 19193 13863 19227
rect 13863 19193 13872 19227
rect 13820 19184 13872 19193
rect 17040 19184 17092 19236
rect 19524 19252 19576 19304
rect 20076 19252 20128 19304
rect 24216 19320 24268 19372
rect 25596 19320 25648 19372
rect 33048 19320 33100 19372
rect 33600 19363 33652 19372
rect 33600 19329 33609 19363
rect 33609 19329 33643 19363
rect 33643 19329 33652 19363
rect 33600 19320 33652 19329
rect 34060 19388 34112 19440
rect 37556 19456 37608 19508
rect 38660 19456 38712 19508
rect 40500 19456 40552 19508
rect 41144 19456 41196 19508
rect 42708 19499 42760 19508
rect 42708 19465 42717 19499
rect 42717 19465 42751 19499
rect 42751 19465 42760 19499
rect 42708 19456 42760 19465
rect 43444 19456 43496 19508
rect 44088 19499 44140 19508
rect 44088 19465 44097 19499
rect 44097 19465 44131 19499
rect 44131 19465 44140 19499
rect 44088 19456 44140 19465
rect 44916 19499 44968 19508
rect 44916 19465 44925 19499
rect 44925 19465 44959 19499
rect 44959 19465 44968 19499
rect 44916 19456 44968 19465
rect 37280 19431 37332 19440
rect 37280 19397 37289 19431
rect 37289 19397 37323 19431
rect 37323 19397 37332 19431
rect 37280 19388 37332 19397
rect 38568 19388 38620 19440
rect 43720 19388 43772 19440
rect 36912 19320 36964 19372
rect 39488 19320 39540 19372
rect 21640 19252 21692 19304
rect 22008 19295 22060 19304
rect 22008 19261 22017 19295
rect 22017 19261 22051 19295
rect 22051 19261 22060 19295
rect 22008 19252 22060 19261
rect 27896 19295 27948 19304
rect 27896 19261 27905 19295
rect 27905 19261 27939 19295
rect 27939 19261 27948 19295
rect 27896 19252 27948 19261
rect 29828 19295 29880 19304
rect 29828 19261 29837 19295
rect 29837 19261 29871 19295
rect 29871 19261 29880 19295
rect 29828 19252 29880 19261
rect 31760 19252 31812 19304
rect 33140 19252 33192 19304
rect 38568 19252 38620 19304
rect 13084 19159 13136 19168
rect 13084 19125 13093 19159
rect 13093 19125 13127 19159
rect 13127 19125 13136 19159
rect 13084 19116 13136 19125
rect 13268 19116 13320 19168
rect 13636 19116 13688 19168
rect 17776 19159 17828 19168
rect 17776 19125 17785 19159
rect 17785 19125 17819 19159
rect 17819 19125 17828 19159
rect 17776 19116 17828 19125
rect 18788 19159 18840 19168
rect 18788 19125 18797 19159
rect 18797 19125 18831 19159
rect 18831 19125 18840 19159
rect 18788 19116 18840 19125
rect 19064 19116 19116 19168
rect 21180 19184 21232 19236
rect 22192 19159 22244 19168
rect 22192 19125 22201 19159
rect 22201 19125 22235 19159
rect 22235 19125 22244 19159
rect 22192 19116 22244 19125
rect 23388 19159 23440 19168
rect 23388 19125 23397 19159
rect 23397 19125 23431 19159
rect 23431 19125 23440 19159
rect 23388 19116 23440 19125
rect 23572 19184 23624 19236
rect 24400 19227 24452 19236
rect 24400 19193 24409 19227
rect 24409 19193 24443 19227
rect 24443 19193 24452 19227
rect 24400 19184 24452 19193
rect 25412 19227 25464 19236
rect 25412 19193 25421 19227
rect 25421 19193 25455 19227
rect 25455 19193 25464 19227
rect 25412 19184 25464 19193
rect 25504 19227 25556 19236
rect 25504 19193 25513 19227
rect 25513 19193 25547 19227
rect 25547 19193 25556 19227
rect 25504 19184 25556 19193
rect 26884 19116 26936 19168
rect 27436 19116 27488 19168
rect 29920 19116 29972 19168
rect 32864 19184 32916 19236
rect 33692 19184 33744 19236
rect 36728 19227 36780 19236
rect 36728 19193 36737 19227
rect 36737 19193 36771 19227
rect 36771 19193 36780 19227
rect 36728 19184 36780 19193
rect 30564 19116 30616 19168
rect 30840 19116 30892 19168
rect 34704 19116 34756 19168
rect 37096 19184 37148 19236
rect 38476 19184 38528 19236
rect 40132 19252 40184 19304
rect 41788 19363 41840 19372
rect 41788 19329 41797 19363
rect 41797 19329 41831 19363
rect 41831 19329 41840 19363
rect 41788 19320 41840 19329
rect 37924 19159 37976 19168
rect 37924 19125 37933 19159
rect 37933 19125 37967 19159
rect 37967 19125 37976 19159
rect 37924 19116 37976 19125
rect 41604 19159 41656 19168
rect 41604 19125 41613 19159
rect 41613 19125 41647 19159
rect 41647 19125 41656 19159
rect 41604 19116 41656 19125
rect 42524 19116 42576 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 10968 18955 11020 18964
rect 10968 18921 10977 18955
rect 10977 18921 11011 18955
rect 11011 18921 11020 18955
rect 10968 18912 11020 18921
rect 11244 18955 11296 18964
rect 11244 18921 11253 18955
rect 11253 18921 11287 18955
rect 11287 18921 11296 18955
rect 11244 18912 11296 18921
rect 13176 18955 13228 18964
rect 13176 18921 13185 18955
rect 13185 18921 13219 18955
rect 13219 18921 13228 18955
rect 13176 18912 13228 18921
rect 13084 18844 13136 18896
rect 13820 18912 13872 18964
rect 18972 18912 19024 18964
rect 19340 18912 19392 18964
rect 20720 18955 20772 18964
rect 20720 18921 20729 18955
rect 20729 18921 20763 18955
rect 20763 18921 20772 18955
rect 20720 18912 20772 18921
rect 20904 18912 20956 18964
rect 22008 18955 22060 18964
rect 22008 18921 22017 18955
rect 22017 18921 22051 18955
rect 22051 18921 22060 18955
rect 22008 18912 22060 18921
rect 23664 18955 23716 18964
rect 23664 18921 23673 18955
rect 23673 18921 23707 18955
rect 23707 18921 23716 18955
rect 23664 18912 23716 18921
rect 25412 18912 25464 18964
rect 32864 18955 32916 18964
rect 32864 18921 32873 18955
rect 32873 18921 32907 18955
rect 32907 18921 32916 18955
rect 32864 18912 32916 18921
rect 33784 18912 33836 18964
rect 13728 18887 13780 18896
rect 13728 18853 13737 18887
rect 13737 18853 13771 18887
rect 13771 18853 13780 18887
rect 13728 18844 13780 18853
rect 14280 18887 14332 18896
rect 14280 18853 14289 18887
rect 14289 18853 14323 18887
rect 14323 18853 14332 18887
rect 14280 18844 14332 18853
rect 18604 18844 18656 18896
rect 19248 18887 19300 18896
rect 19248 18853 19257 18887
rect 19257 18853 19291 18887
rect 19291 18853 19300 18887
rect 19248 18844 19300 18853
rect 23388 18844 23440 18896
rect 23572 18844 23624 18896
rect 29828 18844 29880 18896
rect 30840 18844 30892 18896
rect 31208 18887 31260 18896
rect 31208 18853 31217 18887
rect 31217 18853 31251 18887
rect 31251 18853 31260 18887
rect 31208 18844 31260 18853
rect 33692 18887 33744 18896
rect 33692 18853 33701 18887
rect 33701 18853 33735 18887
rect 33735 18853 33744 18887
rect 33692 18844 33744 18853
rect 34244 18887 34296 18896
rect 34244 18853 34253 18887
rect 34253 18853 34287 18887
rect 34287 18853 34296 18887
rect 34244 18844 34296 18853
rect 34612 18844 34664 18896
rect 35256 18887 35308 18896
rect 35256 18853 35265 18887
rect 35265 18853 35299 18887
rect 35299 18853 35308 18887
rect 38752 18912 38804 18964
rect 40132 18955 40184 18964
rect 40132 18921 40141 18955
rect 40141 18921 40175 18955
rect 40175 18921 40184 18955
rect 40132 18912 40184 18921
rect 41328 18912 41380 18964
rect 35256 18844 35308 18853
rect 37648 18844 37700 18896
rect 41512 18887 41564 18896
rect 41512 18853 41521 18887
rect 41521 18853 41555 18887
rect 41555 18853 41564 18887
rect 41512 18844 41564 18853
rect 41604 18887 41656 18896
rect 41604 18853 41613 18887
rect 41613 18853 41647 18887
rect 41647 18853 41656 18887
rect 41604 18844 41656 18853
rect 10876 18776 10928 18828
rect 11520 18776 11572 18828
rect 12072 18776 12124 18828
rect 12808 18776 12860 18828
rect 15844 18776 15896 18828
rect 17224 18819 17276 18828
rect 17224 18785 17233 18819
rect 17233 18785 17267 18819
rect 17267 18785 17276 18819
rect 17224 18776 17276 18785
rect 17408 18776 17460 18828
rect 21364 18776 21416 18828
rect 23020 18776 23072 18828
rect 24584 18819 24636 18828
rect 13636 18751 13688 18760
rect 13636 18717 13645 18751
rect 13645 18717 13679 18751
rect 13679 18717 13688 18751
rect 13636 18708 13688 18717
rect 16580 18751 16632 18760
rect 16580 18717 16589 18751
rect 16589 18717 16623 18751
rect 16623 18717 16632 18751
rect 16580 18708 16632 18717
rect 19524 18708 19576 18760
rect 19892 18708 19944 18760
rect 20720 18708 20772 18760
rect 22192 18708 22244 18760
rect 24584 18785 24593 18819
rect 24593 18785 24627 18819
rect 24627 18785 24636 18819
rect 24584 18776 24636 18785
rect 25504 18776 25556 18828
rect 27068 18819 27120 18828
rect 27068 18785 27077 18819
rect 27077 18785 27111 18819
rect 27111 18785 27120 18819
rect 27068 18776 27120 18785
rect 29184 18819 29236 18828
rect 29184 18785 29193 18819
rect 29193 18785 29227 18819
rect 29227 18785 29236 18819
rect 29184 18776 29236 18785
rect 29736 18776 29788 18828
rect 32128 18776 32180 18828
rect 36912 18776 36964 18828
rect 40224 18776 40276 18828
rect 43996 18776 44048 18828
rect 24860 18708 24912 18760
rect 28540 18708 28592 18760
rect 33600 18751 33652 18760
rect 33600 18717 33609 18751
rect 33609 18717 33643 18751
rect 33643 18717 33652 18751
rect 33600 18708 33652 18717
rect 34704 18708 34756 18760
rect 38844 18708 38896 18760
rect 40592 18708 40644 18760
rect 44180 18708 44232 18760
rect 8392 18640 8444 18692
rect 9404 18640 9456 18692
rect 11060 18640 11112 18692
rect 14280 18640 14332 18692
rect 16764 18640 16816 18692
rect 17960 18683 18012 18692
rect 17960 18649 17969 18683
rect 17969 18649 18003 18683
rect 18003 18649 18012 18683
rect 17960 18640 18012 18649
rect 8760 18572 8812 18624
rect 16488 18572 16540 18624
rect 18328 18615 18380 18624
rect 18328 18581 18337 18615
rect 18337 18581 18371 18615
rect 18371 18581 18380 18615
rect 18328 18572 18380 18581
rect 19524 18615 19576 18624
rect 19524 18581 19533 18615
rect 19533 18581 19567 18615
rect 19567 18581 19576 18615
rect 19524 18572 19576 18581
rect 25044 18615 25096 18624
rect 25044 18581 25053 18615
rect 25053 18581 25087 18615
rect 25087 18581 25096 18615
rect 25044 18572 25096 18581
rect 26700 18615 26752 18624
rect 26700 18581 26709 18615
rect 26709 18581 26743 18615
rect 26743 18581 26752 18615
rect 26700 18572 26752 18581
rect 31484 18572 31536 18624
rect 36084 18640 36136 18692
rect 38568 18640 38620 18692
rect 39212 18640 39264 18692
rect 36728 18572 36780 18624
rect 43076 18615 43128 18624
rect 43076 18581 43085 18615
rect 43085 18581 43119 18615
rect 43119 18581 43128 18615
rect 43076 18572 43128 18581
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 10876 18411 10928 18420
rect 10876 18377 10885 18411
rect 10885 18377 10919 18411
rect 10919 18377 10928 18411
rect 10876 18368 10928 18377
rect 12072 18411 12124 18420
rect 12072 18377 12081 18411
rect 12081 18377 12115 18411
rect 12115 18377 12124 18411
rect 12072 18368 12124 18377
rect 13636 18368 13688 18420
rect 13084 18300 13136 18352
rect 13728 18300 13780 18352
rect 13360 18275 13412 18284
rect 13360 18241 13369 18275
rect 13369 18241 13403 18275
rect 13403 18241 13412 18275
rect 13360 18232 13412 18241
rect 10048 18207 10100 18216
rect 10048 18173 10057 18207
rect 10057 18173 10091 18207
rect 10091 18173 10100 18207
rect 10048 18164 10100 18173
rect 10324 18207 10376 18216
rect 10324 18173 10333 18207
rect 10333 18173 10367 18207
rect 10367 18173 10376 18207
rect 10324 18164 10376 18173
rect 10508 18139 10560 18148
rect 10508 18105 10517 18139
rect 10517 18105 10551 18139
rect 10551 18105 10560 18139
rect 10508 18096 10560 18105
rect 9220 18071 9272 18080
rect 9220 18037 9229 18071
rect 9229 18037 9263 18071
rect 9263 18037 9272 18071
rect 9220 18028 9272 18037
rect 10876 18028 10928 18080
rect 12992 18139 13044 18148
rect 12992 18105 13001 18139
rect 13001 18105 13035 18139
rect 13035 18105 13044 18139
rect 12992 18096 13044 18105
rect 13084 18139 13136 18148
rect 13084 18105 13093 18139
rect 13093 18105 13127 18139
rect 13127 18105 13136 18139
rect 17224 18368 17276 18420
rect 18328 18368 18380 18420
rect 18604 18411 18656 18420
rect 18604 18377 18613 18411
rect 18613 18377 18647 18411
rect 18647 18377 18656 18411
rect 18604 18368 18656 18377
rect 18972 18411 19024 18420
rect 18972 18377 18981 18411
rect 18981 18377 19015 18411
rect 19015 18377 19024 18411
rect 18972 18368 19024 18377
rect 19892 18368 19944 18420
rect 21364 18411 21416 18420
rect 21364 18377 21373 18411
rect 21373 18377 21407 18411
rect 21407 18377 21416 18411
rect 21364 18368 21416 18377
rect 23020 18411 23072 18420
rect 23020 18377 23029 18411
rect 23029 18377 23063 18411
rect 23063 18377 23072 18411
rect 23020 18368 23072 18377
rect 23848 18368 23900 18420
rect 24584 18368 24636 18420
rect 27068 18411 27120 18420
rect 27068 18377 27077 18411
rect 27077 18377 27111 18411
rect 27111 18377 27120 18411
rect 27068 18368 27120 18377
rect 29184 18368 29236 18420
rect 29736 18411 29788 18420
rect 29736 18377 29745 18411
rect 29745 18377 29779 18411
rect 29779 18377 29788 18411
rect 29736 18368 29788 18377
rect 33600 18368 33652 18420
rect 33692 18368 33744 18420
rect 35256 18368 35308 18420
rect 36912 18368 36964 18420
rect 37648 18411 37700 18420
rect 37648 18377 37657 18411
rect 37657 18377 37691 18411
rect 37691 18377 37700 18411
rect 37648 18368 37700 18377
rect 39580 18368 39632 18420
rect 40592 18368 40644 18420
rect 41512 18368 41564 18420
rect 43996 18411 44048 18420
rect 17408 18300 17460 18352
rect 23664 18300 23716 18352
rect 16488 18275 16540 18284
rect 16488 18241 16497 18275
rect 16497 18241 16531 18275
rect 16531 18241 16540 18275
rect 16488 18232 16540 18241
rect 20444 18275 20496 18284
rect 20444 18241 20453 18275
rect 20453 18241 20487 18275
rect 20487 18241 20496 18275
rect 20444 18232 20496 18241
rect 24216 18275 24268 18284
rect 24216 18241 24225 18275
rect 24225 18241 24259 18275
rect 24259 18241 24268 18275
rect 24216 18232 24268 18241
rect 25412 18232 25464 18284
rect 25872 18232 25924 18284
rect 14464 18164 14516 18216
rect 15108 18207 15160 18216
rect 15108 18173 15117 18207
rect 15117 18173 15151 18207
rect 15151 18173 15160 18207
rect 15108 18164 15160 18173
rect 17960 18207 18012 18216
rect 17960 18173 17969 18207
rect 17969 18173 18003 18207
rect 18003 18173 18012 18207
rect 17960 18164 18012 18173
rect 18236 18164 18288 18216
rect 18788 18164 18840 18216
rect 19524 18164 19576 18216
rect 19984 18207 20036 18216
rect 19984 18173 19993 18207
rect 19993 18173 20027 18207
rect 20027 18173 20036 18207
rect 19984 18164 20036 18173
rect 20260 18164 20312 18216
rect 13084 18096 13136 18105
rect 16028 18096 16080 18148
rect 16580 18139 16632 18148
rect 16580 18105 16589 18139
rect 16589 18105 16623 18139
rect 16623 18105 16632 18139
rect 16580 18096 16632 18105
rect 17132 18139 17184 18148
rect 17132 18105 17141 18139
rect 17141 18105 17175 18139
rect 17175 18105 17184 18139
rect 17132 18096 17184 18105
rect 11888 18028 11940 18080
rect 13728 18028 13780 18080
rect 14924 18028 14976 18080
rect 15844 18028 15896 18080
rect 17868 18028 17920 18080
rect 21916 18071 21968 18080
rect 21916 18037 21925 18071
rect 21925 18037 21959 18071
rect 21959 18037 21968 18071
rect 21916 18028 21968 18037
rect 22008 18028 22060 18080
rect 22192 18139 22244 18148
rect 22192 18105 22201 18139
rect 22201 18105 22235 18139
rect 22235 18105 22244 18139
rect 22192 18096 22244 18105
rect 23848 18139 23900 18148
rect 23848 18105 23857 18139
rect 23857 18105 23891 18139
rect 23891 18105 23900 18139
rect 23848 18096 23900 18105
rect 24952 18096 25004 18148
rect 36820 18300 36872 18352
rect 40224 18343 40276 18352
rect 24216 18028 24268 18080
rect 26792 18096 26844 18148
rect 28724 18232 28776 18284
rect 33508 18232 33560 18284
rect 28816 18164 28868 18216
rect 30656 18207 30708 18216
rect 30656 18173 30665 18207
rect 30665 18173 30699 18207
rect 30699 18173 30708 18207
rect 30656 18164 30708 18173
rect 27712 18139 27764 18148
rect 27712 18105 27721 18139
rect 27721 18105 27755 18139
rect 27755 18105 27764 18139
rect 27712 18096 27764 18105
rect 27436 18071 27488 18080
rect 27436 18037 27445 18071
rect 27445 18037 27479 18071
rect 27479 18037 27488 18071
rect 32220 18139 32272 18148
rect 32220 18105 32229 18139
rect 32229 18105 32263 18139
rect 32263 18105 32272 18139
rect 32220 18096 32272 18105
rect 34704 18164 34756 18216
rect 37372 18232 37424 18284
rect 40224 18309 40233 18343
rect 40233 18309 40267 18343
rect 40267 18309 40276 18343
rect 40224 18300 40276 18309
rect 41604 18343 41656 18352
rect 41604 18309 41613 18343
rect 41613 18309 41647 18343
rect 41647 18309 41656 18343
rect 41604 18300 41656 18309
rect 41696 18300 41748 18352
rect 43996 18377 44005 18411
rect 44005 18377 44039 18411
rect 44039 18377 44048 18411
rect 43996 18368 44048 18377
rect 43076 18275 43128 18284
rect 43076 18241 43085 18275
rect 43085 18241 43119 18275
rect 43119 18241 43128 18275
rect 43076 18232 43128 18241
rect 44180 18232 44232 18284
rect 35348 18207 35400 18216
rect 35348 18173 35357 18207
rect 35357 18173 35391 18207
rect 35391 18173 35400 18207
rect 35348 18164 35400 18173
rect 33508 18096 33560 18148
rect 37096 18096 37148 18148
rect 37280 18139 37332 18148
rect 37280 18105 37289 18139
rect 37289 18105 37323 18139
rect 37323 18105 37332 18139
rect 37280 18096 37332 18105
rect 38200 18139 38252 18148
rect 38200 18105 38209 18139
rect 38209 18105 38243 18139
rect 38243 18105 38252 18139
rect 38200 18096 38252 18105
rect 27436 18028 27488 18037
rect 29000 18028 29052 18080
rect 30564 18071 30616 18080
rect 30564 18037 30573 18071
rect 30573 18037 30607 18071
rect 30607 18037 30616 18071
rect 30564 18028 30616 18037
rect 31116 18028 31168 18080
rect 33232 18028 33284 18080
rect 33968 18028 34020 18080
rect 34612 18071 34664 18080
rect 34612 18037 34621 18071
rect 34621 18037 34655 18071
rect 34655 18037 34664 18071
rect 34612 18028 34664 18037
rect 37924 18071 37976 18080
rect 37924 18037 37933 18071
rect 37933 18037 37967 18071
rect 37967 18037 37976 18071
rect 40684 18139 40736 18148
rect 40684 18105 40693 18139
rect 40693 18105 40727 18139
rect 40727 18105 40736 18139
rect 41236 18139 41288 18148
rect 40684 18096 40736 18105
rect 41236 18105 41245 18139
rect 41245 18105 41279 18139
rect 41279 18105 41288 18139
rect 41236 18096 41288 18105
rect 43536 18096 43588 18148
rect 37924 18028 37976 18037
rect 38568 18028 38620 18080
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 9864 17867 9916 17876
rect 9864 17833 9873 17867
rect 9873 17833 9907 17867
rect 9907 17833 9916 17867
rect 9864 17824 9916 17833
rect 9220 17756 9272 17808
rect 10324 17824 10376 17876
rect 10508 17824 10560 17876
rect 12992 17867 13044 17876
rect 12992 17833 13001 17867
rect 13001 17833 13035 17867
rect 13035 17833 13044 17867
rect 12992 17824 13044 17833
rect 16488 17867 16540 17876
rect 16488 17833 16497 17867
rect 16497 17833 16531 17867
rect 16531 17833 16540 17867
rect 16488 17824 16540 17833
rect 19248 17824 19300 17876
rect 19984 17867 20036 17876
rect 19984 17833 19993 17867
rect 19993 17833 20027 17867
rect 20027 17833 20036 17867
rect 19984 17824 20036 17833
rect 21272 17867 21324 17876
rect 21272 17833 21281 17867
rect 21281 17833 21315 17867
rect 21315 17833 21324 17867
rect 21272 17824 21324 17833
rect 11704 17799 11756 17808
rect 11704 17765 11713 17799
rect 11713 17765 11747 17799
rect 11747 17765 11756 17799
rect 11704 17756 11756 17765
rect 11888 17756 11940 17808
rect 13176 17799 13228 17808
rect 13176 17765 13185 17799
rect 13185 17765 13219 17799
rect 13219 17765 13228 17799
rect 13176 17756 13228 17765
rect 13452 17756 13504 17808
rect 15568 17756 15620 17808
rect 17040 17799 17092 17808
rect 17040 17765 17049 17799
rect 17049 17765 17083 17799
rect 17083 17765 17092 17799
rect 17040 17756 17092 17765
rect 23296 17799 23348 17808
rect 23296 17765 23305 17799
rect 23305 17765 23339 17799
rect 23339 17765 23348 17799
rect 27068 17824 27120 17876
rect 30840 17824 30892 17876
rect 33692 17824 33744 17876
rect 37188 17824 37240 17876
rect 37372 17867 37424 17876
rect 37372 17833 37381 17867
rect 37381 17833 37415 17867
rect 37415 17833 37424 17867
rect 37372 17824 37424 17833
rect 38108 17824 38160 17876
rect 38568 17824 38620 17876
rect 38844 17867 38896 17876
rect 38844 17833 38853 17867
rect 38853 17833 38887 17867
rect 38887 17833 38896 17867
rect 38844 17824 38896 17833
rect 23296 17756 23348 17765
rect 24400 17756 24452 17808
rect 24860 17799 24912 17808
rect 24860 17765 24869 17799
rect 24869 17765 24903 17799
rect 24903 17765 24912 17799
rect 24860 17756 24912 17765
rect 28540 17756 28592 17808
rect 28724 17799 28776 17808
rect 28724 17765 28733 17799
rect 28733 17765 28767 17799
rect 28767 17765 28776 17799
rect 28724 17756 28776 17765
rect 29736 17756 29788 17808
rect 30656 17756 30708 17808
rect 33508 17799 33560 17808
rect 33508 17765 33517 17799
rect 33517 17765 33551 17799
rect 33551 17765 33560 17799
rect 33508 17756 33560 17765
rect 33600 17799 33652 17808
rect 33600 17765 33609 17799
rect 33609 17765 33643 17799
rect 33643 17765 33652 17799
rect 33600 17756 33652 17765
rect 34336 17756 34388 17808
rect 36360 17756 36412 17808
rect 37096 17799 37148 17808
rect 10324 17731 10376 17740
rect 9680 17484 9732 17536
rect 10324 17697 10333 17731
rect 10333 17697 10367 17731
rect 10367 17697 10376 17731
rect 10324 17688 10376 17697
rect 17960 17688 18012 17740
rect 27344 17688 27396 17740
rect 30288 17731 30340 17740
rect 30288 17697 30297 17731
rect 30297 17697 30331 17731
rect 30331 17697 30340 17731
rect 30288 17688 30340 17697
rect 30472 17731 30524 17740
rect 30472 17697 30481 17731
rect 30481 17697 30515 17731
rect 30515 17697 30524 17731
rect 30472 17688 30524 17697
rect 36544 17731 36596 17740
rect 36544 17697 36553 17731
rect 36553 17697 36587 17731
rect 36587 17697 36596 17731
rect 36544 17688 36596 17697
rect 37096 17765 37105 17799
rect 37105 17765 37139 17799
rect 37139 17765 37148 17799
rect 37096 17756 37148 17765
rect 37648 17756 37700 17808
rect 39488 17756 39540 17808
rect 41512 17756 41564 17808
rect 43536 17799 43588 17808
rect 43536 17765 43545 17799
rect 43545 17765 43579 17799
rect 43579 17765 43588 17799
rect 43536 17756 43588 17765
rect 37832 17731 37884 17740
rect 37832 17697 37841 17731
rect 37841 17697 37875 17731
rect 37875 17697 37884 17731
rect 37832 17688 37884 17697
rect 38476 17688 38528 17740
rect 40684 17731 40736 17740
rect 40684 17697 40693 17731
rect 40693 17697 40727 17731
rect 40727 17697 40736 17731
rect 40684 17688 40736 17697
rect 45192 17688 45244 17740
rect 11336 17620 11388 17672
rect 12532 17552 12584 17604
rect 15108 17620 15160 17672
rect 16028 17663 16080 17672
rect 16028 17629 16037 17663
rect 16037 17629 16071 17663
rect 16071 17629 16080 17663
rect 16028 17620 16080 17629
rect 17408 17620 17460 17672
rect 17868 17620 17920 17672
rect 18604 17663 18656 17672
rect 18604 17629 18613 17663
rect 18613 17629 18647 17663
rect 18647 17629 18656 17663
rect 18604 17620 18656 17629
rect 20628 17620 20680 17672
rect 23204 17663 23256 17672
rect 23204 17629 23213 17663
rect 23213 17629 23247 17663
rect 23247 17629 23256 17663
rect 23204 17620 23256 17629
rect 24768 17663 24820 17672
rect 24768 17629 24777 17663
rect 24777 17629 24811 17663
rect 24811 17629 24820 17663
rect 24768 17620 24820 17629
rect 25044 17663 25096 17672
rect 25044 17629 25053 17663
rect 25053 17629 25087 17663
rect 25087 17629 25096 17663
rect 25044 17620 25096 17629
rect 29000 17620 29052 17672
rect 31208 17620 31260 17672
rect 33784 17663 33836 17672
rect 33784 17629 33793 17663
rect 33793 17629 33827 17663
rect 33827 17629 33836 17663
rect 33784 17620 33836 17629
rect 34704 17620 34756 17672
rect 35440 17620 35492 17672
rect 39856 17620 39908 17672
rect 41052 17620 41104 17672
rect 17132 17552 17184 17604
rect 14556 17484 14608 17536
rect 18144 17484 18196 17536
rect 20076 17552 20128 17604
rect 34244 17552 34296 17604
rect 40592 17552 40644 17604
rect 41972 17552 42024 17604
rect 20260 17527 20312 17536
rect 20260 17493 20269 17527
rect 20269 17493 20303 17527
rect 20303 17493 20312 17527
rect 20260 17484 20312 17493
rect 22008 17484 22060 17536
rect 25596 17484 25648 17536
rect 27712 17527 27764 17536
rect 27712 17493 27721 17527
rect 27721 17493 27755 17527
rect 27755 17493 27764 17527
rect 27712 17484 27764 17493
rect 29092 17484 29144 17536
rect 40316 17527 40368 17536
rect 40316 17493 40325 17527
rect 40325 17493 40359 17527
rect 40359 17493 40368 17527
rect 40316 17484 40368 17493
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 9680 17323 9732 17332
rect 9680 17289 9689 17323
rect 9689 17289 9723 17323
rect 9723 17289 9732 17323
rect 9680 17280 9732 17289
rect 13176 17280 13228 17332
rect 14924 17280 14976 17332
rect 17408 17323 17460 17332
rect 13452 17255 13504 17264
rect 13452 17221 13461 17255
rect 13461 17221 13495 17255
rect 13495 17221 13504 17255
rect 13452 17212 13504 17221
rect 10508 17144 10560 17196
rect 12532 17187 12584 17196
rect 12532 17153 12541 17187
rect 12541 17153 12575 17187
rect 12575 17153 12584 17187
rect 12532 17144 12584 17153
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 14280 17119 14332 17128
rect 14280 17085 14289 17119
rect 14289 17085 14323 17119
rect 14323 17085 14332 17119
rect 14280 17076 14332 17085
rect 17408 17289 17417 17323
rect 17417 17289 17451 17323
rect 17451 17289 17460 17323
rect 17408 17280 17460 17289
rect 19248 17323 19300 17332
rect 19248 17289 19257 17323
rect 19257 17289 19291 17323
rect 19291 17289 19300 17323
rect 19248 17280 19300 17289
rect 21456 17280 21508 17332
rect 23296 17280 23348 17332
rect 24860 17280 24912 17332
rect 25688 17280 25740 17332
rect 29000 17323 29052 17332
rect 29000 17289 29009 17323
rect 29009 17289 29043 17323
rect 29043 17289 29052 17323
rect 29000 17280 29052 17289
rect 29092 17280 29144 17332
rect 30472 17323 30524 17332
rect 30472 17289 30481 17323
rect 30481 17289 30515 17323
rect 30515 17289 30524 17323
rect 30472 17280 30524 17289
rect 33140 17280 33192 17332
rect 33876 17280 33928 17332
rect 34336 17323 34388 17332
rect 34336 17289 34345 17323
rect 34345 17289 34379 17323
rect 34379 17289 34388 17323
rect 34336 17280 34388 17289
rect 35992 17280 36044 17332
rect 39488 17323 39540 17332
rect 39488 17289 39497 17323
rect 39497 17289 39531 17323
rect 39531 17289 39540 17323
rect 39488 17280 39540 17289
rect 39856 17323 39908 17332
rect 39856 17289 39865 17323
rect 39865 17289 39899 17323
rect 39899 17289 39908 17323
rect 39856 17280 39908 17289
rect 40316 17323 40368 17332
rect 40316 17289 40325 17323
rect 40325 17289 40359 17323
rect 40359 17289 40368 17323
rect 40316 17280 40368 17289
rect 41512 17323 41564 17332
rect 41512 17289 41521 17323
rect 41521 17289 41555 17323
rect 41555 17289 41564 17323
rect 41512 17280 41564 17289
rect 15844 17212 15896 17264
rect 20812 17212 20864 17264
rect 31116 17212 31168 17264
rect 33600 17212 33652 17264
rect 36544 17255 36596 17264
rect 36544 17221 36553 17255
rect 36553 17221 36587 17255
rect 36587 17221 36596 17255
rect 36544 17212 36596 17221
rect 36820 17212 36872 17264
rect 37832 17255 37884 17264
rect 37832 17221 37841 17255
rect 37841 17221 37875 17255
rect 37875 17221 37884 17255
rect 37832 17212 37884 17221
rect 38384 17255 38436 17264
rect 38384 17221 38393 17255
rect 38393 17221 38427 17255
rect 38427 17221 38436 17255
rect 38384 17212 38436 17221
rect 41236 17212 41288 17264
rect 20444 17187 20496 17196
rect 20444 17153 20453 17187
rect 20453 17153 20487 17187
rect 20487 17153 20496 17187
rect 20444 17144 20496 17153
rect 18144 17076 18196 17128
rect 23112 17144 23164 17196
rect 25044 17144 25096 17196
rect 25872 17187 25924 17196
rect 25872 17153 25881 17187
rect 25881 17153 25915 17187
rect 25915 17153 25924 17187
rect 25872 17144 25924 17153
rect 27344 17144 27396 17196
rect 31208 17187 31260 17196
rect 31208 17153 31217 17187
rect 31217 17153 31251 17187
rect 31251 17153 31260 17187
rect 31208 17144 31260 17153
rect 31300 17144 31352 17196
rect 33048 17144 33100 17196
rect 33968 17144 34020 17196
rect 37096 17144 37148 17196
rect 10324 17008 10376 17060
rect 12624 17051 12676 17060
rect 12624 17017 12633 17051
rect 12633 17017 12667 17051
rect 12667 17017 12676 17051
rect 12624 17008 12676 17017
rect 15476 17008 15528 17060
rect 9220 16983 9272 16992
rect 9220 16949 9229 16983
rect 9229 16949 9263 16983
rect 9263 16949 9272 16983
rect 9220 16940 9272 16949
rect 11060 16983 11112 16992
rect 11060 16949 11069 16983
rect 11069 16949 11103 16983
rect 11103 16949 11112 16983
rect 11060 16940 11112 16949
rect 11704 16940 11756 16992
rect 11888 16940 11940 16992
rect 15568 16940 15620 16992
rect 19248 17008 19300 17060
rect 21272 17008 21324 17060
rect 23756 17051 23808 17060
rect 23756 17017 23765 17051
rect 23765 17017 23799 17051
rect 23799 17017 23808 17051
rect 23756 17008 23808 17017
rect 25596 17051 25648 17060
rect 17040 16983 17092 16992
rect 17040 16949 17049 16983
rect 17049 16949 17083 16983
rect 17083 16949 17092 16983
rect 17040 16940 17092 16949
rect 18328 16940 18380 16992
rect 23572 16940 23624 16992
rect 25596 17017 25605 17051
rect 25605 17017 25639 17051
rect 25639 17017 25648 17051
rect 25596 17008 25648 17017
rect 25688 17051 25740 17060
rect 25688 17017 25697 17051
rect 25697 17017 25731 17051
rect 25731 17017 25740 17051
rect 25688 17008 25740 17017
rect 26792 16940 26844 16992
rect 27160 16940 27212 16992
rect 27620 17076 27672 17128
rect 29184 17076 29236 17128
rect 33140 17076 33192 17128
rect 34428 17076 34480 17128
rect 35256 17076 35308 17128
rect 37556 17076 37608 17128
rect 41052 17144 41104 17196
rect 38568 17076 38620 17128
rect 42432 17119 42484 17128
rect 42432 17085 42441 17119
rect 42441 17085 42475 17119
rect 42475 17085 42484 17119
rect 42432 17076 42484 17085
rect 30288 17008 30340 17060
rect 27804 16983 27856 16992
rect 27804 16949 27813 16983
rect 27813 16949 27847 16983
rect 27847 16949 27856 16983
rect 27804 16940 27856 16949
rect 28632 16983 28684 16992
rect 28632 16949 28641 16983
rect 28641 16949 28675 16983
rect 28675 16949 28684 16983
rect 28632 16940 28684 16949
rect 31208 17008 31260 17060
rect 33324 17051 33376 17060
rect 33324 17017 33333 17051
rect 33333 17017 33367 17051
rect 33367 17017 33376 17051
rect 33324 17008 33376 17017
rect 33600 17008 33652 17060
rect 35808 17051 35860 17060
rect 35808 17017 35817 17051
rect 35817 17017 35851 17051
rect 35851 17017 35860 17051
rect 35808 17008 35860 17017
rect 37004 17008 37056 17060
rect 40592 17051 40644 17060
rect 40592 17017 40601 17051
rect 40601 17017 40635 17051
rect 40635 17017 40644 17051
rect 40592 17008 40644 17017
rect 43260 17280 43312 17332
rect 43536 17280 43588 17332
rect 44364 17280 44416 17332
rect 45192 17323 45244 17332
rect 45192 17289 45201 17323
rect 45201 17289 45235 17323
rect 45235 17289 45244 17323
rect 45192 17280 45244 17289
rect 43720 17144 43772 17196
rect 40316 16940 40368 16992
rect 43812 16940 43864 16992
rect 44364 17051 44416 17060
rect 44364 17017 44373 17051
rect 44373 17017 44407 17051
rect 44407 17017 44416 17051
rect 44364 17008 44416 17017
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 10324 16779 10376 16788
rect 10324 16745 10333 16779
rect 10333 16745 10367 16779
rect 10367 16745 10376 16779
rect 10324 16736 10376 16745
rect 10876 16779 10928 16788
rect 10876 16745 10885 16779
rect 10885 16745 10919 16779
rect 10919 16745 10928 16779
rect 10876 16736 10928 16745
rect 14280 16736 14332 16788
rect 15108 16779 15160 16788
rect 15108 16745 15117 16779
rect 15117 16745 15151 16779
rect 15151 16745 15160 16779
rect 15108 16736 15160 16745
rect 18604 16779 18656 16788
rect 18604 16745 18613 16779
rect 18613 16745 18647 16779
rect 18647 16745 18656 16779
rect 18604 16736 18656 16745
rect 20444 16779 20496 16788
rect 20444 16745 20453 16779
rect 20453 16745 20487 16779
rect 20487 16745 20496 16779
rect 20444 16736 20496 16745
rect 12716 16711 12768 16720
rect 12716 16677 12725 16711
rect 12725 16677 12759 16711
rect 12759 16677 12768 16711
rect 12716 16668 12768 16677
rect 15476 16711 15528 16720
rect 15476 16677 15485 16711
rect 15485 16677 15519 16711
rect 15519 16677 15528 16711
rect 15476 16668 15528 16677
rect 16028 16711 16080 16720
rect 16028 16677 16037 16711
rect 16037 16677 16071 16711
rect 16071 16677 16080 16711
rect 16028 16668 16080 16677
rect 16580 16668 16632 16720
rect 17408 16668 17460 16720
rect 22836 16668 22888 16720
rect 23204 16736 23256 16788
rect 23756 16779 23808 16788
rect 23756 16745 23765 16779
rect 23765 16745 23799 16779
rect 23799 16745 23808 16779
rect 23756 16736 23808 16745
rect 24768 16779 24820 16788
rect 24768 16745 24777 16779
rect 24777 16745 24811 16779
rect 24811 16745 24820 16779
rect 24768 16736 24820 16745
rect 28816 16779 28868 16788
rect 28816 16745 28825 16779
rect 28825 16745 28859 16779
rect 28859 16745 28868 16779
rect 28816 16736 28868 16745
rect 31208 16779 31260 16788
rect 31208 16745 31217 16779
rect 31217 16745 31251 16779
rect 31251 16745 31260 16779
rect 31208 16736 31260 16745
rect 33324 16779 33376 16788
rect 33324 16745 33333 16779
rect 33333 16745 33367 16779
rect 33367 16745 33376 16779
rect 33324 16736 33376 16745
rect 25044 16711 25096 16720
rect 25044 16677 25053 16711
rect 25053 16677 25087 16711
rect 25087 16677 25096 16711
rect 25044 16668 25096 16677
rect 28540 16668 28592 16720
rect 33416 16668 33468 16720
rect 34152 16736 34204 16788
rect 34520 16736 34572 16788
rect 35256 16736 35308 16788
rect 35440 16779 35492 16788
rect 35440 16745 35449 16779
rect 35449 16745 35483 16779
rect 35483 16745 35492 16779
rect 35440 16736 35492 16745
rect 37004 16736 37056 16788
rect 37372 16736 37424 16788
rect 38568 16779 38620 16788
rect 38568 16745 38577 16779
rect 38577 16745 38611 16779
rect 38611 16745 38620 16779
rect 38568 16736 38620 16745
rect 40592 16736 40644 16788
rect 42432 16779 42484 16788
rect 42432 16745 42441 16779
rect 42441 16745 42475 16779
rect 42475 16745 42484 16779
rect 42432 16736 42484 16745
rect 34244 16668 34296 16720
rect 35992 16668 36044 16720
rect 38292 16668 38344 16720
rect 41236 16711 41288 16720
rect 41236 16677 41245 16711
rect 41245 16677 41279 16711
rect 41279 16677 41288 16711
rect 41236 16668 41288 16677
rect 43536 16711 43588 16720
rect 43536 16677 43556 16711
rect 43556 16677 43588 16711
rect 43536 16668 43588 16677
rect 9312 16600 9364 16652
rect 9864 16600 9916 16652
rect 14464 16600 14516 16652
rect 12256 16532 12308 16584
rect 12992 16575 13044 16584
rect 12992 16541 13001 16575
rect 13001 16541 13035 16575
rect 13035 16541 13044 16575
rect 12992 16532 13044 16541
rect 14924 16532 14976 16584
rect 16948 16575 17000 16584
rect 10048 16464 10100 16516
rect 14648 16464 14700 16516
rect 16948 16541 16957 16575
rect 16957 16541 16991 16575
rect 16991 16541 17000 16575
rect 16948 16532 17000 16541
rect 17132 16532 17184 16584
rect 19064 16600 19116 16652
rect 21364 16600 21416 16652
rect 23388 16600 23440 16652
rect 26424 16600 26476 16652
rect 27804 16600 27856 16652
rect 29644 16643 29696 16652
rect 29644 16609 29653 16643
rect 29653 16609 29687 16643
rect 29687 16609 29696 16643
rect 29644 16600 29696 16609
rect 29736 16600 29788 16652
rect 30472 16600 30524 16652
rect 32956 16600 33008 16652
rect 37648 16600 37700 16652
rect 39396 16643 39448 16652
rect 39396 16609 39405 16643
rect 39405 16609 39439 16643
rect 39439 16609 39448 16643
rect 39396 16600 39448 16609
rect 39856 16643 39908 16652
rect 39856 16609 39865 16643
rect 39865 16609 39899 16643
rect 39899 16609 39908 16643
rect 39856 16600 39908 16609
rect 25596 16575 25648 16584
rect 11336 16396 11388 16448
rect 18604 16396 18656 16448
rect 19248 16464 19300 16516
rect 22284 16464 22336 16516
rect 20260 16396 20312 16448
rect 20628 16396 20680 16448
rect 22100 16439 22152 16448
rect 22100 16405 22109 16439
rect 22109 16405 22143 16439
rect 22143 16405 22152 16439
rect 25596 16541 25605 16575
rect 25605 16541 25639 16575
rect 25639 16541 25648 16575
rect 25596 16532 25648 16541
rect 30196 16575 30248 16584
rect 30196 16541 30205 16575
rect 30205 16541 30239 16575
rect 30239 16541 30248 16575
rect 30196 16532 30248 16541
rect 33876 16575 33928 16584
rect 33876 16541 33885 16575
rect 33885 16541 33919 16575
rect 33919 16541 33928 16575
rect 33876 16532 33928 16541
rect 35900 16575 35952 16584
rect 35900 16541 35909 16575
rect 35909 16541 35943 16575
rect 35943 16541 35952 16575
rect 35900 16532 35952 16541
rect 40500 16575 40552 16584
rect 40500 16541 40509 16575
rect 40509 16541 40543 16575
rect 40543 16541 40552 16575
rect 40500 16532 40552 16541
rect 41144 16575 41196 16584
rect 41144 16541 41153 16575
rect 41153 16541 41187 16575
rect 41187 16541 41196 16575
rect 41144 16532 41196 16541
rect 41328 16532 41380 16584
rect 43444 16575 43496 16584
rect 43444 16541 43453 16575
rect 43453 16541 43487 16575
rect 43487 16541 43496 16575
rect 43444 16532 43496 16541
rect 25412 16464 25464 16516
rect 34060 16464 34112 16516
rect 41052 16464 41104 16516
rect 22100 16396 22152 16405
rect 23296 16396 23348 16448
rect 23756 16396 23808 16448
rect 24308 16439 24360 16448
rect 24308 16405 24317 16439
rect 24317 16405 24351 16439
rect 24351 16405 24360 16439
rect 24308 16396 24360 16405
rect 27528 16439 27580 16448
rect 27528 16405 27537 16439
rect 27537 16405 27571 16439
rect 27571 16405 27580 16439
rect 27528 16396 27580 16405
rect 29184 16396 29236 16448
rect 37096 16439 37148 16448
rect 37096 16405 37105 16439
rect 37105 16405 37139 16439
rect 37139 16405 37148 16439
rect 37096 16396 37148 16405
rect 39028 16439 39080 16448
rect 39028 16405 39037 16439
rect 39037 16405 39071 16439
rect 39071 16405 39080 16439
rect 39028 16396 39080 16405
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 9312 16235 9364 16244
rect 9312 16201 9321 16235
rect 9321 16201 9355 16235
rect 9355 16201 9364 16235
rect 9312 16192 9364 16201
rect 11060 16192 11112 16244
rect 11336 16124 11388 16176
rect 11704 16192 11756 16244
rect 12256 16235 12308 16244
rect 12256 16201 12265 16235
rect 12265 16201 12299 16235
rect 12299 16201 12308 16235
rect 12256 16192 12308 16201
rect 12716 16235 12768 16244
rect 12716 16201 12725 16235
rect 12725 16201 12759 16235
rect 12759 16201 12768 16235
rect 12716 16192 12768 16201
rect 13360 16192 13412 16244
rect 14464 16192 14516 16244
rect 14924 16235 14976 16244
rect 14924 16201 14933 16235
rect 14933 16201 14967 16235
rect 14967 16201 14976 16235
rect 14924 16192 14976 16201
rect 13268 16056 13320 16108
rect 10876 15963 10928 15972
rect 10876 15929 10885 15963
rect 10885 15929 10919 15963
rect 10919 15929 10928 15963
rect 10876 15920 10928 15929
rect 10324 15895 10376 15904
rect 10324 15861 10333 15895
rect 10333 15861 10367 15895
rect 10367 15861 10376 15895
rect 10324 15852 10376 15861
rect 11888 15920 11940 15972
rect 13268 15963 13320 15972
rect 13268 15929 13277 15963
rect 13277 15929 13311 15963
rect 13311 15929 13320 15963
rect 13268 15920 13320 15929
rect 13360 15963 13412 15972
rect 13360 15929 13369 15963
rect 13369 15929 13403 15963
rect 13403 15929 13412 15963
rect 13360 15920 13412 15929
rect 14556 15920 14608 15972
rect 15476 16192 15528 16244
rect 17408 16235 17460 16244
rect 17408 16201 17417 16235
rect 17417 16201 17451 16235
rect 17451 16201 17460 16235
rect 17408 16192 17460 16201
rect 19984 16192 20036 16244
rect 24400 16192 24452 16244
rect 24860 16192 24912 16244
rect 25044 16192 25096 16244
rect 27436 16192 27488 16244
rect 29644 16235 29696 16244
rect 29644 16201 29653 16235
rect 29653 16201 29687 16235
rect 29687 16201 29696 16235
rect 29644 16192 29696 16201
rect 33416 16192 33468 16244
rect 34612 16192 34664 16244
rect 37096 16192 37148 16244
rect 37648 16192 37700 16244
rect 39488 16192 39540 16244
rect 18788 16124 18840 16176
rect 22928 16124 22980 16176
rect 32772 16124 32824 16176
rect 35992 16167 36044 16176
rect 16948 16056 17000 16108
rect 17132 16099 17184 16108
rect 17132 16065 17141 16099
rect 17141 16065 17175 16099
rect 17175 16065 17184 16099
rect 17132 16056 17184 16065
rect 20628 16099 20680 16108
rect 20628 16065 20637 16099
rect 20637 16065 20671 16099
rect 20671 16065 20680 16099
rect 20628 16056 20680 16065
rect 22100 16099 22152 16108
rect 22100 16065 22109 16099
rect 22109 16065 22143 16099
rect 22143 16065 22152 16099
rect 22100 16056 22152 16065
rect 23204 16056 23256 16108
rect 25596 16056 25648 16108
rect 30196 16056 30248 16108
rect 31300 16056 31352 16108
rect 31944 16099 31996 16108
rect 31944 16065 31953 16099
rect 31953 16065 31987 16099
rect 31987 16065 31996 16099
rect 31944 16056 31996 16065
rect 33876 16056 33928 16108
rect 34520 16056 34572 16108
rect 18052 16031 18104 16040
rect 18052 15997 18061 16031
rect 18061 15997 18095 16031
rect 18095 15997 18104 16031
rect 18052 15988 18104 15997
rect 18604 16031 18656 16040
rect 18604 15997 18613 16031
rect 18613 15997 18647 16031
rect 18647 15997 18656 16031
rect 18604 15988 18656 15997
rect 19064 15988 19116 16040
rect 19984 16031 20036 16040
rect 19984 15997 19993 16031
rect 19993 15997 20027 16031
rect 20027 15997 20036 16031
rect 19984 15988 20036 15997
rect 20260 15988 20312 16040
rect 16488 15963 16540 15972
rect 16488 15929 16497 15963
rect 16497 15929 16531 15963
rect 16531 15929 16540 15963
rect 16488 15920 16540 15929
rect 21916 15963 21968 15972
rect 21916 15929 21925 15963
rect 21925 15929 21959 15963
rect 21959 15929 21968 15963
rect 21916 15920 21968 15929
rect 22744 15920 22796 15972
rect 24308 15963 24360 15972
rect 24308 15929 24317 15963
rect 24317 15929 24351 15963
rect 24351 15929 24360 15963
rect 24308 15920 24360 15929
rect 24400 15963 24452 15972
rect 24400 15929 24409 15963
rect 24409 15929 24443 15963
rect 24443 15929 24452 15963
rect 24952 15963 25004 15972
rect 24400 15920 24452 15929
rect 24952 15929 24961 15963
rect 24961 15929 24995 15963
rect 24995 15929 25004 15963
rect 24952 15920 25004 15929
rect 25872 15963 25924 15972
rect 25872 15929 25881 15963
rect 25881 15929 25915 15963
rect 25915 15929 25924 15963
rect 25872 15920 25924 15929
rect 17040 15852 17092 15904
rect 18144 15895 18196 15904
rect 18144 15861 18153 15895
rect 18153 15861 18187 15895
rect 18187 15861 18196 15895
rect 18144 15852 18196 15861
rect 18972 15852 19024 15904
rect 19248 15852 19300 15904
rect 21364 15895 21416 15904
rect 21364 15861 21373 15895
rect 21373 15861 21407 15895
rect 21407 15861 21416 15895
rect 21364 15852 21416 15861
rect 22928 15852 22980 15904
rect 23388 15895 23440 15904
rect 23388 15861 23397 15895
rect 23397 15861 23431 15895
rect 23431 15861 23440 15895
rect 23388 15852 23440 15861
rect 26332 15920 26384 15972
rect 26424 15852 26476 15904
rect 27160 15852 27212 15904
rect 28080 16031 28132 16040
rect 28080 15997 28089 16031
rect 28089 15997 28123 16031
rect 28123 15997 28132 16031
rect 28080 15988 28132 15997
rect 34704 16031 34756 16040
rect 34704 15997 34713 16031
rect 34713 15997 34747 16031
rect 34747 15997 34756 16031
rect 34704 15988 34756 15997
rect 35992 16133 36001 16167
rect 36001 16133 36035 16167
rect 36035 16133 36044 16167
rect 35992 16124 36044 16133
rect 39856 16167 39908 16176
rect 39856 16133 39865 16167
rect 39865 16133 39899 16167
rect 39899 16133 39908 16167
rect 39856 16124 39908 16133
rect 35900 16056 35952 16108
rect 39028 16056 39080 16108
rect 35808 15988 35860 16040
rect 28264 15920 28316 15972
rect 28540 15852 28592 15904
rect 30564 15920 30616 15972
rect 31760 15920 31812 15972
rect 35716 15920 35768 15972
rect 38292 15963 38344 15972
rect 38292 15929 38301 15963
rect 38301 15929 38335 15963
rect 38335 15929 38344 15963
rect 38292 15920 38344 15929
rect 38844 15963 38896 15972
rect 38844 15929 38853 15963
rect 38853 15929 38887 15963
rect 38887 15929 38896 15963
rect 38844 15920 38896 15929
rect 41236 16192 41288 16244
rect 43536 16192 43588 16244
rect 41052 16124 41104 16176
rect 40500 16099 40552 16108
rect 40500 16065 40509 16099
rect 40509 16065 40543 16099
rect 40543 16065 40552 16099
rect 40500 16056 40552 16065
rect 43812 16099 43864 16108
rect 43812 16065 43821 16099
rect 43821 16065 43855 16099
rect 43855 16065 43864 16099
rect 43812 16056 43864 16065
rect 42708 16031 42760 16040
rect 42708 15997 42717 16031
rect 42717 15997 42751 16031
rect 42751 15997 42760 16031
rect 42708 15988 42760 15997
rect 41052 15920 41104 15972
rect 43444 15920 43496 15972
rect 32956 15895 33008 15904
rect 32956 15861 32965 15895
rect 32965 15861 32999 15895
rect 32999 15861 33008 15895
rect 32956 15852 33008 15861
rect 34244 15895 34296 15904
rect 34244 15861 34253 15895
rect 34253 15861 34287 15895
rect 34287 15861 34296 15895
rect 34244 15852 34296 15861
rect 37004 15895 37056 15904
rect 37004 15861 37013 15895
rect 37013 15861 37047 15895
rect 37047 15861 37056 15895
rect 37004 15852 37056 15861
rect 38384 15852 38436 15904
rect 39396 15895 39448 15904
rect 39396 15861 39405 15895
rect 39405 15861 39439 15895
rect 39439 15861 39448 15895
rect 39396 15852 39448 15861
rect 42432 15852 42484 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 13268 15648 13320 15700
rect 16948 15648 17000 15700
rect 18788 15691 18840 15700
rect 18788 15657 18797 15691
rect 18797 15657 18831 15691
rect 18831 15657 18840 15691
rect 18788 15648 18840 15657
rect 21272 15691 21324 15700
rect 21272 15657 21281 15691
rect 21281 15657 21315 15691
rect 21315 15657 21324 15691
rect 21272 15648 21324 15657
rect 21364 15648 21416 15700
rect 22284 15691 22336 15700
rect 22284 15657 22293 15691
rect 22293 15657 22327 15691
rect 22327 15657 22336 15691
rect 22284 15648 22336 15657
rect 25412 15691 25464 15700
rect 25412 15657 25421 15691
rect 25421 15657 25455 15691
rect 25455 15657 25464 15691
rect 25412 15648 25464 15657
rect 27804 15648 27856 15700
rect 28540 15648 28592 15700
rect 29184 15691 29236 15700
rect 29184 15657 29193 15691
rect 29193 15657 29227 15691
rect 29227 15657 29236 15691
rect 29184 15648 29236 15657
rect 29736 15691 29788 15700
rect 29736 15657 29745 15691
rect 29745 15657 29779 15691
rect 29779 15657 29788 15691
rect 29736 15648 29788 15657
rect 30196 15691 30248 15700
rect 30196 15657 30205 15691
rect 30205 15657 30239 15691
rect 30239 15657 30248 15691
rect 30196 15648 30248 15657
rect 31944 15691 31996 15700
rect 31944 15657 31953 15691
rect 31953 15657 31987 15691
rect 31987 15657 31996 15691
rect 31944 15648 31996 15657
rect 34244 15648 34296 15700
rect 35900 15648 35952 15700
rect 38292 15648 38344 15700
rect 41144 15648 41196 15700
rect 43444 15648 43496 15700
rect 11152 15623 11204 15632
rect 11152 15589 11161 15623
rect 11161 15589 11195 15623
rect 11195 15589 11204 15623
rect 11152 15580 11204 15589
rect 11704 15623 11756 15632
rect 11704 15589 11713 15623
rect 11713 15589 11747 15623
rect 11747 15589 11756 15623
rect 11704 15580 11756 15589
rect 12624 15580 12676 15632
rect 15568 15580 15620 15632
rect 18328 15580 18380 15632
rect 24676 15580 24728 15632
rect 26792 15580 26844 15632
rect 9956 15555 10008 15564
rect 9956 15521 9965 15555
rect 9965 15521 9999 15555
rect 9999 15521 10008 15555
rect 9956 15512 10008 15521
rect 17224 15512 17276 15564
rect 19800 15512 19852 15564
rect 22560 15512 22612 15564
rect 26424 15512 26476 15564
rect 31760 15580 31812 15632
rect 32772 15580 32824 15632
rect 33968 15623 34020 15632
rect 33968 15589 33977 15623
rect 33977 15589 34011 15623
rect 34011 15589 34020 15623
rect 33968 15580 34020 15589
rect 34336 15623 34388 15632
rect 34336 15589 34345 15623
rect 34345 15589 34379 15623
rect 34379 15589 34388 15623
rect 34336 15580 34388 15589
rect 35808 15580 35860 15632
rect 37004 15580 37056 15632
rect 37924 15580 37976 15632
rect 39120 15580 39172 15632
rect 11520 15444 11572 15496
rect 12164 15444 12216 15496
rect 16028 15444 16080 15496
rect 17500 15444 17552 15496
rect 20904 15487 20956 15496
rect 20904 15453 20913 15487
rect 20913 15453 20947 15487
rect 20947 15453 20956 15487
rect 20904 15444 20956 15453
rect 24216 15444 24268 15496
rect 26608 15487 26660 15496
rect 26608 15453 26617 15487
rect 26617 15453 26651 15487
rect 26651 15453 26660 15487
rect 26608 15444 26660 15453
rect 26884 15444 26936 15496
rect 28080 15444 28132 15496
rect 28264 15487 28316 15496
rect 28264 15453 28273 15487
rect 28273 15453 28307 15487
rect 28307 15453 28316 15487
rect 28264 15444 28316 15453
rect 13176 15419 13228 15428
rect 13176 15385 13185 15419
rect 13185 15385 13219 15419
rect 13219 15385 13228 15419
rect 13176 15376 13228 15385
rect 15936 15419 15988 15428
rect 15936 15385 15945 15419
rect 15945 15385 15979 15419
rect 15979 15385 15988 15419
rect 15936 15376 15988 15385
rect 16488 15419 16540 15428
rect 16488 15385 16497 15419
rect 16497 15385 16531 15419
rect 16531 15385 16540 15419
rect 16488 15376 16540 15385
rect 24952 15376 25004 15428
rect 26700 15376 26752 15428
rect 30288 15376 30340 15428
rect 31116 15512 31168 15564
rect 33876 15444 33928 15496
rect 36084 15512 36136 15564
rect 40500 15555 40552 15564
rect 34520 15487 34572 15496
rect 34520 15453 34529 15487
rect 34529 15453 34563 15487
rect 34563 15453 34572 15487
rect 34520 15444 34572 15453
rect 35256 15444 35308 15496
rect 40500 15521 40509 15555
rect 40509 15521 40543 15555
rect 40543 15521 40552 15555
rect 40500 15512 40552 15521
rect 36268 15444 36320 15496
rect 38476 15444 38528 15496
rect 38844 15487 38896 15496
rect 38844 15453 38853 15487
rect 38853 15453 38887 15487
rect 38887 15453 38896 15487
rect 38844 15444 38896 15453
rect 39856 15444 39908 15496
rect 42708 15512 42760 15564
rect 43352 15512 43404 15564
rect 41144 15487 41196 15496
rect 41144 15453 41153 15487
rect 41153 15453 41187 15487
rect 41187 15453 41196 15487
rect 41144 15444 41196 15453
rect 35348 15376 35400 15428
rect 37556 15376 37608 15428
rect 10876 15351 10928 15360
rect 10876 15317 10885 15351
rect 10885 15317 10919 15351
rect 10919 15317 10928 15351
rect 10876 15308 10928 15317
rect 15660 15308 15712 15360
rect 19064 15351 19116 15360
rect 19064 15317 19073 15351
rect 19073 15317 19107 15351
rect 19107 15317 19116 15351
rect 19064 15308 19116 15317
rect 22652 15308 22704 15360
rect 25872 15351 25924 15360
rect 25872 15317 25881 15351
rect 25881 15317 25915 15351
rect 25915 15317 25924 15351
rect 25872 15308 25924 15317
rect 27344 15308 27396 15360
rect 37188 15351 37240 15360
rect 37188 15317 37197 15351
rect 37197 15317 37231 15351
rect 37231 15317 37240 15351
rect 37188 15308 37240 15317
rect 41880 15351 41932 15360
rect 41880 15317 41889 15351
rect 41889 15317 41923 15351
rect 41923 15317 41932 15351
rect 41880 15308 41932 15317
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 9956 15104 10008 15156
rect 11520 15147 11572 15156
rect 11520 15113 11529 15147
rect 11529 15113 11563 15147
rect 11563 15113 11572 15147
rect 11520 15104 11572 15113
rect 12624 15147 12676 15156
rect 12624 15113 12633 15147
rect 12633 15113 12667 15147
rect 12667 15113 12676 15147
rect 12624 15104 12676 15113
rect 14556 15147 14608 15156
rect 14556 15113 14565 15147
rect 14565 15113 14599 15147
rect 14599 15113 14608 15147
rect 14556 15104 14608 15113
rect 15568 15104 15620 15156
rect 16028 15147 16080 15156
rect 16028 15113 16037 15147
rect 16037 15113 16071 15147
rect 16071 15113 16080 15147
rect 16028 15104 16080 15113
rect 18328 15147 18380 15156
rect 18328 15113 18337 15147
rect 18337 15113 18371 15147
rect 18371 15113 18380 15147
rect 18328 15104 18380 15113
rect 19800 15104 19852 15156
rect 23388 15104 23440 15156
rect 24676 15147 24728 15156
rect 24676 15113 24685 15147
rect 24685 15113 24719 15147
rect 24719 15113 24728 15147
rect 24676 15104 24728 15113
rect 14096 14968 14148 15020
rect 15936 14968 15988 15020
rect 18696 14968 18748 15020
rect 20904 14968 20956 15020
rect 24216 15011 24268 15020
rect 24216 14977 24225 15011
rect 24225 14977 24259 15011
rect 24259 14977 24268 15011
rect 24216 14968 24268 14977
rect 26608 15104 26660 15156
rect 27252 15104 27304 15156
rect 27344 15104 27396 15156
rect 28264 15104 28316 15156
rect 29736 15104 29788 15156
rect 30288 15147 30340 15156
rect 30288 15113 30297 15147
rect 30297 15113 30331 15147
rect 30331 15113 30340 15147
rect 30288 15104 30340 15113
rect 31760 15147 31812 15156
rect 31760 15113 31769 15147
rect 31769 15113 31803 15147
rect 31803 15113 31812 15147
rect 31760 15104 31812 15113
rect 33876 15147 33928 15156
rect 33876 15113 33885 15147
rect 33885 15113 33919 15147
rect 33919 15113 33928 15147
rect 33876 15104 33928 15113
rect 34060 15104 34112 15156
rect 36084 15104 36136 15156
rect 36268 15147 36320 15156
rect 36268 15113 36277 15147
rect 36277 15113 36311 15147
rect 36311 15113 36320 15147
rect 36268 15104 36320 15113
rect 37188 15104 37240 15156
rect 39028 15104 39080 15156
rect 39856 15104 39908 15156
rect 40500 15104 40552 15156
rect 43352 15147 43404 15156
rect 43352 15113 43361 15147
rect 43361 15113 43395 15147
rect 43395 15113 43404 15147
rect 43352 15104 43404 15113
rect 26792 15079 26844 15088
rect 26792 15045 26801 15079
rect 26801 15045 26835 15079
rect 26835 15045 26844 15079
rect 26792 15036 26844 15045
rect 9864 14900 9916 14952
rect 12164 14832 12216 14884
rect 10324 14807 10376 14816
rect 10324 14773 10333 14807
rect 10333 14773 10367 14807
rect 10367 14773 10376 14807
rect 10324 14764 10376 14773
rect 11152 14764 11204 14816
rect 11980 14764 12032 14816
rect 13360 14764 13412 14816
rect 15844 14900 15896 14952
rect 20996 14943 21048 14952
rect 20996 14909 21005 14943
rect 21005 14909 21039 14943
rect 21039 14909 21048 14943
rect 20996 14900 21048 14909
rect 21088 14900 21140 14952
rect 23388 14943 23440 14952
rect 23388 14909 23397 14943
rect 23397 14909 23431 14943
rect 23431 14909 23440 14943
rect 23388 14900 23440 14909
rect 23756 14900 23808 14952
rect 25136 14943 25188 14952
rect 25136 14909 25145 14943
rect 25145 14909 25179 14943
rect 25179 14909 25188 14943
rect 25136 14900 25188 14909
rect 14740 14875 14792 14884
rect 14740 14841 14749 14875
rect 14749 14841 14783 14875
rect 14783 14841 14792 14875
rect 14740 14832 14792 14841
rect 14096 14764 14148 14816
rect 14556 14764 14608 14816
rect 18328 14832 18380 14884
rect 21272 14832 21324 14884
rect 28540 14968 28592 15020
rect 29184 14900 29236 14952
rect 36360 14968 36412 15020
rect 39120 15079 39172 15088
rect 39120 15045 39129 15079
rect 39129 15045 39163 15079
rect 39163 15045 39172 15079
rect 39120 15036 39172 15045
rect 40776 15036 40828 15088
rect 40960 15079 41012 15088
rect 40960 15045 40969 15079
rect 40969 15045 41003 15079
rect 41003 15045 41012 15079
rect 40960 15036 41012 15045
rect 41328 15036 41380 15088
rect 38476 14968 38528 15020
rect 31116 14900 31168 14952
rect 35256 14900 35308 14952
rect 32496 14832 32548 14884
rect 33140 14832 33192 14884
rect 35624 14875 35676 14884
rect 16212 14764 16264 14816
rect 17224 14764 17276 14816
rect 17500 14807 17552 14816
rect 17500 14773 17509 14807
rect 17509 14773 17543 14807
rect 17543 14773 17552 14807
rect 17500 14764 17552 14773
rect 22560 14764 22612 14816
rect 28356 14764 28408 14816
rect 33232 14807 33284 14816
rect 33232 14773 33241 14807
rect 33241 14773 33275 14807
rect 33275 14773 33284 14807
rect 33232 14764 33284 14773
rect 34244 14807 34296 14816
rect 34244 14773 34253 14807
rect 34253 14773 34287 14807
rect 34287 14773 34296 14807
rect 34244 14764 34296 14773
rect 35624 14841 35633 14875
rect 35633 14841 35667 14875
rect 35667 14841 35676 14875
rect 35624 14832 35676 14841
rect 36912 14875 36964 14884
rect 36912 14841 36921 14875
rect 36921 14841 36955 14875
rect 36955 14841 36964 14875
rect 36912 14832 36964 14841
rect 37280 14832 37332 14884
rect 37924 14832 37976 14884
rect 43720 15036 43772 15088
rect 41236 14900 41288 14952
rect 41696 14832 41748 14884
rect 41880 14832 41932 14884
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 10324 14560 10376 14612
rect 13360 14560 13412 14612
rect 11980 14535 12032 14544
rect 11980 14501 11989 14535
rect 11989 14501 12023 14535
rect 12023 14501 12032 14535
rect 11980 14492 12032 14501
rect 17500 14560 17552 14612
rect 20996 14603 21048 14612
rect 20996 14569 21005 14603
rect 21005 14569 21039 14603
rect 21039 14569 21048 14603
rect 20996 14560 21048 14569
rect 23756 14603 23808 14612
rect 23756 14569 23765 14603
rect 23765 14569 23799 14603
rect 23799 14569 23808 14603
rect 23756 14560 23808 14569
rect 24216 14603 24268 14612
rect 24216 14569 24225 14603
rect 24225 14569 24259 14603
rect 24259 14569 24268 14603
rect 24216 14560 24268 14569
rect 25136 14603 25188 14612
rect 25136 14569 25145 14603
rect 25145 14569 25179 14603
rect 25179 14569 25188 14603
rect 25136 14560 25188 14569
rect 27528 14560 27580 14612
rect 13544 14535 13596 14544
rect 13544 14501 13553 14535
rect 13553 14501 13587 14535
rect 13587 14501 13596 14535
rect 15660 14535 15712 14544
rect 13544 14492 13596 14501
rect 15660 14501 15669 14535
rect 15669 14501 15703 14535
rect 15703 14501 15712 14535
rect 15660 14492 15712 14501
rect 15752 14535 15804 14544
rect 15752 14501 15761 14535
rect 15761 14501 15795 14535
rect 15795 14501 15804 14535
rect 15752 14492 15804 14501
rect 16580 14492 16632 14544
rect 22744 14492 22796 14544
rect 23296 14492 23348 14544
rect 26424 14492 26476 14544
rect 27252 14535 27304 14544
rect 27252 14501 27261 14535
rect 27261 14501 27295 14535
rect 27295 14501 27304 14535
rect 27252 14492 27304 14501
rect 28356 14535 28408 14544
rect 28356 14501 28365 14535
rect 28365 14501 28399 14535
rect 28399 14501 28408 14535
rect 28356 14492 28408 14501
rect 17868 14424 17920 14476
rect 18236 14424 18288 14476
rect 9680 14220 9732 14272
rect 11152 14356 11204 14408
rect 12164 14399 12216 14408
rect 12164 14365 12173 14399
rect 12173 14365 12207 14399
rect 12207 14365 12216 14399
rect 12164 14356 12216 14365
rect 13268 14356 13320 14408
rect 13544 14356 13596 14408
rect 15936 14399 15988 14408
rect 15936 14365 15945 14399
rect 15945 14365 15979 14399
rect 15979 14365 15988 14399
rect 15936 14356 15988 14365
rect 17592 14356 17644 14408
rect 19064 14424 19116 14476
rect 19984 14424 20036 14476
rect 21088 14424 21140 14476
rect 21732 14424 21784 14476
rect 23388 14424 23440 14476
rect 24952 14424 25004 14476
rect 25320 14467 25372 14476
rect 25320 14433 25329 14467
rect 25329 14433 25363 14467
rect 25363 14433 25372 14467
rect 25320 14424 25372 14433
rect 30748 14467 30800 14476
rect 30748 14433 30757 14467
rect 30757 14433 30791 14467
rect 30791 14433 30800 14467
rect 30748 14424 30800 14433
rect 31116 14560 31168 14612
rect 32496 14603 32548 14612
rect 32496 14569 32505 14603
rect 32505 14569 32539 14603
rect 32539 14569 32548 14603
rect 32496 14560 32548 14569
rect 34244 14560 34296 14612
rect 35256 14560 35308 14612
rect 35532 14560 35584 14612
rect 41880 14560 41932 14612
rect 33232 14492 33284 14544
rect 34152 14492 34204 14544
rect 36912 14492 36964 14544
rect 38476 14492 38528 14544
rect 41052 14492 41104 14544
rect 36820 14467 36872 14476
rect 36820 14433 36829 14467
rect 36829 14433 36863 14467
rect 36863 14433 36872 14467
rect 41144 14467 41196 14476
rect 36820 14424 36872 14433
rect 41144 14433 41153 14467
rect 41153 14433 41187 14467
rect 41187 14433 41196 14467
rect 41144 14424 41196 14433
rect 22284 14356 22336 14408
rect 22744 14356 22796 14408
rect 23204 14356 23256 14408
rect 26608 14399 26660 14408
rect 26608 14365 26617 14399
rect 26617 14365 26651 14399
rect 26651 14365 26660 14399
rect 26608 14356 26660 14365
rect 14740 14331 14792 14340
rect 14740 14297 14749 14331
rect 14749 14297 14783 14331
rect 14783 14297 14792 14331
rect 14740 14288 14792 14297
rect 24308 14288 24360 14340
rect 29644 14356 29696 14408
rect 31668 14356 31720 14408
rect 33600 14356 33652 14408
rect 33784 14356 33836 14408
rect 36176 14399 36228 14408
rect 36176 14365 36185 14399
rect 36185 14365 36219 14399
rect 36219 14365 36228 14399
rect 36176 14356 36228 14365
rect 38476 14399 38528 14408
rect 38476 14365 38485 14399
rect 38485 14365 38519 14399
rect 38519 14365 38528 14399
rect 38476 14356 38528 14365
rect 39212 14356 39264 14408
rect 34520 14331 34572 14340
rect 34520 14297 34529 14331
rect 34529 14297 34563 14331
rect 34563 14297 34572 14331
rect 34520 14288 34572 14297
rect 10968 14263 11020 14272
rect 10968 14229 10977 14263
rect 10977 14229 11011 14263
rect 11011 14229 11020 14263
rect 10968 14220 11020 14229
rect 13268 14263 13320 14272
rect 13268 14229 13277 14263
rect 13277 14229 13311 14263
rect 13311 14229 13320 14263
rect 13268 14220 13320 14229
rect 16396 14220 16448 14272
rect 16856 14220 16908 14272
rect 18696 14220 18748 14272
rect 29368 14263 29420 14272
rect 29368 14229 29377 14263
rect 29377 14229 29411 14263
rect 29411 14229 29420 14263
rect 29368 14220 29420 14229
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 10876 14016 10928 14068
rect 13360 14016 13412 14068
rect 13452 14016 13504 14068
rect 15752 14059 15804 14068
rect 15752 14025 15761 14059
rect 15761 14025 15795 14059
rect 15795 14025 15804 14059
rect 15752 14016 15804 14025
rect 19984 14016 20036 14068
rect 11980 13948 12032 14000
rect 15936 13948 15988 14000
rect 16028 13948 16080 14000
rect 9220 13880 9272 13932
rect 10232 13855 10284 13864
rect 10232 13821 10241 13855
rect 10241 13821 10275 13855
rect 10275 13821 10284 13855
rect 10232 13812 10284 13821
rect 10968 13812 11020 13864
rect 11980 13812 12032 13864
rect 13360 13880 13412 13932
rect 13544 13923 13596 13932
rect 13544 13889 13553 13923
rect 13553 13889 13587 13923
rect 13587 13889 13596 13923
rect 13544 13880 13596 13889
rect 14832 13923 14884 13932
rect 14832 13889 14841 13923
rect 14841 13889 14875 13923
rect 14875 13889 14884 13923
rect 14832 13880 14884 13889
rect 16212 13880 16264 13932
rect 18880 13948 18932 14000
rect 19432 13948 19484 14000
rect 17132 13880 17184 13932
rect 20260 14016 20312 14068
rect 24952 14059 25004 14068
rect 21088 13948 21140 14000
rect 24952 14025 24961 14059
rect 24961 14025 24995 14059
rect 24995 14025 25004 14059
rect 24952 14016 25004 14025
rect 26608 14016 26660 14068
rect 28356 14016 28408 14068
rect 31116 14016 31168 14068
rect 31668 14059 31720 14068
rect 31668 14025 31677 14059
rect 31677 14025 31711 14059
rect 31711 14025 31720 14059
rect 31668 14016 31720 14025
rect 32496 14016 32548 14068
rect 33600 14059 33652 14068
rect 33600 14025 33609 14059
rect 33609 14025 33643 14059
rect 33643 14025 33652 14059
rect 33600 14016 33652 14025
rect 34152 14059 34204 14068
rect 34152 14025 34161 14059
rect 34161 14025 34195 14059
rect 34195 14025 34204 14059
rect 34152 14016 34204 14025
rect 34520 14059 34572 14068
rect 34520 14025 34529 14059
rect 34529 14025 34563 14059
rect 34563 14025 34572 14059
rect 34520 14016 34572 14025
rect 35716 14016 35768 14068
rect 35992 14016 36044 14068
rect 36176 14016 36228 14068
rect 36912 14016 36964 14068
rect 41144 14016 41196 14068
rect 25320 13991 25372 14000
rect 25320 13957 25329 13991
rect 25329 13957 25363 13991
rect 25363 13957 25372 13991
rect 25320 13948 25372 13957
rect 26424 13991 26476 14000
rect 26424 13957 26433 13991
rect 26433 13957 26467 13991
rect 26467 13957 26476 13991
rect 26424 13948 26476 13957
rect 20904 13923 20956 13932
rect 20904 13889 20913 13923
rect 20913 13889 20947 13923
rect 20947 13889 20956 13923
rect 20904 13880 20956 13889
rect 24768 13880 24820 13932
rect 26700 13880 26752 13932
rect 27252 13923 27304 13932
rect 27252 13889 27261 13923
rect 27261 13889 27295 13923
rect 27295 13889 27304 13923
rect 27252 13880 27304 13889
rect 10140 13744 10192 13796
rect 10324 13744 10376 13796
rect 13268 13787 13320 13796
rect 9864 13719 9916 13728
rect 9864 13685 9873 13719
rect 9873 13685 9907 13719
rect 9907 13685 9916 13719
rect 9864 13676 9916 13685
rect 11152 13719 11204 13728
rect 11152 13685 11161 13719
rect 11161 13685 11195 13719
rect 11195 13685 11204 13719
rect 11152 13676 11204 13685
rect 13268 13753 13277 13787
rect 13277 13753 13311 13787
rect 13311 13753 13320 13787
rect 13268 13744 13320 13753
rect 13360 13787 13412 13796
rect 13360 13753 13369 13787
rect 13369 13753 13403 13787
rect 13403 13753 13412 13787
rect 13360 13744 13412 13753
rect 16212 13744 16264 13796
rect 16396 13787 16448 13796
rect 16396 13753 16405 13787
rect 16405 13753 16439 13787
rect 16439 13753 16448 13787
rect 16396 13744 16448 13753
rect 16580 13744 16632 13796
rect 13636 13676 13688 13728
rect 17408 13719 17460 13728
rect 17408 13685 17417 13719
rect 17417 13685 17451 13719
rect 17451 13685 17460 13719
rect 17408 13676 17460 13685
rect 17592 13676 17644 13728
rect 18236 13676 18288 13728
rect 18696 13719 18748 13728
rect 18696 13685 18705 13719
rect 18705 13685 18739 13719
rect 18739 13685 18748 13719
rect 18696 13676 18748 13685
rect 18972 13744 19024 13796
rect 20536 13812 20588 13864
rect 22744 13812 22796 13864
rect 25412 13812 25464 13864
rect 26424 13812 26476 13864
rect 28264 13812 28316 13864
rect 30748 13948 30800 14000
rect 38292 13948 38344 14000
rect 29644 13923 29696 13932
rect 29644 13889 29653 13923
rect 29653 13889 29687 13923
rect 29687 13889 29696 13923
rect 29644 13880 29696 13889
rect 28632 13812 28684 13864
rect 29092 13855 29144 13864
rect 29092 13821 29101 13855
rect 29101 13821 29135 13855
rect 29135 13821 29144 13855
rect 29092 13812 29144 13821
rect 31208 13812 31260 13864
rect 35624 13923 35676 13932
rect 35624 13889 35633 13923
rect 35633 13889 35667 13923
rect 35667 13889 35676 13923
rect 35624 13880 35676 13889
rect 38844 13923 38896 13932
rect 38844 13889 38853 13923
rect 38853 13889 38887 13923
rect 38887 13889 38896 13923
rect 38844 13880 38896 13889
rect 34520 13812 34572 13864
rect 41328 13948 41380 14000
rect 41052 13880 41104 13932
rect 41604 13880 41656 13932
rect 24032 13787 24084 13796
rect 24032 13753 24041 13787
rect 24041 13753 24075 13787
rect 24075 13753 24084 13787
rect 24032 13744 24084 13753
rect 24124 13787 24176 13796
rect 24124 13753 24133 13787
rect 24133 13753 24167 13787
rect 24167 13753 24176 13787
rect 24124 13744 24176 13753
rect 19248 13676 19300 13728
rect 20260 13676 20312 13728
rect 21732 13719 21784 13728
rect 21732 13685 21741 13719
rect 21741 13685 21775 13719
rect 21775 13685 21784 13719
rect 21732 13676 21784 13685
rect 22284 13676 22336 13728
rect 23020 13676 23072 13728
rect 23204 13676 23256 13728
rect 26332 13676 26384 13728
rect 26700 13787 26752 13796
rect 26700 13753 26709 13787
rect 26709 13753 26743 13787
rect 26743 13753 26752 13787
rect 26700 13744 26752 13753
rect 27528 13744 27580 13796
rect 29368 13787 29420 13796
rect 29368 13753 29377 13787
rect 29377 13753 29411 13787
rect 29411 13753 29420 13787
rect 29368 13744 29420 13753
rect 29092 13676 29144 13728
rect 32680 13676 32732 13728
rect 33600 13676 33652 13728
rect 35992 13719 36044 13728
rect 35992 13685 36001 13719
rect 36001 13685 36035 13719
rect 36035 13685 36044 13719
rect 35992 13676 36044 13685
rect 38384 13676 38436 13728
rect 38660 13676 38712 13728
rect 39580 13676 39632 13728
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 9680 13472 9732 13524
rect 13268 13472 13320 13524
rect 14096 13515 14148 13524
rect 11520 13404 11572 13456
rect 11980 13404 12032 13456
rect 12164 13447 12216 13456
rect 12164 13413 12173 13447
rect 12173 13413 12207 13447
rect 12207 13413 12216 13447
rect 12164 13404 12216 13413
rect 13636 13404 13688 13456
rect 14096 13481 14105 13515
rect 14105 13481 14139 13515
rect 14139 13481 14148 13515
rect 14096 13472 14148 13481
rect 14832 13515 14884 13524
rect 14832 13481 14841 13515
rect 14841 13481 14875 13515
rect 14875 13481 14884 13515
rect 14832 13472 14884 13481
rect 15660 13472 15712 13524
rect 19248 13472 19300 13524
rect 20996 13515 21048 13524
rect 20996 13481 21005 13515
rect 21005 13481 21039 13515
rect 21039 13481 21048 13515
rect 20996 13472 21048 13481
rect 22652 13472 22704 13524
rect 16212 13404 16264 13456
rect 17040 13404 17092 13456
rect 22836 13447 22888 13456
rect 22836 13413 22845 13447
rect 22845 13413 22879 13447
rect 22879 13413 22888 13447
rect 22836 13404 22888 13413
rect 23020 13404 23072 13456
rect 24124 13472 24176 13524
rect 26332 13515 26384 13524
rect 26332 13481 26341 13515
rect 26341 13481 26375 13515
rect 26375 13481 26384 13515
rect 26332 13472 26384 13481
rect 28264 13472 28316 13524
rect 28632 13515 28684 13524
rect 28632 13481 28641 13515
rect 28641 13481 28675 13515
rect 28675 13481 28684 13515
rect 28632 13472 28684 13481
rect 29368 13472 29420 13524
rect 35624 13515 35676 13524
rect 35624 13481 35633 13515
rect 35633 13481 35667 13515
rect 35667 13481 35676 13515
rect 35624 13472 35676 13481
rect 38384 13472 38436 13524
rect 10048 13379 10100 13388
rect 10048 13345 10057 13379
rect 10057 13345 10091 13379
rect 10091 13345 10100 13379
rect 10048 13336 10100 13345
rect 10232 13379 10284 13388
rect 10232 13345 10241 13379
rect 10241 13345 10275 13379
rect 10275 13345 10284 13379
rect 10232 13336 10284 13345
rect 15200 13379 15252 13388
rect 15200 13345 15209 13379
rect 15209 13345 15243 13379
rect 15243 13345 15252 13379
rect 15200 13336 15252 13345
rect 18696 13336 18748 13388
rect 19248 13336 19300 13388
rect 20444 13336 20496 13388
rect 21088 13336 21140 13388
rect 21180 13336 21232 13388
rect 11336 13268 11388 13320
rect 13912 13268 13964 13320
rect 16120 13268 16172 13320
rect 16856 13311 16908 13320
rect 16856 13277 16865 13311
rect 16865 13277 16899 13311
rect 16899 13277 16908 13311
rect 16856 13268 16908 13277
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 23112 13311 23164 13320
rect 23112 13277 23121 13311
rect 23121 13277 23155 13311
rect 23155 13277 23164 13311
rect 23112 13268 23164 13277
rect 26976 13404 27028 13456
rect 35532 13404 35584 13456
rect 35992 13404 36044 13456
rect 37648 13404 37700 13456
rect 39488 13447 39540 13456
rect 39488 13413 39497 13447
rect 39497 13413 39531 13447
rect 39531 13413 39540 13447
rect 39488 13404 39540 13413
rect 30472 13336 30524 13388
rect 33140 13379 33192 13388
rect 33140 13345 33149 13379
rect 33149 13345 33183 13379
rect 33183 13345 33192 13379
rect 33140 13336 33192 13345
rect 34704 13336 34756 13388
rect 24584 13268 24636 13320
rect 24768 13311 24820 13320
rect 24768 13277 24777 13311
rect 24777 13277 24811 13311
rect 24811 13277 24820 13311
rect 24768 13268 24820 13277
rect 26516 13311 26568 13320
rect 26516 13277 26525 13311
rect 26525 13277 26559 13311
rect 26559 13277 26568 13311
rect 26516 13268 26568 13277
rect 28264 13311 28316 13320
rect 28264 13277 28273 13311
rect 28273 13277 28307 13311
rect 28307 13277 28316 13311
rect 28264 13268 28316 13277
rect 35808 13311 35860 13320
rect 35808 13277 35817 13311
rect 35817 13277 35851 13311
rect 35851 13277 35860 13311
rect 35808 13268 35860 13277
rect 37924 13268 37976 13320
rect 39212 13268 39264 13320
rect 40224 13268 40276 13320
rect 38108 13200 38160 13252
rect 38384 13243 38436 13252
rect 38384 13209 38393 13243
rect 38393 13209 38427 13243
rect 38427 13209 38436 13243
rect 38384 13200 38436 13209
rect 10140 13132 10192 13184
rect 16580 13175 16632 13184
rect 16580 13141 16589 13175
rect 16589 13141 16623 13175
rect 16623 13141 16632 13175
rect 16580 13132 16632 13141
rect 17868 13175 17920 13184
rect 17868 13141 17877 13175
rect 17877 13141 17911 13175
rect 17911 13141 17920 13175
rect 17868 13132 17920 13141
rect 20536 13132 20588 13184
rect 22744 13132 22796 13184
rect 22928 13132 22980 13184
rect 25596 13175 25648 13184
rect 25596 13141 25605 13175
rect 25605 13141 25639 13175
rect 25639 13141 25648 13175
rect 25596 13132 25648 13141
rect 27804 13175 27856 13184
rect 27804 13141 27813 13175
rect 27813 13141 27847 13175
rect 27847 13141 27856 13175
rect 27804 13132 27856 13141
rect 29460 13175 29512 13184
rect 29460 13141 29469 13175
rect 29469 13141 29503 13175
rect 29503 13141 29512 13175
rect 29460 13132 29512 13141
rect 31024 13175 31076 13184
rect 31024 13141 31033 13175
rect 31033 13141 31067 13175
rect 31067 13141 31076 13175
rect 31024 13132 31076 13141
rect 32588 13132 32640 13184
rect 33324 13175 33376 13184
rect 33324 13141 33333 13175
rect 33333 13141 33367 13175
rect 33367 13141 33376 13175
rect 33324 13132 33376 13141
rect 37648 13132 37700 13184
rect 37832 13132 37884 13184
rect 40408 13132 40460 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 11336 12928 11388 12980
rect 11520 12971 11572 12980
rect 11520 12937 11529 12971
rect 11529 12937 11563 12971
rect 11563 12937 11572 12971
rect 11520 12928 11572 12937
rect 13636 12928 13688 12980
rect 16120 12971 16172 12980
rect 16120 12937 16129 12971
rect 16129 12937 16163 12971
rect 16163 12937 16172 12971
rect 16120 12928 16172 12937
rect 16212 12928 16264 12980
rect 17868 12928 17920 12980
rect 22652 12928 22704 12980
rect 24032 12928 24084 12980
rect 24584 12971 24636 12980
rect 24584 12937 24593 12971
rect 24593 12937 24627 12971
rect 24627 12937 24636 12971
rect 24584 12928 24636 12937
rect 25596 12928 25648 12980
rect 29184 12928 29236 12980
rect 30472 12971 30524 12980
rect 30472 12937 30481 12971
rect 30481 12937 30515 12971
rect 30515 12937 30524 12971
rect 30472 12928 30524 12937
rect 32588 12971 32640 12980
rect 32588 12937 32597 12971
rect 32597 12937 32631 12971
rect 32631 12937 32640 12971
rect 32588 12928 32640 12937
rect 36912 12928 36964 12980
rect 37648 12971 37700 12980
rect 37648 12937 37657 12971
rect 37657 12937 37691 12971
rect 37691 12937 37700 12971
rect 37648 12928 37700 12937
rect 38200 12928 38252 12980
rect 39488 12928 39540 12980
rect 39948 12928 40000 12980
rect 40224 12971 40276 12980
rect 40224 12937 40233 12971
rect 40233 12937 40267 12971
rect 40267 12937 40276 12971
rect 40224 12928 40276 12937
rect 11152 12860 11204 12912
rect 10048 12792 10100 12844
rect 14096 12860 14148 12912
rect 18328 12903 18380 12912
rect 18328 12869 18337 12903
rect 18337 12869 18371 12903
rect 18371 12869 18380 12903
rect 18328 12860 18380 12869
rect 22836 12860 22888 12912
rect 13912 12835 13964 12844
rect 13912 12801 13921 12835
rect 13921 12801 13955 12835
rect 13955 12801 13964 12835
rect 13912 12792 13964 12801
rect 18236 12792 18288 12844
rect 20996 12792 21048 12844
rect 9036 12767 9088 12776
rect 9036 12733 9045 12767
rect 9045 12733 9079 12767
rect 9079 12733 9088 12767
rect 9036 12724 9088 12733
rect 9680 12724 9732 12776
rect 10140 12767 10192 12776
rect 10140 12733 10149 12767
rect 10149 12733 10183 12767
rect 10183 12733 10192 12767
rect 10140 12724 10192 12733
rect 10232 12724 10284 12776
rect 12900 12724 12952 12776
rect 14188 12767 14240 12776
rect 12808 12656 12860 12708
rect 14188 12733 14197 12767
rect 14197 12733 14231 12767
rect 14231 12733 14240 12767
rect 14188 12724 14240 12733
rect 15384 12767 15436 12776
rect 15384 12733 15393 12767
rect 15393 12733 15427 12767
rect 15427 12733 15436 12767
rect 15384 12724 15436 12733
rect 15752 12656 15804 12708
rect 16580 12699 16632 12708
rect 16580 12665 16589 12699
rect 16589 12665 16623 12699
rect 16623 12665 16632 12699
rect 16580 12656 16632 12665
rect 18512 12724 18564 12776
rect 23940 12724 23992 12776
rect 25136 12767 25188 12776
rect 25136 12733 25145 12767
rect 25145 12733 25179 12767
rect 25179 12733 25188 12767
rect 25136 12724 25188 12733
rect 8668 12631 8720 12640
rect 8668 12597 8677 12631
rect 8677 12597 8711 12631
rect 8711 12597 8720 12631
rect 8668 12588 8720 12597
rect 10232 12631 10284 12640
rect 10232 12597 10241 12631
rect 10241 12597 10275 12631
rect 10275 12597 10284 12631
rect 10232 12588 10284 12597
rect 15016 12631 15068 12640
rect 15016 12597 15025 12631
rect 15025 12597 15059 12631
rect 15059 12597 15068 12631
rect 15016 12588 15068 12597
rect 17500 12631 17552 12640
rect 17500 12597 17509 12631
rect 17509 12597 17543 12631
rect 17543 12597 17552 12631
rect 17500 12588 17552 12597
rect 21272 12656 21324 12708
rect 26976 12860 27028 12912
rect 28632 12860 28684 12912
rect 33140 12860 33192 12912
rect 37832 12860 37884 12912
rect 38476 12860 38528 12912
rect 29460 12792 29512 12844
rect 35808 12835 35860 12844
rect 35808 12801 35817 12835
rect 35817 12801 35851 12835
rect 35851 12801 35860 12835
rect 35808 12792 35860 12801
rect 38384 12792 38436 12844
rect 27160 12724 27212 12776
rect 27804 12724 27856 12776
rect 28724 12724 28776 12776
rect 30472 12724 30524 12776
rect 31024 12767 31076 12776
rect 31024 12733 31033 12767
rect 31033 12733 31067 12767
rect 31067 12733 31076 12767
rect 31024 12724 31076 12733
rect 32588 12724 32640 12776
rect 35348 12767 35400 12776
rect 35348 12733 35357 12767
rect 35357 12733 35391 12767
rect 35391 12733 35400 12767
rect 35348 12724 35400 12733
rect 35532 12767 35584 12776
rect 35532 12733 35541 12767
rect 35541 12733 35575 12767
rect 35575 12733 35584 12767
rect 35532 12724 35584 12733
rect 28632 12699 28684 12708
rect 28632 12665 28641 12699
rect 28641 12665 28675 12699
rect 28675 12665 28684 12699
rect 28632 12656 28684 12665
rect 30932 12699 30984 12708
rect 30932 12665 30941 12699
rect 30941 12665 30975 12699
rect 30975 12665 30984 12699
rect 30932 12656 30984 12665
rect 32404 12656 32456 12708
rect 32772 12699 32824 12708
rect 32772 12665 32781 12699
rect 32781 12665 32815 12699
rect 32815 12665 32824 12699
rect 32772 12656 32824 12665
rect 35440 12656 35492 12708
rect 38200 12724 38252 12776
rect 38936 12699 38988 12708
rect 38936 12665 38945 12699
rect 38945 12665 38979 12699
rect 38979 12665 38988 12699
rect 38936 12656 38988 12665
rect 19248 12588 19300 12640
rect 20444 12631 20496 12640
rect 20444 12597 20453 12631
rect 20453 12597 20487 12631
rect 20487 12597 20496 12631
rect 20444 12588 20496 12597
rect 21824 12631 21876 12640
rect 21824 12597 21833 12631
rect 21833 12597 21867 12631
rect 21867 12597 21876 12631
rect 21824 12588 21876 12597
rect 27436 12631 27488 12640
rect 27436 12597 27445 12631
rect 27445 12597 27479 12631
rect 27479 12597 27488 12631
rect 27436 12588 27488 12597
rect 31944 12631 31996 12640
rect 31944 12597 31953 12631
rect 31953 12597 31987 12631
rect 31987 12597 31996 12631
rect 31944 12588 31996 12597
rect 34704 12631 34756 12640
rect 34704 12597 34713 12631
rect 34713 12597 34747 12631
rect 34747 12597 34756 12631
rect 34704 12588 34756 12597
rect 36544 12588 36596 12640
rect 41696 12588 41748 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 9036 12384 9088 12436
rect 13912 12384 13964 12436
rect 14188 12384 14240 12436
rect 15384 12384 15436 12436
rect 17224 12384 17276 12436
rect 22008 12384 22060 12436
rect 22560 12384 22612 12436
rect 23388 12427 23440 12436
rect 23388 12393 23397 12427
rect 23397 12393 23431 12427
rect 23431 12393 23440 12427
rect 23388 12384 23440 12393
rect 23940 12427 23992 12436
rect 23940 12393 23949 12427
rect 23949 12393 23983 12427
rect 23983 12393 23992 12427
rect 23940 12384 23992 12393
rect 25136 12427 25188 12436
rect 25136 12393 25145 12427
rect 25145 12393 25179 12427
rect 25179 12393 25188 12427
rect 25136 12384 25188 12393
rect 31208 12427 31260 12436
rect 31208 12393 31217 12427
rect 31217 12393 31251 12427
rect 31251 12393 31260 12427
rect 31208 12384 31260 12393
rect 35348 12384 35400 12436
rect 37924 12427 37976 12436
rect 37924 12393 37933 12427
rect 37933 12393 37967 12427
rect 37967 12393 37976 12427
rect 37924 12384 37976 12393
rect 38936 12427 38988 12436
rect 38936 12393 38945 12427
rect 38945 12393 38979 12427
rect 38979 12393 38988 12427
rect 38936 12384 38988 12393
rect 39396 12427 39448 12436
rect 39396 12393 39405 12427
rect 39405 12393 39439 12427
rect 39439 12393 39448 12427
rect 39396 12384 39448 12393
rect 39948 12427 40000 12436
rect 39948 12393 39957 12427
rect 39957 12393 39991 12427
rect 39991 12393 40000 12427
rect 39948 12384 40000 12393
rect 41696 12427 41748 12436
rect 41696 12393 41705 12427
rect 41705 12393 41739 12427
rect 41739 12393 41748 12427
rect 41696 12384 41748 12393
rect 9956 12359 10008 12368
rect 9956 12325 9965 12359
rect 9965 12325 9999 12359
rect 9999 12325 10008 12359
rect 9956 12316 10008 12325
rect 10324 12316 10376 12368
rect 10508 12359 10560 12368
rect 10508 12325 10517 12359
rect 10517 12325 10551 12359
rect 10551 12325 10560 12359
rect 10508 12316 10560 12325
rect 13636 12316 13688 12368
rect 16212 12316 16264 12368
rect 18328 12316 18380 12368
rect 21272 12316 21324 12368
rect 28264 12359 28316 12368
rect 28264 12325 28273 12359
rect 28273 12325 28307 12359
rect 28307 12325 28316 12359
rect 28264 12316 28316 12325
rect 30472 12316 30524 12368
rect 30932 12316 30984 12368
rect 32588 12316 32640 12368
rect 33784 12316 33836 12368
rect 40868 12316 40920 12368
rect 41604 12316 41656 12368
rect 10232 12291 10284 12300
rect 10232 12257 10241 12291
rect 10241 12257 10275 12291
rect 10275 12257 10284 12291
rect 10232 12248 10284 12257
rect 15200 12248 15252 12300
rect 20076 12248 20128 12300
rect 24860 12291 24912 12300
rect 24860 12257 24869 12291
rect 24869 12257 24903 12291
rect 24903 12257 24912 12291
rect 24860 12248 24912 12257
rect 25228 12248 25280 12300
rect 26792 12248 26844 12300
rect 27436 12248 27488 12300
rect 27712 12291 27764 12300
rect 27712 12257 27721 12291
rect 27721 12257 27755 12291
rect 27755 12257 27764 12291
rect 27712 12248 27764 12257
rect 28724 12291 28776 12300
rect 28724 12257 28733 12291
rect 28733 12257 28767 12291
rect 28767 12257 28776 12291
rect 28724 12248 28776 12257
rect 32404 12291 32456 12300
rect 12532 12223 12584 12232
rect 12532 12189 12541 12223
rect 12541 12189 12575 12223
rect 12575 12189 12584 12223
rect 12532 12180 12584 12189
rect 16028 12223 16080 12232
rect 16028 12189 16037 12223
rect 16037 12189 16071 12223
rect 16071 12189 16080 12223
rect 16028 12180 16080 12189
rect 17776 12223 17828 12232
rect 17776 12189 17785 12223
rect 17785 12189 17819 12223
rect 17819 12189 17828 12223
rect 17776 12180 17828 12189
rect 20996 12180 21048 12232
rect 22744 12180 22796 12232
rect 14004 12112 14056 12164
rect 18696 12112 18748 12164
rect 16948 12087 17000 12096
rect 16948 12053 16957 12087
rect 16957 12053 16991 12087
rect 16991 12053 17000 12087
rect 16948 12044 17000 12053
rect 17224 12044 17276 12096
rect 20812 12044 20864 12096
rect 21088 12087 21140 12096
rect 21088 12053 21097 12087
rect 21097 12053 21131 12087
rect 21131 12053 21140 12087
rect 21088 12044 21140 12053
rect 24216 12087 24268 12096
rect 24216 12053 24225 12087
rect 24225 12053 24259 12087
rect 24259 12053 24268 12087
rect 24216 12044 24268 12053
rect 26516 12044 26568 12096
rect 32404 12257 32413 12291
rect 32413 12257 32447 12291
rect 32447 12257 32456 12291
rect 32404 12248 32456 12257
rect 33324 12248 33376 12300
rect 34796 12248 34848 12300
rect 36176 12248 36228 12300
rect 30564 12180 30616 12232
rect 33968 12223 34020 12232
rect 33968 12189 33977 12223
rect 33977 12189 34011 12223
rect 34011 12189 34020 12223
rect 33968 12180 34020 12189
rect 34244 12223 34296 12232
rect 34244 12189 34253 12223
rect 34253 12189 34287 12223
rect 34287 12189 34296 12223
rect 34244 12180 34296 12189
rect 35624 12180 35676 12232
rect 38844 12180 38896 12232
rect 39028 12223 39080 12232
rect 39028 12189 39037 12223
rect 39037 12189 39071 12223
rect 39071 12189 39080 12223
rect 39028 12180 39080 12189
rect 41144 12180 41196 12232
rect 30288 12044 30340 12096
rect 35256 12044 35308 12096
rect 36636 12087 36688 12096
rect 36636 12053 36645 12087
rect 36645 12053 36679 12087
rect 36679 12053 36688 12087
rect 36636 12044 36688 12053
rect 36912 12087 36964 12096
rect 36912 12053 36921 12087
rect 36921 12053 36955 12087
rect 36955 12053 36964 12087
rect 36912 12044 36964 12053
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 10232 11840 10284 11892
rect 15844 11883 15896 11892
rect 15844 11849 15853 11883
rect 15853 11849 15887 11883
rect 15887 11849 15896 11883
rect 15844 11840 15896 11849
rect 16028 11840 16080 11892
rect 16948 11840 17000 11892
rect 18328 11840 18380 11892
rect 20076 11840 20128 11892
rect 21272 11840 21324 11892
rect 8668 11772 8720 11824
rect 13636 11772 13688 11824
rect 16212 11815 16264 11824
rect 10324 11679 10376 11688
rect 10324 11645 10333 11679
rect 10333 11645 10367 11679
rect 10367 11645 10376 11679
rect 10324 11636 10376 11645
rect 10508 11568 10560 11620
rect 12532 11704 12584 11756
rect 15016 11704 15068 11756
rect 12716 11679 12768 11688
rect 12716 11645 12725 11679
rect 12725 11645 12759 11679
rect 12759 11645 12768 11679
rect 12716 11636 12768 11645
rect 12808 11636 12860 11688
rect 16212 11781 16221 11815
rect 16221 11781 16255 11815
rect 16255 11781 16264 11815
rect 16212 11772 16264 11781
rect 16396 11772 16448 11824
rect 16948 11636 17000 11688
rect 21088 11772 21140 11824
rect 22928 11840 22980 11892
rect 30932 11883 30984 11892
rect 30932 11849 30941 11883
rect 30941 11849 30975 11883
rect 30975 11849 30984 11883
rect 30932 11840 30984 11849
rect 22560 11772 22612 11824
rect 23388 11815 23440 11824
rect 23388 11781 23397 11815
rect 23397 11781 23431 11815
rect 23431 11781 23440 11815
rect 23388 11772 23440 11781
rect 20996 11747 21048 11756
rect 20996 11713 21005 11747
rect 21005 11713 21039 11747
rect 21039 11713 21048 11747
rect 20996 11704 21048 11713
rect 18972 11636 19024 11688
rect 20444 11636 20496 11688
rect 20812 11636 20864 11688
rect 23572 11704 23624 11756
rect 24216 11704 24268 11756
rect 26516 11747 26568 11756
rect 26516 11713 26525 11747
rect 26525 11713 26559 11747
rect 26559 11713 26568 11747
rect 26516 11704 26568 11713
rect 28356 11704 28408 11756
rect 22468 11679 22520 11688
rect 22468 11645 22477 11679
rect 22477 11645 22511 11679
rect 22511 11645 22520 11679
rect 22468 11636 22520 11645
rect 23020 11636 23072 11688
rect 24860 11679 24912 11688
rect 24860 11645 24869 11679
rect 24869 11645 24903 11679
rect 24903 11645 24912 11679
rect 24860 11636 24912 11645
rect 22744 11611 22796 11620
rect 22744 11577 22753 11611
rect 22753 11577 22787 11611
rect 22787 11577 22796 11611
rect 22744 11568 22796 11577
rect 24676 11568 24728 11620
rect 25872 11636 25924 11688
rect 30288 11679 30340 11688
rect 26792 11611 26844 11620
rect 26792 11577 26801 11611
rect 26801 11577 26835 11611
rect 26835 11577 26844 11611
rect 26792 11568 26844 11577
rect 27528 11611 27580 11620
rect 27528 11577 27537 11611
rect 27537 11577 27571 11611
rect 27571 11577 27580 11611
rect 27528 11568 27580 11577
rect 27896 11568 27948 11620
rect 28264 11568 28316 11620
rect 30288 11645 30297 11679
rect 30297 11645 30331 11679
rect 30331 11645 30340 11679
rect 30288 11636 30340 11645
rect 31944 11840 31996 11892
rect 32404 11840 32456 11892
rect 33968 11840 34020 11892
rect 36176 11883 36228 11892
rect 36176 11849 36185 11883
rect 36185 11849 36219 11883
rect 36219 11849 36228 11883
rect 36176 11840 36228 11849
rect 38292 11883 38344 11892
rect 38292 11849 38301 11883
rect 38301 11849 38335 11883
rect 38335 11849 38344 11883
rect 38292 11840 38344 11849
rect 39396 11840 39448 11892
rect 40868 11883 40920 11892
rect 40868 11849 40877 11883
rect 40877 11849 40911 11883
rect 40911 11849 40920 11883
rect 40868 11840 40920 11849
rect 33784 11772 33836 11824
rect 32680 11747 32732 11756
rect 32680 11713 32689 11747
rect 32689 11713 32723 11747
rect 32723 11713 32732 11747
rect 32680 11704 32732 11713
rect 34244 11704 34296 11756
rect 36912 11704 36964 11756
rect 39028 11704 39080 11756
rect 36636 11636 36688 11688
rect 38292 11636 38344 11688
rect 38844 11636 38896 11688
rect 30380 11568 30432 11620
rect 30564 11611 30616 11620
rect 30564 11577 30573 11611
rect 30573 11577 30607 11611
rect 30607 11577 30616 11611
rect 30564 11568 30616 11577
rect 32772 11611 32824 11620
rect 32772 11577 32781 11611
rect 32781 11577 32815 11611
rect 32815 11577 32824 11611
rect 32772 11568 32824 11577
rect 34336 11568 34388 11620
rect 36544 11611 36596 11620
rect 36544 11577 36553 11611
rect 36553 11577 36587 11611
rect 36587 11577 36596 11611
rect 36544 11568 36596 11577
rect 39396 11568 39448 11620
rect 18512 11500 18564 11552
rect 25228 11543 25280 11552
rect 25228 11509 25237 11543
rect 25237 11509 25271 11543
rect 25271 11509 25280 11543
rect 25228 11500 25280 11509
rect 27988 11500 28040 11552
rect 28724 11543 28776 11552
rect 28724 11509 28733 11543
rect 28733 11509 28767 11543
rect 28767 11509 28776 11543
rect 28724 11500 28776 11509
rect 37648 11543 37700 11552
rect 37648 11509 37657 11543
rect 37657 11509 37691 11543
rect 37691 11509 37700 11543
rect 37648 11500 37700 11509
rect 41144 11543 41196 11552
rect 41144 11509 41153 11543
rect 41153 11509 41187 11543
rect 41187 11509 41196 11543
rect 41144 11500 41196 11509
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 9956 11339 10008 11348
rect 9956 11305 9965 11339
rect 9965 11305 9999 11339
rect 9999 11305 10008 11339
rect 9956 11296 10008 11305
rect 10324 11339 10376 11348
rect 10324 11305 10333 11339
rect 10333 11305 10367 11339
rect 10367 11305 10376 11339
rect 10324 11296 10376 11305
rect 11796 11296 11848 11348
rect 12440 11296 12492 11348
rect 15016 11339 15068 11348
rect 15016 11305 15025 11339
rect 15025 11305 15059 11339
rect 15059 11305 15068 11339
rect 15016 11296 15068 11305
rect 16028 11339 16080 11348
rect 16028 11305 16037 11339
rect 16037 11305 16071 11339
rect 16071 11305 16080 11339
rect 16028 11296 16080 11305
rect 17776 11339 17828 11348
rect 17776 11305 17785 11339
rect 17785 11305 17819 11339
rect 17819 11305 17828 11339
rect 17776 11296 17828 11305
rect 18972 11296 19024 11348
rect 22744 11296 22796 11348
rect 24584 11296 24636 11348
rect 26608 11339 26660 11348
rect 26608 11305 26617 11339
rect 26617 11305 26651 11339
rect 26651 11305 26660 11339
rect 26608 11296 26660 11305
rect 27712 11296 27764 11348
rect 28264 11296 28316 11348
rect 30564 11339 30616 11348
rect 30564 11305 30573 11339
rect 30573 11305 30607 11339
rect 30607 11305 30616 11339
rect 30564 11296 30616 11305
rect 32680 11339 32732 11348
rect 32680 11305 32689 11339
rect 32689 11305 32723 11339
rect 32723 11305 32732 11339
rect 32680 11296 32732 11305
rect 36176 11296 36228 11348
rect 11888 11228 11940 11280
rect 17684 11228 17736 11280
rect 19340 11228 19392 11280
rect 20352 11228 20404 11280
rect 20720 11228 20772 11280
rect 23572 11271 23624 11280
rect 23572 11237 23581 11271
rect 23581 11237 23615 11271
rect 23615 11237 23624 11271
rect 23572 11228 23624 11237
rect 12532 11203 12584 11212
rect 12532 11169 12541 11203
rect 12541 11169 12575 11203
rect 12575 11169 12584 11203
rect 12532 11160 12584 11169
rect 12900 11203 12952 11212
rect 12900 11169 12909 11203
rect 12909 11169 12943 11203
rect 12943 11169 12952 11203
rect 12900 11160 12952 11169
rect 13728 11203 13780 11212
rect 13728 11169 13737 11203
rect 13737 11169 13771 11203
rect 13771 11169 13780 11203
rect 13728 11160 13780 11169
rect 13820 11160 13872 11212
rect 16212 11203 16264 11212
rect 16212 11169 16221 11203
rect 16221 11169 16255 11203
rect 16255 11169 16264 11203
rect 16212 11160 16264 11169
rect 10324 11092 10376 11144
rect 14280 11135 14332 11144
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 15384 11092 15436 11144
rect 18236 11160 18288 11212
rect 17408 11092 17460 11144
rect 18972 11160 19024 11212
rect 19892 11160 19944 11212
rect 23020 11203 23072 11212
rect 23020 11169 23029 11203
rect 23029 11169 23063 11203
rect 23063 11169 23072 11203
rect 23020 11160 23072 11169
rect 23204 11160 23256 11212
rect 23664 11160 23716 11212
rect 24308 11160 24360 11212
rect 29184 11228 29236 11280
rect 25044 11160 25096 11212
rect 25320 11160 25372 11212
rect 26056 11160 26108 11212
rect 26700 11160 26752 11212
rect 27988 11160 28040 11212
rect 28264 11160 28316 11212
rect 30288 11228 30340 11280
rect 35532 11228 35584 11280
rect 36912 11228 36964 11280
rect 37648 11228 37700 11280
rect 25780 11135 25832 11144
rect 25780 11101 25789 11135
rect 25789 11101 25823 11135
rect 25823 11101 25832 11135
rect 31852 11160 31904 11212
rect 35256 11160 35308 11212
rect 36268 11203 36320 11212
rect 36268 11169 36277 11203
rect 36277 11169 36311 11203
rect 36311 11169 36320 11203
rect 36268 11160 36320 11169
rect 36544 11203 36596 11212
rect 36544 11169 36553 11203
rect 36553 11169 36587 11203
rect 36587 11169 36596 11203
rect 36544 11160 36596 11169
rect 39396 11160 39448 11212
rect 40500 11296 40552 11348
rect 41144 11228 41196 11280
rect 39764 11203 39816 11212
rect 39764 11169 39773 11203
rect 39773 11169 39807 11203
rect 39807 11169 39816 11203
rect 39764 11160 39816 11169
rect 25780 11092 25832 11101
rect 29736 11092 29788 11144
rect 30564 11092 30616 11144
rect 36728 11092 36780 11144
rect 38292 11135 38344 11144
rect 38292 11101 38301 11135
rect 38301 11101 38335 11135
rect 38335 11101 38344 11135
rect 38292 11092 38344 11101
rect 15752 11024 15804 11076
rect 22468 11024 22520 11076
rect 27252 11024 27304 11076
rect 16212 10956 16264 11008
rect 17132 10956 17184 11008
rect 20812 10956 20864 11008
rect 22836 10956 22888 11008
rect 28356 10956 28408 11008
rect 29276 10999 29328 11008
rect 29276 10965 29285 10999
rect 29285 10965 29319 10999
rect 29319 10965 29328 10999
rect 29276 10956 29328 10965
rect 32496 10956 32548 11008
rect 34704 10956 34756 11008
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 10784 10795 10836 10804
rect 10784 10761 10793 10795
rect 10793 10761 10827 10795
rect 10827 10761 10836 10795
rect 10784 10752 10836 10761
rect 11888 10795 11940 10804
rect 11888 10761 11897 10795
rect 11897 10761 11931 10795
rect 11931 10761 11940 10795
rect 11888 10752 11940 10761
rect 12716 10795 12768 10804
rect 12716 10761 12725 10795
rect 12725 10761 12759 10795
rect 12759 10761 12768 10795
rect 12716 10752 12768 10761
rect 14648 10752 14700 10804
rect 18420 10752 18472 10804
rect 19064 10795 19116 10804
rect 16856 10684 16908 10736
rect 17132 10727 17184 10736
rect 17132 10693 17141 10727
rect 17141 10693 17175 10727
rect 17175 10693 17184 10727
rect 17132 10684 17184 10693
rect 17408 10727 17460 10736
rect 17408 10693 17417 10727
rect 17417 10693 17451 10727
rect 17451 10693 17460 10727
rect 17408 10684 17460 10693
rect 9680 10659 9732 10668
rect 9680 10625 9689 10659
rect 9689 10625 9723 10659
rect 9723 10625 9732 10659
rect 9680 10616 9732 10625
rect 13636 10616 13688 10668
rect 15568 10659 15620 10668
rect 10692 10591 10744 10600
rect 10692 10557 10701 10591
rect 10701 10557 10735 10591
rect 10735 10557 10744 10591
rect 12440 10591 12492 10600
rect 10692 10548 10744 10557
rect 9772 10480 9824 10532
rect 10508 10523 10560 10532
rect 10508 10489 10517 10523
rect 10517 10489 10551 10523
rect 10551 10489 10560 10523
rect 10508 10480 10560 10489
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 12440 10548 12492 10557
rect 12532 10480 12584 10532
rect 9220 10412 9272 10464
rect 12716 10412 12768 10464
rect 13728 10480 13780 10532
rect 14280 10523 14332 10532
rect 14280 10489 14289 10523
rect 14289 10489 14323 10523
rect 14323 10489 14332 10523
rect 14280 10480 14332 10489
rect 15568 10625 15577 10659
rect 15577 10625 15611 10659
rect 15611 10625 15620 10659
rect 15568 10616 15620 10625
rect 17684 10616 17736 10668
rect 15660 10548 15712 10600
rect 19064 10761 19073 10795
rect 19073 10761 19107 10795
rect 19107 10761 19116 10795
rect 19064 10752 19116 10761
rect 20720 10752 20772 10804
rect 23020 10795 23072 10804
rect 23020 10761 23029 10795
rect 23029 10761 23063 10795
rect 23063 10761 23072 10795
rect 23020 10752 23072 10761
rect 24308 10795 24360 10804
rect 24308 10761 24317 10795
rect 24317 10761 24351 10795
rect 24351 10761 24360 10795
rect 24308 10752 24360 10761
rect 28264 10752 28316 10804
rect 28356 10752 28408 10804
rect 29736 10795 29788 10804
rect 29736 10761 29745 10795
rect 29745 10761 29779 10795
rect 29779 10761 29788 10795
rect 29736 10752 29788 10761
rect 30932 10752 30984 10804
rect 35256 10752 35308 10804
rect 36268 10752 36320 10804
rect 36544 10795 36596 10804
rect 36544 10761 36553 10795
rect 36553 10761 36587 10795
rect 36587 10761 36596 10795
rect 36544 10752 36596 10761
rect 36728 10752 36780 10804
rect 37648 10752 37700 10804
rect 39396 10795 39448 10804
rect 39396 10761 39405 10795
rect 39405 10761 39439 10795
rect 39439 10761 39448 10795
rect 39396 10752 39448 10761
rect 27988 10684 28040 10736
rect 29184 10684 29236 10736
rect 34704 10727 34756 10736
rect 34704 10693 34713 10727
rect 34713 10693 34747 10727
rect 34747 10693 34756 10727
rect 34704 10684 34756 10693
rect 37740 10684 37792 10736
rect 38844 10684 38896 10736
rect 38936 10684 38988 10736
rect 39764 10684 39816 10736
rect 19892 10480 19944 10532
rect 20904 10548 20956 10600
rect 26608 10659 26660 10668
rect 26608 10625 26617 10659
rect 26617 10625 26651 10659
rect 26651 10625 26660 10659
rect 26608 10616 26660 10625
rect 30564 10659 30616 10668
rect 30564 10625 30573 10659
rect 30573 10625 30607 10659
rect 30607 10625 30616 10659
rect 30564 10616 30616 10625
rect 33508 10616 33560 10668
rect 22836 10548 22888 10600
rect 23572 10591 23624 10600
rect 23572 10557 23581 10591
rect 23581 10557 23615 10591
rect 23615 10557 23624 10591
rect 23572 10548 23624 10557
rect 24860 10591 24912 10600
rect 24860 10557 24869 10591
rect 24869 10557 24903 10591
rect 24903 10557 24912 10591
rect 24860 10548 24912 10557
rect 29276 10591 29328 10600
rect 29276 10557 29320 10591
rect 29320 10557 29328 10591
rect 29276 10548 29328 10557
rect 20996 10480 21048 10532
rect 21548 10523 21600 10532
rect 21548 10489 21557 10523
rect 21557 10489 21591 10523
rect 21591 10489 21600 10523
rect 21548 10480 21600 10489
rect 23296 10480 23348 10532
rect 24676 10480 24728 10532
rect 32588 10523 32640 10532
rect 32588 10489 32597 10523
rect 32597 10489 32631 10523
rect 32631 10489 32640 10523
rect 32588 10480 32640 10489
rect 33140 10523 33192 10532
rect 33140 10489 33149 10523
rect 33149 10489 33183 10523
rect 33183 10489 33192 10523
rect 34980 10523 35032 10532
rect 33140 10480 33192 10489
rect 34980 10489 34989 10523
rect 34989 10489 35023 10523
rect 35023 10489 35032 10523
rect 34980 10480 35032 10489
rect 13820 10455 13872 10464
rect 13820 10421 13829 10455
rect 13829 10421 13863 10455
rect 13863 10421 13872 10455
rect 15200 10455 15252 10464
rect 13820 10412 13872 10421
rect 15200 10421 15209 10455
rect 15209 10421 15243 10455
rect 15243 10421 15252 10455
rect 15200 10412 15252 10421
rect 18328 10455 18380 10464
rect 18328 10421 18337 10455
rect 18337 10421 18371 10455
rect 18371 10421 18380 10455
rect 18328 10412 18380 10421
rect 19432 10412 19484 10464
rect 22928 10412 22980 10464
rect 23204 10412 23256 10464
rect 26056 10455 26108 10464
rect 26056 10421 26065 10455
rect 26065 10421 26099 10455
rect 26099 10421 26108 10455
rect 26056 10412 26108 10421
rect 30932 10455 30984 10464
rect 30932 10421 30941 10455
rect 30941 10421 30975 10455
rect 30975 10421 30984 10455
rect 30932 10412 30984 10421
rect 31484 10455 31536 10464
rect 31484 10421 31493 10455
rect 31493 10421 31527 10455
rect 31527 10421 31536 10455
rect 31484 10412 31536 10421
rect 31852 10455 31904 10464
rect 31852 10421 31861 10455
rect 31861 10421 31895 10455
rect 31895 10421 31904 10455
rect 31852 10412 31904 10421
rect 33508 10455 33560 10464
rect 33508 10421 33517 10455
rect 33517 10421 33551 10455
rect 33551 10421 33560 10455
rect 33508 10412 33560 10421
rect 34704 10412 34756 10464
rect 36176 10480 36228 10532
rect 37832 10412 37884 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 10324 10208 10376 10260
rect 10600 10140 10652 10192
rect 11244 10140 11296 10192
rect 12440 10208 12492 10260
rect 14280 10251 14332 10260
rect 14280 10217 14289 10251
rect 14289 10217 14323 10251
rect 14323 10217 14332 10251
rect 14280 10208 14332 10217
rect 19340 10251 19392 10260
rect 19340 10217 19349 10251
rect 19349 10217 19383 10251
rect 19383 10217 19392 10251
rect 19340 10208 19392 10217
rect 22284 10208 22336 10260
rect 22560 10208 22612 10260
rect 23572 10208 23624 10260
rect 26608 10208 26660 10260
rect 10692 10115 10744 10124
rect 10692 10081 10701 10115
rect 10701 10081 10735 10115
rect 10735 10081 10744 10115
rect 10692 10072 10744 10081
rect 11888 10115 11940 10124
rect 11888 10081 11897 10115
rect 11897 10081 11931 10115
rect 11931 10081 11940 10115
rect 11888 10072 11940 10081
rect 12164 10072 12216 10124
rect 14556 10140 14608 10192
rect 16120 10140 16172 10192
rect 17684 10140 17736 10192
rect 18328 10140 18380 10192
rect 13268 10115 13320 10124
rect 13268 10081 13277 10115
rect 13277 10081 13311 10115
rect 13311 10081 13320 10115
rect 13268 10072 13320 10081
rect 13498 10115 13550 10124
rect 13498 10081 13507 10115
rect 13507 10081 13541 10115
rect 13541 10081 13550 10115
rect 13498 10072 13550 10081
rect 17500 10072 17552 10124
rect 18236 10115 18288 10124
rect 18236 10081 18245 10115
rect 18245 10081 18279 10115
rect 18279 10081 18288 10115
rect 18236 10072 18288 10081
rect 19432 10115 19484 10124
rect 19432 10081 19441 10115
rect 19441 10081 19475 10115
rect 19475 10081 19484 10115
rect 19432 10072 19484 10081
rect 19616 10115 19668 10124
rect 19616 10081 19625 10115
rect 19625 10081 19659 10115
rect 19659 10081 19668 10115
rect 19616 10072 19668 10081
rect 21456 10072 21508 10124
rect 21824 10072 21876 10124
rect 23480 10140 23532 10192
rect 23204 10072 23256 10124
rect 24308 10115 24360 10124
rect 24308 10081 24317 10115
rect 24317 10081 24351 10115
rect 24351 10081 24360 10115
rect 24308 10072 24360 10081
rect 24860 10140 24912 10192
rect 27252 10183 27304 10192
rect 27252 10149 27261 10183
rect 27261 10149 27295 10183
rect 27295 10149 27304 10183
rect 27252 10140 27304 10149
rect 27344 10183 27396 10192
rect 27344 10149 27353 10183
rect 27353 10149 27387 10183
rect 27387 10149 27396 10183
rect 27896 10183 27948 10192
rect 27344 10140 27396 10149
rect 27896 10149 27905 10183
rect 27905 10149 27939 10183
rect 27939 10149 27948 10183
rect 27896 10140 27948 10149
rect 31852 10208 31904 10260
rect 32496 10183 32548 10192
rect 29184 10115 29236 10124
rect 15200 10004 15252 10056
rect 16028 10004 16080 10056
rect 22100 10047 22152 10056
rect 22100 10013 22109 10047
rect 22109 10013 22143 10047
rect 22143 10013 22152 10047
rect 22100 10004 22152 10013
rect 10508 9936 10560 9988
rect 10876 9868 10928 9920
rect 11888 9868 11940 9920
rect 12624 9868 12676 9920
rect 15568 9936 15620 9988
rect 20996 9936 21048 9988
rect 21732 9936 21784 9988
rect 22928 9936 22980 9988
rect 23388 9936 23440 9988
rect 25228 9936 25280 9988
rect 28724 9936 28776 9988
rect 29184 10081 29193 10115
rect 29193 10081 29227 10115
rect 29227 10081 29236 10115
rect 29184 10072 29236 10081
rect 32496 10149 32505 10183
rect 32505 10149 32539 10183
rect 32539 10149 32548 10183
rect 32496 10140 32548 10149
rect 34980 10208 35032 10260
rect 32772 10140 32824 10192
rect 33140 10183 33192 10192
rect 33140 10149 33149 10183
rect 33149 10149 33183 10183
rect 33183 10149 33192 10183
rect 33140 10140 33192 10149
rect 34244 10140 34296 10192
rect 34336 10183 34388 10192
rect 34336 10149 34345 10183
rect 34345 10149 34379 10183
rect 34379 10149 34388 10183
rect 35164 10183 35216 10192
rect 34336 10140 34388 10149
rect 35164 10149 35173 10183
rect 35173 10149 35207 10183
rect 35207 10149 35216 10183
rect 35164 10140 35216 10149
rect 36268 10183 36320 10192
rect 36268 10149 36277 10183
rect 36277 10149 36311 10183
rect 36311 10149 36320 10183
rect 36268 10140 36320 10149
rect 30932 10072 30984 10124
rect 37832 10115 37884 10124
rect 37832 10081 37841 10115
rect 37841 10081 37875 10115
rect 37875 10081 37884 10115
rect 37832 10072 37884 10081
rect 31208 10004 31260 10056
rect 34244 10047 34296 10056
rect 34244 10013 34253 10047
rect 34253 10013 34287 10047
rect 34287 10013 34296 10047
rect 34244 10004 34296 10013
rect 36176 10047 36228 10056
rect 36176 10013 36185 10047
rect 36185 10013 36219 10047
rect 36219 10013 36228 10047
rect 36176 10004 36228 10013
rect 36820 10047 36872 10056
rect 36820 10013 36829 10047
rect 36829 10013 36863 10047
rect 36863 10013 36872 10047
rect 36820 10004 36872 10013
rect 14188 9868 14240 9920
rect 15660 9868 15712 9920
rect 21088 9868 21140 9920
rect 21916 9911 21968 9920
rect 21916 9877 21925 9911
rect 21925 9877 21959 9911
rect 21959 9877 21968 9911
rect 21916 9868 21968 9877
rect 26608 9868 26660 9920
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 8392 9664 8444 9716
rect 10692 9664 10744 9716
rect 13636 9639 13688 9648
rect 13636 9605 13645 9639
rect 13645 9605 13679 9639
rect 13679 9605 13688 9639
rect 13636 9596 13688 9605
rect 9220 9435 9272 9444
rect 9220 9401 9229 9435
rect 9229 9401 9263 9435
rect 9263 9401 9272 9435
rect 9220 9392 9272 9401
rect 9772 9435 9824 9444
rect 9772 9401 9781 9435
rect 9781 9401 9815 9435
rect 9815 9401 9824 9435
rect 9772 9392 9824 9401
rect 15200 9664 15252 9716
rect 15660 9596 15712 9648
rect 17684 9664 17736 9716
rect 18052 9664 18104 9716
rect 20904 9707 20956 9716
rect 20904 9673 20913 9707
rect 20913 9673 20947 9707
rect 20947 9673 20956 9707
rect 20904 9664 20956 9673
rect 21732 9664 21784 9716
rect 22560 9707 22612 9716
rect 22560 9673 22569 9707
rect 22569 9673 22603 9707
rect 22603 9673 22612 9707
rect 22560 9664 22612 9673
rect 24308 9664 24360 9716
rect 27344 9664 27396 9716
rect 28724 9707 28776 9716
rect 28724 9673 28733 9707
rect 28733 9673 28767 9707
rect 28767 9673 28776 9707
rect 28724 9664 28776 9673
rect 15936 9639 15988 9648
rect 15936 9605 15945 9639
rect 15945 9605 15979 9639
rect 15979 9605 15988 9639
rect 15936 9596 15988 9605
rect 16120 9639 16172 9648
rect 16120 9605 16129 9639
rect 16129 9605 16163 9639
rect 16163 9605 16172 9639
rect 16120 9596 16172 9605
rect 14096 9503 14148 9512
rect 9956 9392 10008 9444
rect 10876 9392 10928 9444
rect 11336 9435 11388 9444
rect 11336 9401 11345 9435
rect 11345 9401 11379 9435
rect 11379 9401 11388 9435
rect 11336 9392 11388 9401
rect 13360 9435 13412 9444
rect 13360 9401 13369 9435
rect 13369 9401 13403 9435
rect 13403 9401 13412 9435
rect 13360 9392 13412 9401
rect 12072 9324 12124 9376
rect 13268 9367 13320 9376
rect 13268 9333 13277 9367
rect 13277 9333 13311 9367
rect 13311 9333 13320 9367
rect 14096 9469 14105 9503
rect 14105 9469 14139 9503
rect 14139 9469 14148 9503
rect 14096 9460 14148 9469
rect 16028 9571 16080 9580
rect 16028 9537 16037 9571
rect 16037 9537 16071 9571
rect 16071 9537 16080 9571
rect 16028 9528 16080 9537
rect 16672 9460 16724 9512
rect 18880 9528 18932 9580
rect 18236 9503 18288 9512
rect 18236 9469 18245 9503
rect 18245 9469 18279 9503
rect 18279 9469 18288 9503
rect 20260 9528 20312 9580
rect 21916 9528 21968 9580
rect 23388 9528 23440 9580
rect 18236 9460 18288 9469
rect 19984 9460 20036 9512
rect 20904 9460 20956 9512
rect 13268 9324 13320 9333
rect 14096 9324 14148 9376
rect 15108 9367 15160 9376
rect 15108 9333 15117 9367
rect 15117 9333 15151 9367
rect 15151 9333 15160 9367
rect 15108 9324 15160 9333
rect 15476 9367 15528 9376
rect 15476 9333 15485 9367
rect 15485 9333 15519 9367
rect 15519 9333 15528 9367
rect 15476 9324 15528 9333
rect 15936 9324 15988 9376
rect 18236 9324 18288 9376
rect 19616 9392 19668 9444
rect 23112 9460 23164 9512
rect 25964 9503 26016 9512
rect 25964 9469 25973 9503
rect 25973 9469 26007 9503
rect 26007 9469 26016 9503
rect 25964 9460 26016 9469
rect 26608 9503 26660 9512
rect 26608 9469 26617 9503
rect 26617 9469 26651 9503
rect 26651 9469 26660 9503
rect 26608 9460 26660 9469
rect 22100 9392 22152 9444
rect 24860 9435 24912 9444
rect 20996 9324 21048 9376
rect 21732 9367 21784 9376
rect 21732 9333 21741 9367
rect 21741 9333 21775 9367
rect 21775 9333 21784 9367
rect 21732 9324 21784 9333
rect 21824 9324 21876 9376
rect 23480 9367 23532 9376
rect 23480 9333 23489 9367
rect 23489 9333 23523 9367
rect 23523 9333 23532 9367
rect 23480 9324 23532 9333
rect 24860 9401 24869 9435
rect 24869 9401 24903 9435
rect 24903 9401 24912 9435
rect 24860 9392 24912 9401
rect 26884 9435 26936 9444
rect 26884 9401 26893 9435
rect 26893 9401 26927 9435
rect 26927 9401 26936 9435
rect 26884 9392 26936 9401
rect 29644 9503 29696 9512
rect 29644 9469 29653 9503
rect 29653 9469 29687 9503
rect 29687 9469 29696 9503
rect 29644 9460 29696 9469
rect 30288 9664 30340 9716
rect 30932 9707 30984 9716
rect 30932 9673 30941 9707
rect 30941 9673 30975 9707
rect 30975 9673 30984 9707
rect 30932 9664 30984 9673
rect 31208 9707 31260 9716
rect 31208 9673 31217 9707
rect 31217 9673 31251 9707
rect 31251 9673 31260 9707
rect 31208 9664 31260 9673
rect 33508 9664 33560 9716
rect 34336 9707 34388 9716
rect 34336 9673 34345 9707
rect 34345 9673 34379 9707
rect 34379 9673 34388 9707
rect 34336 9664 34388 9673
rect 32496 9596 32548 9648
rect 31484 9528 31536 9580
rect 33784 9503 33836 9512
rect 33784 9469 33828 9503
rect 33828 9469 33836 9503
rect 33784 9460 33836 9469
rect 32128 9392 32180 9444
rect 24400 9324 24452 9376
rect 25872 9324 25924 9376
rect 27620 9367 27672 9376
rect 27620 9333 27629 9367
rect 27629 9333 27663 9367
rect 27663 9333 27672 9367
rect 27620 9324 27672 9333
rect 27988 9324 28040 9376
rect 30564 9367 30616 9376
rect 30564 9333 30573 9367
rect 30573 9333 30607 9367
rect 30607 9333 30616 9367
rect 30564 9324 30616 9333
rect 32772 9392 32824 9444
rect 32956 9435 33008 9444
rect 32956 9401 32965 9435
rect 32965 9401 32999 9435
rect 32999 9401 33008 9435
rect 32956 9392 33008 9401
rect 36176 9664 36228 9716
rect 37832 9664 37884 9716
rect 35256 9528 35308 9580
rect 36268 9528 36320 9580
rect 38844 9503 38896 9512
rect 38844 9469 38853 9503
rect 38853 9469 38887 9503
rect 38887 9469 38896 9503
rect 38844 9460 38896 9469
rect 34704 9392 34756 9444
rect 35072 9435 35124 9444
rect 35072 9401 35081 9435
rect 35081 9401 35115 9435
rect 35115 9401 35124 9435
rect 35072 9392 35124 9401
rect 35164 9392 35216 9444
rect 37832 9392 37884 9444
rect 37924 9324 37976 9376
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 9956 9163 10008 9172
rect 9956 9129 9965 9163
rect 9965 9129 9999 9163
rect 9999 9129 10008 9163
rect 9956 9120 10008 9129
rect 10876 9120 10928 9172
rect 11244 9163 11296 9172
rect 11244 9129 11253 9163
rect 11253 9129 11287 9163
rect 11287 9129 11296 9163
rect 11244 9120 11296 9129
rect 18880 9163 18932 9172
rect 18880 9129 18889 9163
rect 18889 9129 18923 9163
rect 18923 9129 18932 9163
rect 18880 9120 18932 9129
rect 20260 9163 20312 9172
rect 20260 9129 20269 9163
rect 20269 9129 20303 9163
rect 20303 9129 20312 9163
rect 20260 9120 20312 9129
rect 21456 9163 21508 9172
rect 21456 9129 21465 9163
rect 21465 9129 21499 9163
rect 21499 9129 21508 9163
rect 21456 9120 21508 9129
rect 21824 9163 21876 9172
rect 21824 9129 21833 9163
rect 21833 9129 21867 9163
rect 21867 9129 21876 9163
rect 21824 9120 21876 9129
rect 22836 9163 22888 9172
rect 22836 9129 22845 9163
rect 22845 9129 22879 9163
rect 22879 9129 22888 9163
rect 22836 9120 22888 9129
rect 27160 9163 27212 9172
rect 27160 9129 27169 9163
rect 27169 9129 27203 9163
rect 27203 9129 27212 9163
rect 27160 9120 27212 9129
rect 27252 9120 27304 9172
rect 33784 9163 33836 9172
rect 33784 9129 33793 9163
rect 33793 9129 33827 9163
rect 33827 9129 33836 9163
rect 33784 9120 33836 9129
rect 9864 9052 9916 9104
rect 14004 9095 14056 9104
rect 14004 9061 14013 9095
rect 14013 9061 14047 9095
rect 14047 9061 14056 9095
rect 14004 9052 14056 9061
rect 17868 9052 17920 9104
rect 19340 9052 19392 9104
rect 19984 9095 20036 9104
rect 19984 9061 19993 9095
rect 19993 9061 20027 9095
rect 20027 9061 20036 9095
rect 19984 9052 20036 9061
rect 8760 8984 8812 9036
rect 11888 9027 11940 9036
rect 11888 8993 11897 9027
rect 11897 8993 11931 9027
rect 11931 8993 11940 9027
rect 11888 8984 11940 8993
rect 12072 9027 12124 9036
rect 12072 8993 12081 9027
rect 12081 8993 12115 9027
rect 12115 8993 12124 9027
rect 13268 9027 13320 9036
rect 12072 8984 12124 8993
rect 13268 8993 13277 9027
rect 13277 8993 13311 9027
rect 13311 8993 13320 9027
rect 13268 8984 13320 8993
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 13360 8959 13412 8968
rect 8576 8848 8628 8900
rect 13360 8925 13369 8959
rect 13369 8925 13403 8959
rect 13403 8925 13412 8959
rect 13360 8916 13412 8925
rect 10416 8780 10468 8832
rect 12624 8780 12676 8832
rect 13176 8823 13228 8832
rect 13176 8789 13185 8823
rect 13185 8789 13219 8823
rect 13219 8789 13228 8823
rect 13636 8984 13688 9036
rect 13728 8984 13780 9036
rect 15660 9027 15712 9036
rect 15660 8993 15669 9027
rect 15669 8993 15703 9027
rect 15703 8993 15712 9027
rect 15660 8984 15712 8993
rect 15844 8984 15896 9036
rect 18236 9027 18288 9036
rect 18236 8993 18245 9027
rect 18245 8993 18279 9027
rect 18279 8993 18288 9027
rect 18236 8984 18288 8993
rect 19156 8984 19208 9036
rect 19892 8984 19944 9036
rect 22284 9095 22336 9104
rect 22284 9061 22287 9095
rect 22287 9061 22321 9095
rect 22321 9061 22336 9095
rect 22284 9052 22336 9061
rect 22560 9052 22612 9104
rect 24308 9095 24360 9104
rect 24308 9061 24317 9095
rect 24317 9061 24351 9095
rect 24351 9061 24360 9095
rect 24308 9052 24360 9061
rect 29644 9095 29696 9104
rect 29644 9061 29653 9095
rect 29653 9061 29687 9095
rect 29687 9061 29696 9095
rect 29644 9052 29696 9061
rect 32588 9052 32640 9104
rect 32956 9052 33008 9104
rect 34244 9120 34296 9172
rect 34612 9120 34664 9172
rect 26884 8984 26936 9036
rect 26976 8984 27028 9036
rect 28632 9027 28684 9036
rect 28632 8993 28641 9027
rect 28641 8993 28675 9027
rect 28675 8993 28684 9027
rect 28632 8984 28684 8993
rect 29000 8984 29052 9036
rect 30656 9027 30708 9036
rect 14188 8916 14240 8968
rect 16580 8916 16632 8968
rect 21548 8916 21600 8968
rect 22560 8916 22612 8968
rect 24216 8959 24268 8968
rect 24216 8925 24225 8959
rect 24225 8925 24259 8959
rect 24259 8925 24268 8959
rect 24216 8916 24268 8925
rect 24952 8916 25004 8968
rect 28724 8916 28776 8968
rect 29920 8916 29972 8968
rect 30656 8993 30665 9027
rect 30665 8993 30699 9027
rect 30699 8993 30708 9027
rect 30656 8984 30708 8993
rect 30932 8959 30984 8968
rect 30932 8925 30941 8959
rect 30941 8925 30975 8959
rect 30975 8925 30984 8959
rect 30932 8916 30984 8925
rect 31760 8916 31812 8968
rect 35072 9052 35124 9104
rect 37924 9095 37976 9104
rect 37924 9061 37933 9095
rect 37933 9061 37967 9095
rect 37967 9061 37976 9095
rect 37924 9052 37976 9061
rect 35164 8984 35216 9036
rect 34060 8959 34112 8968
rect 34060 8925 34069 8959
rect 34069 8925 34103 8959
rect 34103 8925 34112 8959
rect 34060 8916 34112 8925
rect 13176 8780 13228 8789
rect 14280 8780 14332 8832
rect 15568 8780 15620 8832
rect 35532 8848 35584 8900
rect 35808 8916 35860 8968
rect 37832 8959 37884 8968
rect 37832 8925 37841 8959
rect 37841 8925 37875 8959
rect 37875 8925 37884 8959
rect 37832 8916 37884 8925
rect 38108 8959 38160 8968
rect 38108 8925 38117 8959
rect 38117 8925 38151 8959
rect 38151 8925 38160 8959
rect 38108 8916 38160 8925
rect 16028 8780 16080 8832
rect 23940 8780 23992 8832
rect 26608 8780 26660 8832
rect 27896 8780 27948 8832
rect 34796 8780 34848 8832
rect 36544 8823 36596 8832
rect 36544 8789 36553 8823
rect 36553 8789 36587 8823
rect 36587 8789 36596 8823
rect 36544 8780 36596 8789
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 8760 8576 8812 8628
rect 12072 8576 12124 8628
rect 13360 8576 13412 8628
rect 14280 8619 14332 8628
rect 14280 8585 14289 8619
rect 14289 8585 14323 8619
rect 14323 8585 14332 8619
rect 14280 8576 14332 8585
rect 17868 8619 17920 8628
rect 17868 8585 17877 8619
rect 17877 8585 17911 8619
rect 17911 8585 17920 8619
rect 17868 8576 17920 8585
rect 19156 8576 19208 8628
rect 20536 8576 20588 8628
rect 20904 8576 20956 8628
rect 22284 8619 22336 8628
rect 22284 8585 22293 8619
rect 22293 8585 22327 8619
rect 22327 8585 22336 8619
rect 22284 8576 22336 8585
rect 22560 8619 22612 8628
rect 22560 8585 22569 8619
rect 22569 8585 22603 8619
rect 22603 8585 22612 8619
rect 22560 8576 22612 8585
rect 24216 8576 24268 8628
rect 25872 8576 25924 8628
rect 27344 8576 27396 8628
rect 28632 8619 28684 8628
rect 28632 8585 28641 8619
rect 28641 8585 28675 8619
rect 28675 8585 28684 8619
rect 28632 8576 28684 8585
rect 29920 8619 29972 8628
rect 29920 8585 29929 8619
rect 29929 8585 29963 8619
rect 29963 8585 29972 8619
rect 29920 8576 29972 8585
rect 30288 8619 30340 8628
rect 30288 8585 30297 8619
rect 30297 8585 30331 8619
rect 30331 8585 30340 8619
rect 30288 8576 30340 8585
rect 31760 8619 31812 8628
rect 31760 8585 31769 8619
rect 31769 8585 31803 8619
rect 31803 8585 31812 8619
rect 31760 8576 31812 8585
rect 32588 8576 32640 8628
rect 34244 8619 34296 8628
rect 34244 8585 34253 8619
rect 34253 8585 34287 8619
rect 34287 8585 34296 8619
rect 34244 8576 34296 8585
rect 34704 8619 34756 8628
rect 34704 8585 34713 8619
rect 34713 8585 34747 8619
rect 34747 8585 34756 8619
rect 34704 8576 34756 8585
rect 36268 8619 36320 8628
rect 36268 8585 36277 8619
rect 36277 8585 36311 8619
rect 36311 8585 36320 8619
rect 36268 8576 36320 8585
rect 37832 8576 37884 8628
rect 15660 8508 15712 8560
rect 16212 8508 16264 8560
rect 13176 8440 13228 8492
rect 15108 8440 15160 8492
rect 15844 8440 15896 8492
rect 16672 8483 16724 8492
rect 10508 8415 10560 8424
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 13544 8372 13596 8424
rect 14096 8372 14148 8424
rect 16672 8449 16681 8483
rect 16681 8449 16715 8483
rect 16715 8449 16724 8483
rect 16672 8440 16724 8449
rect 24308 8508 24360 8560
rect 27160 8508 27212 8560
rect 35808 8508 35860 8560
rect 21364 8440 21416 8492
rect 18788 8415 18840 8424
rect 10416 8304 10468 8356
rect 11888 8304 11940 8356
rect 9864 8279 9916 8288
rect 9864 8245 9873 8279
rect 9873 8245 9907 8279
rect 9907 8245 9916 8279
rect 9864 8236 9916 8245
rect 10048 8236 10100 8288
rect 13268 8236 13320 8288
rect 13636 8236 13688 8288
rect 15476 8236 15528 8288
rect 18788 8381 18797 8415
rect 18797 8381 18831 8415
rect 18831 8381 18840 8415
rect 18788 8372 18840 8381
rect 18972 8415 19024 8424
rect 18972 8381 18981 8415
rect 18981 8381 19015 8415
rect 19015 8381 19024 8415
rect 18972 8372 19024 8381
rect 20444 8372 20496 8424
rect 21272 8372 21324 8424
rect 22100 8440 22152 8492
rect 23296 8440 23348 8492
rect 24032 8440 24084 8492
rect 28356 8483 28408 8492
rect 28356 8449 28365 8483
rect 28365 8449 28399 8483
rect 28399 8449 28408 8483
rect 28356 8440 28408 8449
rect 32128 8440 32180 8492
rect 33140 8440 33192 8492
rect 34980 8483 35032 8492
rect 34980 8449 34989 8483
rect 34989 8449 35023 8483
rect 35023 8449 35032 8483
rect 34980 8440 35032 8449
rect 35256 8483 35308 8492
rect 35256 8449 35265 8483
rect 35265 8449 35299 8483
rect 35299 8449 35308 8483
rect 36544 8483 36596 8492
rect 35256 8440 35308 8449
rect 36544 8449 36553 8483
rect 36553 8449 36587 8483
rect 36587 8449 36596 8483
rect 36544 8440 36596 8449
rect 37188 8483 37240 8492
rect 37188 8449 37197 8483
rect 37197 8449 37231 8483
rect 37231 8449 37240 8483
rect 37188 8440 37240 8449
rect 38108 8440 38160 8492
rect 23480 8372 23532 8424
rect 23940 8372 23992 8424
rect 18236 8304 18288 8356
rect 19892 8304 19944 8356
rect 24308 8347 24360 8356
rect 24308 8313 24317 8347
rect 24317 8313 24351 8347
rect 24351 8313 24360 8347
rect 24308 8304 24360 8313
rect 24860 8347 24912 8356
rect 24860 8313 24869 8347
rect 24869 8313 24903 8347
rect 24903 8313 24912 8347
rect 24860 8304 24912 8313
rect 16120 8236 16172 8288
rect 19064 8279 19116 8288
rect 19064 8245 19073 8279
rect 19073 8245 19107 8279
rect 19107 8245 19116 8279
rect 19064 8236 19116 8245
rect 25136 8236 25188 8288
rect 25688 8236 25740 8288
rect 25872 8347 25924 8356
rect 25872 8313 25881 8347
rect 25881 8313 25915 8347
rect 25915 8313 25924 8347
rect 25872 8304 25924 8313
rect 27252 8304 27304 8356
rect 27712 8347 27764 8356
rect 27712 8313 27721 8347
rect 27721 8313 27755 8347
rect 27755 8313 27764 8347
rect 27712 8304 27764 8313
rect 27344 8236 27396 8288
rect 38016 8415 38068 8424
rect 38016 8381 38025 8415
rect 38025 8381 38059 8415
rect 38059 8381 38068 8415
rect 38476 8415 38528 8424
rect 38016 8372 38068 8381
rect 38476 8381 38485 8415
rect 38485 8381 38519 8415
rect 38519 8381 38528 8415
rect 38476 8372 38528 8381
rect 30288 8304 30340 8356
rect 31668 8304 31720 8356
rect 34244 8304 34296 8356
rect 34704 8304 34756 8356
rect 36268 8304 36320 8356
rect 29000 8279 29052 8288
rect 29000 8245 29009 8279
rect 29009 8245 29043 8279
rect 29043 8245 29052 8279
rect 29000 8236 29052 8245
rect 29552 8279 29604 8288
rect 29552 8245 29561 8279
rect 29561 8245 29595 8279
rect 29595 8245 29604 8279
rect 29552 8236 29604 8245
rect 36360 8236 36412 8288
rect 37924 8236 37976 8288
rect 38200 8279 38252 8288
rect 38200 8245 38209 8279
rect 38209 8245 38243 8279
rect 38243 8245 38252 8279
rect 38200 8236 38252 8245
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 13544 8032 13596 8084
rect 10600 8007 10652 8016
rect 10600 7973 10609 8007
rect 10609 7973 10643 8007
rect 10643 7973 10652 8007
rect 10600 7964 10652 7973
rect 12164 8007 12216 8016
rect 12164 7973 12173 8007
rect 12173 7973 12207 8007
rect 12207 7973 12216 8007
rect 12164 7964 12216 7973
rect 13728 8032 13780 8084
rect 17500 8075 17552 8084
rect 17500 8041 17509 8075
rect 17509 8041 17543 8075
rect 17543 8041 17552 8075
rect 17500 8032 17552 8041
rect 18788 8075 18840 8084
rect 18788 8041 18797 8075
rect 18797 8041 18831 8075
rect 18831 8041 18840 8075
rect 24032 8075 24084 8084
rect 18788 8032 18840 8041
rect 24032 8041 24041 8075
rect 24041 8041 24075 8075
rect 24075 8041 24084 8075
rect 24032 8032 24084 8041
rect 17132 7964 17184 8016
rect 19432 8007 19484 8016
rect 19432 7973 19441 8007
rect 19441 7973 19475 8007
rect 19475 7973 19484 8007
rect 19432 7964 19484 7973
rect 21456 7964 21508 8016
rect 13728 7939 13780 7948
rect 13728 7905 13737 7939
rect 13737 7905 13771 7939
rect 13771 7905 13780 7939
rect 13728 7896 13780 7905
rect 15844 7939 15896 7948
rect 15844 7905 15853 7939
rect 15853 7905 15887 7939
rect 15887 7905 15896 7939
rect 15844 7896 15896 7905
rect 17408 7939 17460 7948
rect 17408 7905 17417 7939
rect 17417 7905 17451 7939
rect 17451 7905 17460 7939
rect 17408 7896 17460 7905
rect 17868 7896 17920 7948
rect 19064 7896 19116 7948
rect 19616 7939 19668 7948
rect 19616 7905 19625 7939
rect 19625 7905 19659 7939
rect 19659 7905 19668 7939
rect 19616 7896 19668 7905
rect 19892 7896 19944 7948
rect 21088 7939 21140 7948
rect 21088 7905 21097 7939
rect 21097 7905 21131 7939
rect 21131 7905 21140 7939
rect 21088 7896 21140 7905
rect 21364 7939 21416 7948
rect 21364 7905 21373 7939
rect 21373 7905 21407 7939
rect 21407 7905 21416 7939
rect 21364 7896 21416 7905
rect 11152 7828 11204 7880
rect 12072 7871 12124 7880
rect 12072 7837 12081 7871
rect 12081 7837 12115 7871
rect 12115 7837 12124 7871
rect 12072 7828 12124 7837
rect 16212 7871 16264 7880
rect 11336 7760 11388 7812
rect 16212 7837 16221 7871
rect 16221 7837 16255 7871
rect 16255 7837 16264 7871
rect 16212 7828 16264 7837
rect 21824 7828 21876 7880
rect 23020 7964 23072 8016
rect 26056 8032 26108 8084
rect 26884 8032 26936 8084
rect 27712 8075 27764 8084
rect 27712 8041 27721 8075
rect 27721 8041 27755 8075
rect 27755 8041 27764 8075
rect 27712 8032 27764 8041
rect 29552 8075 29604 8084
rect 29552 8041 29561 8075
rect 29561 8041 29595 8075
rect 29595 8041 29604 8075
rect 29552 8032 29604 8041
rect 31760 8032 31812 8084
rect 32220 8075 32272 8084
rect 32220 8041 32229 8075
rect 32229 8041 32263 8075
rect 32263 8041 32272 8075
rect 32220 8032 32272 8041
rect 34060 8075 34112 8084
rect 34060 8041 34069 8075
rect 34069 8041 34103 8075
rect 34103 8041 34112 8075
rect 34060 8032 34112 8041
rect 35532 8075 35584 8084
rect 35532 8041 35541 8075
rect 35541 8041 35575 8075
rect 35575 8041 35584 8075
rect 35532 8032 35584 8041
rect 36360 8032 36412 8084
rect 37188 8032 37240 8084
rect 24400 8007 24452 8016
rect 24400 7973 24409 8007
rect 24409 7973 24443 8007
rect 24443 7973 24452 8007
rect 24952 8007 25004 8016
rect 24400 7964 24452 7973
rect 24952 7973 24961 8007
rect 24961 7973 24995 8007
rect 24995 7973 25004 8007
rect 24952 7964 25004 7973
rect 25136 7964 25188 8016
rect 26424 7964 26476 8016
rect 27528 7964 27580 8016
rect 29000 7964 29052 8016
rect 22836 7828 22888 7880
rect 27896 7896 27948 7948
rect 28264 7896 28316 7948
rect 29460 7896 29512 7948
rect 33140 7964 33192 8016
rect 34244 7964 34296 8016
rect 35256 7964 35308 8016
rect 36268 8007 36320 8016
rect 36268 7973 36277 8007
rect 36277 7973 36311 8007
rect 36311 7973 36320 8007
rect 36268 7964 36320 7973
rect 36820 8007 36872 8016
rect 36820 7973 36829 8007
rect 36829 7973 36863 8007
rect 36863 7973 36872 8007
rect 36820 7964 36872 7973
rect 37924 8007 37976 8016
rect 37924 7973 37933 8007
rect 37933 7973 37967 8007
rect 37967 7973 37976 8007
rect 37924 7964 37976 7973
rect 30564 7896 30616 7948
rect 32128 7939 32180 7948
rect 32128 7905 32137 7939
rect 32137 7905 32171 7939
rect 32171 7905 32180 7939
rect 32128 7896 32180 7905
rect 23388 7871 23440 7880
rect 23388 7837 23397 7871
rect 23397 7837 23431 7871
rect 23431 7837 23440 7871
rect 23388 7828 23440 7837
rect 24308 7871 24360 7880
rect 24308 7837 24317 7871
rect 24317 7837 24351 7871
rect 24351 7837 24360 7871
rect 24308 7828 24360 7837
rect 26608 7871 26660 7880
rect 26608 7837 26617 7871
rect 26617 7837 26651 7871
rect 26651 7837 26660 7871
rect 26608 7828 26660 7837
rect 27252 7871 27304 7880
rect 27252 7837 27261 7871
rect 27261 7837 27295 7871
rect 27295 7837 27304 7871
rect 27252 7828 27304 7837
rect 15936 7760 15988 7812
rect 25044 7760 25096 7812
rect 30564 7760 30616 7812
rect 33140 7828 33192 7880
rect 34520 7828 34572 7880
rect 35808 7828 35860 7880
rect 36176 7871 36228 7880
rect 36176 7837 36185 7871
rect 36185 7837 36219 7871
rect 36219 7837 36228 7871
rect 36176 7828 36228 7837
rect 38476 7896 38528 7948
rect 39304 7939 39356 7948
rect 39304 7905 39348 7939
rect 39348 7905 39356 7939
rect 39304 7896 39356 7905
rect 37832 7871 37884 7880
rect 37832 7837 37841 7871
rect 37841 7837 37875 7871
rect 37875 7837 37884 7871
rect 37832 7828 37884 7837
rect 38108 7871 38160 7880
rect 38108 7837 38117 7871
rect 38117 7837 38151 7871
rect 38151 7837 38160 7871
rect 38108 7828 38160 7837
rect 10416 7692 10468 7744
rect 15568 7735 15620 7744
rect 15568 7701 15577 7735
rect 15577 7701 15611 7735
rect 15611 7701 15620 7735
rect 15568 7692 15620 7701
rect 16120 7735 16172 7744
rect 16120 7701 16129 7735
rect 16129 7701 16163 7735
rect 16163 7701 16172 7735
rect 16948 7735 17000 7744
rect 16120 7692 16172 7701
rect 16948 7701 16957 7735
rect 16957 7701 16991 7735
rect 16991 7701 17000 7735
rect 16948 7692 17000 7701
rect 23664 7735 23716 7744
rect 23664 7701 23673 7735
rect 23673 7701 23707 7735
rect 23707 7701 23716 7735
rect 23664 7692 23716 7701
rect 25688 7735 25740 7744
rect 25688 7701 25697 7735
rect 25697 7701 25731 7735
rect 25731 7701 25740 7735
rect 25688 7692 25740 7701
rect 38476 7692 38528 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 9864 7531 9916 7540
rect 9864 7497 9873 7531
rect 9873 7497 9907 7531
rect 9907 7497 9916 7531
rect 9864 7488 9916 7497
rect 10600 7488 10652 7540
rect 11152 7531 11204 7540
rect 11152 7497 11161 7531
rect 11161 7497 11195 7531
rect 11195 7497 11204 7531
rect 11152 7488 11204 7497
rect 14280 7488 14332 7540
rect 15476 7531 15528 7540
rect 15476 7497 15500 7531
rect 15500 7497 15528 7531
rect 8576 7327 8628 7336
rect 8576 7293 8585 7327
rect 8585 7293 8619 7327
rect 8619 7293 8628 7327
rect 8576 7284 8628 7293
rect 10232 7352 10284 7404
rect 12164 7420 12216 7472
rect 15476 7488 15528 7497
rect 15752 7531 15804 7540
rect 15752 7497 15761 7531
rect 15761 7497 15795 7531
rect 15795 7497 15804 7531
rect 15752 7488 15804 7497
rect 17960 7488 18012 7540
rect 21180 7488 21232 7540
rect 21364 7488 21416 7540
rect 22284 7488 22336 7540
rect 23020 7531 23072 7540
rect 23020 7497 23029 7531
rect 23029 7497 23063 7531
rect 23063 7497 23072 7531
rect 23020 7488 23072 7497
rect 14740 7420 14792 7472
rect 17408 7463 17460 7472
rect 17408 7429 17417 7463
rect 17417 7429 17451 7463
rect 17451 7429 17460 7463
rect 17408 7420 17460 7429
rect 17868 7463 17920 7472
rect 17868 7429 17877 7463
rect 17877 7429 17911 7463
rect 17911 7429 17920 7463
rect 17868 7420 17920 7429
rect 13728 7352 13780 7404
rect 19616 7420 19668 7472
rect 9956 7327 10008 7336
rect 9956 7293 9965 7327
rect 9965 7293 9999 7327
rect 9999 7293 10008 7327
rect 9956 7284 10008 7293
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 14096 7284 14148 7336
rect 15844 7284 15896 7336
rect 9864 7216 9916 7268
rect 10784 7216 10836 7268
rect 15752 7216 15804 7268
rect 16120 7216 16172 7268
rect 13268 7148 13320 7200
rect 16948 7284 17000 7336
rect 18972 7216 19024 7268
rect 24308 7488 24360 7540
rect 24400 7488 24452 7540
rect 26424 7488 26476 7540
rect 27160 7488 27212 7540
rect 27620 7488 27672 7540
rect 27896 7488 27948 7540
rect 29460 7531 29512 7540
rect 29460 7497 29469 7531
rect 29469 7497 29503 7531
rect 29503 7497 29512 7531
rect 29460 7488 29512 7497
rect 29736 7488 29788 7540
rect 32128 7488 32180 7540
rect 33140 7531 33192 7540
rect 33140 7497 33149 7531
rect 33149 7497 33183 7531
rect 33183 7497 33192 7531
rect 33140 7488 33192 7497
rect 33416 7488 33468 7540
rect 33600 7488 33652 7540
rect 34244 7531 34296 7540
rect 34244 7497 34253 7531
rect 34253 7497 34287 7531
rect 34287 7497 34296 7531
rect 34244 7488 34296 7497
rect 36268 7488 36320 7540
rect 37832 7488 37884 7540
rect 39304 7531 39356 7540
rect 39304 7497 39313 7531
rect 39313 7497 39347 7531
rect 39347 7497 39356 7531
rect 39304 7488 39356 7497
rect 23756 7420 23808 7472
rect 26608 7420 26660 7472
rect 28816 7420 28868 7472
rect 31668 7463 31720 7472
rect 21088 7352 21140 7404
rect 21640 7352 21692 7404
rect 21824 7395 21876 7404
rect 21824 7361 21833 7395
rect 21833 7361 21867 7395
rect 21867 7361 21876 7395
rect 21824 7352 21876 7361
rect 23664 7395 23716 7404
rect 23664 7361 23673 7395
rect 23673 7361 23707 7395
rect 23707 7361 23716 7395
rect 23664 7352 23716 7361
rect 20812 7327 20864 7336
rect 20812 7293 20821 7327
rect 20821 7293 20855 7327
rect 20855 7293 20864 7327
rect 20812 7284 20864 7293
rect 24492 7284 24544 7336
rect 26792 7327 26844 7336
rect 26792 7293 26801 7327
rect 26801 7293 26835 7327
rect 26835 7293 26844 7327
rect 26792 7284 26844 7293
rect 31668 7429 31677 7463
rect 31677 7429 31711 7463
rect 31711 7429 31720 7463
rect 31668 7420 31720 7429
rect 35808 7420 35860 7472
rect 37280 7420 37332 7472
rect 38108 7420 38160 7472
rect 36360 7352 36412 7404
rect 37924 7352 37976 7404
rect 30564 7327 30616 7336
rect 30564 7293 30573 7327
rect 30573 7293 30607 7327
rect 30607 7293 30616 7327
rect 30564 7284 30616 7293
rect 31852 7327 31904 7336
rect 31852 7293 31861 7327
rect 31861 7293 31895 7327
rect 31895 7293 31904 7327
rect 31852 7284 31904 7293
rect 33600 7327 33652 7336
rect 33600 7293 33609 7327
rect 33609 7293 33643 7327
rect 33643 7293 33652 7327
rect 33600 7284 33652 7293
rect 38200 7327 38252 7336
rect 38200 7293 38209 7327
rect 38209 7293 38243 7327
rect 38243 7293 38252 7327
rect 38200 7284 38252 7293
rect 19340 7148 19392 7200
rect 19984 7148 20036 7200
rect 21548 7148 21600 7200
rect 22284 7148 22336 7200
rect 23756 7216 23808 7268
rect 27160 7216 27212 7268
rect 30840 7259 30892 7268
rect 30840 7225 30849 7259
rect 30849 7225 30883 7259
rect 30883 7225 30892 7259
rect 30840 7216 30892 7225
rect 31668 7216 31720 7268
rect 32496 7216 32548 7268
rect 36360 7259 36412 7268
rect 36360 7225 36369 7259
rect 36369 7225 36403 7259
rect 36403 7225 36412 7259
rect 36360 7216 36412 7225
rect 26332 7148 26384 7200
rect 26700 7148 26752 7200
rect 29000 7191 29052 7200
rect 29000 7157 29009 7191
rect 29009 7157 29043 7191
rect 29043 7157 29052 7191
rect 29000 7148 29052 7157
rect 33784 7191 33836 7200
rect 33784 7157 33793 7191
rect 33793 7157 33827 7191
rect 33827 7157 33836 7191
rect 33784 7148 33836 7157
rect 34520 7191 34572 7200
rect 34520 7157 34529 7191
rect 34529 7157 34563 7191
rect 34563 7157 34572 7191
rect 34520 7148 34572 7157
rect 34612 7148 34664 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 9956 6944 10008 6996
rect 10600 6944 10652 6996
rect 12440 6944 12492 6996
rect 14372 6944 14424 6996
rect 15568 6944 15620 6996
rect 16212 6944 16264 6996
rect 19432 6987 19484 6996
rect 19432 6953 19441 6987
rect 19441 6953 19475 6987
rect 19475 6953 19484 6987
rect 19432 6944 19484 6953
rect 22836 6944 22888 6996
rect 23664 6944 23716 6996
rect 24308 6944 24360 6996
rect 25688 6944 25740 6996
rect 26792 6944 26844 6996
rect 27988 6944 28040 6996
rect 30288 6987 30340 6996
rect 30288 6953 30297 6987
rect 30297 6953 30331 6987
rect 30331 6953 30340 6987
rect 30288 6944 30340 6953
rect 31300 6987 31352 6996
rect 31300 6953 31309 6987
rect 31309 6953 31343 6987
rect 31343 6953 31352 6987
rect 31300 6944 31352 6953
rect 32220 6944 32272 6996
rect 32496 6987 32548 6996
rect 32496 6953 32505 6987
rect 32505 6953 32539 6987
rect 32539 6953 32548 6987
rect 32496 6944 32548 6953
rect 16488 6876 16540 6928
rect 17868 6876 17920 6928
rect 18512 6919 18564 6928
rect 18512 6885 18521 6919
rect 18521 6885 18555 6919
rect 18555 6885 18564 6919
rect 18512 6876 18564 6885
rect 22284 6876 22336 6928
rect 28908 6876 28960 6928
rect 34336 6876 34388 6928
rect 10232 6851 10284 6860
rect 10232 6817 10241 6851
rect 10241 6817 10275 6851
rect 10275 6817 10284 6851
rect 10232 6808 10284 6817
rect 10508 6851 10560 6860
rect 10508 6817 10517 6851
rect 10517 6817 10551 6851
rect 10551 6817 10560 6851
rect 10508 6808 10560 6817
rect 12716 6851 12768 6860
rect 12716 6817 12725 6851
rect 12725 6817 12759 6851
rect 12759 6817 12768 6851
rect 12716 6808 12768 6817
rect 12532 6740 12584 6792
rect 13636 6808 13688 6860
rect 16028 6740 16080 6792
rect 16580 6783 16632 6792
rect 16580 6749 16589 6783
rect 16589 6749 16623 6783
rect 16623 6749 16632 6783
rect 16580 6740 16632 6749
rect 20812 6808 20864 6860
rect 23480 6851 23532 6860
rect 23480 6817 23489 6851
rect 23489 6817 23523 6851
rect 23523 6817 23532 6851
rect 23940 6851 23992 6860
rect 23480 6808 23532 6817
rect 23940 6817 23949 6851
rect 23949 6817 23983 6851
rect 23983 6817 23992 6851
rect 23940 6808 23992 6817
rect 24492 6808 24544 6860
rect 25504 6808 25556 6860
rect 26516 6851 26568 6860
rect 26516 6817 26525 6851
rect 26525 6817 26559 6851
rect 26559 6817 26568 6851
rect 26516 6808 26568 6817
rect 26700 6808 26752 6860
rect 29460 6808 29512 6860
rect 30196 6851 30248 6860
rect 30196 6817 30205 6851
rect 30205 6817 30239 6851
rect 30239 6817 30248 6851
rect 30196 6808 30248 6817
rect 30564 6808 30616 6860
rect 30840 6808 30892 6860
rect 31944 6808 31996 6860
rect 36176 6944 36228 6996
rect 35808 6876 35860 6928
rect 36912 6876 36964 6928
rect 35900 6808 35952 6860
rect 38476 6808 38528 6860
rect 19064 6740 19116 6792
rect 28724 6783 28776 6792
rect 16948 6672 17000 6724
rect 11244 6604 11296 6656
rect 12072 6604 12124 6656
rect 21364 6604 21416 6656
rect 28724 6749 28733 6783
rect 28733 6749 28767 6783
rect 28767 6749 28776 6783
rect 28724 6740 28776 6749
rect 30012 6740 30064 6792
rect 36360 6740 36412 6792
rect 34060 6672 34112 6724
rect 29644 6647 29696 6656
rect 29644 6613 29653 6647
rect 29653 6613 29687 6647
rect 29687 6613 29696 6647
rect 29644 6604 29696 6613
rect 31852 6604 31904 6656
rect 32772 6604 32824 6656
rect 33324 6604 33376 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 10508 6400 10560 6452
rect 12716 6400 12768 6452
rect 14740 6443 14792 6452
rect 14740 6409 14749 6443
rect 14749 6409 14783 6443
rect 14783 6409 14792 6443
rect 14740 6400 14792 6409
rect 19064 6443 19116 6452
rect 19064 6409 19073 6443
rect 19073 6409 19107 6443
rect 19107 6409 19116 6443
rect 19064 6400 19116 6409
rect 22284 6400 22336 6452
rect 23480 6400 23532 6452
rect 25504 6443 25556 6452
rect 25504 6409 25513 6443
rect 25513 6409 25547 6443
rect 25547 6409 25556 6443
rect 25504 6400 25556 6409
rect 25964 6443 26016 6452
rect 25964 6409 25973 6443
rect 25973 6409 26007 6443
rect 26007 6409 26016 6443
rect 25964 6400 26016 6409
rect 27528 6443 27580 6452
rect 27528 6409 27537 6443
rect 27537 6409 27571 6443
rect 27571 6409 27580 6443
rect 27528 6400 27580 6409
rect 30196 6400 30248 6452
rect 30840 6443 30892 6452
rect 30840 6409 30849 6443
rect 30849 6409 30883 6443
rect 30883 6409 30892 6443
rect 30840 6400 30892 6409
rect 10232 6332 10284 6384
rect 15384 6332 15436 6384
rect 12808 6264 12860 6316
rect 10692 6128 10744 6180
rect 10876 6171 10928 6180
rect 10876 6137 10885 6171
rect 10885 6137 10919 6171
rect 10919 6137 10928 6171
rect 10876 6128 10928 6137
rect 11796 6103 11848 6112
rect 11796 6069 11805 6103
rect 11805 6069 11839 6103
rect 11839 6069 11848 6103
rect 11796 6060 11848 6069
rect 13636 6128 13688 6180
rect 15752 6196 15804 6248
rect 16856 6332 16908 6384
rect 16580 6264 16632 6316
rect 17868 6264 17920 6316
rect 20168 6239 20220 6248
rect 20168 6205 20177 6239
rect 20177 6205 20211 6239
rect 20211 6205 20220 6239
rect 20168 6196 20220 6205
rect 23572 6332 23624 6384
rect 21364 6307 21416 6316
rect 21364 6273 21373 6307
rect 21373 6273 21407 6307
rect 21407 6273 21416 6307
rect 21364 6264 21416 6273
rect 23940 6264 23992 6316
rect 20904 6196 20956 6248
rect 21180 6239 21232 6248
rect 21180 6205 21189 6239
rect 21189 6205 21223 6239
rect 21223 6205 21232 6239
rect 21180 6196 21232 6205
rect 21548 6196 21600 6248
rect 26516 6332 26568 6384
rect 27988 6264 28040 6316
rect 28356 6307 28408 6316
rect 28356 6273 28365 6307
rect 28365 6273 28399 6307
rect 28399 6273 28408 6307
rect 28356 6264 28408 6273
rect 29644 6264 29696 6316
rect 31300 6264 31352 6316
rect 24768 6196 24820 6248
rect 25044 6239 25096 6248
rect 25044 6205 25053 6239
rect 25053 6205 25087 6239
rect 25087 6205 25096 6239
rect 25044 6196 25096 6205
rect 25964 6196 26016 6248
rect 26516 6239 26568 6248
rect 26516 6205 26525 6239
rect 26525 6205 26559 6239
rect 26559 6205 26568 6239
rect 26516 6196 26568 6205
rect 26792 6239 26844 6248
rect 26792 6205 26801 6239
rect 26801 6205 26835 6239
rect 26835 6205 26844 6239
rect 26792 6196 26844 6205
rect 19892 6128 19944 6180
rect 20536 6128 20588 6180
rect 22192 6171 22244 6180
rect 22192 6137 22201 6171
rect 22201 6137 22235 6171
rect 22235 6137 22244 6171
rect 22192 6128 22244 6137
rect 26976 6128 27028 6180
rect 27528 6128 27580 6180
rect 29460 6171 29512 6180
rect 29460 6137 29469 6171
rect 29469 6137 29503 6171
rect 29503 6137 29512 6171
rect 30012 6171 30064 6180
rect 29460 6128 29512 6137
rect 30012 6137 30021 6171
rect 30021 6137 30055 6171
rect 30055 6137 30064 6171
rect 30012 6128 30064 6137
rect 31668 6400 31720 6452
rect 33784 6400 33836 6452
rect 35900 6443 35952 6452
rect 33324 6307 33376 6316
rect 33324 6273 33333 6307
rect 33333 6273 33367 6307
rect 33367 6273 33376 6307
rect 33324 6264 33376 6273
rect 35900 6409 35909 6443
rect 35909 6409 35943 6443
rect 35943 6409 35952 6443
rect 35900 6400 35952 6409
rect 36912 6443 36964 6452
rect 36912 6409 36921 6443
rect 36921 6409 36955 6443
rect 36955 6409 36964 6443
rect 36912 6400 36964 6409
rect 37280 6443 37332 6452
rect 37280 6409 37289 6443
rect 37289 6409 37323 6443
rect 37323 6409 37332 6443
rect 37280 6400 37332 6409
rect 38476 6400 38528 6452
rect 37280 6196 37332 6248
rect 38292 6239 38344 6248
rect 38292 6205 38301 6239
rect 38301 6205 38335 6239
rect 38335 6205 38344 6239
rect 38292 6196 38344 6205
rect 14372 6103 14424 6112
rect 14372 6069 14381 6103
rect 14381 6069 14415 6103
rect 14415 6069 14424 6103
rect 14372 6060 14424 6069
rect 16488 6060 16540 6112
rect 17868 6103 17920 6112
rect 17868 6069 17877 6103
rect 17877 6069 17911 6103
rect 17911 6069 17920 6103
rect 17868 6060 17920 6069
rect 18144 6103 18196 6112
rect 18144 6069 18153 6103
rect 18153 6069 18187 6103
rect 18187 6069 18196 6103
rect 18144 6060 18196 6069
rect 22468 6103 22520 6112
rect 22468 6069 22477 6103
rect 22477 6069 22511 6103
rect 22511 6069 22520 6103
rect 22468 6060 22520 6069
rect 28908 6060 28960 6112
rect 31852 6103 31904 6112
rect 31852 6069 31861 6103
rect 31861 6069 31895 6103
rect 31895 6069 31904 6103
rect 31852 6060 31904 6069
rect 33140 6103 33192 6112
rect 33140 6069 33149 6103
rect 33149 6069 33183 6103
rect 33183 6069 33192 6103
rect 34060 6128 34112 6180
rect 34336 6103 34388 6112
rect 33140 6060 33192 6069
rect 34336 6069 34345 6103
rect 34345 6069 34379 6103
rect 34379 6069 34388 6103
rect 34336 6060 34388 6069
rect 35256 6060 35308 6112
rect 37832 6060 37884 6112
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 10232 5899 10284 5908
rect 10232 5865 10241 5899
rect 10241 5865 10275 5899
rect 10275 5865 10284 5899
rect 10232 5856 10284 5865
rect 10784 5856 10836 5908
rect 12532 5899 12584 5908
rect 12532 5865 12541 5899
rect 12541 5865 12575 5899
rect 12575 5865 12584 5899
rect 12532 5856 12584 5865
rect 13084 5899 13136 5908
rect 13084 5865 13093 5899
rect 13093 5865 13127 5899
rect 13127 5865 13136 5899
rect 13084 5856 13136 5865
rect 12716 5720 12768 5772
rect 10876 5652 10928 5704
rect 11336 5652 11388 5704
rect 13176 5720 13228 5772
rect 15752 5720 15804 5772
rect 17408 5856 17460 5908
rect 18144 5899 18196 5908
rect 18144 5865 18153 5899
rect 18153 5865 18187 5899
rect 18187 5865 18196 5899
rect 18144 5856 18196 5865
rect 18512 5899 18564 5908
rect 18512 5865 18521 5899
rect 18521 5865 18555 5899
rect 18555 5865 18564 5899
rect 18512 5856 18564 5865
rect 20996 5899 21048 5908
rect 20996 5865 21005 5899
rect 21005 5865 21039 5899
rect 21039 5865 21048 5899
rect 20996 5856 21048 5865
rect 22192 5899 22244 5908
rect 22192 5865 22201 5899
rect 22201 5865 22235 5899
rect 22235 5865 22244 5899
rect 22192 5856 22244 5865
rect 23940 5856 23992 5908
rect 26700 5899 26752 5908
rect 26700 5865 26709 5899
rect 26709 5865 26743 5899
rect 26743 5865 26752 5899
rect 26700 5856 26752 5865
rect 28632 5856 28684 5908
rect 17316 5831 17368 5840
rect 17316 5797 17325 5831
rect 17325 5797 17359 5831
rect 17359 5797 17368 5831
rect 17316 5788 17368 5797
rect 18880 5831 18932 5840
rect 18880 5797 18889 5831
rect 18889 5797 18923 5831
rect 18923 5797 18932 5831
rect 18880 5788 18932 5797
rect 21180 5788 21232 5840
rect 16120 5763 16172 5772
rect 16120 5729 16129 5763
rect 16129 5729 16163 5763
rect 16163 5729 16172 5763
rect 16120 5720 16172 5729
rect 20904 5763 20956 5772
rect 20904 5729 20913 5763
rect 20913 5729 20947 5763
rect 20947 5729 20956 5763
rect 20904 5720 20956 5729
rect 21456 5763 21508 5772
rect 21456 5729 21465 5763
rect 21465 5729 21499 5763
rect 21499 5729 21508 5763
rect 21456 5720 21508 5729
rect 22836 5788 22888 5840
rect 23480 5788 23532 5840
rect 22928 5763 22980 5772
rect 22928 5729 22937 5763
rect 22937 5729 22971 5763
rect 22971 5729 22980 5763
rect 24768 5788 24820 5840
rect 25044 5788 25096 5840
rect 27160 5788 27212 5840
rect 27528 5788 27580 5840
rect 29828 5831 29880 5840
rect 29828 5797 29831 5831
rect 29831 5797 29865 5831
rect 29865 5797 29880 5831
rect 29828 5788 29880 5797
rect 22928 5720 22980 5729
rect 26976 5720 27028 5772
rect 30288 5720 30340 5772
rect 30932 5856 30984 5908
rect 31944 5899 31996 5908
rect 31944 5865 31953 5899
rect 31953 5865 31987 5899
rect 31987 5865 31996 5899
rect 31944 5856 31996 5865
rect 32036 5856 32088 5908
rect 33416 5856 33468 5908
rect 32128 5763 32180 5772
rect 32128 5729 32137 5763
rect 32137 5729 32171 5763
rect 32171 5729 32180 5763
rect 32128 5720 32180 5729
rect 33140 5788 33192 5840
rect 36084 5788 36136 5840
rect 36360 5831 36412 5840
rect 36360 5797 36369 5831
rect 36369 5797 36403 5831
rect 36403 5797 36412 5831
rect 36360 5788 36412 5797
rect 33416 5720 33468 5772
rect 34152 5720 34204 5772
rect 34612 5720 34664 5772
rect 37832 5720 37884 5772
rect 16212 5695 16264 5704
rect 16212 5661 16221 5695
rect 16221 5661 16255 5695
rect 16255 5661 16264 5695
rect 16212 5652 16264 5661
rect 16856 5652 16908 5704
rect 18788 5695 18840 5704
rect 16948 5584 17000 5636
rect 18788 5661 18797 5695
rect 18797 5661 18831 5695
rect 18831 5661 18840 5695
rect 18788 5652 18840 5661
rect 23112 5695 23164 5704
rect 23112 5661 23121 5695
rect 23121 5661 23155 5695
rect 23155 5661 23164 5695
rect 23112 5652 23164 5661
rect 24124 5652 24176 5704
rect 28724 5695 28776 5704
rect 28724 5661 28733 5695
rect 28733 5661 28767 5695
rect 28767 5661 28776 5695
rect 28724 5652 28776 5661
rect 30104 5652 30156 5704
rect 30196 5652 30248 5704
rect 35440 5652 35492 5704
rect 36912 5652 36964 5704
rect 30012 5584 30064 5636
rect 36176 5584 36228 5636
rect 11428 5559 11480 5568
rect 11428 5525 11437 5559
rect 11437 5525 11471 5559
rect 11471 5525 11480 5559
rect 11428 5516 11480 5525
rect 12808 5559 12860 5568
rect 12808 5525 12817 5559
rect 12817 5525 12851 5559
rect 12851 5525 12860 5559
rect 12808 5516 12860 5525
rect 24768 5516 24820 5568
rect 26516 5516 26568 5568
rect 27160 5516 27212 5568
rect 29368 5559 29420 5568
rect 29368 5525 29377 5559
rect 29377 5525 29411 5559
rect 29411 5525 29420 5559
rect 29368 5516 29420 5525
rect 29552 5516 29604 5568
rect 36544 5516 36596 5568
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 10784 5312 10836 5364
rect 11796 5312 11848 5364
rect 12716 5355 12768 5364
rect 12716 5321 12725 5355
rect 12725 5321 12759 5355
rect 12759 5321 12768 5355
rect 12716 5312 12768 5321
rect 15384 5355 15436 5364
rect 15384 5321 15393 5355
rect 15393 5321 15427 5355
rect 15427 5321 15436 5355
rect 15384 5312 15436 5321
rect 16856 5355 16908 5364
rect 16856 5321 16865 5355
rect 16865 5321 16899 5355
rect 16899 5321 16908 5355
rect 16856 5312 16908 5321
rect 17316 5312 17368 5364
rect 18880 5312 18932 5364
rect 20260 5312 20312 5364
rect 20904 5312 20956 5364
rect 22836 5355 22888 5364
rect 22836 5321 22845 5355
rect 22845 5321 22879 5355
rect 22879 5321 22888 5355
rect 22836 5312 22888 5321
rect 22928 5312 22980 5364
rect 23388 5312 23440 5364
rect 24124 5355 24176 5364
rect 24124 5321 24133 5355
rect 24133 5321 24167 5355
rect 24167 5321 24176 5355
rect 24124 5312 24176 5321
rect 26976 5312 27028 5364
rect 29828 5312 29880 5364
rect 30840 5355 30892 5364
rect 30840 5321 30849 5355
rect 30849 5321 30883 5355
rect 30883 5321 30892 5355
rect 30840 5312 30892 5321
rect 32128 5355 32180 5364
rect 32128 5321 32137 5355
rect 32137 5321 32171 5355
rect 32171 5321 32180 5355
rect 32128 5312 32180 5321
rect 34152 5355 34204 5364
rect 34152 5321 34161 5355
rect 34161 5321 34195 5355
rect 34195 5321 34204 5355
rect 34152 5312 34204 5321
rect 36912 5355 36964 5364
rect 36912 5321 36921 5355
rect 36921 5321 36955 5355
rect 36955 5321 36964 5355
rect 36912 5312 36964 5321
rect 37832 5312 37884 5364
rect 10600 5151 10652 5160
rect 10600 5117 10609 5151
rect 10609 5117 10643 5151
rect 10643 5117 10652 5151
rect 10600 5108 10652 5117
rect 10784 5040 10836 5092
rect 13084 5176 13136 5228
rect 16488 5176 16540 5228
rect 15384 5108 15436 5160
rect 16120 5151 16172 5160
rect 16120 5117 16129 5151
rect 16129 5117 16163 5151
rect 16163 5117 16172 5151
rect 16120 5108 16172 5117
rect 15016 5040 15068 5092
rect 18144 5176 18196 5228
rect 20260 5151 20312 5160
rect 20260 5117 20269 5151
rect 20269 5117 20303 5151
rect 20303 5117 20312 5151
rect 20260 5108 20312 5117
rect 20352 5108 20404 5160
rect 21456 5108 21508 5160
rect 21640 5108 21692 5160
rect 22560 5176 22612 5228
rect 26700 5244 26752 5296
rect 27528 5287 27580 5296
rect 27528 5253 27537 5287
rect 27537 5253 27571 5287
rect 27571 5253 27580 5287
rect 27528 5244 27580 5253
rect 22836 5108 22888 5160
rect 24584 5151 24636 5160
rect 24584 5117 24593 5151
rect 24593 5117 24627 5151
rect 24627 5117 24636 5151
rect 24584 5108 24636 5117
rect 29092 5176 29144 5228
rect 29828 5219 29880 5228
rect 29828 5185 29837 5219
rect 29837 5185 29871 5219
rect 29871 5185 29880 5219
rect 29828 5176 29880 5185
rect 30932 5219 30984 5228
rect 30932 5185 30941 5219
rect 30941 5185 30975 5219
rect 30975 5185 30984 5219
rect 30932 5176 30984 5185
rect 30380 5108 30432 5160
rect 33416 5108 33468 5160
rect 36544 5151 36596 5160
rect 36544 5117 36553 5151
rect 36553 5117 36587 5151
rect 36587 5117 36596 5151
rect 36544 5108 36596 5117
rect 37832 5108 37884 5160
rect 20720 5040 20772 5092
rect 21180 5040 21232 5092
rect 23664 5040 23716 5092
rect 24492 5083 24544 5092
rect 24492 5049 24501 5083
rect 24501 5049 24535 5083
rect 24535 5049 24544 5083
rect 24492 5040 24544 5049
rect 26700 5083 26752 5092
rect 26700 5049 26703 5083
rect 26703 5049 26737 5083
rect 26737 5049 26752 5083
rect 26700 5040 26752 5049
rect 28816 5040 28868 5092
rect 29368 5083 29420 5092
rect 29368 5049 29377 5083
rect 29377 5049 29411 5083
rect 29411 5049 29420 5083
rect 29368 5040 29420 5049
rect 9588 5015 9640 5024
rect 9588 4981 9597 5015
rect 9597 4981 9631 5015
rect 9631 4981 9640 5015
rect 9588 4972 9640 4981
rect 14096 5015 14148 5024
rect 14096 4981 14105 5015
rect 14105 4981 14139 5015
rect 14139 4981 14148 5015
rect 14096 4972 14148 4981
rect 15660 5015 15712 5024
rect 15660 4981 15669 5015
rect 15669 4981 15703 5015
rect 15703 4981 15712 5015
rect 15660 4972 15712 4981
rect 25504 5015 25556 5024
rect 25504 4981 25513 5015
rect 25513 4981 25547 5015
rect 25547 4981 25556 5015
rect 25504 4972 25556 4981
rect 26516 4972 26568 5024
rect 28448 4972 28500 5024
rect 28908 4972 28960 5024
rect 31024 5040 31076 5092
rect 36636 5083 36688 5092
rect 30840 4972 30892 5024
rect 36636 5049 36645 5083
rect 36645 5049 36679 5083
rect 36679 5049 36688 5083
rect 36636 5040 36688 5049
rect 32772 5015 32824 5024
rect 32772 4981 32781 5015
rect 32781 4981 32815 5015
rect 32815 4981 32824 5015
rect 32772 4972 32824 4981
rect 34244 4972 34296 5024
rect 36084 4972 36136 5024
rect 37648 5015 37700 5024
rect 37648 4981 37657 5015
rect 37657 4981 37691 5015
rect 37691 4981 37700 5015
rect 37648 4972 37700 4981
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 10600 4811 10652 4820
rect 10600 4777 10609 4811
rect 10609 4777 10643 4811
rect 10643 4777 10652 4811
rect 10600 4768 10652 4777
rect 11336 4811 11388 4820
rect 11336 4777 11345 4811
rect 11345 4777 11379 4811
rect 11379 4777 11388 4811
rect 11336 4768 11388 4777
rect 12808 4768 12860 4820
rect 15752 4768 15804 4820
rect 16120 4768 16172 4820
rect 12440 4743 12492 4752
rect 12440 4709 12449 4743
rect 12449 4709 12483 4743
rect 12483 4709 12492 4743
rect 12440 4700 12492 4709
rect 14096 4700 14148 4752
rect 15016 4700 15068 4752
rect 16488 4700 16540 4752
rect 17316 4768 17368 4820
rect 18788 4768 18840 4820
rect 20352 4811 20404 4820
rect 20352 4777 20361 4811
rect 20361 4777 20395 4811
rect 20395 4777 20404 4811
rect 20352 4768 20404 4777
rect 22560 4811 22612 4820
rect 22560 4777 22569 4811
rect 22569 4777 22603 4811
rect 22603 4777 22612 4811
rect 22560 4768 22612 4777
rect 24584 4768 24636 4820
rect 26792 4768 26844 4820
rect 30288 4811 30340 4820
rect 30288 4777 30297 4811
rect 30297 4777 30331 4811
rect 30331 4777 30340 4811
rect 30288 4768 30340 4777
rect 36544 4768 36596 4820
rect 17592 4700 17644 4752
rect 10508 4675 10560 4684
rect 10508 4641 10517 4675
rect 10517 4641 10551 4675
rect 10551 4641 10560 4675
rect 10508 4632 10560 4641
rect 10692 4632 10744 4684
rect 16028 4632 16080 4684
rect 17500 4632 17552 4684
rect 17868 4675 17920 4684
rect 17868 4641 17877 4675
rect 17877 4641 17911 4675
rect 17911 4641 17920 4675
rect 17868 4632 17920 4641
rect 22468 4700 22520 4752
rect 13176 4564 13228 4616
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 13636 4607 13688 4616
rect 13636 4573 13645 4607
rect 13645 4573 13679 4607
rect 13679 4573 13688 4607
rect 13636 4564 13688 4573
rect 18512 4607 18564 4616
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 19524 4632 19576 4684
rect 19984 4632 20036 4684
rect 21272 4632 21324 4684
rect 24492 4700 24544 4752
rect 25044 4743 25096 4752
rect 25044 4709 25053 4743
rect 25053 4709 25087 4743
rect 25087 4709 25096 4743
rect 25044 4700 25096 4709
rect 27068 4700 27120 4752
rect 29092 4700 29144 4752
rect 30840 4700 30892 4752
rect 32220 4700 32272 4752
rect 33140 4700 33192 4752
rect 34152 4743 34204 4752
rect 34152 4709 34161 4743
rect 34161 4709 34195 4743
rect 34195 4709 34204 4743
rect 34152 4700 34204 4709
rect 36084 4743 36136 4752
rect 36084 4709 36093 4743
rect 36093 4709 36127 4743
rect 36127 4709 36136 4743
rect 36084 4700 36136 4709
rect 23112 4675 23164 4684
rect 23112 4641 23121 4675
rect 23121 4641 23155 4675
rect 23155 4641 23164 4675
rect 23112 4632 23164 4641
rect 28172 4675 28224 4684
rect 28172 4641 28190 4675
rect 28190 4641 28224 4675
rect 28172 4632 28224 4641
rect 29552 4632 29604 4684
rect 30380 4632 30432 4684
rect 31852 4632 31904 4684
rect 35992 4632 36044 4684
rect 37648 4632 37700 4684
rect 20628 4564 20680 4616
rect 22192 4607 22244 4616
rect 22192 4573 22201 4607
rect 22201 4573 22235 4607
rect 22235 4573 22244 4607
rect 22192 4564 22244 4573
rect 25228 4564 25280 4616
rect 26608 4607 26660 4616
rect 26608 4573 26617 4607
rect 26617 4573 26651 4607
rect 26651 4573 26660 4607
rect 26608 4564 26660 4573
rect 27344 4564 27396 4616
rect 32036 4564 32088 4616
rect 33508 4564 33560 4616
rect 34060 4607 34112 4616
rect 34060 4573 34069 4607
rect 34069 4573 34103 4607
rect 34103 4573 34112 4607
rect 34060 4564 34112 4573
rect 34704 4564 34756 4616
rect 13728 4428 13780 4480
rect 15108 4471 15160 4480
rect 15108 4437 15117 4471
rect 15117 4437 15151 4471
rect 15151 4437 15160 4471
rect 15108 4428 15160 4437
rect 17776 4471 17828 4480
rect 17776 4437 17785 4471
rect 17785 4437 17819 4471
rect 17819 4437 17828 4471
rect 17776 4428 17828 4437
rect 25596 4496 25648 4548
rect 29644 4496 29696 4548
rect 33048 4539 33100 4548
rect 33048 4505 33057 4539
rect 33057 4505 33091 4539
rect 33091 4505 33100 4539
rect 33048 4496 33100 4505
rect 34612 4539 34664 4548
rect 34612 4505 34621 4539
rect 34621 4505 34655 4539
rect 34655 4505 34664 4539
rect 34612 4496 34664 4505
rect 22928 4471 22980 4480
rect 22928 4437 22937 4471
rect 22937 4437 22971 4471
rect 22971 4437 22980 4471
rect 22928 4428 22980 4437
rect 28632 4428 28684 4480
rect 30012 4471 30064 4480
rect 30012 4437 30021 4471
rect 30021 4437 30055 4471
rect 30055 4437 30064 4471
rect 30012 4428 30064 4437
rect 30932 4471 30984 4480
rect 30932 4437 30941 4471
rect 30941 4437 30975 4471
rect 30975 4437 30984 4471
rect 30932 4428 30984 4437
rect 32496 4428 32548 4480
rect 34796 4428 34848 4480
rect 35900 4428 35952 4480
rect 38108 4428 38160 4480
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 10692 4224 10744 4276
rect 12348 4224 12400 4276
rect 14372 4224 14424 4276
rect 15752 4224 15804 4276
rect 16488 4267 16540 4276
rect 16488 4233 16497 4267
rect 16497 4233 16531 4267
rect 16531 4233 16540 4267
rect 16488 4224 16540 4233
rect 16856 4224 16908 4276
rect 17592 4224 17644 4276
rect 17868 4267 17920 4276
rect 17868 4233 17877 4267
rect 17877 4233 17911 4267
rect 17911 4233 17920 4267
rect 17868 4224 17920 4233
rect 19524 4267 19576 4276
rect 19524 4233 19533 4267
rect 19533 4233 19567 4267
rect 19567 4233 19576 4267
rect 19524 4224 19576 4233
rect 20628 4224 20680 4276
rect 21272 4224 21324 4276
rect 22560 4224 22612 4276
rect 25412 4224 25464 4276
rect 30380 4267 30432 4276
rect 30380 4233 30389 4267
rect 30389 4233 30423 4267
rect 30423 4233 30432 4267
rect 30380 4224 30432 4233
rect 31024 4224 31076 4276
rect 33324 4224 33376 4276
rect 33508 4267 33560 4276
rect 33508 4233 33517 4267
rect 33517 4233 33551 4267
rect 33551 4233 33560 4267
rect 33508 4224 33560 4233
rect 34244 4224 34296 4276
rect 35992 4267 36044 4276
rect 35992 4233 36001 4267
rect 36001 4233 36035 4267
rect 36035 4233 36044 4267
rect 35992 4224 36044 4233
rect 36636 4224 36688 4276
rect 38200 4224 38252 4276
rect 10508 4156 10560 4208
rect 13636 4156 13688 4208
rect 26700 4199 26752 4208
rect 26700 4165 26709 4199
rect 26709 4165 26743 4199
rect 26743 4165 26752 4199
rect 26700 4156 26752 4165
rect 28172 4199 28224 4208
rect 28172 4165 28181 4199
rect 28181 4165 28215 4199
rect 28215 4165 28224 4199
rect 28172 4156 28224 4165
rect 29092 4199 29144 4208
rect 29092 4165 29101 4199
rect 29101 4165 29135 4199
rect 29135 4165 29144 4199
rect 29092 4156 29144 4165
rect 32220 4199 32272 4208
rect 32220 4165 32229 4199
rect 32229 4165 32263 4199
rect 32263 4165 32272 4199
rect 32220 4156 32272 4165
rect 33048 4199 33100 4208
rect 9588 4088 9640 4140
rect 12716 4088 12768 4140
rect 14188 4131 14240 4140
rect 14188 4097 14197 4131
rect 14197 4097 14231 4131
rect 14231 4097 14240 4131
rect 14188 4088 14240 4097
rect 18420 4131 18472 4140
rect 18420 4097 18429 4131
rect 18429 4097 18463 4131
rect 18463 4097 18472 4131
rect 18420 4088 18472 4097
rect 18788 4088 18840 4140
rect 20996 4088 21048 4140
rect 26792 4131 26844 4140
rect 26792 4097 26801 4131
rect 26801 4097 26835 4131
rect 26835 4097 26844 4131
rect 26792 4088 26844 4097
rect 29828 4088 29880 4140
rect 32496 4131 32548 4140
rect 32496 4097 32505 4131
rect 32505 4097 32539 4131
rect 32539 4097 32548 4131
rect 32496 4088 32548 4097
rect 33048 4165 33057 4199
rect 33057 4165 33091 4199
rect 33091 4165 33100 4199
rect 33048 4156 33100 4165
rect 36360 4156 36412 4208
rect 34796 4088 34848 4140
rect 35900 4088 35952 4140
rect 36268 4088 36320 4140
rect 36820 4131 36872 4140
rect 36820 4097 36829 4131
rect 36829 4097 36863 4131
rect 36863 4097 36872 4131
rect 36820 4088 36872 4097
rect 38108 4131 38160 4140
rect 38108 4097 38117 4131
rect 38117 4097 38151 4131
rect 38151 4097 38160 4131
rect 38108 4088 38160 4097
rect 12348 4020 12400 4072
rect 12624 4063 12676 4072
rect 12624 4029 12633 4063
rect 12633 4029 12667 4063
rect 12667 4029 12676 4063
rect 13268 4063 13320 4072
rect 12624 4020 12676 4029
rect 13268 4029 13277 4063
rect 13277 4029 13311 4063
rect 13311 4029 13320 4063
rect 13268 4020 13320 4029
rect 11336 3952 11388 4004
rect 13636 3927 13688 3936
rect 13636 3893 13645 3927
rect 13645 3893 13679 3927
rect 13679 3893 13688 3927
rect 15476 4020 15528 4072
rect 14556 3952 14608 4004
rect 16120 3927 16172 3936
rect 13636 3884 13688 3893
rect 16120 3893 16129 3927
rect 16129 3893 16163 3927
rect 16163 3893 16172 3927
rect 16120 3884 16172 3893
rect 16580 3884 16632 3936
rect 17776 3952 17828 4004
rect 18236 3995 18288 4004
rect 18236 3961 18245 3995
rect 18245 3961 18279 3995
rect 18279 3961 18288 3995
rect 18236 3952 18288 3961
rect 18880 3884 18932 3936
rect 19892 4020 19944 4072
rect 22928 4020 22980 4072
rect 23664 4063 23716 4072
rect 23664 4029 23673 4063
rect 23673 4029 23707 4063
rect 23707 4029 23716 4063
rect 23664 4020 23716 4029
rect 25504 4020 25556 4072
rect 19156 3952 19208 4004
rect 20536 3952 20588 4004
rect 20720 3995 20772 4004
rect 20720 3961 20729 3995
rect 20729 3961 20763 3995
rect 20763 3961 20772 3995
rect 20720 3952 20772 3961
rect 23848 3952 23900 4004
rect 24492 3952 24544 4004
rect 26700 3952 26752 4004
rect 27344 3952 27396 4004
rect 29460 3995 29512 4004
rect 21732 3927 21784 3936
rect 21732 3893 21741 3927
rect 21741 3893 21775 3927
rect 21775 3893 21784 3927
rect 21732 3884 21784 3893
rect 23296 3884 23348 3936
rect 24584 3927 24636 3936
rect 24584 3893 24593 3927
rect 24593 3893 24627 3927
rect 24627 3893 24636 3927
rect 24584 3884 24636 3893
rect 25044 3884 25096 3936
rect 25228 3927 25280 3936
rect 25228 3893 25237 3927
rect 25237 3893 25271 3927
rect 25271 3893 25280 3927
rect 25228 3884 25280 3893
rect 26056 3884 26108 3936
rect 27068 3884 27120 3936
rect 28264 3884 28316 3936
rect 29460 3961 29469 3995
rect 29469 3961 29503 3995
rect 29503 3961 29512 3995
rect 29460 3952 29512 3961
rect 30932 3995 30984 4004
rect 30932 3961 30941 3995
rect 30941 3961 30975 3995
rect 30975 3961 30984 3995
rect 30932 3952 30984 3961
rect 31024 3995 31076 4004
rect 31024 3961 31033 3995
rect 31033 3961 31067 3995
rect 31067 3961 31076 3995
rect 31024 3952 31076 3961
rect 32312 3952 32364 4004
rect 31944 3927 31996 3936
rect 31944 3893 31953 3927
rect 31953 3893 31987 3927
rect 31987 3893 31996 3927
rect 34336 3952 34388 4004
rect 35072 3995 35124 4004
rect 35072 3961 35081 3995
rect 35081 3961 35115 3995
rect 35115 3961 35124 3995
rect 35072 3952 35124 3961
rect 31944 3884 31996 3893
rect 33324 3884 33376 3936
rect 34152 3884 34204 3936
rect 36360 3927 36412 3936
rect 36360 3893 36369 3927
rect 36369 3893 36403 3927
rect 36403 3893 36412 3927
rect 38200 3995 38252 4004
rect 38200 3961 38209 3995
rect 38209 3961 38243 3995
rect 38243 3961 38252 3995
rect 38200 3952 38252 3961
rect 36360 3884 36412 3893
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 11244 3680 11296 3732
rect 11428 3723 11480 3732
rect 11428 3689 11437 3723
rect 11437 3689 11471 3723
rect 11471 3689 11480 3723
rect 11428 3680 11480 3689
rect 14556 3723 14608 3732
rect 14556 3689 14565 3723
rect 14565 3689 14599 3723
rect 14599 3689 14608 3723
rect 14556 3680 14608 3689
rect 16028 3723 16080 3732
rect 16028 3689 16037 3723
rect 16037 3689 16071 3723
rect 16071 3689 16080 3723
rect 16028 3680 16080 3689
rect 16488 3680 16540 3732
rect 18236 3680 18288 3732
rect 20996 3680 21048 3732
rect 23664 3680 23716 3732
rect 25504 3680 25556 3732
rect 26608 3680 26660 3732
rect 28632 3680 28684 3732
rect 18144 3655 18196 3664
rect 18144 3621 18153 3655
rect 18153 3621 18187 3655
rect 18187 3621 18196 3655
rect 18144 3612 18196 3621
rect 22652 3612 22704 3664
rect 23848 3655 23900 3664
rect 23848 3621 23857 3655
rect 23857 3621 23891 3655
rect 23891 3621 23900 3655
rect 23848 3612 23900 3621
rect 25044 3655 25096 3664
rect 25044 3621 25053 3655
rect 25053 3621 25087 3655
rect 25087 3621 25096 3655
rect 25044 3612 25096 3621
rect 27344 3612 27396 3664
rect 28172 3655 28224 3664
rect 28172 3621 28181 3655
rect 28181 3621 28215 3655
rect 28215 3621 28224 3655
rect 28172 3612 28224 3621
rect 28816 3612 28868 3664
rect 30012 3680 30064 3732
rect 32036 3680 32088 3732
rect 30564 3655 30616 3664
rect 30564 3621 30573 3655
rect 30573 3621 30607 3655
rect 30607 3621 30616 3655
rect 30564 3612 30616 3621
rect 30748 3612 30800 3664
rect 32220 3612 32272 3664
rect 32496 3680 32548 3732
rect 34704 3723 34756 3732
rect 34704 3689 34713 3723
rect 34713 3689 34747 3723
rect 34747 3689 34756 3723
rect 34704 3680 34756 3689
rect 36268 3680 36320 3732
rect 11520 3544 11572 3596
rect 13728 3587 13780 3596
rect 13728 3553 13737 3587
rect 13737 3553 13771 3587
rect 13771 3553 13780 3587
rect 13728 3544 13780 3553
rect 19156 3544 19208 3596
rect 19892 3544 19944 3596
rect 20904 3587 20956 3596
rect 20904 3553 20913 3587
rect 20913 3553 20947 3587
rect 20947 3553 20956 3587
rect 20904 3544 20956 3553
rect 21364 3587 21416 3596
rect 21364 3553 21373 3587
rect 21373 3553 21407 3587
rect 21407 3553 21416 3587
rect 21364 3544 21416 3553
rect 22192 3544 22244 3596
rect 26424 3587 26476 3596
rect 26424 3553 26433 3587
rect 26433 3553 26467 3587
rect 26467 3553 26476 3587
rect 26424 3544 26476 3553
rect 29460 3544 29512 3596
rect 33048 3612 33100 3664
rect 33508 3612 33560 3664
rect 33876 3655 33928 3664
rect 33876 3621 33885 3655
rect 33885 3621 33919 3655
rect 33919 3621 33928 3655
rect 33876 3612 33928 3621
rect 35072 3612 35124 3664
rect 35256 3612 35308 3664
rect 35440 3544 35492 3596
rect 37740 3587 37792 3596
rect 37740 3553 37749 3587
rect 37749 3553 37783 3587
rect 37783 3553 37792 3587
rect 37740 3544 37792 3553
rect 11888 3519 11940 3528
rect 11888 3485 11897 3519
rect 11897 3485 11931 3519
rect 11931 3485 11940 3519
rect 11888 3476 11940 3485
rect 12440 3476 12492 3528
rect 16212 3519 16264 3528
rect 16212 3485 16221 3519
rect 16221 3485 16255 3519
rect 16255 3485 16264 3519
rect 16212 3476 16264 3485
rect 16764 3476 16816 3528
rect 18236 3476 18288 3528
rect 13360 3408 13412 3460
rect 15568 3408 15620 3460
rect 18420 3476 18472 3528
rect 21456 3519 21508 3528
rect 21456 3485 21465 3519
rect 21465 3485 21499 3519
rect 21499 3485 21508 3519
rect 21456 3476 21508 3485
rect 26056 3476 26108 3528
rect 26976 3476 27028 3528
rect 29000 3476 29052 3528
rect 31208 3519 31260 3528
rect 31208 3485 31217 3519
rect 31217 3485 31251 3519
rect 31251 3485 31260 3519
rect 32220 3519 32272 3528
rect 31208 3476 31260 3485
rect 32220 3485 32229 3519
rect 32229 3485 32263 3519
rect 32263 3485 32272 3519
rect 32220 3476 32272 3485
rect 32312 3476 32364 3528
rect 21180 3408 21232 3460
rect 33508 3476 33560 3528
rect 33784 3519 33836 3528
rect 33784 3485 33793 3519
rect 33793 3485 33827 3519
rect 33827 3485 33836 3519
rect 33784 3476 33836 3485
rect 37188 3476 37240 3528
rect 34336 3451 34388 3460
rect 34336 3417 34345 3451
rect 34345 3417 34379 3451
rect 34379 3417 34388 3451
rect 34336 3408 34388 3417
rect 34612 3408 34664 3460
rect 1676 3340 1728 3392
rect 9956 3340 10008 3392
rect 11520 3340 11572 3392
rect 14188 3383 14240 3392
rect 14188 3349 14197 3383
rect 14197 3349 14231 3383
rect 14231 3349 14240 3383
rect 14188 3340 14240 3349
rect 14280 3340 14332 3392
rect 18880 3340 18932 3392
rect 18972 3340 19024 3392
rect 23480 3383 23532 3392
rect 23480 3349 23489 3383
rect 23489 3349 23523 3383
rect 23523 3349 23532 3383
rect 24768 3383 24820 3392
rect 23480 3340 23532 3349
rect 24768 3349 24777 3383
rect 24777 3349 24811 3383
rect 24811 3349 24820 3383
rect 24768 3340 24820 3349
rect 27712 3383 27764 3392
rect 27712 3349 27721 3383
rect 27721 3349 27755 3383
rect 27755 3349 27764 3383
rect 27712 3340 27764 3349
rect 36176 3340 36228 3392
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 8668 3179 8720 3188
rect 8668 3145 8677 3179
rect 8677 3145 8711 3179
rect 8711 3145 8720 3179
rect 8668 3136 8720 3145
rect 11520 3179 11572 3188
rect 11520 3145 11529 3179
rect 11529 3145 11563 3179
rect 11563 3145 11572 3179
rect 11520 3136 11572 3145
rect 13360 3136 13412 3188
rect 13728 3136 13780 3188
rect 15476 3136 15528 3188
rect 11888 3000 11940 3052
rect 13636 3043 13688 3052
rect 13636 3009 13645 3043
rect 13645 3009 13679 3043
rect 13679 3009 13688 3043
rect 13636 3000 13688 3009
rect 10876 2932 10928 2984
rect 12716 2932 12768 2984
rect 12900 2932 12952 2984
rect 14280 2932 14332 2984
rect 16580 3136 16632 3188
rect 16764 3179 16816 3188
rect 16764 3145 16773 3179
rect 16773 3145 16807 3179
rect 16807 3145 16816 3179
rect 16764 3136 16816 3145
rect 17776 3136 17828 3188
rect 18144 3136 18196 3188
rect 19892 3179 19944 3188
rect 19892 3145 19901 3179
rect 19901 3145 19935 3179
rect 19935 3145 19944 3179
rect 19892 3136 19944 3145
rect 20904 3136 20956 3188
rect 22192 3136 22244 3188
rect 23112 3136 23164 3188
rect 24032 3136 24084 3188
rect 26056 3179 26108 3188
rect 26056 3145 26065 3179
rect 26065 3145 26099 3179
rect 26099 3145 26108 3179
rect 26056 3136 26108 3145
rect 26516 3179 26568 3188
rect 26516 3145 26525 3179
rect 26525 3145 26559 3179
rect 26559 3145 26568 3179
rect 26516 3136 26568 3145
rect 26976 3136 27028 3188
rect 27160 3179 27212 3188
rect 27160 3145 27169 3179
rect 27169 3145 27203 3179
rect 27203 3145 27212 3179
rect 27160 3136 27212 3145
rect 29000 3179 29052 3188
rect 29000 3145 29009 3179
rect 29009 3145 29043 3179
rect 29043 3145 29052 3179
rect 29000 3136 29052 3145
rect 29920 3136 29972 3188
rect 30748 3136 30800 3188
rect 32036 3179 32088 3188
rect 32036 3145 32045 3179
rect 32045 3145 32079 3179
rect 32079 3145 32088 3179
rect 32036 3136 32088 3145
rect 32220 3136 32272 3188
rect 33876 3136 33928 3188
rect 37740 3136 37792 3188
rect 39488 3136 39540 3188
rect 16488 3111 16540 3120
rect 16488 3077 16497 3111
rect 16497 3077 16531 3111
rect 16531 3077 16540 3111
rect 16488 3068 16540 3077
rect 18420 3068 18472 3120
rect 18972 3043 19024 3052
rect 18972 3009 18981 3043
rect 18981 3009 19015 3043
rect 19015 3009 19024 3043
rect 18972 3000 19024 3009
rect 21364 3068 21416 3120
rect 22652 3111 22704 3120
rect 22652 3077 22661 3111
rect 22661 3077 22695 3111
rect 22695 3077 22704 3111
rect 22652 3068 22704 3077
rect 21180 3043 21232 3052
rect 21180 3009 21189 3043
rect 21189 3009 21223 3043
rect 21223 3009 21232 3043
rect 21180 3000 21232 3009
rect 25412 3043 25464 3052
rect 25412 3009 25421 3043
rect 25421 3009 25455 3043
rect 25455 3009 25464 3043
rect 25412 3000 25464 3009
rect 27712 3043 27764 3052
rect 27712 3009 27721 3043
rect 27721 3009 27755 3043
rect 27755 3009 27764 3043
rect 27712 3000 27764 3009
rect 28816 3000 28868 3052
rect 31208 3043 31260 3052
rect 31208 3009 31217 3043
rect 31217 3009 31251 3043
rect 31251 3009 31260 3043
rect 31208 3000 31260 3009
rect 36360 3000 36412 3052
rect 37188 3043 37240 3052
rect 16120 2932 16172 2984
rect 23480 2932 23532 2984
rect 27160 2932 27212 2984
rect 30012 2932 30064 2984
rect 31760 2975 31812 2984
rect 31760 2941 31769 2975
rect 31769 2941 31803 2975
rect 31803 2941 31812 2975
rect 31760 2932 31812 2941
rect 9956 2864 10008 2916
rect 11980 2864 12032 2916
rect 9036 2839 9088 2848
rect 9036 2805 9045 2839
rect 9045 2805 9079 2839
rect 9079 2805 9088 2839
rect 11888 2839 11940 2848
rect 9036 2796 9088 2805
rect 11888 2805 11897 2839
rect 11897 2805 11931 2839
rect 11931 2805 11940 2839
rect 11888 2796 11940 2805
rect 14556 2864 14608 2916
rect 19432 2864 19484 2916
rect 20720 2864 20772 2916
rect 20996 2864 21048 2916
rect 22652 2864 22704 2916
rect 24768 2907 24820 2916
rect 24768 2873 24777 2907
rect 24777 2873 24811 2907
rect 24811 2873 24820 2907
rect 24768 2864 24820 2873
rect 18236 2839 18288 2848
rect 18236 2805 18245 2839
rect 18245 2805 18279 2839
rect 18279 2805 18288 2839
rect 18236 2796 18288 2805
rect 22100 2839 22152 2848
rect 22100 2805 22109 2839
rect 22109 2805 22143 2839
rect 22143 2805 22152 2839
rect 22100 2796 22152 2805
rect 27068 2864 27120 2916
rect 28356 2864 28408 2916
rect 30564 2907 30616 2916
rect 30564 2873 30573 2907
rect 30573 2873 30607 2907
rect 30607 2873 30616 2907
rect 30564 2864 30616 2873
rect 25044 2796 25096 2848
rect 28172 2796 28224 2848
rect 31944 2864 31996 2916
rect 36176 2975 36228 2984
rect 36176 2941 36185 2975
rect 36185 2941 36219 2975
rect 36219 2941 36228 2975
rect 36176 2932 36228 2941
rect 37188 3009 37197 3043
rect 37197 3009 37231 3043
rect 37231 3009 37240 3043
rect 37188 3000 37240 3009
rect 38108 3000 38160 3052
rect 33600 2839 33652 2848
rect 33600 2805 33609 2839
rect 33609 2805 33643 2839
rect 33643 2805 33652 2839
rect 33600 2796 33652 2805
rect 33692 2796 33744 2848
rect 35440 2839 35492 2848
rect 35440 2805 35449 2839
rect 35449 2805 35483 2839
rect 35483 2805 35492 2839
rect 35440 2796 35492 2805
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 9956 2592 10008 2644
rect 11980 2635 12032 2644
rect 11980 2601 11989 2635
rect 11989 2601 12023 2635
rect 12023 2601 12032 2635
rect 11980 2592 12032 2601
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12440 2592 12492 2601
rect 12900 2635 12952 2644
rect 12900 2601 12909 2635
rect 12909 2601 12943 2635
rect 12943 2601 12952 2635
rect 12900 2592 12952 2601
rect 14188 2592 14240 2644
rect 14280 2635 14332 2644
rect 14280 2601 14289 2635
rect 14289 2601 14323 2635
rect 14323 2601 14332 2635
rect 15660 2635 15712 2644
rect 14280 2592 14332 2601
rect 15660 2601 15669 2635
rect 15669 2601 15703 2635
rect 15703 2601 15712 2635
rect 15660 2592 15712 2601
rect 16488 2592 16540 2644
rect 16396 2524 16448 2576
rect 18144 2592 18196 2644
rect 19432 2635 19484 2644
rect 19432 2601 19441 2635
rect 19441 2601 19475 2635
rect 19475 2601 19484 2635
rect 19432 2592 19484 2601
rect 20996 2635 21048 2644
rect 20996 2601 21005 2635
rect 21005 2601 21039 2635
rect 21039 2601 21048 2635
rect 20996 2592 21048 2601
rect 22836 2592 22888 2644
rect 23296 2592 23348 2644
rect 27712 2592 27764 2644
rect 30564 2592 30616 2644
rect 31760 2592 31812 2644
rect 25136 2567 25188 2576
rect 25136 2533 25145 2567
rect 25145 2533 25179 2567
rect 25179 2533 25188 2567
rect 25136 2524 25188 2533
rect 27068 2567 27120 2576
rect 27068 2533 27077 2567
rect 27077 2533 27111 2567
rect 27111 2533 27120 2567
rect 27068 2524 27120 2533
rect 28264 2567 28316 2576
rect 28264 2533 28273 2567
rect 28273 2533 28307 2567
rect 28307 2533 28316 2567
rect 28264 2524 28316 2533
rect 28356 2524 28408 2576
rect 29920 2567 29972 2576
rect 29920 2533 29929 2567
rect 29929 2533 29963 2567
rect 29963 2533 29972 2567
rect 29920 2524 29972 2533
rect 30656 2524 30708 2576
rect 11060 2456 11112 2508
rect 11428 2456 11480 2508
rect 12716 2456 12768 2508
rect 13728 2456 13780 2508
rect 15568 2456 15620 2508
rect 15660 2456 15712 2508
rect 18512 2499 18564 2508
rect 18512 2465 18521 2499
rect 18521 2465 18555 2499
rect 18555 2465 18564 2499
rect 18512 2456 18564 2465
rect 21456 2456 21508 2508
rect 31576 2499 31628 2508
rect 31576 2465 31594 2499
rect 31594 2465 31628 2499
rect 31576 2456 31628 2465
rect 35256 2635 35308 2644
rect 35256 2601 35265 2635
rect 35265 2601 35299 2635
rect 35299 2601 35308 2635
rect 35256 2592 35308 2601
rect 35440 2592 35492 2644
rect 33784 2567 33836 2576
rect 33784 2533 33793 2567
rect 33793 2533 33827 2567
rect 33827 2533 33836 2567
rect 33784 2524 33836 2533
rect 36820 2524 36872 2576
rect 37740 2592 37792 2644
rect 16672 2388 16724 2440
rect 25136 2388 25188 2440
rect 25412 2431 25464 2440
rect 25412 2397 25421 2431
rect 25421 2397 25455 2431
rect 25455 2397 25464 2431
rect 25412 2388 25464 2397
rect 26240 2388 26292 2440
rect 18236 2320 18288 2372
rect 25596 2320 25648 2372
rect 30104 2431 30156 2440
rect 28448 2320 28500 2372
rect 30104 2397 30113 2431
rect 30113 2397 30147 2431
rect 30147 2397 30156 2431
rect 30104 2388 30156 2397
rect 33324 2431 33376 2440
rect 33324 2397 33333 2431
rect 33333 2397 33367 2431
rect 33367 2397 33376 2431
rect 33324 2388 33376 2397
rect 34336 2388 34388 2440
rect 5632 2252 5684 2304
rect 10876 2252 10928 2304
rect 11060 2295 11112 2304
rect 11060 2261 11069 2295
rect 11069 2261 11103 2295
rect 11103 2261 11112 2295
rect 11060 2252 11112 2261
rect 11428 2295 11480 2304
rect 11428 2261 11437 2295
rect 11437 2261 11471 2295
rect 11471 2261 11480 2295
rect 11428 2252 11480 2261
rect 11888 2252 11940 2304
rect 26240 2295 26292 2304
rect 26240 2261 26249 2295
rect 26249 2261 26283 2295
rect 26283 2261 26292 2295
rect 26240 2252 26292 2261
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
rect 33232 76 33284 128
rect 33876 76 33928 128
rect 40040 76 40092 128
rect 40960 76 41012 128
rect 41328 76 41380 128
rect 48136 76 48188 128
<< metal2 >>
rect 2778 49586 2834 50000
rect 8298 49586 8354 50000
rect 2778 49558 2912 49586
rect 2778 49520 2834 49558
rect 2884 42794 2912 49558
rect 8298 49558 8432 49586
rect 8298 49520 8354 49558
rect 4220 46812 4516 46832
rect 4276 46810 4300 46812
rect 4356 46810 4380 46812
rect 4436 46810 4460 46812
rect 4298 46758 4300 46810
rect 4362 46758 4374 46810
rect 4436 46758 4438 46810
rect 4276 46756 4300 46758
rect 4356 46756 4380 46758
rect 4436 46756 4460 46758
rect 4220 46736 4516 46756
rect 4220 45724 4516 45744
rect 4276 45722 4300 45724
rect 4356 45722 4380 45724
rect 4436 45722 4460 45724
rect 4298 45670 4300 45722
rect 4362 45670 4374 45722
rect 4436 45670 4438 45722
rect 4276 45668 4300 45670
rect 4356 45668 4380 45670
rect 4436 45668 4460 45670
rect 4220 45648 4516 45668
rect 4220 44636 4516 44656
rect 4276 44634 4300 44636
rect 4356 44634 4380 44636
rect 4436 44634 4460 44636
rect 4298 44582 4300 44634
rect 4362 44582 4374 44634
rect 4436 44582 4438 44634
rect 4276 44580 4300 44582
rect 4356 44580 4380 44582
rect 4436 44580 4460 44582
rect 4220 44560 4516 44580
rect 4220 43548 4516 43568
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4298 43494 4300 43546
rect 4362 43494 4374 43546
rect 4436 43494 4438 43546
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4220 43472 4516 43492
rect 8404 42794 8432 49558
rect 13818 49564 13874 50000
rect 13818 49520 13820 49564
rect 13872 49520 13874 49564
rect 16120 49564 16172 49570
rect 13820 49506 13872 49512
rect 19430 49564 19486 50000
rect 19430 49520 19432 49564
rect 16120 49506 16172 49512
rect 19484 49520 19486 49564
rect 20260 49564 20312 49570
rect 19432 49506 19484 49512
rect 20260 49506 20312 49512
rect 24216 49564 24268 49570
rect 24950 49564 25006 50000
rect 30470 49586 30526 50000
rect 36082 49586 36138 50000
rect 41602 49586 41658 50000
rect 47122 49586 47178 50000
rect 24950 49520 24952 49564
rect 24216 49506 24268 49512
rect 25004 49520 25006 49564
rect 30392 49558 30526 49586
rect 24952 49506 25004 49512
rect 13832 49475 13860 49506
rect 2792 42766 2912 42794
rect 8312 42766 8432 42794
rect 2792 23089 2820 42766
rect 4220 42460 4516 42480
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4298 42406 4300 42458
rect 4362 42406 4374 42458
rect 4436 42406 4438 42458
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4220 42384 4516 42404
rect 4220 41372 4516 41392
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4298 41318 4300 41370
rect 4362 41318 4374 41370
rect 4436 41318 4438 41370
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4220 41296 4516 41316
rect 4220 40284 4516 40304
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4298 40230 4300 40282
rect 4362 40230 4374 40282
rect 4436 40230 4438 40282
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4220 40208 4516 40228
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4220 39120 4516 39140
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 8312 30977 8340 42766
rect 14188 42152 14240 42158
rect 14188 42094 14240 42100
rect 11426 41576 11482 41585
rect 11426 41511 11482 41520
rect 11440 39953 11468 41511
rect 14200 40526 14228 42094
rect 14556 41132 14608 41138
rect 14556 41074 14608 41080
rect 14280 41064 14332 41070
rect 14280 41006 14332 41012
rect 14188 40520 14240 40526
rect 14188 40462 14240 40468
rect 14200 40186 14228 40462
rect 14188 40180 14240 40186
rect 14188 40122 14240 40128
rect 13360 40044 13412 40050
rect 13360 39986 13412 39992
rect 12992 39976 13044 39982
rect 11426 39944 11482 39953
rect 13372 39953 13400 39986
rect 12992 39918 13044 39924
rect 13358 39944 13414 39953
rect 11426 39879 11482 39888
rect 11888 39500 11940 39506
rect 11888 39442 11940 39448
rect 10508 38888 10560 38894
rect 10508 38830 10560 38836
rect 11336 38888 11388 38894
rect 11336 38830 11388 38836
rect 10232 37664 10284 37670
rect 10232 37606 10284 37612
rect 9680 35828 9732 35834
rect 9680 35770 9732 35776
rect 9692 31890 9720 35770
rect 10140 32904 10192 32910
rect 10140 32846 10192 32852
rect 10152 32570 10180 32846
rect 10140 32564 10192 32570
rect 10140 32506 10192 32512
rect 9680 31884 9732 31890
rect 9680 31826 9732 31832
rect 9954 31512 10010 31521
rect 9954 31447 10010 31456
rect 8298 30968 8354 30977
rect 8298 30903 8354 30912
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 9496 30048 9548 30054
rect 9496 29990 9548 29996
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 9508 29034 9536 29990
rect 9864 29640 9916 29646
rect 9864 29582 9916 29588
rect 9496 29028 9548 29034
rect 9496 28970 9548 28976
rect 9876 28762 9904 29582
rect 9864 28756 9916 28762
rect 9864 28698 9916 28704
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 9864 27872 9916 27878
rect 9864 27814 9916 27820
rect 9876 27577 9904 27814
rect 9862 27568 9918 27577
rect 9862 27503 9918 27512
rect 9968 27334 9996 31447
rect 10048 30048 10100 30054
rect 10048 29990 10100 29996
rect 9956 27328 10008 27334
rect 9956 27270 10008 27276
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 9864 26920 9916 26926
rect 9864 26862 9916 26868
rect 9876 26246 9904 26862
rect 9968 26790 9996 27270
rect 9956 26784 10008 26790
rect 9956 26726 10008 26732
rect 9864 26240 9916 26246
rect 9864 26182 9916 26188
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 9404 25696 9456 25702
rect 9404 25638 9456 25644
rect 9416 25265 9444 25638
rect 9402 25256 9458 25265
rect 9402 25191 9458 25200
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 2778 23080 2834 23089
rect 2778 23015 2834 23024
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 9416 18737 9444 25191
rect 9876 23474 9904 26182
rect 9968 23594 9996 26726
rect 10060 26450 10088 29990
rect 10140 29504 10192 29510
rect 10140 29446 10192 29452
rect 10048 26444 10100 26450
rect 10048 26386 10100 26392
rect 10048 25152 10100 25158
rect 10048 25094 10100 25100
rect 10060 24818 10088 25094
rect 10048 24812 10100 24818
rect 10048 24754 10100 24760
rect 9956 23588 10008 23594
rect 9956 23530 10008 23536
rect 9876 23446 10088 23474
rect 10060 22098 10088 23446
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 10152 20602 10180 29446
rect 10244 29306 10272 37606
rect 10416 36236 10468 36242
rect 10416 36178 10468 36184
rect 10428 35834 10456 36178
rect 10416 35828 10468 35834
rect 10416 35770 10468 35776
rect 10520 33658 10548 38830
rect 11348 38729 11376 38830
rect 11704 38820 11756 38826
rect 11704 38762 11756 38768
rect 11334 38720 11390 38729
rect 11334 38655 11390 38664
rect 11348 38554 11376 38655
rect 11716 38554 11744 38762
rect 11900 38758 11928 39442
rect 12624 38888 12676 38894
rect 12624 38830 12676 38836
rect 11888 38752 11940 38758
rect 11888 38694 11940 38700
rect 11336 38548 11388 38554
rect 11336 38490 11388 38496
rect 11704 38548 11756 38554
rect 11704 38490 11756 38496
rect 11348 37806 11376 38490
rect 11520 38344 11572 38350
rect 11520 38286 11572 38292
rect 11336 37800 11388 37806
rect 11336 37742 11388 37748
rect 11348 37466 11376 37742
rect 11532 37738 11560 38286
rect 11520 37732 11572 37738
rect 11520 37674 11572 37680
rect 11532 37466 11560 37674
rect 11716 37670 11744 38490
rect 11704 37664 11756 37670
rect 11704 37606 11756 37612
rect 10876 37460 10928 37466
rect 10876 37402 10928 37408
rect 11336 37460 11388 37466
rect 11336 37402 11388 37408
rect 11520 37460 11572 37466
rect 11520 37402 11572 37408
rect 10888 36242 10916 37402
rect 11900 37369 11928 38694
rect 12636 38554 12664 38830
rect 12624 38548 12676 38554
rect 12624 38490 12676 38496
rect 12624 38344 12676 38350
rect 12624 38286 12676 38292
rect 12348 38208 12400 38214
rect 12348 38150 12400 38156
rect 12532 38208 12584 38214
rect 12532 38150 12584 38156
rect 12360 37670 12388 38150
rect 12544 37874 12572 38150
rect 12636 37874 12664 38286
rect 12532 37868 12584 37874
rect 12532 37810 12584 37816
rect 12624 37868 12676 37874
rect 12624 37810 12676 37816
rect 11980 37664 12032 37670
rect 11980 37606 12032 37612
rect 12348 37664 12400 37670
rect 12348 37606 12400 37612
rect 11886 37360 11942 37369
rect 11886 37295 11942 37304
rect 11244 37256 11296 37262
rect 11244 37198 11296 37204
rect 11256 36689 11284 37198
rect 11242 36680 11298 36689
rect 11242 36615 11298 36624
rect 11256 36582 11284 36615
rect 11244 36576 11296 36582
rect 11244 36518 11296 36524
rect 11612 36576 11664 36582
rect 11612 36518 11664 36524
rect 10876 36236 10928 36242
rect 10876 36178 10928 36184
rect 10888 35834 10916 36178
rect 10968 36168 11020 36174
rect 10968 36110 11020 36116
rect 10876 35828 10928 35834
rect 10876 35770 10928 35776
rect 10888 35290 10916 35770
rect 10876 35284 10928 35290
rect 10876 35226 10928 35232
rect 10888 34542 10916 35226
rect 10980 35154 11008 36110
rect 10968 35148 11020 35154
rect 10968 35090 11020 35096
rect 10876 34536 10928 34542
rect 10876 34478 10928 34484
rect 10600 34400 10652 34406
rect 10600 34342 10652 34348
rect 10508 33652 10560 33658
rect 10508 33594 10560 33600
rect 10520 33454 10548 33594
rect 10508 33448 10560 33454
rect 10508 33390 10560 33396
rect 10520 33134 10548 33390
rect 10336 33106 10548 33134
rect 10232 29300 10284 29306
rect 10232 29242 10284 29248
rect 10244 29102 10272 29242
rect 10232 29096 10284 29102
rect 10232 29038 10284 29044
rect 10244 26042 10272 29038
rect 10336 28626 10364 33106
rect 10508 32360 10560 32366
rect 10508 32302 10560 32308
rect 10520 32026 10548 32302
rect 10508 32020 10560 32026
rect 10508 31962 10560 31968
rect 10416 31884 10468 31890
rect 10416 31826 10468 31832
rect 10428 31249 10456 31826
rect 10414 31240 10470 31249
rect 10414 31175 10470 31184
rect 10428 31142 10456 31175
rect 10416 31136 10468 31142
rect 10416 31078 10468 31084
rect 10506 31104 10562 31113
rect 10324 28620 10376 28626
rect 10324 28562 10376 28568
rect 10336 27606 10364 28562
rect 10324 27600 10376 27606
rect 10324 27542 10376 27548
rect 10428 26926 10456 31078
rect 10612 31090 10640 34342
rect 10888 34134 10916 34478
rect 10980 34202 11008 35090
rect 10968 34196 11020 34202
rect 10968 34138 11020 34144
rect 10876 34128 10928 34134
rect 10876 34070 10928 34076
rect 10968 33448 11020 33454
rect 10968 33390 11020 33396
rect 10980 32774 11008 33390
rect 10692 32768 10744 32774
rect 10692 32710 10744 32716
rect 10968 32768 11020 32774
rect 10968 32710 11020 32716
rect 10704 31890 10732 32710
rect 10692 31884 10744 31890
rect 10692 31826 10744 31832
rect 10704 31142 10732 31826
rect 10562 31062 10640 31090
rect 10692 31136 10744 31142
rect 10692 31078 10744 31084
rect 10506 31039 10562 31048
rect 10520 30802 10548 31039
rect 10704 30802 10732 31078
rect 10508 30796 10560 30802
rect 10508 30738 10560 30744
rect 10692 30796 10744 30802
rect 10692 30738 10744 30744
rect 10520 29850 10548 30738
rect 10508 29844 10560 29850
rect 10508 29786 10560 29792
rect 10704 29034 10732 30738
rect 10784 30728 10836 30734
rect 10784 30670 10836 30676
rect 10796 30258 10824 30670
rect 10784 30252 10836 30258
rect 10784 30194 10836 30200
rect 10796 29850 10824 30194
rect 11256 30190 11284 36518
rect 11336 35828 11388 35834
rect 11336 35770 11388 35776
rect 11348 35630 11376 35770
rect 11336 35624 11388 35630
rect 11336 35566 11388 35572
rect 11428 33380 11480 33386
rect 11428 33322 11480 33328
rect 11440 32910 11468 33322
rect 11428 32904 11480 32910
rect 11428 32846 11480 32852
rect 11440 32026 11468 32846
rect 11428 32020 11480 32026
rect 11428 31962 11480 31968
rect 11244 30184 11296 30190
rect 11244 30126 11296 30132
rect 11336 30116 11388 30122
rect 11336 30058 11388 30064
rect 10784 29844 10836 29850
rect 10784 29786 10836 29792
rect 11348 29782 11376 30058
rect 11336 29776 11388 29782
rect 11336 29718 11388 29724
rect 10876 29640 10928 29646
rect 10876 29582 10928 29588
rect 10888 29170 10916 29582
rect 11348 29238 11376 29718
rect 11336 29232 11388 29238
rect 11336 29174 11388 29180
rect 10876 29164 10928 29170
rect 10876 29106 10928 29112
rect 10692 29028 10744 29034
rect 10692 28970 10744 28976
rect 10600 28620 10652 28626
rect 10600 28562 10652 28568
rect 10508 28416 10560 28422
rect 10508 28358 10560 28364
rect 10520 28082 10548 28358
rect 10508 28076 10560 28082
rect 10508 28018 10560 28024
rect 10520 27062 10548 28018
rect 10612 27334 10640 28562
rect 10876 28552 10928 28558
rect 10876 28494 10928 28500
rect 10888 27538 10916 28494
rect 11348 28014 11376 29174
rect 11336 28008 11388 28014
rect 11336 27950 11388 27956
rect 11348 27606 11376 27950
rect 11428 27872 11480 27878
rect 11428 27814 11480 27820
rect 11440 27674 11468 27814
rect 11428 27668 11480 27674
rect 11428 27610 11480 27616
rect 11336 27600 11388 27606
rect 11336 27542 11388 27548
rect 10876 27532 10928 27538
rect 10876 27474 10928 27480
rect 10600 27328 10652 27334
rect 10600 27270 10652 27276
rect 10508 27056 10560 27062
rect 10508 26998 10560 27004
rect 10416 26920 10468 26926
rect 10416 26862 10468 26868
rect 10612 26858 10640 27270
rect 10888 27130 10916 27474
rect 10876 27124 10928 27130
rect 10876 27066 10928 27072
rect 11348 27062 11376 27542
rect 11152 27056 11204 27062
rect 11152 26998 11204 27004
rect 11336 27056 11388 27062
rect 11336 26998 11388 27004
rect 10600 26852 10652 26858
rect 10600 26794 10652 26800
rect 10508 26444 10560 26450
rect 10508 26386 10560 26392
rect 10232 26036 10284 26042
rect 10232 25978 10284 25984
rect 10244 25838 10272 25978
rect 10232 25832 10284 25838
rect 10232 25774 10284 25780
rect 10244 25362 10272 25774
rect 10520 25702 10548 26386
rect 10612 25838 10640 26794
rect 10600 25832 10652 25838
rect 10600 25774 10652 25780
rect 11058 25800 11114 25809
rect 10508 25696 10560 25702
rect 10508 25638 10560 25644
rect 10324 25424 10376 25430
rect 10324 25366 10376 25372
rect 10232 25356 10284 25362
rect 10232 25298 10284 25304
rect 10336 24954 10364 25366
rect 10324 24948 10376 24954
rect 10324 24890 10376 24896
rect 10612 24818 10640 25774
rect 10784 25764 10836 25770
rect 11058 25735 11114 25744
rect 10784 25706 10836 25712
rect 10796 25294 10824 25706
rect 11072 25702 11100 25735
rect 11060 25696 11112 25702
rect 11060 25638 11112 25644
rect 11164 25430 11192 26998
rect 11336 26512 11388 26518
rect 11336 26454 11388 26460
rect 11348 25974 11376 26454
rect 11336 25968 11388 25974
rect 11336 25910 11388 25916
rect 11348 25702 11376 25910
rect 11336 25696 11388 25702
rect 11336 25638 11388 25644
rect 11348 25498 11376 25638
rect 11336 25492 11388 25498
rect 11336 25434 11388 25440
rect 11152 25424 11204 25430
rect 11204 25384 11284 25412
rect 11152 25366 11204 25372
rect 10784 25288 10836 25294
rect 10784 25230 10836 25236
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 10416 24744 10468 24750
rect 10416 24686 10468 24692
rect 10428 24410 10456 24686
rect 10796 24410 10824 25230
rect 11256 24886 11284 25384
rect 11244 24880 11296 24886
rect 11244 24822 11296 24828
rect 11152 24676 11204 24682
rect 11152 24618 11204 24624
rect 10416 24404 10468 24410
rect 10784 24404 10836 24410
rect 10468 24364 10548 24392
rect 10416 24346 10468 24352
rect 10416 23656 10468 23662
rect 10416 23598 10468 23604
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 10152 19922 10180 20538
rect 10140 19916 10192 19922
rect 10140 19858 10192 19864
rect 10152 19514 10180 19858
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 9402 18728 9458 18737
rect 8392 18692 8444 18698
rect 9402 18663 9404 18672
rect 8392 18634 8444 18640
rect 9456 18663 9458 18672
rect 9404 18634 9456 18640
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 8404 9722 8432 18634
rect 8760 18624 8812 18630
rect 9416 18603 9444 18634
rect 8760 18566 8812 18572
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8680 11830 8708 12582
rect 8668 11824 8720 11830
rect 8668 11766 8720 11772
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8772 9042 8800 18566
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9232 17814 9260 18022
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9220 17808 9272 17814
rect 9220 17750 9272 17756
rect 9232 16998 9260 17750
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9692 17338 9720 17478
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 9232 13938 9260 16934
rect 9876 16658 9904 17818
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9324 16250 9352 16594
rect 10060 16522 10088 18158
rect 10336 17882 10364 18158
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10336 17746 10364 17818
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 10324 17060 10376 17066
rect 10324 17002 10376 17008
rect 10336 16794 10364 17002
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 10048 16516 10100 16522
rect 10048 16458 10100 16464
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 10336 15910 10364 16730
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9968 15162 9996 15506
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9692 13530 9720 14214
rect 9876 13734 9904 14894
rect 10336 14822 10364 15846
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10336 14618 10364 14758
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 10140 13796 10192 13802
rect 10140 13738 10192 13744
rect 9864 13728 9916 13734
rect 10152 13705 10180 13738
rect 9864 13670 9916 13676
rect 10138 13696 10194 13705
rect 10138 13631 10194 13640
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 10244 13394 10272 13806
rect 10336 13802 10364 14554
rect 10324 13796 10376 13802
rect 10324 13738 10376 13744
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10060 12850 10088 13330
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10152 12782 10180 13126
rect 10244 12782 10272 13330
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10232 12776 10284 12782
rect 10284 12736 10364 12764
rect 10232 12718 10284 12724
rect 9048 12442 9076 12718
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 9692 10985 9720 12718
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 9956 12368 10008 12374
rect 9956 12310 10008 12316
rect 9968 11354 9996 12310
rect 10244 12306 10272 12582
rect 10336 12374 10364 12736
rect 10324 12368 10376 12374
rect 10324 12310 10376 12316
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 10244 11898 10272 12242
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10336 11354 10364 11630
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10322 11248 10378 11257
rect 10322 11183 10378 11192
rect 10336 11150 10364 11183
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 9678 10976 9734 10985
rect 9678 10911 9734 10920
rect 9692 10674 9720 10911
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9232 9450 9260 10406
rect 9784 10033 9812 10474
rect 10336 10266 10364 11086
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10428 10033 10456 23598
rect 10520 22681 10548 24364
rect 10784 24346 10836 24352
rect 11164 24206 11192 24618
rect 11256 24342 11284 24822
rect 11244 24336 11296 24342
rect 11244 24278 11296 24284
rect 11152 24200 11204 24206
rect 11152 24142 11204 24148
rect 11164 23866 11192 24142
rect 11152 23860 11204 23866
rect 11152 23802 11204 23808
rect 11256 23798 11284 24278
rect 11244 23792 11296 23798
rect 11244 23734 11296 23740
rect 10506 22672 10562 22681
rect 10506 22607 10562 22616
rect 10508 22500 10560 22506
rect 10508 22442 10560 22448
rect 10520 19938 10548 22442
rect 11244 22432 11296 22438
rect 11244 22374 11296 22380
rect 11256 21962 11284 22374
rect 11244 21956 11296 21962
rect 11244 21898 11296 21904
rect 11256 21690 11284 21898
rect 11244 21684 11296 21690
rect 11244 21626 11296 21632
rect 11624 21078 11652 36518
rect 11900 34066 11928 37295
rect 11992 35562 12020 37606
rect 12544 37466 12572 37810
rect 12532 37460 12584 37466
rect 12532 37402 12584 37408
rect 12164 37392 12216 37398
rect 12084 37352 12164 37380
rect 12084 36038 12112 37352
rect 12164 37334 12216 37340
rect 12636 37262 12664 37810
rect 12164 37256 12216 37262
rect 12164 37198 12216 37204
rect 12624 37256 12676 37262
rect 12624 37198 12676 37204
rect 12176 36922 12204 37198
rect 12164 36916 12216 36922
rect 12164 36858 12216 36864
rect 12636 36174 12664 37198
rect 12716 36304 12768 36310
rect 12716 36246 12768 36252
rect 12164 36168 12216 36174
rect 12164 36110 12216 36116
rect 12624 36168 12676 36174
rect 12624 36110 12676 36116
rect 12072 36032 12124 36038
rect 12072 35974 12124 35980
rect 11980 35556 12032 35562
rect 11980 35498 12032 35504
rect 11992 35222 12020 35498
rect 11980 35216 12032 35222
rect 11980 35158 12032 35164
rect 11992 34746 12020 35158
rect 12084 35154 12112 35974
rect 12176 35290 12204 36110
rect 12532 35760 12584 35766
rect 12532 35702 12584 35708
rect 12164 35284 12216 35290
rect 12164 35226 12216 35232
rect 12072 35148 12124 35154
rect 12072 35090 12124 35096
rect 12440 35080 12492 35086
rect 12440 35022 12492 35028
rect 11980 34740 12032 34746
rect 11980 34682 12032 34688
rect 11888 34060 11940 34066
rect 11888 34002 11940 34008
rect 11900 33658 11928 34002
rect 11888 33652 11940 33658
rect 11888 33594 11940 33600
rect 11992 33046 12020 34682
rect 12452 34610 12480 35022
rect 12440 34604 12492 34610
rect 12440 34546 12492 34552
rect 12544 34490 12572 35702
rect 12728 35290 12756 36246
rect 12716 35284 12768 35290
rect 12716 35226 12768 35232
rect 12452 34462 12572 34490
rect 11980 33040 12032 33046
rect 11980 32982 12032 32988
rect 11992 32502 12020 32982
rect 11980 32496 12032 32502
rect 11980 32438 12032 32444
rect 12348 31884 12400 31890
rect 12348 31826 12400 31832
rect 12360 31142 12388 31826
rect 11704 31136 11756 31142
rect 11704 31078 11756 31084
rect 12348 31136 12400 31142
rect 12348 31078 12400 31084
rect 11716 27946 11744 31078
rect 11980 30864 12032 30870
rect 11980 30806 12032 30812
rect 11888 30728 11940 30734
rect 11888 30670 11940 30676
rect 11900 30326 11928 30670
rect 11888 30320 11940 30326
rect 11888 30262 11940 30268
rect 11992 30258 12020 30806
rect 11796 30252 11848 30258
rect 11796 30194 11848 30200
rect 11980 30252 12032 30258
rect 11980 30194 12032 30200
rect 11808 29850 11836 30194
rect 11796 29844 11848 29850
rect 11796 29786 11848 29792
rect 12452 29306 12480 34462
rect 12900 34400 12952 34406
rect 12900 34342 12952 34348
rect 12532 33856 12584 33862
rect 12532 33798 12584 33804
rect 12544 33522 12572 33798
rect 12532 33516 12584 33522
rect 12532 33458 12584 33464
rect 12716 33380 12768 33386
rect 12716 33322 12768 33328
rect 12532 32768 12584 32774
rect 12728 32756 12756 33322
rect 12912 33046 12940 34342
rect 12900 33040 12952 33046
rect 12900 32982 12952 32988
rect 12584 32728 12756 32756
rect 12532 32710 12584 32716
rect 12544 31958 12572 32710
rect 12624 32292 12676 32298
rect 12624 32234 12676 32240
rect 12636 32026 12664 32234
rect 12624 32020 12676 32026
rect 12624 31962 12676 31968
rect 12532 31952 12584 31958
rect 12532 31894 12584 31900
rect 13004 31890 13032 39918
rect 13358 39879 13414 39888
rect 13176 39840 13228 39846
rect 13176 39782 13228 39788
rect 13188 39574 13216 39782
rect 13176 39568 13228 39574
rect 13176 39510 13228 39516
rect 14004 39568 14056 39574
rect 14004 39510 14056 39516
rect 13188 39098 13216 39510
rect 13268 39296 13320 39302
rect 13268 39238 13320 39244
rect 13634 39264 13690 39273
rect 13176 39092 13228 39098
rect 13176 39034 13228 39040
rect 13280 38486 13308 39238
rect 13634 39199 13690 39208
rect 13452 38752 13504 38758
rect 13452 38694 13504 38700
rect 13464 38486 13492 38694
rect 13268 38480 13320 38486
rect 13268 38422 13320 38428
rect 13452 38480 13504 38486
rect 13452 38422 13504 38428
rect 13280 37942 13308 38422
rect 13464 38010 13492 38422
rect 13452 38004 13504 38010
rect 13452 37946 13504 37952
rect 13268 37936 13320 37942
rect 13268 37878 13320 37884
rect 13452 37324 13504 37330
rect 13452 37266 13504 37272
rect 13464 36922 13492 37266
rect 13452 36916 13504 36922
rect 13452 36858 13504 36864
rect 13268 36848 13320 36854
rect 13268 36790 13320 36796
rect 13280 36310 13308 36790
rect 13268 36304 13320 36310
rect 13268 36246 13320 36252
rect 13360 35556 13412 35562
rect 13360 35498 13412 35504
rect 13372 35222 13400 35498
rect 13360 35216 13412 35222
rect 13360 35158 13412 35164
rect 13372 34678 13400 35158
rect 13464 34746 13492 36858
rect 13452 34740 13504 34746
rect 13452 34682 13504 34688
rect 13360 34672 13412 34678
rect 13360 34614 13412 34620
rect 13084 34536 13136 34542
rect 13084 34478 13136 34484
rect 12992 31884 13044 31890
rect 12992 31826 13044 31832
rect 12992 31680 13044 31686
rect 12992 31622 13044 31628
rect 13004 31482 13032 31622
rect 13096 31521 13124 34478
rect 13176 33380 13228 33386
rect 13176 33322 13228 33328
rect 13188 32434 13216 33322
rect 13452 33040 13504 33046
rect 13452 32982 13504 32988
rect 13544 33040 13596 33046
rect 13544 32982 13596 32988
rect 13464 32570 13492 32982
rect 13452 32564 13504 32570
rect 13452 32506 13504 32512
rect 13556 32502 13584 32982
rect 13544 32496 13596 32502
rect 13544 32438 13596 32444
rect 13176 32428 13228 32434
rect 13176 32370 13228 32376
rect 13188 32026 13216 32370
rect 13556 32298 13584 32438
rect 13544 32292 13596 32298
rect 13544 32234 13596 32240
rect 13176 32020 13228 32026
rect 13176 31962 13228 31968
rect 13082 31512 13138 31521
rect 12992 31476 13044 31482
rect 13082 31447 13138 31456
rect 12992 31418 13044 31424
rect 13188 31346 13216 31962
rect 13452 31952 13504 31958
rect 13452 31894 13504 31900
rect 13464 31482 13492 31894
rect 13452 31476 13504 31482
rect 13452 31418 13504 31424
rect 13648 31414 13676 39199
rect 13728 38956 13780 38962
rect 13728 38898 13780 38904
rect 13740 38554 13768 38898
rect 13728 38548 13780 38554
rect 13728 38490 13780 38496
rect 13820 36780 13872 36786
rect 14016 36768 14044 39510
rect 14292 39273 14320 41006
rect 14372 40928 14424 40934
rect 14372 40870 14424 40876
rect 14278 39264 14334 39273
rect 14278 39199 14334 39208
rect 14384 38962 14412 40870
rect 14372 38956 14424 38962
rect 14372 38898 14424 38904
rect 14568 38729 14596 41074
rect 14648 40384 14700 40390
rect 14648 40326 14700 40332
rect 14660 40050 14688 40326
rect 16028 40112 16080 40118
rect 16028 40054 16080 40060
rect 14648 40044 14700 40050
rect 14648 39986 14700 39992
rect 14740 39908 14792 39914
rect 14740 39850 14792 39856
rect 15292 39908 15344 39914
rect 15292 39850 15344 39856
rect 14752 39642 14780 39850
rect 14740 39636 14792 39642
rect 14740 39578 14792 39584
rect 14752 39098 14780 39578
rect 15304 39438 15332 39850
rect 16040 39574 16068 40054
rect 16028 39568 16080 39574
rect 16028 39510 16080 39516
rect 15660 39500 15712 39506
rect 15660 39442 15712 39448
rect 15292 39432 15344 39438
rect 15292 39374 15344 39380
rect 15672 39098 15700 39442
rect 15936 39432 15988 39438
rect 15936 39374 15988 39380
rect 14740 39092 14792 39098
rect 14740 39034 14792 39040
rect 15660 39092 15712 39098
rect 15660 39034 15712 39040
rect 14752 38826 14780 39034
rect 15384 38888 15436 38894
rect 15384 38830 15436 38836
rect 14740 38820 14792 38826
rect 14740 38762 14792 38768
rect 14554 38720 14610 38729
rect 14554 38655 14610 38664
rect 14280 37392 14332 37398
rect 14280 37334 14332 37340
rect 13872 36740 14044 36768
rect 13820 36722 13872 36728
rect 13728 36644 13780 36650
rect 13728 36586 13780 36592
rect 13740 36378 13768 36586
rect 14016 36378 14044 36740
rect 13728 36372 13780 36378
rect 13728 36314 13780 36320
rect 14004 36372 14056 36378
rect 14004 36314 14056 36320
rect 13740 35834 13768 36314
rect 13728 35828 13780 35834
rect 13728 35770 13780 35776
rect 14016 35766 14044 36314
rect 14096 36236 14148 36242
rect 14096 36178 14148 36184
rect 14004 35760 14056 35766
rect 14004 35702 14056 35708
rect 14108 35698 14136 36178
rect 14096 35692 14148 35698
rect 14096 35634 14148 35640
rect 14108 34746 14136 35634
rect 14096 34740 14148 34746
rect 14096 34682 14148 34688
rect 14108 34542 14136 34682
rect 14096 34536 14148 34542
rect 14094 34504 14096 34513
rect 14148 34504 14150 34513
rect 14094 34439 14150 34448
rect 13912 34400 13964 34406
rect 13912 34342 13964 34348
rect 13728 34060 13780 34066
rect 13728 34002 13780 34008
rect 13740 33658 13768 34002
rect 13728 33652 13780 33658
rect 13728 33594 13780 33600
rect 13924 33522 13952 34342
rect 14096 34060 14148 34066
rect 14096 34002 14148 34008
rect 14108 33658 14136 34002
rect 14096 33652 14148 33658
rect 14096 33594 14148 33600
rect 13912 33516 13964 33522
rect 13912 33458 13964 33464
rect 13728 32904 13780 32910
rect 13728 32846 13780 32852
rect 13740 31754 13768 32846
rect 13820 31816 13872 31822
rect 13820 31758 13872 31764
rect 13728 31748 13780 31754
rect 13728 31690 13780 31696
rect 13636 31408 13688 31414
rect 13636 31350 13688 31356
rect 12532 31340 12584 31346
rect 12532 31282 12584 31288
rect 13176 31340 13228 31346
rect 13176 31282 13228 31288
rect 12544 30870 12572 31282
rect 12808 31204 12860 31210
rect 12808 31146 12860 31152
rect 12900 31204 12952 31210
rect 12900 31146 12952 31152
rect 12532 30864 12584 30870
rect 12532 30806 12584 30812
rect 12820 30598 12848 31146
rect 12808 30592 12860 30598
rect 12808 30534 12860 30540
rect 12820 30394 12848 30534
rect 12808 30388 12860 30394
rect 12808 30330 12860 30336
rect 12912 29714 12940 31146
rect 13084 31136 13136 31142
rect 13136 31096 13216 31124
rect 13084 31078 13136 31084
rect 12900 29708 12952 29714
rect 12900 29650 12952 29656
rect 12992 29640 13044 29646
rect 12992 29582 13044 29588
rect 12532 29504 12584 29510
rect 12532 29446 12584 29452
rect 12440 29300 12492 29306
rect 12440 29242 12492 29248
rect 12452 29102 12480 29242
rect 12544 29102 12572 29446
rect 13004 29170 13032 29582
rect 12992 29164 13044 29170
rect 12992 29106 13044 29112
rect 12440 29096 12492 29102
rect 12440 29038 12492 29044
rect 12532 29096 12584 29102
rect 12532 29038 12584 29044
rect 12164 28688 12216 28694
rect 12164 28630 12216 28636
rect 12072 28552 12124 28558
rect 12072 28494 12124 28500
rect 11796 28076 11848 28082
rect 11796 28018 11848 28024
rect 11704 27940 11756 27946
rect 11704 27882 11756 27888
rect 11808 27538 11836 28018
rect 11796 27532 11848 27538
rect 11796 27474 11848 27480
rect 12084 27334 12112 28494
rect 12176 28082 12204 28630
rect 12164 28076 12216 28082
rect 12164 28018 12216 28024
rect 12164 27396 12216 27402
rect 12164 27338 12216 27344
rect 12256 27396 12308 27402
rect 12256 27338 12308 27344
rect 12072 27328 12124 27334
rect 12072 27270 12124 27276
rect 12084 26518 12112 27270
rect 12176 27130 12204 27338
rect 12164 27124 12216 27130
rect 12164 27066 12216 27072
rect 12072 26512 12124 26518
rect 12072 26454 12124 26460
rect 11888 26376 11940 26382
rect 11888 26318 11940 26324
rect 11900 26042 11928 26318
rect 11888 26036 11940 26042
rect 11888 25978 11940 25984
rect 11886 25936 11942 25945
rect 11886 25871 11942 25880
rect 11900 25362 11928 25871
rect 11888 25356 11940 25362
rect 11888 25298 11940 25304
rect 11900 23186 11928 25298
rect 12072 25152 12124 25158
rect 12072 25094 12124 25100
rect 12084 24410 12112 25094
rect 12072 24404 12124 24410
rect 12072 24346 12124 24352
rect 12268 23866 12296 27338
rect 12452 24274 12480 29038
rect 12808 28552 12860 28558
rect 12808 28494 12860 28500
rect 12532 28212 12584 28218
rect 12532 28154 12584 28160
rect 12544 27946 12572 28154
rect 12532 27940 12584 27946
rect 12532 27882 12584 27888
rect 12544 24290 12572 27882
rect 12624 27668 12676 27674
rect 12624 27610 12676 27616
rect 12636 26858 12664 27610
rect 12716 27056 12768 27062
rect 12716 26998 12768 27004
rect 12624 26852 12676 26858
rect 12624 26794 12676 26800
rect 12624 24744 12676 24750
rect 12624 24686 12676 24692
rect 12636 24410 12664 24686
rect 12624 24404 12676 24410
rect 12624 24346 12676 24352
rect 12440 24268 12492 24274
rect 12544 24262 12664 24290
rect 12440 24210 12492 24216
rect 12348 24064 12400 24070
rect 12348 24006 12400 24012
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 12268 23662 12296 23802
rect 12360 23730 12388 24006
rect 12348 23724 12400 23730
rect 12348 23666 12400 23672
rect 12256 23656 12308 23662
rect 12256 23598 12308 23604
rect 12360 23186 12388 23666
rect 12636 23474 12664 24262
rect 12544 23446 12664 23474
rect 11888 23180 11940 23186
rect 11888 23122 11940 23128
rect 12348 23180 12400 23186
rect 12348 23122 12400 23128
rect 11900 22506 11928 23122
rect 11888 22500 11940 22506
rect 11888 22442 11940 22448
rect 11796 22092 11848 22098
rect 11796 22034 11848 22040
rect 11808 21350 11836 22034
rect 12360 21962 12388 23122
rect 12440 23112 12492 23118
rect 12440 23054 12492 23060
rect 12452 22642 12480 23054
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12452 22234 12480 22578
rect 12440 22228 12492 22234
rect 12440 22170 12492 22176
rect 12348 21956 12400 21962
rect 12348 21898 12400 21904
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11612 21072 11664 21078
rect 11612 21014 11664 21020
rect 10600 21004 10652 21010
rect 10600 20946 10652 20952
rect 10612 20058 10640 20946
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10692 20324 10744 20330
rect 10692 20266 10744 20272
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 10520 19910 10640 19938
rect 10508 18148 10560 18154
rect 10508 18090 10560 18096
rect 10520 17882 10548 18090
rect 10508 17876 10560 17882
rect 10508 17818 10560 17824
rect 10520 17202 10548 17818
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10508 12368 10560 12374
rect 10508 12310 10560 12316
rect 10520 11626 10548 12310
rect 10508 11620 10560 11626
rect 10508 11562 10560 11568
rect 10508 10532 10560 10538
rect 10508 10474 10560 10480
rect 9770 10024 9826 10033
rect 9770 9959 9826 9968
rect 10414 10024 10470 10033
rect 10520 9994 10548 10474
rect 10612 10198 10640 19910
rect 10704 19514 10732 20266
rect 10980 19990 11008 20742
rect 10968 19984 11020 19990
rect 10968 19926 11020 19932
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10704 19174 10732 19450
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10980 18970 11008 19926
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 10968 18964 11020 18970
rect 10968 18906 11020 18912
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 10888 18426 10916 18770
rect 11072 18698 11100 19314
rect 11256 18970 11284 19790
rect 11520 19780 11572 19786
rect 11520 19722 11572 19728
rect 11532 19378 11560 19722
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11532 18834 11560 19314
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11060 18692 11112 18698
rect 11060 18634 11112 18640
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 10888 16794 10916 18022
rect 11704 17808 11756 17814
rect 11704 17750 11756 17756
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 11072 16250 11100 16934
rect 11348 16454 11376 17614
rect 11716 16998 11744 17750
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11336 16448 11388 16454
rect 11336 16390 11388 16396
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11348 16182 11376 16390
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11336 16176 11388 16182
rect 11336 16118 11388 16124
rect 10876 15972 10928 15978
rect 10876 15914 10928 15920
rect 10888 15366 10916 15914
rect 11716 15638 11744 16186
rect 11152 15632 11204 15638
rect 11152 15574 11204 15580
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10888 14074 10916 15302
rect 11164 14822 11192 15574
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11532 15162 11560 15438
rect 11520 15156 11572 15162
rect 11520 15098 11572 15104
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10980 13870 11008 14214
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 11164 13734 11192 14350
rect 11152 13728 11204 13734
rect 10782 13696 10838 13705
rect 11152 13670 11204 13676
rect 10782 13631 10838 13640
rect 10796 10810 10824 13631
rect 11164 12918 11192 13670
rect 11520 13456 11572 13462
rect 11520 13398 11572 13404
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11348 12986 11376 13262
rect 11532 12986 11560 13398
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11152 12912 11204 12918
rect 11152 12854 11204 12860
rect 11808 11354 11836 21286
rect 12164 21072 12216 21078
rect 12164 21014 12216 21020
rect 12176 19514 12204 21014
rect 12544 21010 12572 23446
rect 12728 21690 12756 26998
rect 12820 26994 12848 28494
rect 13084 27872 13136 27878
rect 13084 27814 13136 27820
rect 13096 27334 13124 27814
rect 13084 27328 13136 27334
rect 13084 27270 13136 27276
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 12820 26450 12848 26930
rect 13096 26586 13124 27270
rect 13084 26580 13136 26586
rect 13084 26522 13136 26528
rect 13188 26450 13216 31096
rect 13740 30938 13768 31690
rect 13832 31482 13860 31758
rect 13820 31476 13872 31482
rect 13820 31418 13872 31424
rect 13728 30932 13780 30938
rect 13728 30874 13780 30880
rect 13636 30796 13688 30802
rect 13636 30738 13688 30744
rect 13360 30388 13412 30394
rect 13360 30330 13412 30336
rect 13372 30190 13400 30330
rect 13360 30184 13412 30190
rect 13360 30126 13412 30132
rect 13268 28076 13320 28082
rect 13268 28018 13320 28024
rect 13280 27946 13308 28018
rect 13268 27940 13320 27946
rect 13268 27882 13320 27888
rect 13280 26858 13308 27882
rect 13268 26852 13320 26858
rect 13268 26794 13320 26800
rect 12808 26444 12860 26450
rect 12808 26386 12860 26392
rect 13176 26444 13228 26450
rect 13176 26386 13228 26392
rect 12820 25294 12848 26386
rect 13188 25702 13216 26386
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 13176 25696 13228 25702
rect 13176 25638 13228 25644
rect 12808 25288 12860 25294
rect 12808 25230 12860 25236
rect 12820 24954 12848 25230
rect 12808 24948 12860 24954
rect 12808 24890 12860 24896
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 12808 22500 12860 22506
rect 12808 22442 12860 22448
rect 12820 22166 12848 22442
rect 12808 22160 12860 22166
rect 12808 22102 12860 22108
rect 12820 21690 12848 22102
rect 13004 22098 13032 23666
rect 12992 22092 13044 22098
rect 12992 22034 13044 22040
rect 12900 22024 12952 22030
rect 12900 21966 12952 21972
rect 12716 21684 12768 21690
rect 12716 21626 12768 21632
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 12820 21418 12848 21626
rect 12912 21486 12940 21966
rect 13004 21690 13032 22034
rect 12992 21684 13044 21690
rect 12992 21626 13044 21632
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 12808 21412 12860 21418
rect 12808 21354 12860 21360
rect 12820 21078 12848 21354
rect 12912 21146 12940 21422
rect 12900 21140 12952 21146
rect 12900 21082 12952 21088
rect 12808 21072 12860 21078
rect 12808 21014 12860 21020
rect 12532 21004 12584 21010
rect 12532 20946 12584 20952
rect 12544 20602 12572 20946
rect 12808 20868 12860 20874
rect 12808 20810 12860 20816
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 12636 19514 12664 20334
rect 12164 19508 12216 19514
rect 12164 19450 12216 19456
rect 12624 19508 12676 19514
rect 12624 19450 12676 19456
rect 12176 19310 12204 19450
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12820 18834 12848 20810
rect 13188 20398 13216 25638
rect 13280 25430 13308 25842
rect 13268 25424 13320 25430
rect 13268 25366 13320 25372
rect 13372 24410 13400 30126
rect 13452 29776 13504 29782
rect 13452 29718 13504 29724
rect 13464 29306 13492 29718
rect 13452 29300 13504 29306
rect 13452 29242 13504 29248
rect 13544 25764 13596 25770
rect 13544 25706 13596 25712
rect 13556 24954 13584 25706
rect 13648 25362 13676 30738
rect 13740 30122 13768 30874
rect 14292 30394 14320 37334
rect 14372 37120 14424 37126
rect 14372 37062 14424 37068
rect 14384 35698 14412 37062
rect 14464 36576 14516 36582
rect 14464 36518 14516 36524
rect 14372 35692 14424 35698
rect 14372 35634 14424 35640
rect 14384 35290 14412 35634
rect 14476 35562 14504 36518
rect 14464 35556 14516 35562
rect 14464 35498 14516 35504
rect 14372 35284 14424 35290
rect 14372 35226 14424 35232
rect 14476 35154 14504 35498
rect 14464 35148 14516 35154
rect 14464 35090 14516 35096
rect 14476 34746 14504 35090
rect 14568 34746 14596 38655
rect 14740 37800 14792 37806
rect 14740 37742 14792 37748
rect 14752 37670 14780 37742
rect 15292 37732 15344 37738
rect 15292 37674 15344 37680
rect 14740 37664 14792 37670
rect 14740 37606 14792 37612
rect 14752 37233 14780 37606
rect 15304 37466 15332 37674
rect 15292 37460 15344 37466
rect 15292 37402 15344 37408
rect 14738 37224 14794 37233
rect 14738 37159 14794 37168
rect 14648 36032 14700 36038
rect 14648 35974 14700 35980
rect 14464 34740 14516 34746
rect 14464 34682 14516 34688
rect 14556 34740 14608 34746
rect 14556 34682 14608 34688
rect 14476 34474 14504 34682
rect 14464 34468 14516 34474
rect 14464 34410 14516 34416
rect 14568 34066 14596 34682
rect 14660 34610 14688 35974
rect 14648 34604 14700 34610
rect 14648 34546 14700 34552
rect 14660 34202 14688 34546
rect 14648 34196 14700 34202
rect 14648 34138 14700 34144
rect 14752 34082 14780 37159
rect 15200 36644 15252 36650
rect 15200 36586 15252 36592
rect 15212 36378 15240 36586
rect 15200 36372 15252 36378
rect 15200 36314 15252 36320
rect 15292 36236 15344 36242
rect 15292 36178 15344 36184
rect 15304 35494 15332 36178
rect 15292 35488 15344 35494
rect 15292 35430 15344 35436
rect 14556 34060 14608 34066
rect 14556 34002 14608 34008
rect 14660 34054 14780 34082
rect 14556 33312 14608 33318
rect 14554 33280 14556 33289
rect 14608 33280 14610 33289
rect 14554 33215 14610 33224
rect 14568 33046 14596 33215
rect 14556 33040 14608 33046
rect 14556 32982 14608 32988
rect 14660 30802 14688 34054
rect 14740 33516 14792 33522
rect 14740 33458 14792 33464
rect 14752 33114 14780 33458
rect 14924 33312 14976 33318
rect 14844 33272 14924 33300
rect 14740 33108 14792 33114
rect 14740 33050 14792 33056
rect 14844 32298 14872 33272
rect 14924 33254 14976 33260
rect 14740 32292 14792 32298
rect 14740 32234 14792 32240
rect 14832 32292 14884 32298
rect 14832 32234 14884 32240
rect 14752 31686 14780 32234
rect 14844 31958 14872 32234
rect 14832 31952 14884 31958
rect 14832 31894 14884 31900
rect 14740 31680 14792 31686
rect 14740 31622 14792 31628
rect 15304 31278 15332 35430
rect 15396 34610 15424 38830
rect 15476 38480 15528 38486
rect 15476 38422 15528 38428
rect 15488 37738 15516 38422
rect 15844 38344 15896 38350
rect 15844 38286 15896 38292
rect 15856 37942 15884 38286
rect 15844 37936 15896 37942
rect 15844 37878 15896 37884
rect 15476 37732 15528 37738
rect 15476 37674 15528 37680
rect 15856 37466 15884 37878
rect 15948 37806 15976 39374
rect 16040 38350 16068 39510
rect 16028 38344 16080 38350
rect 16028 38286 16080 38292
rect 15936 37800 15988 37806
rect 15936 37742 15988 37748
rect 15844 37460 15896 37466
rect 15844 37402 15896 37408
rect 15948 36854 15976 37742
rect 16028 37324 16080 37330
rect 16028 37266 16080 37272
rect 16040 36922 16068 37266
rect 16028 36916 16080 36922
rect 16028 36858 16080 36864
rect 15936 36848 15988 36854
rect 15936 36790 15988 36796
rect 15948 35562 15976 36790
rect 16040 36145 16068 36858
rect 16026 36136 16082 36145
rect 16026 36071 16082 36080
rect 15936 35556 15988 35562
rect 15936 35498 15988 35504
rect 15660 35216 15712 35222
rect 15660 35158 15712 35164
rect 15568 35080 15620 35086
rect 15568 35022 15620 35028
rect 15384 34604 15436 34610
rect 15384 34546 15436 34552
rect 15580 34202 15608 35022
rect 15672 34678 15700 35158
rect 15660 34672 15712 34678
rect 15660 34614 15712 34620
rect 15568 34196 15620 34202
rect 15568 34138 15620 34144
rect 15476 34128 15528 34134
rect 15476 34070 15528 34076
rect 15384 33992 15436 33998
rect 15384 33934 15436 33940
rect 15396 33658 15424 33934
rect 15384 33652 15436 33658
rect 15384 33594 15436 33600
rect 15384 33380 15436 33386
rect 15384 33322 15436 33328
rect 15396 32434 15424 33322
rect 15488 33318 15516 34070
rect 15936 33924 15988 33930
rect 15936 33866 15988 33872
rect 15476 33312 15528 33318
rect 15476 33254 15528 33260
rect 15566 33280 15622 33289
rect 15566 33215 15622 33224
rect 15580 33134 15608 33215
rect 15488 33106 15608 33134
rect 15384 32428 15436 32434
rect 15384 32370 15436 32376
rect 15488 31958 15516 33106
rect 15752 32972 15804 32978
rect 15752 32914 15804 32920
rect 15764 32230 15792 32914
rect 15844 32428 15896 32434
rect 15844 32370 15896 32376
rect 15752 32224 15804 32230
rect 15752 32166 15804 32172
rect 15476 31952 15528 31958
rect 15476 31894 15528 31900
rect 15384 31816 15436 31822
rect 15384 31758 15436 31764
rect 15396 31346 15424 31758
rect 15488 31482 15516 31894
rect 15476 31476 15528 31482
rect 15476 31418 15528 31424
rect 15384 31340 15436 31346
rect 15384 31282 15436 31288
rect 15292 31272 15344 31278
rect 15292 31214 15344 31220
rect 14924 31136 14976 31142
rect 14924 31078 14976 31084
rect 14648 30796 14700 30802
rect 14648 30738 14700 30744
rect 14372 30592 14424 30598
rect 14372 30534 14424 30540
rect 14280 30388 14332 30394
rect 14280 30330 14332 30336
rect 14384 30190 14412 30534
rect 14660 30394 14688 30738
rect 14648 30388 14700 30394
rect 14648 30330 14700 30336
rect 14372 30184 14424 30190
rect 14372 30126 14424 30132
rect 13728 30116 13780 30122
rect 13728 30058 13780 30064
rect 13820 30116 13872 30122
rect 13820 30058 13872 30064
rect 13832 29850 13860 30058
rect 13820 29844 13872 29850
rect 13820 29786 13872 29792
rect 14384 29714 14412 30126
rect 14372 29708 14424 29714
rect 14372 29650 14424 29656
rect 14648 29640 14700 29646
rect 14648 29582 14700 29588
rect 14660 29306 14688 29582
rect 14648 29300 14700 29306
rect 14648 29242 14700 29248
rect 14936 29102 14964 31078
rect 15476 30864 15528 30870
rect 15476 30806 15528 30812
rect 15016 30728 15068 30734
rect 15016 30670 15068 30676
rect 15028 29850 15056 30670
rect 15488 30122 15516 30806
rect 15476 30116 15528 30122
rect 15476 30058 15528 30064
rect 15016 29844 15068 29850
rect 15016 29786 15068 29792
rect 15488 29782 15516 30058
rect 15476 29776 15528 29782
rect 15476 29718 15528 29724
rect 15488 29306 15516 29718
rect 15476 29300 15528 29306
rect 15476 29242 15528 29248
rect 14464 29096 14516 29102
rect 14464 29038 14516 29044
rect 14924 29096 14976 29102
rect 14924 29038 14976 29044
rect 14280 28620 14332 28626
rect 14280 28562 14332 28568
rect 14292 28257 14320 28562
rect 14278 28248 14334 28257
rect 14278 28183 14334 28192
rect 14188 28076 14240 28082
rect 14188 28018 14240 28024
rect 13728 27872 13780 27878
rect 13728 27814 13780 27820
rect 13740 27674 13768 27814
rect 13728 27668 13780 27674
rect 13728 27610 13780 27616
rect 14200 27606 14228 28018
rect 14292 28014 14320 28183
rect 14280 28008 14332 28014
rect 14280 27950 14332 27956
rect 14188 27600 14240 27606
rect 14188 27542 14240 27548
rect 13820 27464 13872 27470
rect 13820 27406 13872 27412
rect 13832 27130 13860 27406
rect 13820 27124 13872 27130
rect 13820 27066 13872 27072
rect 13912 25764 13964 25770
rect 13912 25706 13964 25712
rect 13636 25356 13688 25362
rect 13636 25298 13688 25304
rect 13924 25226 13952 25706
rect 14188 25356 14240 25362
rect 14188 25298 14240 25304
rect 13912 25220 13964 25226
rect 13912 25162 13964 25168
rect 13544 24948 13596 24954
rect 13544 24890 13596 24896
rect 13452 24676 13504 24682
rect 13452 24618 13504 24624
rect 13360 24404 13412 24410
rect 13360 24346 13412 24352
rect 13464 24274 13492 24618
rect 14200 24614 14228 25298
rect 14188 24608 14240 24614
rect 14188 24550 14240 24556
rect 13268 24268 13320 24274
rect 13268 24210 13320 24216
rect 13452 24268 13504 24274
rect 13452 24210 13504 24216
rect 13280 23866 13308 24210
rect 13268 23860 13320 23866
rect 13268 23802 13320 23808
rect 13464 23322 13492 24210
rect 13452 23316 13504 23322
rect 13452 23258 13504 23264
rect 14200 22137 14228 24550
rect 14292 23186 14320 27950
rect 14372 26444 14424 26450
rect 14372 26386 14424 26392
rect 14384 26042 14412 26386
rect 14372 26036 14424 26042
rect 14372 25978 14424 25984
rect 14372 24744 14424 24750
rect 14372 24686 14424 24692
rect 14384 24410 14412 24686
rect 14372 24404 14424 24410
rect 14372 24346 14424 24352
rect 14384 24138 14412 24346
rect 14372 24132 14424 24138
rect 14372 24074 14424 24080
rect 14372 23724 14424 23730
rect 14372 23666 14424 23672
rect 14280 23180 14332 23186
rect 14280 23122 14332 23128
rect 14292 22778 14320 23122
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 14186 22128 14242 22137
rect 14186 22063 14242 22072
rect 14004 21004 14056 21010
rect 14004 20946 14056 20952
rect 14016 20602 14044 20946
rect 14004 20596 14056 20602
rect 14004 20538 14056 20544
rect 13176 20392 13228 20398
rect 13176 20334 13228 20340
rect 13728 20324 13780 20330
rect 13728 20266 13780 20272
rect 13268 19984 13320 19990
rect 13268 19926 13320 19932
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 13096 18902 13124 19110
rect 13188 18970 13216 19790
rect 13280 19174 13308 19926
rect 13360 19780 13412 19786
rect 13360 19722 13412 19728
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13176 18964 13228 18970
rect 13228 18924 13308 18952
rect 13176 18906 13228 18912
rect 13084 18896 13136 18902
rect 13084 18838 13136 18844
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12808 18828 12860 18834
rect 12808 18770 12860 18776
rect 12084 18426 12112 18770
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 13084 18352 13136 18358
rect 13084 18294 13136 18300
rect 13096 18154 13124 18294
rect 12992 18148 13044 18154
rect 12992 18090 13044 18096
rect 13084 18148 13136 18154
rect 13084 18090 13136 18096
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 11900 17814 11928 18022
rect 13004 17882 13032 18090
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 11888 17808 11940 17814
rect 11888 17750 11940 17756
rect 12532 17604 12584 17610
rect 12532 17546 12584 17552
rect 12544 17202 12572 17546
rect 13004 17202 13032 17818
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 13188 17338 13216 17750
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11900 15978 11928 16934
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12268 16250 12296 16526
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 11888 15972 11940 15978
rect 11888 15914 11940 15920
rect 11900 13852 11928 15914
rect 12636 15638 12664 17002
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 12728 16250 12756 16662
rect 13004 16590 13032 17138
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 13280 16114 13308 18924
rect 13372 18290 13400 19722
rect 13634 19272 13690 19281
rect 13634 19207 13690 19216
rect 13648 19174 13676 19207
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13740 18902 13768 20266
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14108 19281 14136 19654
rect 14280 19440 14332 19446
rect 14280 19382 14332 19388
rect 14094 19272 14150 19281
rect 13820 19236 13872 19242
rect 14094 19207 14150 19216
rect 13820 19178 13872 19184
rect 13832 18970 13860 19178
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13728 18896 13780 18902
rect 13728 18838 13780 18844
rect 13636 18760 13688 18766
rect 13636 18702 13688 18708
rect 13648 18426 13676 18702
rect 13636 18420 13688 18426
rect 13636 18362 13688 18368
rect 13740 18358 13768 18838
rect 13728 18352 13780 18358
rect 13728 18294 13780 18300
rect 13360 18284 13412 18290
rect 13360 18226 13412 18232
rect 13740 18086 13768 18294
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13452 17808 13504 17814
rect 13452 17750 13504 17756
rect 13464 17270 13492 17750
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 13360 16244 13412 16250
rect 13360 16186 13412 16192
rect 13268 16108 13320 16114
rect 13188 16068 13268 16096
rect 12624 15632 12676 15638
rect 12624 15574 12676 15580
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12176 14890 12204 15438
rect 12636 15162 12664 15574
rect 13188 15434 13216 16068
rect 13268 16050 13320 16056
rect 13372 15978 13400 16186
rect 13268 15972 13320 15978
rect 13268 15914 13320 15920
rect 13360 15972 13412 15978
rect 13360 15914 13412 15920
rect 13280 15706 13308 15914
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 13176 15428 13228 15434
rect 13176 15370 13228 15376
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12164 14884 12216 14890
rect 12164 14826 12216 14832
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11992 14550 12020 14758
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 11992 14006 12020 14486
rect 12176 14414 12204 14826
rect 13280 14414 13308 15642
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 13372 14618 13400 14758
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 11980 14000 12032 14006
rect 11980 13942 12032 13948
rect 11980 13864 12032 13870
rect 11900 13824 11980 13852
rect 11980 13806 12032 13812
rect 11992 13462 12020 13806
rect 12176 13462 12204 14350
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13280 13802 13308 14214
rect 13372 14074 13400 14554
rect 13464 14532 13492 17206
rect 14108 15026 14136 19207
rect 14292 18902 14320 19382
rect 14280 18896 14332 18902
rect 14280 18838 14332 18844
rect 14292 18698 14320 18838
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 14292 16794 14320 17070
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 13544 14544 13596 14550
rect 13464 14504 13544 14532
rect 13464 14074 13492 14504
rect 13544 14486 13596 14492
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13556 13938 13584 14350
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13372 13802 13400 13874
rect 13268 13796 13320 13802
rect 13268 13738 13320 13744
rect 13360 13796 13412 13802
rect 13360 13738 13412 13744
rect 13280 13530 13308 13738
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13648 13462 13676 13670
rect 14108 13530 14136 14758
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 12164 13456 12216 13462
rect 12164 13398 12216 13404
rect 13636 13456 13688 13462
rect 13636 13398 13688 13404
rect 13648 12986 13676 13398
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12808 12708 12860 12714
rect 12808 12650 12860 12656
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12544 11762 12572 12174
rect 12714 11792 12770 11801
rect 12532 11756 12584 11762
rect 12714 11727 12770 11736
rect 12532 11698 12584 11704
rect 12728 11694 12756 11727
rect 12820 11694 12848 12650
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 11888 11280 11940 11286
rect 11888 11222 11940 11228
rect 11900 10810 11928 11222
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 12452 10606 12480 11290
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10704 10130 10732 10542
rect 12452 10266 12480 10542
rect 12544 10538 12572 11154
rect 12728 10810 12756 11630
rect 12912 11218 12940 12718
rect 13648 12374 13676 12922
rect 13924 12850 13952 13262
rect 14096 12912 14148 12918
rect 14096 12854 14148 12860
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 13924 12442 13952 12786
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 13648 11830 13676 12310
rect 14004 12164 14056 12170
rect 14004 12106 14056 12112
rect 13636 11824 13688 11830
rect 13636 11766 13688 11772
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 12912 11121 12940 11154
rect 12898 11112 12954 11121
rect 12898 11047 12954 11056
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 11244 10192 11296 10198
rect 11244 10134 11296 10140
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10414 9959 10470 9968
rect 10508 9988 10560 9994
rect 9784 9450 9812 9959
rect 10508 9930 10560 9936
rect 10704 9722 10732 10066
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10888 9450 10916 9862
rect 9220 9444 9272 9450
rect 9220 9386 9272 9392
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9956 9444 10008 9450
rect 9956 9386 10008 9392
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 9968 9178 9996 9386
rect 10888 9178 10916 9386
rect 11256 9178 11284 10134
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 11900 9926 11928 10066
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 12176 9674 12204 10066
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12084 9646 12204 9674
rect 11336 9444 11388 9450
rect 11336 9386 11388 9392
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 8588 7342 8616 8842
rect 8772 8634 8800 8978
rect 8760 8628 8812 8634
rect 8680 8588 8760 8616
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1688 82 1716 3334
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 8680 3194 8708 8588
rect 8760 8570 8812 8576
rect 9876 8294 9904 9046
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10060 8294 10088 8910
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10428 8362 10456 8774
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 9876 7546 9904 8230
rect 10428 7750 10456 8298
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9876 7274 9904 7482
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9968 7002 9996 7278
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 10244 6866 10272 7346
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10244 6390 10272 6802
rect 10232 6384 10284 6390
rect 10232 6326 10284 6332
rect 10244 5914 10272 6326
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9600 4146 9628 4966
rect 10428 4842 10456 7686
rect 10520 6866 10548 8366
rect 10600 8016 10652 8022
rect 10600 7958 10652 7964
rect 10612 7546 10640 7958
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11164 7546 11192 7822
rect 11348 7818 11376 9386
rect 12084 9382 12112 9646
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 11900 8362 11928 8978
rect 12084 8634 12112 8978
rect 12636 8838 12664 9862
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 10612 7002 10640 7482
rect 10784 7268 10836 7274
rect 10784 7210 10836 7216
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10520 6458 10548 6802
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10506 4856 10562 4865
rect 10428 4814 10506 4842
rect 10612 4826 10640 5102
rect 10506 4791 10562 4800
rect 10600 4820 10652 4826
rect 10520 4690 10548 4791
rect 10600 4762 10652 4768
rect 10704 4690 10732 6122
rect 10796 5914 10824 7210
rect 12084 6662 12112 7822
rect 12176 7478 12204 7958
rect 12164 7472 12216 7478
rect 12164 7414 12216 7420
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12452 7002 12480 7278
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12728 6866 12756 10406
rect 13648 10146 13676 10610
rect 13740 10538 13768 11154
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 13832 10470 13860 11154
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13510 10130 13676 10146
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13498 10124 13676 10130
rect 13550 10118 13676 10124
rect 13498 10066 13550 10072
rect 13280 9382 13308 10066
rect 13648 9738 13676 10118
rect 13556 9710 13676 9738
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13280 9042 13308 9318
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13188 8498 13216 8774
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13280 8294 13308 8978
rect 13372 8974 13400 9386
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13372 8634 13400 8910
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13556 8430 13584 9710
rect 13832 9674 13860 10406
rect 13648 9654 13860 9674
rect 13636 9648 13860 9654
rect 13688 9646 13860 9648
rect 13636 9590 13688 9596
rect 13648 9042 13676 9590
rect 14016 9110 14044 12106
rect 14108 9518 14136 12854
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14200 12442 14228 12718
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14292 10538 14320 11086
rect 14280 10532 14332 10538
rect 14280 10474 14332 10480
rect 14292 10266 14320 10474
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14004 9104 14056 9110
rect 14004 9046 14056 9052
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13556 8090 13584 8366
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13648 7936 13676 8230
rect 13740 8090 13768 8978
rect 14108 8430 14136 9318
rect 14200 8974 14228 9862
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14292 8634 14320 8774
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13728 7948 13780 7954
rect 13648 7908 13728 7936
rect 13728 7890 13780 7896
rect 13740 7410 13768 7890
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 14108 7342 14136 8366
rect 14292 7546 14320 8570
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10796 5370 10824 5850
rect 10888 5710 10916 6122
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10796 5098 10824 5306
rect 10784 5092 10836 5098
rect 10784 5034 10836 5040
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10520 4214 10548 4626
rect 10704 4282 10732 4626
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 11256 3738 11284 6598
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11348 4826 11376 5646
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11336 4004 11388 4010
rect 11440 3992 11468 5510
rect 11808 5370 11836 6054
rect 12544 5914 12572 6734
rect 12728 6458 12756 6802
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 12728 5778 12756 6394
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12728 5370 12756 5714
rect 12820 5574 12848 6258
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12438 5264 12494 5273
rect 12438 5199 12494 5208
rect 12452 4758 12480 5199
rect 12440 4752 12492 4758
rect 12440 4694 12492 4700
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 12360 4078 12388 4218
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 11388 3964 11468 3992
rect 11336 3946 11388 3952
rect 11440 3738 11468 3964
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11532 3398 11560 3538
rect 12452 3534 12480 4694
rect 12728 4146 12756 5306
rect 12820 4826 12848 5510
rect 13096 5234 13124 5850
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 13188 4622 13216 5714
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 13280 4078 13308 7142
rect 14384 7002 14412 23666
rect 14476 23662 14504 29038
rect 15016 28960 15068 28966
rect 15016 28902 15068 28908
rect 15028 28762 15056 28902
rect 15016 28756 15068 28762
rect 15016 28698 15068 28704
rect 15476 28688 15528 28694
rect 15476 28630 15528 28636
rect 15016 28416 15068 28422
rect 15016 28358 15068 28364
rect 15028 26994 15056 28358
rect 15292 28076 15344 28082
rect 15292 28018 15344 28024
rect 15108 27940 15160 27946
rect 15108 27882 15160 27888
rect 15120 27334 15148 27882
rect 15108 27328 15160 27334
rect 15108 27270 15160 27276
rect 15120 27130 15148 27270
rect 15108 27124 15160 27130
rect 15108 27066 15160 27072
rect 15016 26988 15068 26994
rect 15016 26930 15068 26936
rect 15028 26586 15056 26930
rect 15016 26580 15068 26586
rect 15016 26522 15068 26528
rect 15200 26376 15252 26382
rect 15200 26318 15252 26324
rect 14924 25968 14976 25974
rect 14924 25910 14976 25916
rect 14936 25770 14964 25910
rect 14832 25764 14884 25770
rect 14832 25706 14884 25712
rect 14924 25764 14976 25770
rect 14924 25706 14976 25712
rect 14844 25498 14872 25706
rect 14832 25492 14884 25498
rect 14832 25434 14884 25440
rect 15108 25288 15160 25294
rect 15108 25230 15160 25236
rect 14556 24948 14608 24954
rect 14556 24890 14608 24896
rect 14464 23656 14516 23662
rect 14464 23598 14516 23604
rect 14568 23474 14596 24890
rect 15120 24682 15148 25230
rect 15212 25158 15240 26318
rect 15304 25906 15332 28018
rect 15488 27946 15516 28630
rect 15660 28552 15712 28558
rect 15660 28494 15712 28500
rect 15476 27940 15528 27946
rect 15476 27882 15528 27888
rect 15476 27600 15528 27606
rect 15382 27568 15438 27577
rect 15476 27542 15528 27548
rect 15382 27503 15438 27512
rect 15396 27470 15424 27503
rect 15384 27464 15436 27470
rect 15384 27406 15436 27412
rect 15396 26586 15424 27406
rect 15488 26790 15516 27542
rect 15672 26994 15700 28494
rect 15764 28257 15792 32166
rect 15856 30326 15884 32370
rect 15948 31754 15976 33866
rect 16028 33652 16080 33658
rect 16028 33594 16080 33600
rect 16040 33114 16068 33594
rect 16028 33108 16080 33114
rect 16028 33050 16080 33056
rect 15936 31748 15988 31754
rect 15936 31690 15988 31696
rect 15844 30320 15896 30326
rect 15844 30262 15896 30268
rect 15948 29578 15976 31690
rect 16132 31414 16160 49506
rect 19444 49475 19472 49506
rect 19580 47356 19876 47376
rect 19636 47354 19660 47356
rect 19716 47354 19740 47356
rect 19796 47354 19820 47356
rect 19658 47302 19660 47354
rect 19722 47302 19734 47354
rect 19796 47302 19798 47354
rect 19636 47300 19660 47302
rect 19716 47300 19740 47302
rect 19796 47300 19820 47302
rect 19580 47280 19876 47300
rect 19580 46268 19876 46288
rect 19636 46266 19660 46268
rect 19716 46266 19740 46268
rect 19796 46266 19820 46268
rect 19658 46214 19660 46266
rect 19722 46214 19734 46266
rect 19796 46214 19798 46266
rect 19636 46212 19660 46214
rect 19716 46212 19740 46214
rect 19796 46212 19820 46214
rect 19580 46192 19876 46212
rect 19580 45180 19876 45200
rect 19636 45178 19660 45180
rect 19716 45178 19740 45180
rect 19796 45178 19820 45180
rect 19658 45126 19660 45178
rect 19722 45126 19734 45178
rect 19796 45126 19798 45178
rect 19636 45124 19660 45126
rect 19716 45124 19740 45126
rect 19796 45124 19820 45126
rect 19580 45104 19876 45124
rect 19580 44092 19876 44112
rect 19636 44090 19660 44092
rect 19716 44090 19740 44092
rect 19796 44090 19820 44092
rect 19658 44038 19660 44090
rect 19722 44038 19734 44090
rect 19796 44038 19798 44090
rect 19636 44036 19660 44038
rect 19716 44036 19740 44038
rect 19796 44036 19820 44038
rect 19580 44016 19876 44036
rect 19580 43004 19876 43024
rect 19636 43002 19660 43004
rect 19716 43002 19740 43004
rect 19796 43002 19820 43004
rect 19658 42950 19660 43002
rect 19722 42950 19734 43002
rect 19796 42950 19798 43002
rect 19636 42948 19660 42950
rect 19716 42948 19740 42950
rect 19796 42948 19820 42950
rect 19580 42928 19876 42948
rect 19580 41916 19876 41936
rect 19636 41914 19660 41916
rect 19716 41914 19740 41916
rect 19796 41914 19820 41916
rect 19658 41862 19660 41914
rect 19722 41862 19734 41914
rect 19796 41862 19798 41914
rect 19636 41860 19660 41862
rect 19716 41860 19740 41862
rect 19796 41860 19820 41862
rect 19580 41840 19876 41860
rect 19062 41712 19118 41721
rect 17500 41676 17552 41682
rect 19062 41647 19064 41656
rect 17500 41618 17552 41624
rect 19116 41647 19118 41656
rect 19064 41618 19116 41624
rect 16488 41472 16540 41478
rect 16488 41414 16540 41420
rect 16580 41472 16632 41478
rect 16580 41414 16632 41420
rect 16500 41138 16528 41414
rect 16488 41132 16540 41138
rect 16488 41074 16540 41080
rect 16488 40928 16540 40934
rect 16488 40870 16540 40876
rect 16212 40384 16264 40390
rect 16212 40326 16264 40332
rect 16224 39642 16252 40326
rect 16396 39840 16448 39846
rect 16396 39782 16448 39788
rect 16212 39636 16264 39642
rect 16212 39578 16264 39584
rect 16408 39574 16436 39782
rect 16500 39642 16528 40870
rect 16592 40050 16620 41414
rect 17512 41070 17540 41618
rect 19076 41274 19104 41618
rect 19156 41472 19208 41478
rect 19156 41414 19208 41420
rect 19432 41472 19484 41478
rect 19432 41414 19484 41420
rect 19708 41472 19760 41478
rect 19708 41414 19760 41420
rect 19064 41268 19116 41274
rect 19064 41210 19116 41216
rect 17500 41064 17552 41070
rect 17500 41006 17552 41012
rect 18604 41064 18656 41070
rect 18788 41064 18840 41070
rect 18604 41006 18656 41012
rect 18786 41032 18788 41041
rect 18840 41032 18842 41041
rect 18420 40996 18472 41002
rect 18420 40938 18472 40944
rect 16764 40656 16816 40662
rect 16764 40598 16816 40604
rect 16672 40384 16724 40390
rect 16672 40326 16724 40332
rect 16580 40044 16632 40050
rect 16580 39986 16632 39992
rect 16488 39636 16540 39642
rect 16488 39578 16540 39584
rect 16396 39568 16448 39574
rect 16396 39510 16448 39516
rect 16500 38962 16528 39578
rect 16684 39574 16712 40326
rect 16776 39914 16804 40598
rect 17868 40588 17920 40594
rect 17868 40530 17920 40536
rect 17224 40520 17276 40526
rect 17224 40462 17276 40468
rect 16764 39908 16816 39914
rect 16764 39850 16816 39856
rect 16776 39574 16804 39850
rect 16672 39568 16724 39574
rect 16672 39510 16724 39516
rect 16764 39568 16816 39574
rect 16764 39510 16816 39516
rect 16488 38956 16540 38962
rect 16488 38898 16540 38904
rect 16684 38554 16712 39510
rect 16776 39098 16804 39510
rect 16764 39092 16816 39098
rect 16764 39034 16816 39040
rect 17236 38894 17264 40462
rect 17880 40186 17908 40530
rect 17868 40180 17920 40186
rect 17920 40140 18000 40168
rect 17868 40122 17920 40128
rect 17500 39908 17552 39914
rect 17500 39850 17552 39856
rect 17224 38888 17276 38894
rect 17224 38830 17276 38836
rect 16672 38548 16724 38554
rect 16672 38490 16724 38496
rect 17236 38350 17264 38830
rect 16948 38344 17000 38350
rect 16948 38286 17000 38292
rect 17224 38344 17276 38350
rect 17224 38286 17276 38292
rect 16960 37738 16988 38286
rect 17224 37936 17276 37942
rect 17224 37878 17276 37884
rect 17236 37806 17264 37878
rect 17224 37800 17276 37806
rect 17224 37742 17276 37748
rect 16948 37732 17000 37738
rect 16948 37674 17000 37680
rect 17236 37398 17264 37742
rect 17224 37392 17276 37398
rect 17224 37334 17276 37340
rect 16488 37324 16540 37330
rect 16488 37266 16540 37272
rect 17040 37324 17092 37330
rect 17040 37266 17092 37272
rect 16500 36582 16528 37266
rect 17052 36922 17080 37266
rect 17316 37256 17368 37262
rect 17316 37198 17368 37204
rect 17040 36916 17092 36922
rect 17040 36858 17092 36864
rect 16764 36780 16816 36786
rect 16764 36722 16816 36728
rect 16488 36576 16540 36582
rect 16488 36518 16540 36524
rect 16304 36372 16356 36378
rect 16304 36314 16356 36320
rect 16316 35834 16344 36314
rect 16396 36168 16448 36174
rect 16396 36110 16448 36116
rect 16304 35828 16356 35834
rect 16304 35770 16356 35776
rect 16316 35222 16344 35770
rect 16408 35290 16436 36110
rect 16500 36106 16528 36518
rect 16488 36100 16540 36106
rect 16488 36042 16540 36048
rect 16500 35977 16528 36042
rect 16580 36032 16632 36038
rect 16580 35974 16632 35980
rect 16592 35698 16620 35974
rect 16776 35698 16804 36722
rect 17328 36242 17356 37198
rect 17408 36576 17460 36582
rect 17408 36518 17460 36524
rect 17316 36236 17368 36242
rect 17316 36178 17368 36184
rect 17222 36136 17278 36145
rect 17222 36071 17278 36080
rect 16580 35692 16632 35698
rect 16580 35634 16632 35640
rect 16764 35692 16816 35698
rect 16764 35634 16816 35640
rect 16592 35562 16620 35634
rect 16580 35556 16632 35562
rect 16580 35498 16632 35504
rect 16396 35284 16448 35290
rect 16396 35226 16448 35232
rect 16304 35216 16356 35222
rect 16304 35158 16356 35164
rect 16488 34944 16540 34950
rect 16488 34886 16540 34892
rect 16500 34474 16528 34886
rect 16776 34678 16804 35634
rect 16764 34672 16816 34678
rect 16764 34614 16816 34620
rect 16672 34604 16724 34610
rect 16672 34546 16724 34552
rect 16488 34468 16540 34474
rect 16488 34410 16540 34416
rect 16580 34400 16632 34406
rect 16580 34342 16632 34348
rect 16488 32428 16540 32434
rect 16488 32370 16540 32376
rect 16500 32026 16528 32370
rect 16488 32020 16540 32026
rect 16488 31962 16540 31968
rect 16120 31408 16172 31414
rect 16120 31350 16172 31356
rect 16488 31272 16540 31278
rect 16408 31232 16488 31260
rect 16408 30598 16436 31232
rect 16488 31214 16540 31220
rect 16396 30592 16448 30598
rect 16396 30534 16448 30540
rect 16304 30048 16356 30054
rect 16304 29990 16356 29996
rect 16316 29646 16344 29990
rect 16304 29640 16356 29646
rect 16304 29582 16356 29588
rect 15936 29572 15988 29578
rect 15936 29514 15988 29520
rect 16408 29492 16436 30534
rect 16316 29464 16436 29492
rect 16212 29096 16264 29102
rect 16212 29038 16264 29044
rect 15750 28248 15806 28257
rect 15750 28183 15806 28192
rect 15752 27940 15804 27946
rect 15752 27882 15804 27888
rect 15764 27470 15792 27882
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 15660 26988 15712 26994
rect 15660 26930 15712 26936
rect 15476 26784 15528 26790
rect 15476 26726 15528 26732
rect 15384 26580 15436 26586
rect 15384 26522 15436 26528
rect 15672 26314 15700 26930
rect 16224 26518 16252 29038
rect 16316 29034 16344 29464
rect 16592 29102 16620 34342
rect 16684 34202 16712 34546
rect 16672 34196 16724 34202
rect 16672 34138 16724 34144
rect 16764 33924 16816 33930
rect 16764 33866 16816 33872
rect 16580 29096 16632 29102
rect 16580 29038 16632 29044
rect 16304 29028 16356 29034
rect 16304 28970 16356 28976
rect 16316 28762 16344 28970
rect 16304 28756 16356 28762
rect 16304 28698 16356 28704
rect 16028 26512 16080 26518
rect 16028 26454 16080 26460
rect 16212 26512 16264 26518
rect 16212 26454 16264 26460
rect 15660 26308 15712 26314
rect 15660 26250 15712 26256
rect 16040 25974 16068 26454
rect 16028 25968 16080 25974
rect 16028 25910 16080 25916
rect 15292 25900 15344 25906
rect 15292 25842 15344 25848
rect 15304 25430 15332 25842
rect 16040 25770 16068 25910
rect 16028 25764 16080 25770
rect 16028 25706 16080 25712
rect 16488 25764 16540 25770
rect 16488 25706 16540 25712
rect 16500 25498 16528 25706
rect 16488 25492 16540 25498
rect 16488 25434 16540 25440
rect 15292 25424 15344 25430
rect 15292 25366 15344 25372
rect 15476 25424 15528 25430
rect 15476 25366 15528 25372
rect 15200 25152 15252 25158
rect 15200 25094 15252 25100
rect 15108 24676 15160 24682
rect 15108 24618 15160 24624
rect 15120 24410 15148 24618
rect 15108 24404 15160 24410
rect 15108 24346 15160 24352
rect 15212 24206 15240 25094
rect 15488 24954 15516 25366
rect 16304 25220 16356 25226
rect 16304 25162 16356 25168
rect 16212 25152 16264 25158
rect 16212 25094 16264 25100
rect 15476 24948 15528 24954
rect 15476 24890 15528 24896
rect 16120 24812 16172 24818
rect 16120 24754 16172 24760
rect 16132 24342 16160 24754
rect 16224 24682 16252 25094
rect 16316 24682 16344 25162
rect 16212 24676 16264 24682
rect 16212 24618 16264 24624
rect 16304 24676 16356 24682
rect 16304 24618 16356 24624
rect 16120 24336 16172 24342
rect 16120 24278 16172 24284
rect 16028 24268 16080 24274
rect 16028 24210 16080 24216
rect 15200 24200 15252 24206
rect 15200 24142 15252 24148
rect 15568 23792 15620 23798
rect 15568 23734 15620 23740
rect 15580 23594 15608 23734
rect 16040 23594 16068 24210
rect 14740 23588 14792 23594
rect 14740 23530 14792 23536
rect 15108 23588 15160 23594
rect 15108 23530 15160 23536
rect 15568 23588 15620 23594
rect 15568 23530 15620 23536
rect 15844 23588 15896 23594
rect 15844 23530 15896 23536
rect 16028 23588 16080 23594
rect 16028 23530 16080 23536
rect 14476 23446 14596 23474
rect 14476 22166 14504 23446
rect 14464 22160 14516 22166
rect 14464 22102 14516 22108
rect 14752 22030 14780 23530
rect 15120 23322 15148 23530
rect 15580 23322 15608 23530
rect 15108 23316 15160 23322
rect 15108 23258 15160 23264
rect 15568 23316 15620 23322
rect 15568 23258 15620 23264
rect 15856 23118 15884 23530
rect 16120 23520 16172 23526
rect 16120 23462 16172 23468
rect 15936 23316 15988 23322
rect 15936 23258 15988 23264
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 15844 23112 15896 23118
rect 15844 23054 15896 23060
rect 15108 22636 15160 22642
rect 15108 22578 15160 22584
rect 14832 22228 14884 22234
rect 14832 22170 14884 22176
rect 14740 22024 14792 22030
rect 14740 21966 14792 21972
rect 14844 20602 14872 22170
rect 15120 22166 15148 22578
rect 15396 22234 15424 23054
rect 15660 22976 15712 22982
rect 15660 22918 15712 22924
rect 15672 22710 15700 22918
rect 15476 22704 15528 22710
rect 15476 22646 15528 22652
rect 15660 22704 15712 22710
rect 15660 22646 15712 22652
rect 15488 22506 15516 22646
rect 15476 22500 15528 22506
rect 15476 22442 15528 22448
rect 15752 22432 15804 22438
rect 15752 22374 15804 22380
rect 15384 22228 15436 22234
rect 15384 22170 15436 22176
rect 15764 22166 15792 22374
rect 15856 22166 15884 23054
rect 15948 22438 15976 23258
rect 16132 22642 16160 23462
rect 16394 22672 16450 22681
rect 16120 22636 16172 22642
rect 16394 22607 16450 22616
rect 16120 22578 16172 22584
rect 15936 22432 15988 22438
rect 15936 22374 15988 22380
rect 15108 22160 15160 22166
rect 15108 22102 15160 22108
rect 15752 22160 15804 22166
rect 15752 22102 15804 22108
rect 15844 22160 15896 22166
rect 15844 22102 15896 22108
rect 15764 21418 15792 22102
rect 15948 21894 15976 22374
rect 15936 21888 15988 21894
rect 15936 21830 15988 21836
rect 15752 21412 15804 21418
rect 15752 21354 15804 21360
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 15212 19990 15240 20878
rect 15764 20330 15792 21354
rect 15844 21072 15896 21078
rect 15948 21060 15976 21830
rect 16028 21412 16080 21418
rect 16028 21354 16080 21360
rect 15896 21032 15976 21060
rect 15844 21014 15896 21020
rect 15856 20466 15884 21014
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15752 20324 15804 20330
rect 15752 20266 15804 20272
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15200 19984 15252 19990
rect 15200 19926 15252 19932
rect 15212 19514 15240 19926
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15396 19378 15424 20198
rect 15856 19990 15884 20402
rect 16040 20262 16068 21354
rect 16212 20868 16264 20874
rect 16212 20810 16264 20816
rect 16224 20534 16252 20810
rect 16408 20806 16436 22607
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 16592 21690 16620 21966
rect 16580 21684 16632 21690
rect 16580 21626 16632 21632
rect 16396 20800 16448 20806
rect 16396 20742 16448 20748
rect 16212 20528 16264 20534
rect 16212 20470 16264 20476
rect 16304 20324 16356 20330
rect 16304 20266 16356 20272
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 16040 19990 16068 20198
rect 16316 20058 16344 20266
rect 16304 20052 16356 20058
rect 16304 19994 16356 20000
rect 15844 19984 15896 19990
rect 15844 19926 15896 19932
rect 16028 19984 16080 19990
rect 16028 19926 16080 19932
rect 15856 19514 15884 19926
rect 15844 19508 15896 19514
rect 15844 19450 15896 19456
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15844 18828 15896 18834
rect 15844 18770 15896 18776
rect 15106 18320 15162 18329
rect 15106 18255 15162 18264
rect 15120 18222 15148 18255
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 14476 16658 14504 18158
rect 15856 18086 15884 18770
rect 16028 18148 16080 18154
rect 16028 18090 16080 18096
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14476 16250 14504 16594
rect 14464 16244 14516 16250
rect 14464 16186 14516 16192
rect 14568 16130 14596 17478
rect 14936 17338 14964 18022
rect 15568 17808 15620 17814
rect 15568 17750 15620 17756
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 14924 17332 14976 17338
rect 14924 17274 14976 17280
rect 15120 16794 15148 17614
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15108 16788 15160 16794
rect 15108 16730 15160 16736
rect 15488 16726 15516 17002
rect 15580 16998 15608 17750
rect 15856 17270 15884 18022
rect 16040 17678 16068 18090
rect 16028 17672 16080 17678
rect 16028 17614 16080 17620
rect 15844 17264 15896 17270
rect 15844 17206 15896 17212
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 15476 16720 15528 16726
rect 15476 16662 15528 16668
rect 14924 16584 14976 16590
rect 14924 16526 14976 16532
rect 14648 16516 14700 16522
rect 14648 16458 14700 16464
rect 14476 16102 14596 16130
rect 14476 13814 14504 16102
rect 14556 15972 14608 15978
rect 14556 15914 14608 15920
rect 14568 15162 14596 15914
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14568 14822 14596 15098
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14476 13786 14596 13814
rect 14568 10198 14596 13786
rect 14660 10810 14688 16458
rect 14936 16250 14964 16526
rect 15488 16250 15516 16662
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15580 15638 15608 16934
rect 16040 16726 16068 17614
rect 16028 16720 16080 16726
rect 16028 16662 16080 16668
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 15580 15162 15608 15574
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 15936 15428 15988 15434
rect 15936 15370 15988 15376
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 14752 14346 14780 14826
rect 15672 14550 15700 15302
rect 15948 15026 15976 15370
rect 16040 15162 16068 15438
rect 16408 15314 16436 20742
rect 16776 19922 16804 33866
rect 16948 33312 17000 33318
rect 16948 33254 17000 33260
rect 16960 31958 16988 33254
rect 17236 33134 17264 36071
rect 17316 35148 17368 35154
rect 17420 35136 17448 36518
rect 17368 35108 17448 35136
rect 17316 35090 17368 35096
rect 17328 34678 17356 35090
rect 17316 34672 17368 34678
rect 17316 34614 17368 34620
rect 17328 34406 17356 34614
rect 17316 34400 17368 34406
rect 17316 34342 17368 34348
rect 17512 34066 17540 39850
rect 17868 38752 17920 38758
rect 17868 38694 17920 38700
rect 17880 38554 17908 38694
rect 17868 38548 17920 38554
rect 17868 38490 17920 38496
rect 17684 38004 17736 38010
rect 17684 37946 17736 37952
rect 17592 37732 17644 37738
rect 17592 37674 17644 37680
rect 17604 37466 17632 37674
rect 17592 37460 17644 37466
rect 17592 37402 17644 37408
rect 17500 34060 17552 34066
rect 17500 34002 17552 34008
rect 17512 33658 17540 34002
rect 17500 33652 17552 33658
rect 17500 33594 17552 33600
rect 17696 33134 17724 37946
rect 17776 35148 17828 35154
rect 17776 35090 17828 35096
rect 17788 34746 17816 35090
rect 17776 34740 17828 34746
rect 17776 34682 17828 34688
rect 17788 34610 17816 34682
rect 17776 34604 17828 34610
rect 17776 34546 17828 34552
rect 17776 34400 17828 34406
rect 17776 34342 17828 34348
rect 17236 33106 17356 33134
rect 17040 32904 17092 32910
rect 17040 32846 17092 32852
rect 16948 31952 17000 31958
rect 16948 31894 17000 31900
rect 16960 30938 16988 31894
rect 17052 31686 17080 32846
rect 17132 32292 17184 32298
rect 17132 32234 17184 32240
rect 17040 31680 17092 31686
rect 17040 31622 17092 31628
rect 17052 31346 17080 31622
rect 17040 31340 17092 31346
rect 17040 31282 17092 31288
rect 16948 30932 17000 30938
rect 16948 30874 17000 30880
rect 17144 30870 17172 32234
rect 17224 32224 17276 32230
rect 17224 32166 17276 32172
rect 17236 31958 17264 32166
rect 17224 31952 17276 31958
rect 17224 31894 17276 31900
rect 17236 31482 17264 31894
rect 17224 31476 17276 31482
rect 17224 31418 17276 31424
rect 17132 30864 17184 30870
rect 17132 30806 17184 30812
rect 17328 30394 17356 33106
rect 17420 33106 17724 33134
rect 17420 31210 17448 33106
rect 17500 33040 17552 33046
rect 17500 32982 17552 32988
rect 17512 32570 17540 32982
rect 17684 32768 17736 32774
rect 17684 32710 17736 32716
rect 17500 32564 17552 32570
rect 17500 32506 17552 32512
rect 17696 32298 17724 32710
rect 17788 32434 17816 34342
rect 17868 33856 17920 33862
rect 17868 33798 17920 33804
rect 17776 32428 17828 32434
rect 17776 32370 17828 32376
rect 17880 32298 17908 33798
rect 17972 33658 18000 40140
rect 18432 38457 18460 40938
rect 18512 39432 18564 39438
rect 18512 39374 18564 39380
rect 18524 38554 18552 39374
rect 18512 38548 18564 38554
rect 18512 38490 18564 38496
rect 18418 38448 18474 38457
rect 18418 38383 18420 38392
rect 18472 38383 18474 38392
rect 18420 38354 18472 38360
rect 18432 38010 18460 38354
rect 18420 38004 18472 38010
rect 18420 37946 18472 37952
rect 18144 37324 18196 37330
rect 18144 37266 18196 37272
rect 18156 36582 18184 37266
rect 18420 37120 18472 37126
rect 18420 37062 18472 37068
rect 18144 36576 18196 36582
rect 18144 36518 18196 36524
rect 18328 36236 18380 36242
rect 18328 36178 18380 36184
rect 18340 35834 18368 36178
rect 18432 36038 18460 37062
rect 18420 36032 18472 36038
rect 18420 35974 18472 35980
rect 18328 35828 18380 35834
rect 18328 35770 18380 35776
rect 18052 35012 18104 35018
rect 18052 34954 18104 34960
rect 18064 34066 18092 34954
rect 18052 34060 18104 34066
rect 18052 34002 18104 34008
rect 17960 33652 18012 33658
rect 17960 33594 18012 33600
rect 17972 33454 18000 33594
rect 17960 33448 18012 33454
rect 17960 33390 18012 33396
rect 17684 32292 17736 32298
rect 17684 32234 17736 32240
rect 17868 32292 17920 32298
rect 17868 32234 17920 32240
rect 17500 31748 17552 31754
rect 17500 31690 17552 31696
rect 17408 31204 17460 31210
rect 17408 31146 17460 31152
rect 17512 30734 17540 31690
rect 17868 31204 17920 31210
rect 17868 31146 17920 31152
rect 17592 30864 17644 30870
rect 17592 30806 17644 30812
rect 17500 30728 17552 30734
rect 17500 30670 17552 30676
rect 17316 30388 17368 30394
rect 17316 30330 17368 30336
rect 17328 30190 17356 30330
rect 17316 30184 17368 30190
rect 17368 30144 17448 30172
rect 17316 30126 17368 30132
rect 17316 29844 17368 29850
rect 17316 29786 17368 29792
rect 16948 29640 17000 29646
rect 16948 29582 17000 29588
rect 16960 29170 16988 29582
rect 16948 29164 17000 29170
rect 16948 29106 17000 29112
rect 17328 29034 17356 29786
rect 17316 29028 17368 29034
rect 17316 28970 17368 28976
rect 17224 28688 17276 28694
rect 17224 28630 17276 28636
rect 17236 27946 17264 28630
rect 17224 27940 17276 27946
rect 17224 27882 17276 27888
rect 16948 27872 17000 27878
rect 16948 27814 17000 27820
rect 16960 27606 16988 27814
rect 17236 27606 17264 27882
rect 16948 27600 17000 27606
rect 16948 27542 17000 27548
rect 17224 27600 17276 27606
rect 17224 27542 17276 27548
rect 16960 26586 16988 27542
rect 17132 27464 17184 27470
rect 17132 27406 17184 27412
rect 16948 26580 17000 26586
rect 16948 26522 17000 26528
rect 17144 25906 17172 27406
rect 17236 27130 17264 27542
rect 17224 27124 17276 27130
rect 17224 27066 17276 27072
rect 17420 26081 17448 30144
rect 17512 29782 17540 30670
rect 17604 30394 17632 30806
rect 17592 30388 17644 30394
rect 17592 30330 17644 30336
rect 17604 29850 17632 30330
rect 17684 30184 17736 30190
rect 17684 30126 17736 30132
rect 17592 29844 17644 29850
rect 17592 29786 17644 29792
rect 17500 29776 17552 29782
rect 17500 29718 17552 29724
rect 17500 28960 17552 28966
rect 17500 28902 17552 28908
rect 17512 28558 17540 28902
rect 17500 28552 17552 28558
rect 17500 28494 17552 28500
rect 17592 28552 17644 28558
rect 17592 28494 17644 28500
rect 17512 28218 17540 28494
rect 17500 28212 17552 28218
rect 17500 28154 17552 28160
rect 17604 28082 17632 28494
rect 17592 28076 17644 28082
rect 17592 28018 17644 28024
rect 17696 28014 17724 30126
rect 17684 28008 17736 28014
rect 17684 27950 17736 27956
rect 17880 26790 17908 31146
rect 17972 28626 18000 33390
rect 18064 33114 18092 34002
rect 18432 33862 18460 35974
rect 18616 34746 18644 41006
rect 18786 40967 18842 40976
rect 18800 40934 18828 40967
rect 18788 40928 18840 40934
rect 18788 40870 18840 40876
rect 19076 40594 19104 41210
rect 19064 40588 19116 40594
rect 19064 40530 19116 40536
rect 19168 40526 19196 41414
rect 19444 41002 19472 41414
rect 19720 41138 19748 41414
rect 19892 41200 19944 41206
rect 19892 41142 19944 41148
rect 19708 41132 19760 41138
rect 19708 41074 19760 41080
rect 19432 40996 19484 41002
rect 19432 40938 19484 40944
rect 19444 40662 19472 40938
rect 19580 40828 19876 40848
rect 19636 40826 19660 40828
rect 19716 40826 19740 40828
rect 19796 40826 19820 40828
rect 19658 40774 19660 40826
rect 19722 40774 19734 40826
rect 19796 40774 19798 40826
rect 19636 40772 19660 40774
rect 19716 40772 19740 40774
rect 19796 40772 19820 40774
rect 19580 40752 19876 40772
rect 19432 40656 19484 40662
rect 19432 40598 19484 40604
rect 19156 40520 19208 40526
rect 19156 40462 19208 40468
rect 18788 39840 18840 39846
rect 18788 39782 18840 39788
rect 18696 39568 18748 39574
rect 18800 39545 18828 39782
rect 19168 39574 19196 40462
rect 19444 40186 19472 40598
rect 19432 40180 19484 40186
rect 19432 40122 19484 40128
rect 19444 39914 19472 40122
rect 19432 39908 19484 39914
rect 19432 39850 19484 39856
rect 19444 39642 19472 39850
rect 19580 39740 19876 39760
rect 19636 39738 19660 39740
rect 19716 39738 19740 39740
rect 19796 39738 19820 39740
rect 19658 39686 19660 39738
rect 19722 39686 19734 39738
rect 19796 39686 19798 39738
rect 19636 39684 19660 39686
rect 19716 39684 19740 39686
rect 19796 39684 19820 39686
rect 19580 39664 19876 39684
rect 19432 39636 19484 39642
rect 19432 39578 19484 39584
rect 19156 39568 19208 39574
rect 18696 39510 18748 39516
rect 18786 39536 18842 39545
rect 18708 39098 18736 39510
rect 19156 39510 19208 39516
rect 18786 39471 18842 39480
rect 19432 39364 19484 39370
rect 19432 39306 19484 39312
rect 18696 39092 18748 39098
rect 18696 39034 18748 39040
rect 18708 38826 18736 39034
rect 19248 38888 19300 38894
rect 19168 38848 19248 38876
rect 18696 38820 18748 38826
rect 18748 38780 18828 38808
rect 18696 38762 18748 38768
rect 18696 37256 18748 37262
rect 18696 37198 18748 37204
rect 18708 36786 18736 37198
rect 18800 36922 18828 38780
rect 19168 38418 19196 38848
rect 19248 38830 19300 38836
rect 19156 38412 19208 38418
rect 19156 38354 19208 38360
rect 19168 38214 19196 38354
rect 19156 38208 19208 38214
rect 19156 38150 19208 38156
rect 19168 37738 19196 38150
rect 19340 37800 19392 37806
rect 19340 37742 19392 37748
rect 19156 37732 19208 37738
rect 19156 37674 19208 37680
rect 19168 37126 19196 37674
rect 19246 37224 19302 37233
rect 19246 37159 19302 37168
rect 19260 37126 19288 37159
rect 19156 37120 19208 37126
rect 19156 37062 19208 37068
rect 19248 37120 19300 37126
rect 19352 37097 19380 37742
rect 19248 37062 19300 37068
rect 19338 37088 19394 37097
rect 19338 37023 19394 37032
rect 18788 36916 18840 36922
rect 18788 36858 18840 36864
rect 18696 36780 18748 36786
rect 18696 36722 18748 36728
rect 18800 36650 18828 36858
rect 18788 36644 18840 36650
rect 18788 36586 18840 36592
rect 18800 36310 18828 36586
rect 18788 36304 18840 36310
rect 18788 36246 18840 36252
rect 18800 35834 18828 36246
rect 18788 35828 18840 35834
rect 18788 35770 18840 35776
rect 18800 34746 18828 35770
rect 19340 35216 19392 35222
rect 19340 35158 19392 35164
rect 18604 34740 18656 34746
rect 18604 34682 18656 34688
rect 18788 34740 18840 34746
rect 18788 34682 18840 34688
rect 18616 34542 18644 34682
rect 19156 34604 19208 34610
rect 19156 34546 19208 34552
rect 18604 34536 18656 34542
rect 18604 34478 18656 34484
rect 18420 33856 18472 33862
rect 18420 33798 18472 33804
rect 18432 33454 18460 33798
rect 18328 33448 18380 33454
rect 18328 33390 18380 33396
rect 18420 33448 18472 33454
rect 18420 33390 18472 33396
rect 18052 33108 18104 33114
rect 18052 33050 18104 33056
rect 18340 32774 18368 33390
rect 18616 33134 18644 34478
rect 18880 33992 18932 33998
rect 18880 33934 18932 33940
rect 18892 33522 18920 33934
rect 18880 33516 18932 33522
rect 18880 33458 18932 33464
rect 18432 33106 18644 33134
rect 18328 32768 18380 32774
rect 18328 32710 18380 32716
rect 18144 32292 18196 32298
rect 18144 32234 18196 32240
rect 18156 30938 18184 32234
rect 18236 32020 18288 32026
rect 18236 31962 18288 31968
rect 18248 31278 18276 31962
rect 18236 31272 18288 31278
rect 18236 31214 18288 31220
rect 18144 30932 18196 30938
rect 18144 30874 18196 30880
rect 18340 30802 18368 32710
rect 18328 30796 18380 30802
rect 18328 30738 18380 30744
rect 18340 30054 18368 30738
rect 18328 30048 18380 30054
rect 18328 29990 18380 29996
rect 17960 28620 18012 28626
rect 17960 28562 18012 28568
rect 18144 28416 18196 28422
rect 18144 28358 18196 28364
rect 18156 28014 18184 28358
rect 18144 28008 18196 28014
rect 18144 27950 18196 27956
rect 18156 26790 18184 27950
rect 18236 27328 18288 27334
rect 18236 27270 18288 27276
rect 18248 26926 18276 27270
rect 18236 26920 18288 26926
rect 18236 26862 18288 26868
rect 17868 26784 17920 26790
rect 17868 26726 17920 26732
rect 18144 26784 18196 26790
rect 18144 26726 18196 26732
rect 17500 26444 17552 26450
rect 17500 26386 17552 26392
rect 17406 26072 17462 26081
rect 17406 26007 17462 26016
rect 16856 25900 16908 25906
rect 16856 25842 16908 25848
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 16868 25158 16896 25842
rect 16856 25152 16908 25158
rect 16856 25094 16908 25100
rect 16868 24410 16896 25094
rect 17144 24818 17172 25842
rect 17132 24812 17184 24818
rect 17132 24754 17184 24760
rect 16856 24404 16908 24410
rect 16856 24346 16908 24352
rect 17420 24274 17448 26007
rect 17512 25974 17540 26386
rect 17776 26308 17828 26314
rect 17776 26250 17828 26256
rect 17684 26036 17736 26042
rect 17684 25978 17736 25984
rect 17500 25968 17552 25974
rect 17500 25910 17552 25916
rect 17696 24698 17724 25978
rect 17788 25906 17816 26250
rect 17776 25900 17828 25906
rect 17776 25842 17828 25848
rect 17788 25498 17816 25842
rect 17776 25492 17828 25498
rect 17776 25434 17828 25440
rect 17880 24750 17908 26726
rect 18248 26450 18276 26862
rect 18236 26444 18288 26450
rect 18236 26386 18288 26392
rect 18052 26376 18104 26382
rect 18052 26318 18104 26324
rect 18064 25362 18092 26318
rect 18248 25702 18276 26386
rect 18236 25696 18288 25702
rect 18236 25638 18288 25644
rect 18052 25356 18104 25362
rect 18052 25298 18104 25304
rect 18064 24954 18092 25298
rect 18052 24948 18104 24954
rect 18052 24890 18104 24896
rect 18248 24886 18276 25638
rect 18236 24880 18288 24886
rect 18236 24822 18288 24828
rect 17868 24744 17920 24750
rect 17774 24712 17830 24721
rect 17696 24670 17774 24698
rect 17868 24686 17920 24692
rect 18052 24744 18104 24750
rect 18052 24686 18104 24692
rect 17774 24647 17830 24656
rect 17408 24268 17460 24274
rect 17408 24210 17460 24216
rect 17420 23866 17448 24210
rect 17408 23860 17460 23866
rect 17408 23802 17460 23808
rect 17420 23474 17448 23802
rect 17328 23446 17448 23474
rect 17224 23248 17276 23254
rect 17224 23190 17276 23196
rect 17040 23112 17092 23118
rect 17040 23054 17092 23060
rect 17052 22778 17080 23054
rect 17040 22772 17092 22778
rect 17040 22714 17092 22720
rect 17236 22506 17264 23190
rect 17328 22778 17356 23446
rect 17788 23066 17816 24647
rect 18064 24313 18092 24686
rect 18144 24608 18196 24614
rect 18144 24550 18196 24556
rect 18050 24304 18106 24313
rect 18156 24274 18184 24550
rect 18050 24239 18106 24248
rect 18144 24268 18196 24274
rect 17788 23038 17908 23066
rect 17776 22976 17828 22982
rect 17776 22918 17828 22924
rect 17316 22772 17368 22778
rect 17316 22714 17368 22720
rect 17788 22710 17816 22918
rect 17776 22704 17828 22710
rect 17776 22646 17828 22652
rect 17224 22500 17276 22506
rect 17224 22442 17276 22448
rect 17236 22166 17264 22442
rect 17788 22166 17816 22646
rect 17224 22160 17276 22166
rect 17776 22160 17828 22166
rect 17224 22102 17276 22108
rect 17314 22128 17370 22137
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17144 21690 17172 21966
rect 17236 21690 17264 22102
rect 17776 22102 17828 22108
rect 17314 22063 17370 22072
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 17224 21684 17276 21690
rect 17224 21626 17276 21632
rect 17144 21146 17172 21626
rect 17328 21622 17356 22063
rect 17592 21684 17644 21690
rect 17592 21626 17644 21632
rect 17316 21616 17368 21622
rect 17316 21558 17368 21564
rect 17132 21140 17184 21146
rect 17132 21082 17184 21088
rect 17604 21078 17632 21626
rect 17592 21072 17644 21078
rect 17592 21014 17644 21020
rect 16948 20936 17000 20942
rect 16948 20878 17000 20884
rect 17500 20936 17552 20942
rect 17500 20878 17552 20884
rect 16960 20602 16988 20878
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 16960 20058 16988 20538
rect 17512 20058 17540 20878
rect 17604 20602 17632 21014
rect 17592 20596 17644 20602
rect 17592 20538 17644 20544
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 16776 19514 16804 19858
rect 16948 19712 17000 19718
rect 16948 19654 17000 19660
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 16960 19310 16988 19654
rect 17512 19514 17540 19994
rect 17880 19904 17908 23038
rect 17960 19916 18012 19922
rect 17880 19876 17960 19904
rect 17960 19858 18012 19864
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17500 19508 17552 19514
rect 17500 19450 17552 19456
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 17040 19236 17092 19242
rect 17040 19178 17092 19184
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 16488 18624 16540 18630
rect 16488 18566 16540 18572
rect 16500 18290 16528 18566
rect 16488 18284 16540 18290
rect 16488 18226 16540 18232
rect 16500 17882 16528 18226
rect 16592 18154 16620 18702
rect 16764 18692 16816 18698
rect 16764 18634 16816 18640
rect 16580 18148 16632 18154
rect 16580 18090 16632 18096
rect 16488 17876 16540 17882
rect 16488 17818 16540 17824
rect 16592 16726 16620 18090
rect 16580 16720 16632 16726
rect 16580 16662 16632 16668
rect 16488 15972 16540 15978
rect 16488 15914 16540 15920
rect 16500 15434 16528 15914
rect 16488 15428 16540 15434
rect 16488 15370 16540 15376
rect 16408 15286 16528 15314
rect 16028 15156 16080 15162
rect 16028 15098 16080 15104
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 15844 14952 15896 14958
rect 15844 14894 15896 14900
rect 15660 14544 15712 14550
rect 15660 14486 15712 14492
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 14740 14340 14792 14346
rect 14740 14282 14792 14288
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 14844 13530 14872 13874
rect 15672 13530 15700 14486
rect 15764 14074 15792 14486
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 15028 11762 15056 12582
rect 15212 12306 15240 13330
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15396 12442 15424 12718
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 15028 11354 15056 11698
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 15396 11150 15424 12378
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15764 11082 15792 12650
rect 15856 11898 15884 14894
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15948 14006 15976 14350
rect 16040 14006 16068 15098
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 15936 14000 15988 14006
rect 15936 13942 15988 13948
rect 16028 14000 16080 14006
rect 16028 13942 16080 13948
rect 16224 13938 16252 14758
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 16408 13802 16436 14214
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16224 13462 16252 13738
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 16132 12986 16160 13262
rect 16224 12986 16252 13398
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16212 12980 16264 12986
rect 16212 12922 16264 12928
rect 16212 12368 16264 12374
rect 16212 12310 16264 12316
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16040 11898 16068 12174
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 16040 11354 16068 11834
rect 16224 11830 16252 12310
rect 16408 11830 16436 13738
rect 16500 13172 16528 15286
rect 16592 14550 16620 16662
rect 16580 14544 16632 14550
rect 16580 14486 16632 14492
rect 16592 13802 16620 14486
rect 16580 13796 16632 13802
rect 16580 13738 16632 13744
rect 16580 13184 16632 13190
rect 16500 13144 16580 13172
rect 16580 13126 16632 13132
rect 16592 12714 16620 13126
rect 16580 12708 16632 12714
rect 16580 12650 16632 12656
rect 16212 11824 16264 11830
rect 16212 11766 16264 11772
rect 16396 11824 16448 11830
rect 16396 11766 16448 11772
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 15752 11076 15804 11082
rect 15752 11018 15804 11024
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 14556 10192 14608 10198
rect 14556 10134 14608 10140
rect 15212 10062 15240 10406
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15212 9722 15240 9998
rect 15580 9994 15608 10610
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15568 9988 15620 9994
rect 15568 9930 15620 9936
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 15108 9376 15160 9382
rect 15108 9318 15160 9324
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15120 8498 15148 9318
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15488 8294 15516 9318
rect 15580 8838 15608 9930
rect 15672 9926 15700 10542
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 15672 9654 15700 9862
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15672 9042 15700 9590
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15672 8566 15700 8978
rect 15660 8560 15712 8566
rect 15660 8502 15712 8508
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15476 7540 15528 7546
rect 15580 7528 15608 7686
rect 15764 7546 15792 11018
rect 16224 11014 16252 11154
rect 16212 11008 16264 11014
rect 16212 10950 16264 10956
rect 16120 10192 16172 10198
rect 16120 10134 16172 10140
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 15936 9648 15988 9654
rect 15856 9608 15936 9636
rect 15856 9042 15884 9608
rect 15936 9590 15988 9596
rect 16040 9586 16068 9998
rect 16132 9654 16160 10134
rect 16120 9648 16172 9654
rect 16120 9590 16172 9596
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15844 9036 15896 9042
rect 15844 8978 15896 8984
rect 15856 8498 15884 8978
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15528 7500 15608 7528
rect 15476 7482 15528 7488
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13648 6186 13676 6802
rect 14752 6458 14780 7414
rect 15580 7002 15608 7500
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15856 7342 15884 7890
rect 15948 7818 15976 9318
rect 16592 8974 16620 12650
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 15936 7812 15988 7818
rect 15936 7754 15988 7760
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 15752 7268 15804 7274
rect 15752 7210 15804 7216
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 15384 6384 15436 6390
rect 15384 6326 15436 6332
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13648 4622 13676 6122
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 14108 4758 14136 4966
rect 14096 4752 14148 4758
rect 14096 4694 14148 4700
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 9968 2922 9996 3334
rect 11532 3194 11560 3334
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11900 3058 11928 3470
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 9956 2916 10008 2922
rect 9956 2858 10008 2864
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 5632 2304 5684 2310
rect 5632 2246 5684 2252
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 1766 82 1822 480
rect 1688 54 1822 82
rect 1766 0 1822 54
rect 5262 82 5318 480
rect 5644 82 5672 2246
rect 5262 54 5672 82
rect 8850 82 8906 480
rect 9048 82 9076 2790
rect 9968 2650 9996 2858
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 10888 2310 10916 2926
rect 11900 2854 11928 2994
rect 11980 2916 12032 2922
rect 11980 2858 12032 2864
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 11992 2650 12020 2858
rect 12452 2650 12480 3470
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 11072 2310 11100 2450
rect 11440 2310 11468 2450
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11428 2304 11480 2310
rect 11428 2246 11480 2252
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11072 1737 11100 2246
rect 11440 2145 11468 2246
rect 11426 2136 11482 2145
rect 11426 2071 11482 2080
rect 11900 1873 11928 2246
rect 11886 1864 11942 1873
rect 11886 1799 11942 1808
rect 11058 1728 11114 1737
rect 11058 1663 11114 1672
rect 8850 54 9076 82
rect 12438 82 12494 480
rect 12636 82 12664 4014
rect 13372 3466 13400 4558
rect 13648 4214 13676 4558
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 13636 4208 13688 4214
rect 13636 4150 13688 4156
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13360 3460 13412 3466
rect 13360 3402 13412 3408
rect 13372 3194 13400 3402
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13648 3058 13676 3878
rect 13740 3602 13768 4422
rect 14384 4282 14412 6054
rect 15396 5370 15424 6326
rect 15764 6254 15792 7210
rect 16040 6798 16068 8774
rect 16212 8560 16264 8566
rect 16212 8502 16264 8508
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16132 7750 16160 8230
rect 16224 7886 16252 8502
rect 16684 8498 16712 9454
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16120 7744 16172 7750
rect 16120 7686 16172 7692
rect 16132 7274 16160 7686
rect 16120 7268 16172 7274
rect 16120 7210 16172 7216
rect 16224 7002 16252 7822
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 16488 6928 16540 6934
rect 16488 6870 16540 6876
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 15752 6248 15804 6254
rect 15752 6190 15804 6196
rect 16500 6118 16528 6870
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 16592 6322 16620 6734
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15396 5166 15424 5306
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15016 5092 15068 5098
rect 15016 5034 15068 5040
rect 15028 4758 15056 5034
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 15016 4752 15068 4758
rect 15016 4694 15068 4700
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 15120 4185 15148 4422
rect 14186 4176 14242 4185
rect 14186 4111 14188 4120
rect 14240 4111 14242 4120
rect 15106 4176 15162 4185
rect 15106 4111 15162 4120
rect 14188 4082 14240 4088
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 14556 4004 14608 4010
rect 14556 3946 14608 3952
rect 14568 3738 14596 3946
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13740 3194 13768 3538
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12728 2514 12756 2926
rect 12912 2650 12940 2926
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 13740 2514 13768 3130
rect 14200 2650 14228 3334
rect 14292 2990 14320 3334
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14292 2650 14320 2926
rect 14568 2922 14596 3674
rect 15488 3194 15516 4014
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 14556 2916 14608 2922
rect 14556 2858 14608 2864
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 15580 2514 15608 3402
rect 15672 2650 15700 4966
rect 15764 4826 15792 5714
rect 16132 5166 16160 5714
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 16132 4826 16160 5102
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 16120 4820 16172 4826
rect 16120 4762 16172 4768
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15660 2644 15712 2650
rect 15660 2586 15712 2592
rect 15672 2514 15700 2586
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15660 2508 15712 2514
rect 15660 2450 15712 2456
rect 12438 54 12664 82
rect 15764 82 15792 4218
rect 16040 3738 16068 4626
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 16132 2990 16160 3878
rect 16224 3534 16252 5646
rect 16500 5234 16528 6054
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16500 4758 16528 5170
rect 16488 4752 16540 4758
rect 16488 4694 16540 4700
rect 16500 4282 16528 4694
rect 16488 4276 16540 4282
rect 16488 4218 16540 4224
rect 16500 3738 16528 4218
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 16500 3126 16528 3674
rect 16592 3194 16620 3878
rect 16776 3618 16804 18634
rect 17052 17814 17080 19178
rect 17420 18834 17448 19450
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 17408 18828 17460 18834
rect 17408 18770 17460 18776
rect 17236 18426 17264 18770
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17420 18358 17448 18770
rect 17788 18737 17816 19110
rect 17774 18728 17830 18737
rect 17972 18698 18000 19858
rect 17774 18663 17830 18672
rect 17960 18692 18012 18698
rect 17960 18634 18012 18640
rect 17408 18352 17460 18358
rect 18064 18306 18092 24239
rect 18144 24210 18196 24216
rect 18156 23866 18184 24210
rect 18340 24120 18368 29990
rect 18432 29306 18460 33106
rect 19064 32972 19116 32978
rect 19064 32914 19116 32920
rect 18788 32428 18840 32434
rect 18788 32370 18840 32376
rect 18694 30968 18750 30977
rect 18694 30903 18750 30912
rect 18512 30116 18564 30122
rect 18512 30058 18564 30064
rect 18420 29300 18472 29306
rect 18420 29242 18472 29248
rect 18432 29102 18460 29242
rect 18420 29096 18472 29102
rect 18420 29038 18472 29044
rect 18524 29034 18552 30058
rect 18708 29170 18736 30903
rect 18800 29646 18828 32370
rect 18880 32360 18932 32366
rect 18880 32302 18932 32308
rect 18892 32026 18920 32302
rect 19076 32230 19104 32914
rect 19064 32224 19116 32230
rect 19064 32166 19116 32172
rect 18880 32020 18932 32026
rect 18880 31962 18932 31968
rect 18972 31136 19024 31142
rect 19076 31113 19104 32166
rect 19168 31482 19196 34546
rect 19248 34468 19300 34474
rect 19248 34410 19300 34416
rect 19260 34202 19288 34410
rect 19352 34406 19380 35158
rect 19444 35086 19472 39306
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19580 38576 19876 38596
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 19706 37360 19762 37369
rect 19706 37295 19762 37304
rect 19720 37262 19748 37295
rect 19708 37256 19760 37262
rect 19708 37198 19760 37204
rect 19720 36922 19748 37198
rect 19708 36916 19760 36922
rect 19708 36858 19760 36864
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 19904 36310 19932 41142
rect 19984 39908 20036 39914
rect 19984 39850 20036 39856
rect 19996 39370 20024 39850
rect 19984 39364 20036 39370
rect 19984 39306 20036 39312
rect 19984 38752 20036 38758
rect 19984 38694 20036 38700
rect 19996 38214 20024 38694
rect 19984 38208 20036 38214
rect 19984 38150 20036 38156
rect 19892 36304 19944 36310
rect 19892 36246 19944 36252
rect 19524 36032 19576 36038
rect 19524 35974 19576 35980
rect 19536 35834 19564 35974
rect 19904 35834 19932 36246
rect 19524 35828 19576 35834
rect 19524 35770 19576 35776
rect 19892 35828 19944 35834
rect 19892 35770 19944 35776
rect 19536 35544 19564 35770
rect 19892 35692 19944 35698
rect 19892 35634 19944 35640
rect 19708 35556 19760 35562
rect 19536 35516 19708 35544
rect 19708 35498 19760 35504
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 19432 35080 19484 35086
rect 19432 35022 19484 35028
rect 19444 34610 19472 35022
rect 19904 35018 19932 35634
rect 19892 35012 19944 35018
rect 19892 34954 19944 34960
rect 19432 34604 19484 34610
rect 19432 34546 19484 34552
rect 20076 34536 20128 34542
rect 20076 34478 20128 34484
rect 19432 34468 19484 34474
rect 19432 34410 19484 34416
rect 19340 34400 19392 34406
rect 19340 34342 19392 34348
rect 19352 34202 19380 34342
rect 19248 34196 19300 34202
rect 19248 34138 19300 34144
rect 19340 34196 19392 34202
rect 19340 34138 19392 34144
rect 19444 33658 19472 34410
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 20088 34202 20116 34478
rect 20076 34196 20128 34202
rect 20076 34138 20128 34144
rect 19432 33652 19484 33658
rect 19432 33594 19484 33600
rect 19248 33380 19300 33386
rect 19248 33322 19300 33328
rect 19260 33046 19288 33322
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 20088 33046 20116 34138
rect 19248 33040 19300 33046
rect 19248 32982 19300 32988
rect 20076 33040 20128 33046
rect 20076 32982 20128 32988
rect 19892 32428 19944 32434
rect 19892 32370 19944 32376
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19340 31884 19392 31890
rect 19340 31826 19392 31832
rect 19156 31476 19208 31482
rect 19156 31418 19208 31424
rect 19156 31204 19208 31210
rect 19156 31146 19208 31152
rect 18972 31078 19024 31084
rect 19062 31104 19118 31113
rect 18984 30802 19012 31078
rect 19062 31039 19118 31048
rect 19064 30932 19116 30938
rect 19064 30874 19116 30880
rect 18972 30796 19024 30802
rect 18972 30738 19024 30744
rect 18972 30660 19024 30666
rect 18972 30602 19024 30608
rect 18880 30048 18932 30054
rect 18880 29990 18932 29996
rect 18892 29782 18920 29990
rect 18880 29776 18932 29782
rect 18880 29718 18932 29724
rect 18788 29640 18840 29646
rect 18788 29582 18840 29588
rect 18800 29238 18828 29582
rect 18892 29306 18920 29718
rect 18984 29646 19012 30602
rect 19076 30258 19104 30874
rect 19064 30252 19116 30258
rect 19064 30194 19116 30200
rect 19076 29850 19104 30194
rect 19064 29844 19116 29850
rect 19064 29786 19116 29792
rect 18972 29640 19024 29646
rect 18972 29582 19024 29588
rect 19168 29306 19196 31146
rect 19352 30784 19380 31826
rect 19616 31816 19668 31822
rect 19616 31758 19668 31764
rect 19432 31680 19484 31686
rect 19432 31622 19484 31628
rect 19444 31278 19472 31622
rect 19628 31414 19656 31758
rect 19904 31754 19932 32370
rect 20272 32366 20300 49506
rect 21824 42764 21876 42770
rect 21824 42706 21876 42712
rect 21640 42560 21692 42566
rect 21640 42502 21692 42508
rect 21652 41614 21680 42502
rect 21836 42022 21864 42706
rect 21732 42016 21784 42022
rect 21732 41958 21784 41964
rect 21824 42016 21876 42022
rect 21824 41958 21876 41964
rect 21640 41608 21692 41614
rect 21640 41550 21692 41556
rect 21652 41274 21680 41550
rect 21640 41268 21692 41274
rect 21640 41210 21692 41216
rect 21744 40662 21772 41958
rect 21732 40656 21784 40662
rect 21732 40598 21784 40604
rect 20536 40520 20588 40526
rect 20536 40462 20588 40468
rect 20444 38888 20496 38894
rect 20444 38830 20496 38836
rect 20456 38554 20484 38830
rect 20444 38548 20496 38554
rect 20444 38490 20496 38496
rect 20548 36786 20576 40462
rect 21744 40186 21772 40598
rect 21732 40180 21784 40186
rect 21732 40122 21784 40128
rect 21836 39522 21864 41958
rect 21916 41744 21968 41750
rect 21916 41686 21968 41692
rect 21928 41002 21956 41686
rect 24228 41682 24256 49506
rect 24964 49475 24992 49506
rect 24308 42152 24360 42158
rect 24308 42094 24360 42100
rect 24860 42152 24912 42158
rect 24860 42094 24912 42100
rect 24216 41676 24268 41682
rect 24216 41618 24268 41624
rect 22284 41608 22336 41614
rect 22284 41550 22336 41556
rect 22296 41206 22324 41550
rect 23204 41540 23256 41546
rect 23204 41482 23256 41488
rect 22284 41200 22336 41206
rect 22284 41142 22336 41148
rect 21916 40996 21968 41002
rect 21916 40938 21968 40944
rect 22100 40996 22152 41002
rect 22100 40938 22152 40944
rect 21744 39494 21864 39522
rect 20628 38820 20680 38826
rect 20628 38762 20680 38768
rect 20640 38010 20668 38762
rect 20628 38004 20680 38010
rect 20680 37964 20760 37992
rect 20628 37946 20680 37952
rect 20628 37800 20680 37806
rect 20628 37742 20680 37748
rect 20640 37466 20668 37742
rect 20732 37738 20760 37964
rect 20720 37732 20772 37738
rect 20720 37674 20772 37680
rect 20628 37460 20680 37466
rect 20628 37402 20680 37408
rect 21744 37126 21772 39494
rect 21824 39432 21876 39438
rect 21824 39374 21876 39380
rect 21836 39098 21864 39374
rect 21824 39092 21876 39098
rect 21824 39034 21876 39040
rect 21824 38480 21876 38486
rect 21928 38468 21956 40938
rect 22008 40656 22060 40662
rect 22008 40598 22060 40604
rect 22020 39846 22048 40598
rect 22112 40526 22140 40938
rect 22100 40520 22152 40526
rect 22100 40462 22152 40468
rect 22296 40118 22324 41142
rect 23020 40928 23072 40934
rect 23020 40870 23072 40876
rect 22744 40384 22796 40390
rect 22744 40326 22796 40332
rect 22756 40186 22784 40326
rect 22744 40180 22796 40186
rect 22744 40122 22796 40128
rect 22284 40112 22336 40118
rect 22284 40054 22336 40060
rect 22008 39840 22060 39846
rect 22008 39782 22060 39788
rect 22020 39574 22048 39782
rect 22008 39568 22060 39574
rect 22008 39510 22060 39516
rect 22020 38826 22048 39510
rect 22284 39364 22336 39370
rect 22284 39306 22336 39312
rect 22008 38820 22060 38826
rect 22008 38762 22060 38768
rect 21876 38440 21956 38468
rect 21824 38422 21876 38428
rect 21836 37670 21864 38422
rect 22296 38350 22324 39306
rect 22650 39264 22706 39273
rect 22650 39199 22706 39208
rect 22664 38894 22692 39199
rect 22652 38888 22704 38894
rect 22652 38830 22704 38836
rect 22192 38344 22244 38350
rect 22192 38286 22244 38292
rect 22284 38344 22336 38350
rect 22284 38286 22336 38292
rect 22204 38010 22232 38286
rect 22192 38004 22244 38010
rect 22192 37946 22244 37952
rect 22560 37800 22612 37806
rect 22560 37742 22612 37748
rect 21824 37664 21876 37670
rect 21824 37606 21876 37612
rect 21836 37398 21864 37606
rect 21824 37392 21876 37398
rect 21824 37334 21876 37340
rect 21732 37120 21784 37126
rect 21732 37062 21784 37068
rect 21836 36922 21864 37334
rect 21824 36916 21876 36922
rect 21824 36858 21876 36864
rect 22572 36786 22600 37742
rect 20536 36780 20588 36786
rect 20536 36722 20588 36728
rect 22560 36780 22612 36786
rect 22560 36722 22612 36728
rect 20548 36378 20576 36722
rect 21732 36712 21784 36718
rect 21732 36654 21784 36660
rect 21180 36644 21232 36650
rect 21180 36586 21232 36592
rect 20536 36372 20588 36378
rect 20536 36314 20588 36320
rect 20996 36168 21048 36174
rect 20996 36110 21048 36116
rect 21008 35834 21036 36110
rect 20996 35828 21048 35834
rect 20996 35770 21048 35776
rect 21088 35216 21140 35222
rect 21088 35158 21140 35164
rect 20996 35080 21048 35086
rect 20996 35022 21048 35028
rect 21008 34202 21036 35022
rect 21100 34746 21128 35158
rect 21192 35018 21220 36586
rect 21744 36281 21772 36654
rect 21916 36576 21968 36582
rect 21916 36518 21968 36524
rect 21730 36272 21786 36281
rect 21730 36207 21732 36216
rect 21784 36207 21786 36216
rect 21732 36178 21784 36184
rect 21744 36147 21772 36178
rect 21928 36174 21956 36518
rect 22100 36304 22152 36310
rect 22100 36246 22152 36252
rect 21916 36168 21968 36174
rect 21916 36110 21968 36116
rect 22008 35692 22060 35698
rect 22008 35634 22060 35640
rect 22020 35290 22048 35634
rect 22112 35562 22140 36246
rect 22100 35556 22152 35562
rect 22100 35498 22152 35504
rect 22008 35284 22060 35290
rect 22008 35226 22060 35232
rect 22112 35222 22140 35498
rect 22376 35488 22428 35494
rect 22376 35430 22428 35436
rect 22100 35216 22152 35222
rect 22100 35158 22152 35164
rect 21180 35012 21232 35018
rect 21180 34954 21232 34960
rect 21088 34740 21140 34746
rect 21088 34682 21140 34688
rect 21086 34504 21142 34513
rect 22112 34474 22140 35158
rect 22388 35086 22416 35430
rect 22376 35080 22428 35086
rect 22376 35022 22428 35028
rect 22388 34746 22416 35022
rect 22376 34740 22428 34746
rect 22376 34682 22428 34688
rect 21086 34439 21142 34448
rect 22008 34468 22060 34474
rect 20996 34196 21048 34202
rect 20996 34138 21048 34144
rect 20352 33652 20404 33658
rect 20352 33594 20404 33600
rect 20364 33046 20392 33594
rect 20352 33040 20404 33046
rect 20352 32982 20404 32988
rect 20364 32570 20392 32982
rect 20352 32564 20404 32570
rect 20352 32506 20404 32512
rect 20996 32428 21048 32434
rect 20996 32370 21048 32376
rect 20260 32360 20312 32366
rect 20260 32302 20312 32308
rect 21008 32230 21036 32370
rect 19984 32224 20036 32230
rect 19984 32166 20036 32172
rect 20996 32224 21048 32230
rect 20996 32166 21048 32172
rect 19892 31748 19944 31754
rect 19812 31708 19892 31736
rect 19812 31414 19840 31708
rect 19892 31690 19944 31696
rect 19616 31408 19668 31414
rect 19616 31350 19668 31356
rect 19800 31408 19852 31414
rect 19852 31368 19932 31396
rect 19800 31350 19852 31356
rect 19432 31272 19484 31278
rect 19432 31214 19484 31220
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 19904 30802 19932 31368
rect 19996 30977 20024 32166
rect 20076 32020 20128 32026
rect 20076 31962 20128 31968
rect 19982 30968 20038 30977
rect 19982 30903 20038 30912
rect 19432 30796 19484 30802
rect 19352 30756 19432 30784
rect 19432 30738 19484 30744
rect 19892 30796 19944 30802
rect 19892 30738 19944 30744
rect 19444 30394 19472 30738
rect 19432 30388 19484 30394
rect 19432 30330 19484 30336
rect 19892 30184 19944 30190
rect 19892 30126 19944 30132
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 18880 29300 18932 29306
rect 18880 29242 18932 29248
rect 19156 29300 19208 29306
rect 19156 29242 19208 29248
rect 18788 29232 18840 29238
rect 18788 29174 18840 29180
rect 18696 29164 18748 29170
rect 18696 29106 18748 29112
rect 18512 29028 18564 29034
rect 18512 28970 18564 28976
rect 18524 27878 18552 28970
rect 18602 28656 18658 28665
rect 18602 28591 18604 28600
rect 18656 28591 18658 28600
rect 18604 28562 18656 28568
rect 18616 27946 18644 28562
rect 18696 28416 18748 28422
rect 18696 28358 18748 28364
rect 18604 27940 18656 27946
rect 18604 27882 18656 27888
rect 18512 27872 18564 27878
rect 18512 27814 18564 27820
rect 18512 25424 18564 25430
rect 18512 25366 18564 25372
rect 18524 24818 18552 25366
rect 18512 24812 18564 24818
rect 18512 24754 18564 24760
rect 18524 24342 18552 24754
rect 18512 24336 18564 24342
rect 18512 24278 18564 24284
rect 18420 24132 18472 24138
rect 18340 24092 18420 24120
rect 18420 24074 18472 24080
rect 18144 23860 18196 23866
rect 18144 23802 18196 23808
rect 18432 23769 18460 24074
rect 18524 23866 18552 24278
rect 18512 23860 18564 23866
rect 18512 23802 18564 23808
rect 18418 23760 18474 23769
rect 18144 23724 18196 23730
rect 18418 23695 18474 23704
rect 18144 23666 18196 23672
rect 18156 22953 18184 23666
rect 18142 22944 18198 22953
rect 18142 22879 18198 22888
rect 18156 21350 18184 22879
rect 18236 21412 18288 21418
rect 18236 21354 18288 21360
rect 18144 21344 18196 21350
rect 18144 21286 18196 21292
rect 18248 21162 18276 21354
rect 17408 18294 17460 18300
rect 17696 18278 18092 18306
rect 18156 21134 18276 21162
rect 17132 18148 17184 18154
rect 17132 18090 17184 18096
rect 17040 17808 17092 17814
rect 17040 17750 17092 17756
rect 17052 16998 17080 17750
rect 17144 17610 17172 18090
rect 17408 17672 17460 17678
rect 17408 17614 17460 17620
rect 17132 17604 17184 17610
rect 17132 17546 17184 17552
rect 17420 17338 17448 17614
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16960 16114 16988 16526
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16960 15706 16988 16050
rect 17052 15910 17080 16934
rect 17408 16720 17460 16726
rect 17408 16662 17460 16668
rect 17132 16584 17184 16590
rect 17132 16526 17184 16532
rect 17144 16114 17172 16526
rect 17420 16250 17448 16662
rect 17408 16244 17460 16250
rect 17408 16186 17460 16192
rect 17132 16108 17184 16114
rect 17132 16050 17184 16056
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 16868 13326 16896 14214
rect 17052 13462 17080 15846
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 17236 14822 17264 15506
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 17512 14822 17540 15438
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17500 14816 17552 14822
rect 17500 14758 17552 14764
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 17040 13456 17092 13462
rect 17040 13398 17092 13404
rect 17144 13326 17172 13874
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17236 12442 17264 14758
rect 17512 14618 17540 14758
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17604 13734 17632 14350
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 16960 11898 16988 12038
rect 16948 11892 17000 11898
rect 16948 11834 17000 11840
rect 16960 11694 16988 11834
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17144 10742 17172 10950
rect 16856 10736 16908 10742
rect 16856 10678 16908 10684
rect 17132 10736 17184 10742
rect 17132 10678 17184 10684
rect 16868 6390 16896 10678
rect 17144 8022 17172 10678
rect 17132 8016 17184 8022
rect 17132 7958 17184 7964
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16960 7342 16988 7686
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 16960 6730 16988 7278
rect 16948 6724 17000 6730
rect 16948 6666 17000 6672
rect 16856 6384 16908 6390
rect 16856 6326 16908 6332
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16868 5370 16896 5646
rect 16960 5642 16988 6666
rect 16948 5636 17000 5642
rect 16948 5578 17000 5584
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16868 4282 16896 5306
rect 17236 5273 17264 12038
rect 17420 11150 17448 13670
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17420 10742 17448 11086
rect 17408 10736 17460 10742
rect 17408 10678 17460 10684
rect 17512 10130 17540 12582
rect 17696 11286 17724 18278
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17880 17678 17908 18022
rect 17972 17746 18000 18158
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 17868 17672 17920 17678
rect 18156 17626 18184 21134
rect 18432 20058 18460 23695
rect 18616 22098 18644 27882
rect 18708 27606 18736 28358
rect 18788 27872 18840 27878
rect 18788 27814 18840 27820
rect 18800 27606 18828 27814
rect 18696 27600 18748 27606
rect 18696 27542 18748 27548
rect 18788 27600 18840 27606
rect 18788 27542 18840 27548
rect 18800 27130 18828 27542
rect 18880 27464 18932 27470
rect 18880 27406 18932 27412
rect 18788 27124 18840 27130
rect 18788 27066 18840 27072
rect 18800 26586 18828 27066
rect 18788 26580 18840 26586
rect 18788 26522 18840 26528
rect 18892 25906 18920 27406
rect 19168 27130 19196 29242
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19708 28416 19760 28422
rect 19708 28358 19760 28364
rect 19720 28150 19748 28358
rect 19708 28144 19760 28150
rect 19708 28086 19760 28092
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 19156 27124 19208 27130
rect 19156 27066 19208 27072
rect 19168 26382 19196 27066
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19524 26444 19576 26450
rect 19444 26404 19524 26432
rect 19156 26376 19208 26382
rect 19156 26318 19208 26324
rect 18972 26240 19024 26246
rect 18972 26182 19024 26188
rect 18880 25900 18932 25906
rect 18880 25842 18932 25848
rect 18984 25770 19012 26182
rect 18972 25764 19024 25770
rect 18972 25706 19024 25712
rect 19064 25764 19116 25770
rect 19064 25706 19116 25712
rect 18984 25498 19012 25706
rect 18972 25492 19024 25498
rect 18972 25434 19024 25440
rect 19076 24682 19104 25706
rect 19168 25498 19196 26318
rect 19248 25968 19300 25974
rect 19248 25910 19300 25916
rect 19156 25492 19208 25498
rect 19156 25434 19208 25440
rect 19064 24676 19116 24682
rect 19064 24618 19116 24624
rect 18788 24132 18840 24138
rect 18788 24074 18840 24080
rect 18800 23322 18828 24074
rect 18880 24064 18932 24070
rect 18880 24006 18932 24012
rect 19156 24064 19208 24070
rect 19156 24006 19208 24012
rect 18892 23866 18920 24006
rect 18880 23860 18932 23866
rect 18880 23802 18932 23808
rect 18892 23594 18920 23802
rect 19168 23730 19196 24006
rect 19156 23724 19208 23730
rect 19156 23666 19208 23672
rect 18880 23588 18932 23594
rect 18880 23530 18932 23536
rect 18788 23316 18840 23322
rect 18788 23258 18840 23264
rect 18800 22642 18828 23258
rect 18892 23236 18920 23530
rect 19064 23248 19116 23254
rect 18892 23208 19064 23236
rect 18788 22636 18840 22642
rect 18788 22578 18840 22584
rect 18786 22536 18842 22545
rect 18892 22506 18920 23208
rect 19064 23190 19116 23196
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 18786 22471 18842 22480
rect 18880 22500 18932 22506
rect 18604 22092 18656 22098
rect 18604 22034 18656 22040
rect 18616 21690 18644 22034
rect 18604 21684 18656 21690
rect 18604 21626 18656 21632
rect 18800 21486 18828 22471
rect 18880 22442 18932 22448
rect 18984 22234 19012 23054
rect 19064 22636 19116 22642
rect 19064 22578 19116 22584
rect 18972 22228 19024 22234
rect 18972 22170 19024 22176
rect 19076 22030 19104 22578
rect 19168 22166 19196 23666
rect 19260 23322 19288 25910
rect 19444 25430 19472 26404
rect 19524 26386 19576 26392
rect 19616 26376 19668 26382
rect 19616 26318 19668 26324
rect 19628 26042 19656 26318
rect 19616 26036 19668 26042
rect 19616 25978 19668 25984
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19432 25424 19484 25430
rect 19432 25366 19484 25372
rect 19340 25152 19392 25158
rect 19340 25094 19392 25100
rect 19352 24614 19380 25094
rect 19340 24608 19392 24614
rect 19340 24550 19392 24556
rect 19248 23316 19300 23322
rect 19248 23258 19300 23264
rect 19246 22808 19302 22817
rect 19246 22743 19302 22752
rect 19156 22160 19208 22166
rect 19156 22102 19208 22108
rect 19064 22024 19116 22030
rect 19260 22012 19288 22743
rect 19352 22658 19380 24550
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 19904 24274 19932 30126
rect 19984 29164 20036 29170
rect 19984 29106 20036 29112
rect 19996 26382 20024 29106
rect 20088 26926 20116 31962
rect 20812 31884 20864 31890
rect 20812 31826 20864 31832
rect 20352 31680 20404 31686
rect 20352 31622 20404 31628
rect 20364 31210 20392 31622
rect 20824 31521 20852 31826
rect 21008 31822 21036 32166
rect 20996 31816 21048 31822
rect 20996 31758 21048 31764
rect 20810 31512 20866 31521
rect 20810 31447 20866 31456
rect 20824 31414 20852 31447
rect 21008 31414 21036 31758
rect 20812 31408 20864 31414
rect 20812 31350 20864 31356
rect 20996 31408 21048 31414
rect 20996 31350 21048 31356
rect 20444 31272 20496 31278
rect 20904 31272 20956 31278
rect 20444 31214 20496 31220
rect 20626 31240 20682 31249
rect 20352 31204 20404 31210
rect 20352 31146 20404 31152
rect 20364 30666 20392 31146
rect 20456 30938 20484 31214
rect 20904 31214 20956 31220
rect 20626 31175 20682 31184
rect 20444 30932 20496 30938
rect 20444 30874 20496 30880
rect 20640 30802 20668 31175
rect 20628 30796 20680 30802
rect 20628 30738 20680 30744
rect 20352 30660 20404 30666
rect 20352 30602 20404 30608
rect 20364 29034 20392 30602
rect 20640 30394 20668 30738
rect 20628 30388 20680 30394
rect 20628 30330 20680 30336
rect 20444 29504 20496 29510
rect 20444 29446 20496 29452
rect 20456 29238 20484 29446
rect 20444 29232 20496 29238
rect 20916 29209 20944 31214
rect 21100 29714 21128 34439
rect 22008 34410 22060 34416
rect 22100 34468 22152 34474
rect 22100 34410 22152 34416
rect 21824 34196 21876 34202
rect 21824 34138 21876 34144
rect 21456 33992 21508 33998
rect 21456 33934 21508 33940
rect 21468 33522 21496 33934
rect 21836 33658 21864 34138
rect 22020 33658 22048 34410
rect 22112 34202 22140 34410
rect 22100 34196 22152 34202
rect 22100 34138 22152 34144
rect 22192 33924 22244 33930
rect 22192 33866 22244 33872
rect 21824 33652 21876 33658
rect 21824 33594 21876 33600
rect 22008 33652 22060 33658
rect 22008 33594 22060 33600
rect 21456 33516 21508 33522
rect 21456 33458 21508 33464
rect 21180 33448 21232 33454
rect 21180 33390 21232 33396
rect 21732 33448 21784 33454
rect 21732 33390 21784 33396
rect 21192 30802 21220 33390
rect 21548 32768 21600 32774
rect 21548 32710 21600 32716
rect 21560 32502 21588 32710
rect 21744 32570 21772 33390
rect 21732 32564 21784 32570
rect 21732 32506 21784 32512
rect 21548 32496 21600 32502
rect 21548 32438 21600 32444
rect 21364 32224 21416 32230
rect 21364 32166 21416 32172
rect 21376 31686 21404 32166
rect 21560 31958 21588 32438
rect 21732 32360 21784 32366
rect 21732 32302 21784 32308
rect 21548 31952 21600 31958
rect 21548 31894 21600 31900
rect 21364 31680 21416 31686
rect 21364 31622 21416 31628
rect 21744 31482 21772 32302
rect 22204 31890 22232 33866
rect 22284 32972 22336 32978
rect 22284 32914 22336 32920
rect 22468 32972 22520 32978
rect 22468 32914 22520 32920
rect 22296 32337 22324 32914
rect 22480 32570 22508 32914
rect 22468 32564 22520 32570
rect 22468 32506 22520 32512
rect 22282 32328 22338 32337
rect 22282 32263 22338 32272
rect 22296 32230 22324 32263
rect 22284 32224 22336 32230
rect 22284 32166 22336 32172
rect 22192 31884 22244 31890
rect 22192 31826 22244 31832
rect 21732 31476 21784 31482
rect 21732 31418 21784 31424
rect 22296 31142 22324 32166
rect 22284 31136 22336 31142
rect 22284 31078 22336 31084
rect 21180 30796 21232 30802
rect 21180 30738 21232 30744
rect 21640 30796 21692 30802
rect 21640 30738 21692 30744
rect 21362 30288 21418 30297
rect 21362 30223 21418 30232
rect 21376 30190 21404 30223
rect 21364 30184 21416 30190
rect 21364 30126 21416 30132
rect 21088 29708 21140 29714
rect 21088 29650 21140 29656
rect 20444 29174 20496 29180
rect 20902 29200 20958 29209
rect 20352 29028 20404 29034
rect 20352 28970 20404 28976
rect 20364 28422 20392 28970
rect 20352 28416 20404 28422
rect 20352 28358 20404 28364
rect 20260 27872 20312 27878
rect 20260 27814 20312 27820
rect 20272 27674 20300 27814
rect 20260 27668 20312 27674
rect 20260 27610 20312 27616
rect 20364 27554 20392 28358
rect 20456 27606 20484 29174
rect 21100 29170 21128 29650
rect 21652 29510 21680 30738
rect 22192 30728 22244 30734
rect 22192 30670 22244 30676
rect 21824 30592 21876 30598
rect 21824 30534 21876 30540
rect 21836 30190 21864 30534
rect 21824 30184 21876 30190
rect 21824 30126 21876 30132
rect 21640 29504 21692 29510
rect 21640 29446 21692 29452
rect 20902 29135 20904 29144
rect 20956 29135 20958 29144
rect 21088 29164 21140 29170
rect 20904 29106 20956 29112
rect 21088 29106 21140 29112
rect 20916 29075 20944 29106
rect 20904 29028 20956 29034
rect 21100 28994 21128 29106
rect 21548 29096 21600 29102
rect 21548 29038 21600 29044
rect 20904 28970 20956 28976
rect 20916 28014 20944 28970
rect 21008 28966 21128 28994
rect 21560 28966 21588 29038
rect 21652 29034 21680 29446
rect 21640 29028 21692 29034
rect 21640 28970 21692 28976
rect 21836 28966 21864 30126
rect 22204 29646 22232 30670
rect 22468 30116 22520 30122
rect 22468 30058 22520 30064
rect 22480 29850 22508 30058
rect 22468 29844 22520 29850
rect 22468 29786 22520 29792
rect 22192 29640 22244 29646
rect 22192 29582 22244 29588
rect 20904 28008 20956 28014
rect 20904 27950 20956 27956
rect 20272 27526 20392 27554
rect 20444 27600 20496 27606
rect 20444 27542 20496 27548
rect 20076 26920 20128 26926
rect 20076 26862 20128 26868
rect 20088 26586 20116 26862
rect 20076 26580 20128 26586
rect 20076 26522 20128 26528
rect 19984 26376 20036 26382
rect 19984 26318 20036 26324
rect 19892 24268 19944 24274
rect 19892 24210 19944 24216
rect 19904 23866 19932 24210
rect 19892 23860 19944 23866
rect 19892 23802 19944 23808
rect 19432 23792 19484 23798
rect 19432 23734 19484 23740
rect 19444 23050 19472 23734
rect 19996 23474 20024 26318
rect 20076 25832 20128 25838
rect 20076 25774 20128 25780
rect 20088 25498 20116 25774
rect 20168 25696 20220 25702
rect 20168 25638 20220 25644
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 20076 25288 20128 25294
rect 20076 25230 20128 25236
rect 20088 23882 20116 25230
rect 20180 24818 20208 25638
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20180 24410 20208 24754
rect 20168 24404 20220 24410
rect 20168 24346 20220 24352
rect 20088 23854 20208 23882
rect 20076 23792 20128 23798
rect 20076 23734 20128 23740
rect 19904 23446 20024 23474
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19616 23112 19668 23118
rect 19616 23054 19668 23060
rect 19432 23044 19484 23050
rect 19432 22986 19484 22992
rect 19444 22778 19472 22986
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19628 22710 19656 23054
rect 19616 22704 19668 22710
rect 19352 22630 19472 22658
rect 19616 22646 19668 22652
rect 19064 21966 19116 21972
rect 19168 21984 19288 22012
rect 18972 21888 19024 21894
rect 18972 21830 19024 21836
rect 18984 21486 19012 21830
rect 18788 21480 18840 21486
rect 18788 21422 18840 21428
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 18512 21344 18564 21350
rect 18512 21286 18564 21292
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18340 18426 18368 18566
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18236 18216 18288 18222
rect 18236 18158 18288 18164
rect 17868 17614 17920 17620
rect 17972 17598 18184 17626
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17880 13190 17908 14418
rect 17868 13184 17920 13190
rect 17868 13126 17920 13132
rect 17880 12986 17908 13126
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17788 11354 17816 12174
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 17684 11280 17736 11286
rect 17684 11222 17736 11228
rect 17696 10674 17724 11222
rect 17684 10668 17736 10674
rect 17684 10610 17736 10616
rect 17696 10198 17724 10610
rect 17684 10192 17736 10198
rect 17684 10134 17736 10140
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 17696 9722 17724 10134
rect 17684 9716 17736 9722
rect 17684 9658 17736 9664
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 17880 8634 17908 9046
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17420 7478 17448 7890
rect 17408 7472 17460 7478
rect 17408 7414 17460 7420
rect 17420 5914 17448 7414
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17316 5840 17368 5846
rect 17316 5782 17368 5788
rect 17328 5370 17356 5782
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17222 5264 17278 5273
rect 17222 5199 17278 5208
rect 17328 4826 17356 5306
rect 17316 4820 17368 4826
rect 17316 4762 17368 4768
rect 17512 4690 17540 8026
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17880 7478 17908 7890
rect 17972 7546 18000 17598
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 18156 17134 18184 17478
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 18052 16040 18104 16046
rect 18052 15982 18104 15988
rect 18064 11665 18092 15982
rect 18156 15910 18184 17070
rect 18144 15904 18196 15910
rect 18144 15846 18196 15852
rect 18248 15722 18276 18158
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18156 15694 18276 15722
rect 18050 11656 18106 11665
rect 18050 11591 18106 11600
rect 18064 9722 18092 11591
rect 18052 9716 18104 9722
rect 18052 9658 18104 9664
rect 18156 8945 18184 15694
rect 18340 15638 18368 16934
rect 18328 15632 18380 15638
rect 18328 15574 18380 15580
rect 18340 15162 18368 15574
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 18340 14890 18368 15098
rect 18328 14884 18380 14890
rect 18328 14826 18380 14832
rect 18236 14476 18288 14482
rect 18236 14418 18288 14424
rect 18248 13734 18276 14418
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18248 13297 18276 13670
rect 18234 13288 18290 13297
rect 18234 13223 18290 13232
rect 18248 12850 18276 13223
rect 18340 12918 18368 14826
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18340 12374 18368 12854
rect 18328 12368 18380 12374
rect 18328 12310 18380 12316
rect 18340 11898 18368 12310
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 18236 11212 18288 11218
rect 18288 11172 18368 11200
rect 18236 11154 18288 11160
rect 18340 10470 18368 11172
rect 18432 10810 18460 19994
rect 18524 13376 18552 21286
rect 18800 20806 18828 21422
rect 18972 21344 19024 21350
rect 18972 21286 19024 21292
rect 18984 21010 19012 21286
rect 18972 21004 19024 21010
rect 18972 20946 19024 20952
rect 18788 20800 18840 20806
rect 18788 20742 18840 20748
rect 18984 20602 19012 20946
rect 18972 20596 19024 20602
rect 18972 20538 19024 20544
rect 19076 20330 19104 21966
rect 19168 21162 19196 21984
rect 19444 21894 19472 22630
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19616 22092 19668 22098
rect 19616 22034 19668 22040
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19168 21134 19288 21162
rect 19156 21072 19208 21078
rect 19156 21014 19208 21020
rect 19168 20534 19196 21014
rect 19156 20528 19208 20534
rect 19156 20470 19208 20476
rect 19064 20324 19116 20330
rect 19064 20266 19116 20272
rect 19260 19922 19288 21134
rect 19340 19984 19392 19990
rect 19340 19926 19392 19932
rect 19248 19916 19300 19922
rect 19248 19858 19300 19864
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 18880 19508 18932 19514
rect 18880 19450 18932 19456
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 18604 18896 18656 18902
rect 18604 18838 18656 18844
rect 18616 18426 18644 18838
rect 18604 18420 18656 18426
rect 18604 18362 18656 18368
rect 18800 18222 18828 19110
rect 18788 18216 18840 18222
rect 18788 18158 18840 18164
rect 18604 17672 18656 17678
rect 18604 17614 18656 17620
rect 18616 16794 18644 17614
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18616 16046 18644 16390
rect 18788 16176 18840 16182
rect 18788 16118 18840 16124
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 18800 15706 18828 16118
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18696 15020 18748 15026
rect 18696 14962 18748 14968
rect 18708 14278 18736 14962
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18708 13734 18736 14214
rect 18892 14090 18920 19450
rect 19076 19174 19104 19790
rect 19156 19780 19208 19786
rect 19156 19722 19208 19728
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 18972 18964 19024 18970
rect 18972 18906 19024 18912
rect 18984 18426 19012 18906
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 19076 16046 19104 16594
rect 19064 16040 19116 16046
rect 19064 15982 19116 15988
rect 18972 15904 19024 15910
rect 18972 15846 19024 15852
rect 18984 14362 19012 15846
rect 19076 15366 19104 15982
rect 19064 15360 19116 15366
rect 19064 15302 19116 15308
rect 19076 14482 19104 15302
rect 19064 14476 19116 14482
rect 19064 14418 19116 14424
rect 18984 14334 19104 14362
rect 18800 14062 18920 14090
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18694 13424 18750 13433
rect 18524 13368 18694 13376
rect 18524 13348 18696 13368
rect 18748 13359 18750 13368
rect 18696 13330 18748 13336
rect 18512 12776 18564 12782
rect 18512 12718 18564 12724
rect 18524 11558 18552 12718
rect 18708 12170 18736 13330
rect 18696 12164 18748 12170
rect 18696 12106 18748 12112
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18340 10198 18368 10406
rect 18328 10192 18380 10198
rect 18328 10134 18380 10140
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18248 9518 18276 10066
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18248 9382 18276 9454
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18236 9036 18288 9042
rect 18236 8978 18288 8984
rect 18142 8936 18198 8945
rect 18142 8871 18198 8880
rect 18248 8362 18276 8978
rect 18800 8430 18828 14062
rect 18880 14000 18932 14006
rect 18880 13942 18932 13948
rect 18892 9586 18920 13942
rect 18972 13796 19024 13802
rect 18972 13738 19024 13744
rect 18984 11694 19012 13738
rect 18972 11688 19024 11694
rect 18972 11630 19024 11636
rect 18984 11354 19012 11630
rect 18972 11348 19024 11354
rect 18972 11290 19024 11296
rect 18984 11218 19012 11290
rect 18972 11212 19024 11218
rect 18972 11154 19024 11160
rect 19076 10810 19104 14334
rect 19064 10804 19116 10810
rect 19064 10746 19116 10752
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 18892 9178 18920 9522
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 19168 9042 19196 19722
rect 19260 18902 19288 19858
rect 19352 19718 19380 19926
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19352 19446 19380 19654
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19352 18970 19380 19382
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19248 18896 19300 18902
rect 19352 18873 19380 18906
rect 19248 18838 19300 18844
rect 19338 18864 19394 18873
rect 19338 18799 19394 18808
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 19260 17338 19288 17818
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19260 17066 19288 17274
rect 19248 17060 19300 17066
rect 19248 17002 19300 17008
rect 19248 16516 19300 16522
rect 19248 16458 19300 16464
rect 19260 16017 19288 16458
rect 19246 16008 19302 16017
rect 19246 15943 19302 15952
rect 19260 15910 19288 15943
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 19444 14006 19472 21490
rect 19628 21418 19656 22034
rect 19616 21412 19668 21418
rect 19616 21354 19668 21360
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 19536 19310 19564 19654
rect 19904 19378 19932 23446
rect 19984 23316 20036 23322
rect 19984 23258 20036 23264
rect 19996 22642 20024 23258
rect 19984 22636 20036 22642
rect 19984 22578 20036 22584
rect 19996 21554 20024 22578
rect 19984 21548 20036 21554
rect 19984 21490 20036 21496
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19996 19514 20024 20198
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19892 19372 19944 19378
rect 19892 19314 19944 19320
rect 19524 19304 19576 19310
rect 19524 19246 19576 19252
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19522 18864 19578 18873
rect 19522 18799 19578 18808
rect 19536 18766 19564 18799
rect 19904 18766 19932 19314
rect 20088 19310 20116 23734
rect 20180 19990 20208 23854
rect 20272 22817 20300 27526
rect 20456 27130 20484 27542
rect 20444 27124 20496 27130
rect 20444 27066 20496 27072
rect 20456 26314 20484 27066
rect 21008 27062 21036 28966
rect 21548 28960 21600 28966
rect 21548 28902 21600 28908
rect 21824 28960 21876 28966
rect 21824 28902 21876 28908
rect 21456 28756 21508 28762
rect 21456 28698 21508 28704
rect 21180 28552 21232 28558
rect 21180 28494 21232 28500
rect 21192 28082 21220 28494
rect 21180 28076 21232 28082
rect 21180 28018 21232 28024
rect 21468 27878 21496 28698
rect 21456 27872 21508 27878
rect 21456 27814 21508 27820
rect 21088 27532 21140 27538
rect 21088 27474 21140 27480
rect 20996 27056 21048 27062
rect 20996 26998 21048 27004
rect 20904 26988 20956 26994
rect 20904 26930 20956 26936
rect 20536 26784 20588 26790
rect 20536 26726 20588 26732
rect 20444 26308 20496 26314
rect 20444 26250 20496 26256
rect 20456 26042 20484 26250
rect 20444 26036 20496 26042
rect 20444 25978 20496 25984
rect 20548 25838 20576 26726
rect 20536 25832 20588 25838
rect 20536 25774 20588 25780
rect 20352 25356 20404 25362
rect 20352 25298 20404 25304
rect 20364 23322 20392 25298
rect 20548 25158 20576 25774
rect 20628 25696 20680 25702
rect 20628 25638 20680 25644
rect 20536 25152 20588 25158
rect 20536 25094 20588 25100
rect 20548 24342 20576 25094
rect 20536 24336 20588 24342
rect 20536 24278 20588 24284
rect 20536 23860 20588 23866
rect 20536 23802 20588 23808
rect 20352 23316 20404 23322
rect 20352 23258 20404 23264
rect 20548 22953 20576 23802
rect 20640 23769 20668 25638
rect 20720 24608 20772 24614
rect 20720 24550 20772 24556
rect 20626 23760 20682 23769
rect 20626 23695 20682 23704
rect 20732 23526 20760 24550
rect 20720 23520 20772 23526
rect 20720 23462 20772 23468
rect 20534 22944 20590 22953
rect 20534 22879 20590 22888
rect 20258 22808 20314 22817
rect 20258 22743 20314 22752
rect 20272 22234 20300 22743
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20548 20380 20576 21422
rect 20732 21350 20760 23462
rect 20812 23316 20864 23322
rect 20812 23258 20864 23264
rect 20720 21344 20772 21350
rect 20720 21286 20772 21292
rect 20732 21078 20760 21286
rect 20720 21072 20772 21078
rect 20720 21014 20772 21020
rect 20628 20392 20680 20398
rect 20548 20352 20628 20380
rect 20352 20256 20404 20262
rect 20352 20198 20404 20204
rect 20364 20058 20392 20198
rect 20548 20058 20576 20352
rect 20628 20334 20680 20340
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20824 19990 20852 23258
rect 20168 19984 20220 19990
rect 20812 19984 20864 19990
rect 20168 19926 20220 19932
rect 20732 19944 20812 19972
rect 20180 19718 20208 19926
rect 20352 19780 20404 19786
rect 20352 19722 20404 19728
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 19524 18760 19576 18766
rect 19524 18702 19576 18708
rect 19892 18760 19944 18766
rect 19892 18702 19944 18708
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19536 18222 19564 18566
rect 19904 18426 19932 18702
rect 19892 18420 19944 18426
rect 19892 18362 19944 18368
rect 19524 18216 19576 18222
rect 19524 18158 19576 18164
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 20260 18216 20312 18222
rect 20260 18158 20312 18164
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19996 17882 20024 18158
rect 19984 17876 20036 17882
rect 19984 17818 20036 17824
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19996 16250 20024 17818
rect 20076 17604 20128 17610
rect 20076 17546 20128 17552
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 19996 16046 20024 16186
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 19800 15564 19852 15570
rect 19800 15506 19852 15512
rect 19812 15162 19840 15506
rect 19800 15156 19852 15162
rect 19800 15098 19852 15104
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 19996 14482 20024 15982
rect 19984 14476 20036 14482
rect 19984 14418 20036 14424
rect 19996 14074 20024 14418
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 19260 13530 19288 13670
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19260 12646 19288 13330
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 20088 12306 20116 17546
rect 20272 17542 20300 18158
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 20260 16448 20312 16454
rect 20260 16390 20312 16396
rect 20272 16046 20300 16390
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 20272 13734 20300 14010
rect 20260 13728 20312 13734
rect 20260 13670 20312 13676
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 20088 11898 20116 12242
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 20364 11286 20392 19722
rect 20732 18970 20760 19944
rect 20812 19926 20864 19932
rect 20916 19836 20944 26930
rect 21100 26790 21128 27474
rect 21468 26790 21496 27814
rect 21088 26784 21140 26790
rect 21088 26726 21140 26732
rect 21456 26784 21508 26790
rect 21456 26726 21508 26732
rect 21100 26450 21128 26726
rect 21088 26444 21140 26450
rect 21088 26386 21140 26392
rect 21100 25945 21128 26386
rect 21086 25936 21142 25945
rect 21086 25871 21142 25880
rect 21272 24744 21324 24750
rect 21272 24686 21324 24692
rect 20996 24608 21048 24614
rect 20996 24550 21048 24556
rect 21008 23254 21036 24550
rect 21180 24404 21232 24410
rect 21180 24346 21232 24352
rect 21192 23730 21220 24346
rect 21284 24274 21312 24686
rect 21560 24313 21588 28902
rect 22204 28762 22232 29582
rect 22480 29170 22508 29786
rect 22468 29164 22520 29170
rect 22468 29106 22520 29112
rect 22192 28756 22244 28762
rect 22192 28698 22244 28704
rect 22480 28694 22508 29106
rect 22468 28688 22520 28694
rect 22468 28630 22520 28636
rect 22572 28218 22600 36722
rect 23032 36310 23060 40870
rect 23216 40594 23244 41482
rect 24228 40916 24256 41618
rect 24320 41206 24348 42094
rect 24872 42022 24900 42094
rect 30392 42022 30420 49558
rect 30470 49520 30526 49558
rect 35912 49558 36138 49586
rect 34940 46812 35236 46832
rect 34996 46810 35020 46812
rect 35076 46810 35100 46812
rect 35156 46810 35180 46812
rect 35018 46758 35020 46810
rect 35082 46758 35094 46810
rect 35156 46758 35158 46810
rect 34996 46756 35020 46758
rect 35076 46756 35100 46758
rect 35156 46756 35180 46758
rect 34940 46736 35236 46756
rect 34940 45724 35236 45744
rect 34996 45722 35020 45724
rect 35076 45722 35100 45724
rect 35156 45722 35180 45724
rect 35018 45670 35020 45722
rect 35082 45670 35094 45722
rect 35156 45670 35158 45722
rect 34996 45668 35020 45670
rect 35076 45668 35100 45670
rect 35156 45668 35180 45670
rect 34940 45648 35236 45668
rect 34940 44636 35236 44656
rect 34996 44634 35020 44636
rect 35076 44634 35100 44636
rect 35156 44634 35180 44636
rect 35018 44582 35020 44634
rect 35082 44582 35094 44634
rect 35156 44582 35158 44634
rect 34996 44580 35020 44582
rect 35076 44580 35100 44582
rect 35156 44580 35180 44582
rect 34940 44560 35236 44580
rect 34940 43548 35236 43568
rect 34996 43546 35020 43548
rect 35076 43546 35100 43548
rect 35156 43546 35180 43548
rect 35018 43494 35020 43546
rect 35082 43494 35094 43546
rect 35156 43494 35158 43546
rect 34996 43492 35020 43494
rect 35076 43492 35100 43494
rect 35156 43492 35180 43494
rect 34940 43472 35236 43492
rect 34940 42460 35236 42480
rect 34996 42458 35020 42460
rect 35076 42458 35100 42460
rect 35156 42458 35180 42460
rect 35018 42406 35020 42458
rect 35082 42406 35094 42458
rect 35156 42406 35158 42458
rect 34996 42404 35020 42406
rect 35076 42404 35100 42406
rect 35156 42404 35180 42406
rect 34940 42384 35236 42404
rect 24768 42016 24820 42022
rect 24768 41958 24820 41964
rect 24860 42016 24912 42022
rect 24860 41958 24912 41964
rect 30380 42016 30432 42022
rect 30380 41958 30432 41964
rect 24780 41818 24808 41958
rect 24768 41812 24820 41818
rect 24768 41754 24820 41760
rect 24584 41472 24636 41478
rect 24584 41414 24636 41420
rect 24308 41200 24360 41206
rect 24308 41142 24360 41148
rect 24308 40928 24360 40934
rect 24228 40888 24308 40916
rect 24308 40870 24360 40876
rect 23204 40588 23256 40594
rect 23204 40530 23256 40536
rect 23216 40050 23244 40530
rect 24320 40458 24348 40870
rect 24596 40730 24624 41414
rect 24780 41138 24808 41754
rect 24872 41721 24900 41958
rect 24858 41712 24914 41721
rect 24858 41647 24914 41656
rect 25964 41676 26016 41682
rect 25964 41618 26016 41624
rect 30196 41676 30248 41682
rect 30196 41618 30248 41624
rect 24952 41472 25004 41478
rect 24952 41414 25004 41420
rect 24768 41132 24820 41138
rect 24768 41074 24820 41080
rect 24584 40724 24636 40730
rect 24584 40666 24636 40672
rect 24308 40452 24360 40458
rect 24228 40412 24308 40440
rect 23204 40044 23256 40050
rect 23204 39986 23256 39992
rect 23216 39953 23244 39986
rect 23202 39944 23258 39953
rect 23202 39879 23258 39888
rect 24228 39545 24256 40412
rect 24308 40394 24360 40400
rect 24596 40118 24624 40666
rect 24964 40526 24992 41414
rect 25976 41041 26004 41618
rect 27436 41608 27488 41614
rect 27436 41550 27488 41556
rect 26884 41472 26936 41478
rect 26884 41414 26936 41420
rect 25962 41032 26018 41041
rect 25044 40996 25096 41002
rect 25962 40967 25964 40976
rect 25044 40938 25096 40944
rect 26016 40967 26018 40976
rect 25964 40938 26016 40944
rect 25056 40662 25084 40938
rect 25976 40907 26004 40938
rect 26896 40730 26924 41414
rect 27448 41274 27476 41550
rect 30104 41472 30156 41478
rect 30104 41414 30156 41420
rect 27436 41268 27488 41274
rect 27436 41210 27488 41216
rect 27252 41132 27304 41138
rect 27252 41074 27304 41080
rect 26976 40928 27028 40934
rect 26976 40870 27028 40876
rect 26884 40724 26936 40730
rect 26884 40666 26936 40672
rect 25044 40656 25096 40662
rect 25044 40598 25096 40604
rect 24952 40520 25004 40526
rect 24952 40462 25004 40468
rect 24584 40112 24636 40118
rect 24584 40054 24636 40060
rect 24964 39846 24992 40462
rect 25056 40186 25084 40598
rect 26148 40520 26200 40526
rect 26148 40462 26200 40468
rect 25044 40180 25096 40186
rect 25044 40122 25096 40128
rect 25056 39914 25084 40122
rect 25044 39908 25096 39914
rect 25044 39850 25096 39856
rect 24952 39840 25004 39846
rect 24952 39782 25004 39788
rect 25056 39642 25084 39850
rect 24308 39636 24360 39642
rect 24308 39578 24360 39584
rect 25044 39636 25096 39642
rect 25044 39578 25096 39584
rect 24214 39536 24270 39545
rect 24214 39471 24270 39480
rect 23940 39432 23992 39438
rect 23940 39374 23992 39380
rect 23756 39296 23808 39302
rect 23756 39238 23808 39244
rect 23768 38894 23796 39238
rect 23480 38888 23532 38894
rect 23480 38830 23532 38836
rect 23756 38888 23808 38894
rect 23756 38830 23808 38836
rect 23204 38820 23256 38826
rect 23204 38762 23256 38768
rect 23216 38486 23244 38762
rect 23388 38752 23440 38758
rect 23388 38694 23440 38700
rect 23400 38554 23428 38694
rect 23388 38548 23440 38554
rect 23388 38490 23440 38496
rect 23204 38480 23256 38486
rect 23256 38440 23336 38468
rect 23492 38457 23520 38830
rect 23952 38758 23980 39374
rect 24320 38962 24348 39578
rect 25228 39296 25280 39302
rect 25228 39238 25280 39244
rect 25240 38962 25268 39238
rect 24308 38956 24360 38962
rect 24308 38898 24360 38904
rect 24768 38956 24820 38962
rect 24768 38898 24820 38904
rect 25228 38956 25280 38962
rect 25228 38898 25280 38904
rect 23940 38752 23992 38758
rect 23940 38694 23992 38700
rect 23204 38422 23256 38428
rect 23204 38344 23256 38350
rect 23204 38286 23256 38292
rect 23216 37194 23244 38286
rect 23308 38010 23336 38440
rect 23478 38448 23534 38457
rect 23478 38383 23534 38392
rect 23664 38344 23716 38350
rect 23664 38286 23716 38292
rect 23296 38004 23348 38010
rect 23296 37946 23348 37952
rect 23388 37664 23440 37670
rect 23388 37606 23440 37612
rect 23400 37262 23428 37606
rect 23676 37398 23704 38286
rect 24780 38010 24808 38898
rect 25240 38554 25268 38898
rect 25320 38888 25372 38894
rect 25320 38830 25372 38836
rect 25228 38548 25280 38554
rect 25228 38490 25280 38496
rect 25332 38418 25360 38830
rect 25504 38820 25556 38826
rect 25504 38762 25556 38768
rect 25516 38554 25544 38762
rect 25504 38548 25556 38554
rect 25504 38490 25556 38496
rect 25136 38412 25188 38418
rect 25136 38354 25188 38360
rect 25320 38412 25372 38418
rect 25320 38354 25372 38360
rect 25148 38214 25176 38354
rect 25136 38208 25188 38214
rect 25136 38150 25188 38156
rect 24768 38004 24820 38010
rect 24768 37946 24820 37952
rect 25148 37942 25176 38150
rect 25136 37936 25188 37942
rect 25136 37878 25188 37884
rect 24768 37800 24820 37806
rect 24768 37742 24820 37748
rect 24676 37732 24728 37738
rect 24676 37674 24728 37680
rect 24308 37664 24360 37670
rect 24308 37606 24360 37612
rect 23664 37392 23716 37398
rect 23664 37334 23716 37340
rect 23388 37256 23440 37262
rect 23388 37198 23440 37204
rect 23204 37188 23256 37194
rect 23204 37130 23256 37136
rect 23400 36922 23428 37198
rect 23388 36916 23440 36922
rect 23388 36858 23440 36864
rect 23296 36712 23348 36718
rect 23296 36654 23348 36660
rect 23112 36644 23164 36650
rect 23112 36586 23164 36592
rect 22744 36304 22796 36310
rect 22744 36246 22796 36252
rect 23020 36304 23072 36310
rect 23020 36246 23072 36252
rect 22756 36145 22784 36246
rect 22742 36136 22798 36145
rect 22742 36071 22798 36080
rect 23124 35834 23152 36586
rect 23112 35828 23164 35834
rect 23112 35770 23164 35776
rect 23124 35290 23152 35770
rect 23112 35284 23164 35290
rect 23112 35226 23164 35232
rect 22926 34504 22982 34513
rect 22926 34439 22982 34448
rect 22940 33862 22968 34439
rect 23308 33930 23336 36654
rect 23572 36576 23624 36582
rect 23572 36518 23624 36524
rect 23388 36100 23440 36106
rect 23388 36042 23440 36048
rect 23400 35834 23428 36042
rect 23388 35828 23440 35834
rect 23388 35770 23440 35776
rect 23584 35698 23612 36518
rect 23572 35692 23624 35698
rect 23572 35634 23624 35640
rect 23676 35086 23704 37334
rect 24032 37324 24084 37330
rect 24032 37266 24084 37272
rect 24044 37097 24072 37266
rect 24030 37088 24086 37097
rect 24030 37023 24086 37032
rect 24044 36922 24072 37023
rect 24032 36916 24084 36922
rect 24032 36858 24084 36864
rect 24320 36718 24348 37606
rect 24584 37324 24636 37330
rect 24584 37266 24636 37272
rect 24308 36712 24360 36718
rect 24306 36680 24308 36689
rect 24360 36680 24362 36689
rect 24216 36644 24268 36650
rect 24596 36650 24624 37266
rect 24306 36615 24362 36624
rect 24584 36644 24636 36650
rect 24216 36586 24268 36592
rect 24584 36586 24636 36592
rect 24228 36242 24256 36586
rect 24216 36236 24268 36242
rect 24216 36178 24268 36184
rect 24308 36168 24360 36174
rect 24308 36110 24360 36116
rect 23848 35284 23900 35290
rect 23848 35226 23900 35232
rect 23664 35080 23716 35086
rect 23664 35022 23716 35028
rect 23860 34950 23888 35226
rect 24320 35154 24348 36110
rect 24688 35834 24716 37674
rect 24780 37398 24808 37742
rect 25148 37466 25176 37878
rect 25332 37466 25360 38354
rect 25516 37738 25544 38490
rect 25504 37732 25556 37738
rect 25504 37674 25556 37680
rect 25136 37460 25188 37466
rect 25136 37402 25188 37408
rect 25320 37460 25372 37466
rect 25320 37402 25372 37408
rect 24768 37392 24820 37398
rect 24768 37334 24820 37340
rect 24768 37120 24820 37126
rect 24768 37062 24820 37068
rect 24780 36242 24808 37062
rect 24768 36236 24820 36242
rect 24768 36178 24820 36184
rect 25412 36236 25464 36242
rect 25412 36178 25464 36184
rect 24768 36032 24820 36038
rect 24768 35974 24820 35980
rect 24676 35828 24728 35834
rect 24676 35770 24728 35776
rect 24688 35494 24716 35770
rect 24780 35698 24808 35974
rect 25424 35834 25452 36178
rect 25412 35828 25464 35834
rect 25412 35770 25464 35776
rect 26160 35698 26188 40462
rect 26896 40186 26924 40666
rect 26884 40180 26936 40186
rect 26884 40122 26936 40128
rect 26988 40050 27016 40870
rect 27068 40656 27120 40662
rect 27068 40598 27120 40604
rect 26976 40044 27028 40050
rect 26976 39986 27028 39992
rect 27080 39914 27108 40598
rect 27264 40050 27292 41074
rect 29920 40928 29972 40934
rect 29920 40870 29972 40876
rect 29932 40526 29960 40870
rect 29092 40520 29144 40526
rect 29092 40462 29144 40468
rect 29920 40520 29972 40526
rect 29920 40462 29972 40468
rect 27804 40112 27856 40118
rect 27804 40054 27856 40060
rect 27252 40044 27304 40050
rect 27252 39986 27304 39992
rect 27068 39908 27120 39914
rect 27068 39850 27120 39856
rect 27080 39574 27108 39850
rect 27068 39568 27120 39574
rect 27068 39510 27120 39516
rect 26976 39432 27028 39438
rect 26976 39374 27028 39380
rect 26988 39098 27016 39374
rect 26976 39092 27028 39098
rect 26976 39034 27028 39040
rect 27080 38758 27108 39510
rect 27068 38752 27120 38758
rect 27068 38694 27120 38700
rect 27080 38486 27108 38694
rect 27068 38480 27120 38486
rect 27068 38422 27120 38428
rect 26516 37868 26568 37874
rect 26516 37810 26568 37816
rect 26528 36854 26556 37810
rect 26620 37738 26924 37754
rect 26620 37732 26936 37738
rect 26620 37726 26884 37732
rect 26620 37670 26648 37726
rect 26608 37664 26660 37670
rect 26608 37606 26660 37612
rect 26700 37664 26752 37670
rect 26700 37606 26752 37612
rect 26712 37126 26740 37606
rect 26804 37398 26832 37726
rect 26884 37674 26936 37680
rect 26792 37392 26844 37398
rect 26792 37334 26844 37340
rect 26700 37120 26752 37126
rect 26700 37062 26752 37068
rect 26712 36922 26740 37062
rect 26700 36916 26752 36922
rect 26700 36858 26752 36864
rect 26804 36854 26832 37334
rect 27264 37262 27292 39986
rect 27816 39438 27844 40054
rect 29104 39846 29132 40462
rect 29920 40384 29972 40390
rect 29920 40326 29972 40332
rect 29092 39840 29144 39846
rect 29092 39782 29144 39788
rect 29000 39568 29052 39574
rect 29000 39510 29052 39516
rect 27804 39432 27856 39438
rect 27804 39374 27856 39380
rect 27712 38480 27764 38486
rect 27712 38422 27764 38428
rect 27528 38276 27580 38282
rect 27528 38218 27580 38224
rect 26976 37256 27028 37262
rect 26976 37198 27028 37204
rect 27252 37256 27304 37262
rect 27252 37198 27304 37204
rect 26516 36848 26568 36854
rect 26516 36790 26568 36796
rect 26792 36848 26844 36854
rect 26792 36790 26844 36796
rect 26792 36576 26844 36582
rect 26844 36553 26924 36564
rect 26844 36544 26938 36553
rect 26844 36536 26882 36544
rect 26792 36518 26844 36524
rect 26882 36479 26938 36488
rect 26988 36378 27016 37198
rect 27068 36848 27120 36854
rect 27068 36790 27120 36796
rect 27080 36650 27108 36790
rect 27068 36644 27120 36650
rect 27068 36586 27120 36592
rect 27080 36378 27108 36586
rect 26976 36372 27028 36378
rect 26976 36314 27028 36320
rect 27068 36372 27120 36378
rect 27068 36314 27120 36320
rect 26514 36272 26570 36281
rect 26514 36207 26570 36216
rect 27068 36236 27120 36242
rect 24768 35692 24820 35698
rect 24768 35634 24820 35640
rect 26148 35692 26200 35698
rect 26148 35634 26200 35640
rect 26424 35692 26476 35698
rect 26424 35634 26476 35640
rect 24676 35488 24728 35494
rect 24676 35430 24728 35436
rect 24688 35290 24716 35430
rect 24676 35284 24728 35290
rect 24676 35226 24728 35232
rect 24308 35148 24360 35154
rect 24308 35090 24360 35096
rect 23848 34944 23900 34950
rect 23848 34886 23900 34892
rect 23860 34542 23888 34886
rect 23848 34536 23900 34542
rect 23848 34478 23900 34484
rect 24320 34202 24348 35090
rect 24688 34746 24716 35226
rect 24676 34740 24728 34746
rect 24676 34682 24728 34688
rect 24308 34196 24360 34202
rect 24308 34138 24360 34144
rect 23296 33924 23348 33930
rect 23296 33866 23348 33872
rect 22928 33856 22980 33862
rect 22928 33798 22980 33804
rect 22940 33454 22968 33798
rect 24688 33522 24716 34682
rect 24780 34610 24808 35634
rect 25228 35488 25280 35494
rect 25228 35430 25280 35436
rect 25872 35488 25924 35494
rect 25872 35430 25924 35436
rect 25240 34746 25268 35430
rect 25884 35290 25912 35430
rect 26160 35290 26188 35634
rect 25872 35284 25924 35290
rect 25872 35226 25924 35232
rect 26148 35284 26200 35290
rect 26148 35226 26200 35232
rect 25412 35216 25464 35222
rect 25412 35158 25464 35164
rect 25228 34740 25280 34746
rect 25228 34682 25280 34688
rect 24768 34604 24820 34610
rect 24768 34546 24820 34552
rect 24952 34536 25004 34542
rect 24952 34478 25004 34484
rect 24964 34066 24992 34478
rect 25240 34406 25268 34682
rect 25424 34610 25452 35158
rect 26436 34610 26464 35634
rect 26528 35494 26556 36207
rect 27068 36178 27120 36184
rect 27080 35834 27108 36178
rect 27068 35828 27120 35834
rect 27068 35770 27120 35776
rect 26516 35488 26568 35494
rect 26516 35430 26568 35436
rect 25412 34604 25464 34610
rect 25412 34546 25464 34552
rect 26424 34604 26476 34610
rect 26424 34546 26476 34552
rect 25228 34400 25280 34406
rect 25228 34342 25280 34348
rect 25686 34368 25742 34377
rect 25686 34303 25742 34312
rect 25700 34066 25728 34303
rect 24952 34060 25004 34066
rect 24952 34002 25004 34008
rect 25688 34060 25740 34066
rect 25688 34002 25740 34008
rect 24676 33516 24728 33522
rect 24676 33458 24728 33464
rect 22928 33448 22980 33454
rect 22928 33390 22980 33396
rect 24400 33312 24452 33318
rect 24400 33254 24452 33260
rect 24412 33114 24440 33254
rect 24688 33134 24716 33458
rect 24400 33108 24452 33114
rect 24688 33106 24808 33134
rect 24964 33114 24992 34002
rect 25596 33992 25648 33998
rect 25596 33934 25648 33940
rect 25608 33522 25636 33934
rect 25700 33658 25728 34002
rect 25688 33652 25740 33658
rect 25688 33594 25740 33600
rect 25596 33516 25648 33522
rect 25596 33458 25648 33464
rect 26056 33516 26108 33522
rect 26056 33458 26108 33464
rect 25228 33380 25280 33386
rect 25228 33322 25280 33328
rect 25240 33153 25268 33322
rect 25226 33144 25282 33153
rect 24400 33050 24452 33056
rect 24780 33046 24808 33106
rect 24952 33108 25004 33114
rect 26068 33114 26096 33458
rect 26436 33153 26464 34546
rect 26422 33144 26478 33153
rect 25226 33079 25282 33088
rect 26056 33108 26108 33114
rect 24952 33050 25004 33056
rect 23112 33040 23164 33046
rect 23112 32982 23164 32988
rect 24768 33040 24820 33046
rect 24768 32982 24820 32988
rect 23124 32502 23152 32982
rect 23296 32904 23348 32910
rect 23296 32846 23348 32852
rect 23112 32496 23164 32502
rect 23112 32438 23164 32444
rect 22744 32428 22796 32434
rect 22744 32370 22796 32376
rect 22652 31884 22704 31890
rect 22756 31872 22784 32370
rect 23112 32292 23164 32298
rect 23112 32234 23164 32240
rect 23124 32026 23152 32234
rect 23308 32026 23336 32846
rect 23572 32768 23624 32774
rect 23572 32710 23624 32716
rect 23112 32020 23164 32026
rect 23112 31962 23164 31968
rect 23296 32020 23348 32026
rect 23296 31962 23348 31968
rect 23480 31952 23532 31958
rect 23480 31894 23532 31900
rect 22704 31844 22784 31872
rect 22652 31826 22704 31832
rect 22664 31414 22692 31826
rect 23492 31482 23520 31894
rect 23480 31476 23532 31482
rect 23480 31418 23532 31424
rect 22652 31408 22704 31414
rect 22652 31350 22704 31356
rect 22928 30864 22980 30870
rect 22928 30806 22980 30812
rect 22652 30728 22704 30734
rect 22652 30670 22704 30676
rect 22664 30394 22692 30670
rect 22940 30394 22968 30806
rect 23480 30728 23532 30734
rect 23480 30670 23532 30676
rect 22652 30388 22704 30394
rect 22652 30330 22704 30336
rect 22928 30388 22980 30394
rect 22928 30330 22980 30336
rect 22940 30122 22968 30330
rect 22928 30116 22980 30122
rect 22928 30058 22980 30064
rect 23492 29578 23520 30670
rect 23296 29572 23348 29578
rect 23296 29514 23348 29520
rect 23480 29572 23532 29578
rect 23480 29514 23532 29520
rect 23018 29200 23074 29209
rect 23018 29135 23074 29144
rect 23032 28422 23060 29135
rect 23112 28688 23164 28694
rect 23112 28630 23164 28636
rect 23020 28416 23072 28422
rect 23020 28358 23072 28364
rect 23124 28218 23152 28630
rect 23308 28558 23336 29514
rect 23296 28552 23348 28558
rect 23296 28494 23348 28500
rect 22560 28212 22612 28218
rect 22560 28154 22612 28160
rect 23112 28212 23164 28218
rect 23112 28154 23164 28160
rect 22572 28014 22600 28154
rect 21640 28008 21692 28014
rect 21640 27950 21692 27956
rect 21732 28008 21784 28014
rect 21732 27950 21784 27956
rect 22560 28008 22612 28014
rect 22560 27950 22612 27956
rect 21652 27538 21680 27950
rect 21640 27532 21692 27538
rect 21640 27474 21692 27480
rect 21652 26246 21680 27474
rect 21640 26240 21692 26246
rect 21640 26182 21692 26188
rect 21640 25832 21692 25838
rect 21640 25774 21692 25780
rect 21652 25702 21680 25774
rect 21640 25696 21692 25702
rect 21640 25638 21692 25644
rect 21546 24304 21602 24313
rect 21272 24268 21324 24274
rect 21546 24239 21602 24248
rect 21272 24210 21324 24216
rect 21284 23866 21312 24210
rect 21640 24064 21692 24070
rect 21640 24006 21692 24012
rect 21272 23860 21324 23866
rect 21272 23802 21324 23808
rect 21180 23724 21232 23730
rect 21180 23666 21232 23672
rect 21456 23520 21508 23526
rect 21456 23462 21508 23468
rect 20996 23248 21048 23254
rect 20996 23190 21048 23196
rect 21008 22778 21036 23190
rect 20996 22772 21048 22778
rect 20996 22714 21048 22720
rect 21468 22506 21496 23462
rect 21548 23044 21600 23050
rect 21548 22986 21600 22992
rect 21560 22642 21588 22986
rect 21548 22636 21600 22642
rect 21548 22578 21600 22584
rect 21456 22500 21508 22506
rect 21456 22442 21508 22448
rect 21272 22160 21324 22166
rect 21272 22102 21324 22108
rect 21180 22024 21232 22030
rect 21180 21966 21232 21972
rect 21192 21146 21220 21966
rect 21284 21690 21312 22102
rect 21560 22030 21588 22578
rect 21548 22024 21600 22030
rect 21548 21966 21600 21972
rect 21456 21956 21508 21962
rect 21456 21898 21508 21904
rect 21272 21684 21324 21690
rect 21272 21626 21324 21632
rect 21364 21480 21416 21486
rect 21364 21422 21416 21428
rect 21180 21140 21232 21146
rect 21180 21082 21232 21088
rect 21088 21072 21140 21078
rect 21088 21014 21140 21020
rect 21100 20602 21128 21014
rect 21088 20596 21140 20602
rect 21088 20538 21140 20544
rect 21376 20466 21404 21422
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 20996 19848 21048 19854
rect 20916 19808 20996 19836
rect 20812 19440 20864 19446
rect 20916 19428 20944 19808
rect 20996 19790 21048 19796
rect 21088 19712 21140 19718
rect 21088 19654 21140 19660
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 21100 19514 21128 19654
rect 21088 19508 21140 19514
rect 21088 19450 21140 19456
rect 20864 19400 20944 19428
rect 20812 19382 20864 19388
rect 20916 18970 20944 19400
rect 21192 19242 21220 19654
rect 21180 19236 21232 19242
rect 21180 19178 21232 19184
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 21364 18828 21416 18834
rect 21364 18770 21416 18776
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 20456 17202 20484 18226
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20456 16794 20484 17138
rect 20444 16788 20496 16794
rect 20444 16730 20496 16736
rect 20640 16454 20668 17614
rect 20628 16448 20680 16454
rect 20628 16390 20680 16396
rect 20640 16114 20668 16390
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20536 13864 20588 13870
rect 20534 13832 20536 13841
rect 20588 13832 20590 13841
rect 20534 13767 20590 13776
rect 20444 13388 20496 13394
rect 20444 13330 20496 13336
rect 20456 12646 20484 13330
rect 20548 13190 20576 13767
rect 20536 13184 20588 13190
rect 20536 13126 20588 13132
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 20456 11694 20484 12582
rect 20444 11688 20496 11694
rect 20444 11630 20496 11636
rect 19340 11280 19392 11286
rect 19340 11222 19392 11228
rect 20352 11280 20404 11286
rect 20352 11222 20404 11228
rect 19352 10266 19380 11222
rect 19892 11212 19944 11218
rect 19892 11154 19944 11160
rect 19904 10538 19932 11154
rect 19892 10532 19944 10538
rect 19892 10474 19944 10480
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19340 10260 19392 10266
rect 19444 10248 19472 10406
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19444 10220 19564 10248
rect 19340 10202 19392 10208
rect 19352 9110 19380 10202
rect 19432 10124 19484 10130
rect 19536 10112 19564 10220
rect 19616 10124 19668 10130
rect 19536 10084 19616 10112
rect 19432 10066 19484 10072
rect 19616 10066 19668 10072
rect 19444 10033 19472 10066
rect 19430 10024 19486 10033
rect 19430 9959 19486 9968
rect 19628 9450 19656 10066
rect 19616 9444 19668 9450
rect 19616 9386 19668 9392
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19340 9104 19392 9110
rect 19340 9046 19392 9052
rect 19904 9042 19932 10474
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 19984 9512 20036 9518
rect 19984 9454 20036 9460
rect 19996 9110 20024 9454
rect 20272 9178 20300 9522
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 19984 9104 20036 9110
rect 19984 9046 20036 9052
rect 19156 9036 19208 9042
rect 19156 8978 19208 8984
rect 19892 9036 19944 9042
rect 19892 8978 19944 8984
rect 19168 8634 19196 8978
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 18788 8424 18840 8430
rect 18788 8366 18840 8372
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 18800 8090 18828 8366
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17868 7472 17920 7478
rect 17868 7414 17920 7420
rect 17880 6934 17908 7414
rect 18984 7274 19012 8366
rect 19904 8362 19932 8978
rect 19892 8356 19944 8362
rect 19892 8298 19944 8304
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 19076 7954 19104 8230
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 19432 8016 19484 8022
rect 19432 7958 19484 7964
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 18972 7268 19024 7274
rect 18972 7210 19024 7216
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 18512 6928 18564 6934
rect 18512 6870 18564 6876
rect 17880 6322 17908 6870
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 17880 4865 17908 6054
rect 18156 5914 18184 6054
rect 18524 5914 18552 6870
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 19076 6458 19104 6734
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18156 5234 18184 5850
rect 18880 5840 18932 5846
rect 18880 5782 18932 5788
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 17866 4856 17922 4865
rect 18800 4826 18828 5646
rect 18892 5370 18920 5782
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 17866 4791 17922 4800
rect 18788 4820 18840 4826
rect 17592 4752 17644 4758
rect 17592 4694 17644 4700
rect 17500 4684 17552 4690
rect 17500 4626 17552 4632
rect 17604 4282 17632 4694
rect 17880 4690 17908 4791
rect 18788 4762 18840 4768
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 17592 4276 17644 4282
rect 17592 4218 17644 4224
rect 17788 4010 17816 4422
rect 17880 4282 17908 4626
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 17868 4276 17920 4282
rect 17868 4218 17920 4224
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 17776 4004 17828 4010
rect 17776 3946 17828 3952
rect 18236 4004 18288 4010
rect 18236 3946 18288 3952
rect 16684 3590 16804 3618
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16488 3120 16540 3126
rect 16488 3062 16540 3068
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 16500 2650 16528 3062
rect 16488 2644 16540 2650
rect 16488 2586 16540 2592
rect 16396 2576 16448 2582
rect 16396 2518 16448 2524
rect 16408 2417 16436 2518
rect 16684 2446 16712 3590
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16776 3194 16804 3470
rect 17788 3194 17816 3946
rect 18248 3738 18276 3946
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 18156 3194 18184 3606
rect 18432 3534 18460 4082
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18156 2650 18184 3130
rect 18248 2854 18276 3470
rect 18432 3126 18460 3470
rect 18420 3120 18472 3126
rect 18420 3062 18472 3068
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 16672 2440 16724 2446
rect 16394 2408 16450 2417
rect 16672 2382 16724 2388
rect 18248 2378 18276 2790
rect 18524 2514 18552 4558
rect 18800 4146 18828 4762
rect 19154 4176 19210 4185
rect 18788 4140 18840 4146
rect 19154 4111 19210 4120
rect 18788 4082 18840 4088
rect 19168 4010 19196 4111
rect 19156 4004 19208 4010
rect 19156 3946 19208 3952
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18892 3398 18920 3878
rect 19168 3602 19196 3946
rect 19156 3596 19208 3602
rect 19156 3538 19208 3544
rect 18880 3392 18932 3398
rect 18880 3334 18932 3340
rect 18972 3392 19024 3398
rect 18972 3334 19024 3340
rect 18984 3058 19012 3334
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18512 2508 18564 2514
rect 18512 2450 18564 2456
rect 16394 2343 16450 2352
rect 18236 2372 18288 2378
rect 18236 2314 18288 2320
rect 16026 82 16082 480
rect 15764 54 16082 82
rect 19352 82 19380 7142
rect 19444 7002 19472 7958
rect 19904 7954 19932 8298
rect 19616 7948 19668 7954
rect 19616 7890 19668 7896
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 19628 7478 19656 7890
rect 19616 7472 19668 7478
rect 19616 7414 19668 7420
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19892 6180 19944 6186
rect 19892 6122 19944 6128
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 19524 4684 19576 4690
rect 19524 4626 19576 4632
rect 19536 4282 19564 4626
rect 19524 4276 19576 4282
rect 19524 4218 19576 4224
rect 19904 4078 19932 6122
rect 19996 4690 20024 7142
rect 20166 6352 20222 6361
rect 20166 6287 20222 6296
rect 20180 6254 20208 6287
rect 20168 6248 20220 6254
rect 20168 6190 20220 6196
rect 20272 5370 20300 9114
rect 20548 8786 20576 13126
rect 20732 11286 20760 18702
rect 21376 18426 21404 18770
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 21272 17876 21324 17882
rect 21272 17818 21324 17824
rect 20812 17264 20864 17270
rect 20812 17206 20864 17212
rect 20824 12102 20852 17206
rect 21284 17066 21312 17818
rect 21468 17338 21496 21898
rect 21560 20874 21588 21966
rect 21548 20868 21600 20874
rect 21548 20810 21600 20816
rect 21560 20398 21588 20810
rect 21548 20392 21600 20398
rect 21548 20334 21600 20340
rect 21652 19310 21680 24006
rect 21744 23798 21772 27950
rect 22560 27872 22612 27878
rect 22560 27814 22612 27820
rect 22572 27606 22600 27814
rect 22560 27600 22612 27606
rect 22560 27542 22612 27548
rect 23020 27600 23072 27606
rect 23020 27542 23072 27548
rect 21824 27464 21876 27470
rect 21824 27406 21876 27412
rect 21836 26994 21864 27406
rect 22572 27062 22600 27542
rect 23032 27130 23060 27542
rect 23308 27402 23336 28494
rect 23296 27396 23348 27402
rect 23296 27338 23348 27344
rect 23020 27124 23072 27130
rect 23020 27066 23072 27072
rect 22560 27056 22612 27062
rect 22560 26998 22612 27004
rect 21824 26988 21876 26994
rect 21824 26930 21876 26936
rect 21836 26586 21864 26930
rect 22744 26784 22796 26790
rect 22744 26726 22796 26732
rect 21824 26580 21876 26586
rect 21824 26522 21876 26528
rect 22756 26518 22784 26726
rect 22744 26512 22796 26518
rect 22744 26454 22796 26460
rect 22192 26376 22244 26382
rect 22192 26318 22244 26324
rect 22100 26240 22152 26246
rect 22100 26182 22152 26188
rect 22112 25838 22140 26182
rect 22204 25906 22232 26318
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 22100 25832 22152 25838
rect 22100 25774 22152 25780
rect 22112 25158 22140 25774
rect 22204 25498 22232 25842
rect 22284 25764 22336 25770
rect 22284 25706 22336 25712
rect 22192 25492 22244 25498
rect 22192 25434 22244 25440
rect 22100 25152 22152 25158
rect 22100 25094 22152 25100
rect 22296 24274 22324 25706
rect 22756 25702 22784 26454
rect 23020 26240 23072 26246
rect 23020 26182 23072 26188
rect 22744 25696 22796 25702
rect 22744 25638 22796 25644
rect 22652 25152 22704 25158
rect 22652 25094 22704 25100
rect 22664 24750 22692 25094
rect 22652 24744 22704 24750
rect 22652 24686 22704 24692
rect 22664 24342 22692 24686
rect 22756 24682 22784 25638
rect 23032 25430 23060 26182
rect 23020 25424 23072 25430
rect 23020 25366 23072 25372
rect 23032 24954 23060 25366
rect 23308 25294 23336 27338
rect 23296 25288 23348 25294
rect 23296 25230 23348 25236
rect 23020 24948 23072 24954
rect 23020 24890 23072 24896
rect 22744 24676 22796 24682
rect 22744 24618 22796 24624
rect 23308 24410 23336 25230
rect 23296 24404 23348 24410
rect 23296 24346 23348 24352
rect 22652 24336 22704 24342
rect 22652 24278 22704 24284
rect 22192 24268 22244 24274
rect 22192 24210 22244 24216
rect 22284 24268 22336 24274
rect 22284 24210 22336 24216
rect 22928 24268 22980 24274
rect 22928 24210 22980 24216
rect 22204 23866 22232 24210
rect 22940 23866 22968 24210
rect 22192 23860 22244 23866
rect 22192 23802 22244 23808
rect 22928 23860 22980 23866
rect 22928 23802 22980 23808
rect 21732 23792 21784 23798
rect 21732 23734 21784 23740
rect 23584 23474 23612 32710
rect 24032 32564 24084 32570
rect 24032 32506 24084 32512
rect 23940 32496 23992 32502
rect 23940 32438 23992 32444
rect 23952 32026 23980 32438
rect 24044 32026 24072 32506
rect 24780 32230 24808 32982
rect 24964 32570 24992 33050
rect 25240 32978 25268 33079
rect 26422 33079 26478 33088
rect 26056 33050 26108 33056
rect 26424 33040 26476 33046
rect 26424 32982 26476 32988
rect 25228 32972 25280 32978
rect 25228 32914 25280 32920
rect 24952 32564 25004 32570
rect 24952 32506 25004 32512
rect 24768 32224 24820 32230
rect 24768 32166 24820 32172
rect 23940 32020 23992 32026
rect 23940 31962 23992 31968
rect 24032 32020 24084 32026
rect 24032 31962 24084 31968
rect 24860 31952 24912 31958
rect 24860 31894 24912 31900
rect 24492 31884 24544 31890
rect 24492 31826 24544 31832
rect 23940 31136 23992 31142
rect 23940 31078 23992 31084
rect 23952 30938 23980 31078
rect 24504 30938 24532 31826
rect 24872 31362 24900 31894
rect 24964 31890 24992 32506
rect 25136 32428 25188 32434
rect 25136 32370 25188 32376
rect 25148 31958 25176 32370
rect 25240 32026 25268 32914
rect 26332 32836 26384 32842
rect 26332 32778 26384 32784
rect 25688 32768 25740 32774
rect 25688 32710 25740 32716
rect 25700 32434 25728 32710
rect 25688 32428 25740 32434
rect 25688 32370 25740 32376
rect 26344 32026 26372 32778
rect 26436 32230 26464 32982
rect 26424 32224 26476 32230
rect 26424 32166 26476 32172
rect 26436 32026 26464 32166
rect 25228 32020 25280 32026
rect 25228 31962 25280 31968
rect 26332 32020 26384 32026
rect 26332 31962 26384 31968
rect 26424 32020 26476 32026
rect 26424 31962 26476 31968
rect 25136 31952 25188 31958
rect 25136 31894 25188 31900
rect 24952 31884 25004 31890
rect 24952 31826 25004 31832
rect 26424 31884 26476 31890
rect 26424 31826 26476 31832
rect 26332 31748 26384 31754
rect 26332 31690 26384 31696
rect 25412 31680 25464 31686
rect 25412 31622 25464 31628
rect 25872 31680 25924 31686
rect 25872 31622 25924 31628
rect 24950 31376 25006 31385
rect 24872 31334 24950 31362
rect 24950 31311 25006 31320
rect 24964 31278 24992 31311
rect 24952 31272 25004 31278
rect 24952 31214 25004 31220
rect 24964 30977 24992 31214
rect 25424 31210 25452 31622
rect 25780 31340 25832 31346
rect 25780 31282 25832 31288
rect 25412 31204 25464 31210
rect 25412 31146 25464 31152
rect 24950 30968 25006 30977
rect 23940 30932 23992 30938
rect 23940 30874 23992 30880
rect 24492 30932 24544 30938
rect 24950 30903 25006 30912
rect 24492 30874 24544 30880
rect 24952 30864 25004 30870
rect 24952 30806 25004 30812
rect 24124 30728 24176 30734
rect 24124 30670 24176 30676
rect 24136 30394 24164 30670
rect 24124 30388 24176 30394
rect 24124 30330 24176 30336
rect 23756 30184 23808 30190
rect 23756 30126 23808 30132
rect 23768 30054 23796 30126
rect 24964 30122 24992 30806
rect 24952 30116 25004 30122
rect 24952 30058 25004 30064
rect 23756 30048 23808 30054
rect 23756 29990 23808 29996
rect 23768 28665 23796 29990
rect 24964 29850 24992 30058
rect 25424 30054 25452 31146
rect 25792 30598 25820 31282
rect 25780 30592 25832 30598
rect 25780 30534 25832 30540
rect 25596 30184 25648 30190
rect 25596 30126 25648 30132
rect 25412 30048 25464 30054
rect 25412 29990 25464 29996
rect 25424 29850 25452 29990
rect 24952 29844 25004 29850
rect 24952 29786 25004 29792
rect 25412 29844 25464 29850
rect 25412 29786 25464 29792
rect 24124 29776 24176 29782
rect 24124 29718 24176 29724
rect 24032 29640 24084 29646
rect 24032 29582 24084 29588
rect 24044 29306 24072 29582
rect 24032 29300 24084 29306
rect 24032 29242 24084 29248
rect 24136 29170 24164 29718
rect 25228 29572 25280 29578
rect 25228 29514 25280 29520
rect 24124 29164 24176 29170
rect 24124 29106 24176 29112
rect 25240 29034 25268 29514
rect 25228 29028 25280 29034
rect 25228 28970 25280 28976
rect 25424 28966 25452 29786
rect 25412 28960 25464 28966
rect 25412 28902 25464 28908
rect 25608 28694 25636 30126
rect 25792 29850 25820 30534
rect 25884 30394 25912 31622
rect 25964 31204 26016 31210
rect 25964 31146 26016 31152
rect 25976 30870 26004 31146
rect 26240 31136 26292 31142
rect 26240 31078 26292 31084
rect 25964 30864 26016 30870
rect 25964 30806 26016 30812
rect 25872 30388 25924 30394
rect 25872 30330 25924 30336
rect 25780 29844 25832 29850
rect 25780 29786 25832 29792
rect 25044 28688 25096 28694
rect 23754 28656 23810 28665
rect 25044 28630 25096 28636
rect 25596 28688 25648 28694
rect 25648 28648 25728 28676
rect 25596 28630 25648 28636
rect 23754 28591 23810 28600
rect 24768 28552 24820 28558
rect 24768 28494 24820 28500
rect 23664 28484 23716 28490
rect 23664 28426 23716 28432
rect 23676 27674 23704 28426
rect 24780 28218 24808 28494
rect 24768 28212 24820 28218
rect 24768 28154 24820 28160
rect 25056 28150 25084 28630
rect 25044 28144 25096 28150
rect 25044 28086 25096 28092
rect 25596 28076 25648 28082
rect 25596 28018 25648 28024
rect 25320 27872 25372 27878
rect 25320 27814 25372 27820
rect 23664 27668 23716 27674
rect 23664 27610 23716 27616
rect 25136 27600 25188 27606
rect 25136 27542 25188 27548
rect 24860 27532 24912 27538
rect 24860 27474 24912 27480
rect 24872 27130 24900 27474
rect 24952 27328 25004 27334
rect 24952 27270 25004 27276
rect 24492 27124 24544 27130
rect 24492 27066 24544 27072
rect 24860 27124 24912 27130
rect 24860 27066 24912 27072
rect 24400 26920 24452 26926
rect 24400 26862 24452 26868
rect 23940 26444 23992 26450
rect 23940 26386 23992 26392
rect 23952 26081 23980 26386
rect 23938 26072 23994 26081
rect 23938 26007 23994 26016
rect 23952 25974 23980 26007
rect 23940 25968 23992 25974
rect 23940 25910 23992 25916
rect 24412 25809 24440 26862
rect 24398 25800 24454 25809
rect 24398 25735 24454 25744
rect 23940 25152 23992 25158
rect 23940 25094 23992 25100
rect 23952 24818 23980 25094
rect 23940 24812 23992 24818
rect 23940 24754 23992 24760
rect 24216 24676 24268 24682
rect 24216 24618 24268 24624
rect 24228 24410 24256 24618
rect 24216 24404 24268 24410
rect 24216 24346 24268 24352
rect 23848 24200 23900 24206
rect 23848 24142 23900 24148
rect 23492 23446 23612 23474
rect 22928 23180 22980 23186
rect 22928 23122 22980 23128
rect 23388 23180 23440 23186
rect 23388 23122 23440 23128
rect 22940 22778 22968 23122
rect 23400 22778 23428 23122
rect 22928 22772 22980 22778
rect 22928 22714 22980 22720
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 22744 22092 22796 22098
rect 22744 22034 22796 22040
rect 22756 21690 22784 22034
rect 23112 21888 23164 21894
rect 23112 21830 23164 21836
rect 22744 21684 22796 21690
rect 22744 21626 22796 21632
rect 22376 21480 22428 21486
rect 22376 21422 22428 21428
rect 21916 20936 21968 20942
rect 21916 20878 21968 20884
rect 21928 20602 21956 20878
rect 22388 20602 22416 21422
rect 21916 20596 21968 20602
rect 21916 20538 21968 20544
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 23124 19990 23152 21830
rect 23296 20868 23348 20874
rect 23296 20810 23348 20816
rect 23204 20460 23256 20466
rect 23204 20402 23256 20408
rect 23112 19984 23164 19990
rect 23112 19926 23164 19932
rect 23124 19514 23152 19926
rect 23216 19786 23244 20402
rect 23308 19854 23336 20810
rect 23388 20800 23440 20806
rect 23388 20742 23440 20748
rect 23400 20602 23428 20742
rect 23388 20596 23440 20602
rect 23388 20538 23440 20544
rect 23400 20262 23428 20538
rect 23388 20256 23440 20262
rect 23388 20198 23440 20204
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 23204 19780 23256 19786
rect 23204 19722 23256 19728
rect 23112 19508 23164 19514
rect 23112 19450 23164 19456
rect 21640 19304 21692 19310
rect 21640 19246 21692 19252
rect 22008 19304 22060 19310
rect 22008 19246 22060 19252
rect 22020 18970 22048 19246
rect 22192 19168 22244 19174
rect 22192 19110 22244 19116
rect 22008 18964 22060 18970
rect 22008 18906 22060 18912
rect 22204 18766 22232 19110
rect 23020 18828 23072 18834
rect 23020 18770 23072 18776
rect 22192 18760 22244 18766
rect 22192 18702 22244 18708
rect 23032 18426 23060 18770
rect 23020 18420 23072 18426
rect 23020 18362 23072 18368
rect 21928 18154 22232 18170
rect 21928 18148 22244 18154
rect 21928 18142 22192 18148
rect 21928 18086 21956 18142
rect 22192 18090 22244 18096
rect 21916 18080 21968 18086
rect 21916 18022 21968 18028
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 21456 17332 21508 17338
rect 21456 17274 21508 17280
rect 21272 17060 21324 17066
rect 21272 17002 21324 17008
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 21376 15910 21404 16594
rect 21928 15978 21956 18022
rect 22020 17542 22048 18022
rect 23216 17762 23244 19722
rect 23388 19168 23440 19174
rect 23388 19110 23440 19116
rect 23400 18902 23428 19110
rect 23388 18896 23440 18902
rect 23388 18838 23440 18844
rect 23492 18329 23520 23446
rect 23860 23322 23888 24142
rect 24032 24064 24084 24070
rect 24032 24006 24084 24012
rect 24044 23662 24072 24006
rect 24228 23866 24256 24346
rect 24216 23860 24268 23866
rect 24216 23802 24268 23808
rect 23940 23656 23992 23662
rect 23940 23598 23992 23604
rect 24032 23656 24084 23662
rect 24032 23598 24084 23604
rect 23848 23316 23900 23322
rect 23848 23258 23900 23264
rect 23952 22710 23980 23598
rect 24044 23186 24072 23598
rect 24504 23497 24532 27066
rect 24860 26852 24912 26858
rect 24860 26794 24912 26800
rect 24872 26586 24900 26794
rect 24860 26580 24912 26586
rect 24860 26522 24912 26528
rect 24964 26518 24992 27270
rect 25148 26858 25176 27542
rect 25228 27056 25280 27062
rect 25228 26998 25280 27004
rect 25136 26852 25188 26858
rect 25136 26794 25188 26800
rect 25148 26518 25176 26794
rect 24952 26512 25004 26518
rect 24952 26454 25004 26460
rect 25136 26512 25188 26518
rect 25136 26454 25188 26460
rect 24768 25764 24820 25770
rect 24768 25706 24820 25712
rect 24780 24410 24808 25706
rect 24964 25498 24992 26454
rect 25148 26042 25176 26454
rect 25136 26036 25188 26042
rect 25136 25978 25188 25984
rect 25240 25906 25268 26998
rect 25228 25900 25280 25906
rect 25228 25842 25280 25848
rect 25240 25498 25268 25842
rect 24952 25492 25004 25498
rect 24952 25434 25004 25440
rect 25228 25492 25280 25498
rect 25228 25434 25280 25440
rect 25044 25424 25096 25430
rect 25044 25366 25096 25372
rect 25136 25424 25188 25430
rect 25136 25366 25188 25372
rect 25056 24954 25084 25366
rect 25148 25294 25176 25366
rect 25136 25288 25188 25294
rect 25136 25230 25188 25236
rect 25044 24948 25096 24954
rect 25044 24890 25096 24896
rect 25148 24410 25176 25230
rect 24768 24404 24820 24410
rect 24768 24346 24820 24352
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 24490 23488 24546 23497
rect 24412 23446 24490 23474
rect 24032 23180 24084 23186
rect 24032 23122 24084 23128
rect 23940 22704 23992 22710
rect 23940 22646 23992 22652
rect 23572 22568 23624 22574
rect 23952 22545 23980 22646
rect 23572 22510 23624 22516
rect 23938 22536 23994 22545
rect 23584 22234 23612 22510
rect 23938 22471 23994 22480
rect 23664 22432 23716 22438
rect 23664 22374 23716 22380
rect 23572 22228 23624 22234
rect 23572 22170 23624 22176
rect 23584 21962 23612 22170
rect 23572 21956 23624 21962
rect 23572 21898 23624 21904
rect 23572 21344 23624 21350
rect 23572 21286 23624 21292
rect 23584 21010 23612 21286
rect 23572 21004 23624 21010
rect 23572 20946 23624 20952
rect 23584 20534 23612 20946
rect 23572 20528 23624 20534
rect 23572 20470 23624 20476
rect 23572 19236 23624 19242
rect 23572 19178 23624 19184
rect 23584 18902 23612 19178
rect 23676 18970 23704 22374
rect 24412 22137 24440 23446
rect 24490 23423 24546 23432
rect 24492 23180 24544 23186
rect 24492 23122 24544 23128
rect 25228 23180 25280 23186
rect 25228 23122 25280 23128
rect 24504 23089 24532 23122
rect 24490 23080 24546 23089
rect 24490 23015 24546 23024
rect 24504 22778 24532 23015
rect 24492 22772 24544 22778
rect 24492 22714 24544 22720
rect 24398 22128 24454 22137
rect 24504 22098 24532 22714
rect 25240 22574 25268 23122
rect 25332 23050 25360 27814
rect 25608 27674 25636 28018
rect 25596 27668 25648 27674
rect 25596 27610 25648 27616
rect 25700 26518 25728 28648
rect 25976 28490 26004 30806
rect 26056 29164 26108 29170
rect 26056 29106 26108 29112
rect 25964 28484 26016 28490
rect 25964 28426 26016 28432
rect 25976 27062 26004 28426
rect 26068 28014 26096 29106
rect 26252 29102 26280 31078
rect 26344 30258 26372 31690
rect 26436 31482 26464 31826
rect 26424 31476 26476 31482
rect 26424 31418 26476 31424
rect 26332 30252 26384 30258
rect 26332 30194 26384 30200
rect 26344 29782 26372 30194
rect 26332 29776 26384 29782
rect 26332 29718 26384 29724
rect 26240 29096 26292 29102
rect 26240 29038 26292 29044
rect 26056 28008 26108 28014
rect 26056 27950 26108 27956
rect 26068 27062 26096 27950
rect 25964 27056 26016 27062
rect 25964 26998 26016 27004
rect 26056 27056 26108 27062
rect 26056 26998 26108 27004
rect 25688 26512 25740 26518
rect 25688 26454 25740 26460
rect 25412 25900 25464 25906
rect 25412 25842 25464 25848
rect 25424 25294 25452 25842
rect 25700 25430 25728 26454
rect 25688 25424 25740 25430
rect 25688 25366 25740 25372
rect 26436 25362 26464 31418
rect 26528 29696 26556 35430
rect 27160 35216 27212 35222
rect 27264 35204 27292 37198
rect 27540 36718 27568 38218
rect 27724 38010 27752 38422
rect 27712 38004 27764 38010
rect 27712 37946 27764 37952
rect 27816 37738 27844 39374
rect 29012 39098 29040 39510
rect 29000 39092 29052 39098
rect 29000 39034 29052 39040
rect 29012 38758 29040 39034
rect 29000 38752 29052 38758
rect 29000 38694 29052 38700
rect 29012 38554 29040 38694
rect 29000 38548 29052 38554
rect 29000 38490 29052 38496
rect 28448 38412 28500 38418
rect 28448 38354 28500 38360
rect 28080 38344 28132 38350
rect 28080 38286 28132 38292
rect 28092 38010 28120 38286
rect 28080 38004 28132 38010
rect 28080 37946 28132 37952
rect 28460 37874 28488 38354
rect 28448 37868 28500 37874
rect 28448 37810 28500 37816
rect 27804 37732 27856 37738
rect 27804 37674 27856 37680
rect 27528 36712 27580 36718
rect 27528 36654 27580 36660
rect 27344 35284 27396 35290
rect 27344 35226 27396 35232
rect 27212 35176 27292 35204
rect 27160 35158 27212 35164
rect 27160 35080 27212 35086
rect 27160 35022 27212 35028
rect 26976 34400 27028 34406
rect 26976 34342 27028 34348
rect 26988 34134 27016 34342
rect 27172 34202 27200 35022
rect 27264 35018 27292 35176
rect 27252 35012 27304 35018
rect 27252 34954 27304 34960
rect 27356 34610 27384 35226
rect 27540 34610 27568 36654
rect 27712 36032 27764 36038
rect 27712 35974 27764 35980
rect 27724 35562 27752 35974
rect 27712 35556 27764 35562
rect 27712 35498 27764 35504
rect 27724 35290 27752 35498
rect 27712 35284 27764 35290
rect 27712 35226 27764 35232
rect 27344 34604 27396 34610
rect 27528 34604 27580 34610
rect 27344 34546 27396 34552
rect 27448 34564 27528 34592
rect 27356 34474 27384 34546
rect 27344 34468 27396 34474
rect 27344 34410 27396 34416
rect 27160 34196 27212 34202
rect 27160 34138 27212 34144
rect 27356 34134 27384 34410
rect 26976 34128 27028 34134
rect 26976 34070 27028 34076
rect 27344 34128 27396 34134
rect 27344 34070 27396 34076
rect 27356 33658 27384 34070
rect 27344 33652 27396 33658
rect 27344 33594 27396 33600
rect 26882 33144 26938 33153
rect 26882 33079 26938 33088
rect 26896 32910 26924 33079
rect 26884 32904 26936 32910
rect 26884 32846 26936 32852
rect 27448 32842 27476 34564
rect 27528 34546 27580 34552
rect 27712 34468 27764 34474
rect 27712 34410 27764 34416
rect 27620 33992 27672 33998
rect 27620 33934 27672 33940
rect 27528 33856 27580 33862
rect 27528 33798 27580 33804
rect 27540 33454 27568 33798
rect 27632 33658 27660 33934
rect 27724 33930 27752 34410
rect 27816 33930 27844 37674
rect 28460 37233 28488 37810
rect 29012 37466 29040 38490
rect 29104 37913 29132 39782
rect 29184 39432 29236 39438
rect 29184 39374 29236 39380
rect 29196 38758 29224 39374
rect 29276 38888 29328 38894
rect 29276 38830 29328 38836
rect 29184 38752 29236 38758
rect 29184 38694 29236 38700
rect 29288 38214 29316 38830
rect 29552 38480 29604 38486
rect 29552 38422 29604 38428
rect 29276 38208 29328 38214
rect 29276 38150 29328 38156
rect 29564 38010 29592 38422
rect 29932 38350 29960 40326
rect 30116 40050 30144 41414
rect 30208 40934 30236 41618
rect 30392 41070 30420 41958
rect 32128 41676 32180 41682
rect 32128 41618 32180 41624
rect 32140 41206 32168 41618
rect 32772 41472 32824 41478
rect 32772 41414 32824 41420
rect 30932 41200 30984 41206
rect 30932 41142 30984 41148
rect 32128 41200 32180 41206
rect 32128 41142 32180 41148
rect 30380 41064 30432 41070
rect 30380 41006 30432 41012
rect 30196 40928 30248 40934
rect 30196 40870 30248 40876
rect 30208 40769 30236 40870
rect 30194 40760 30250 40769
rect 30194 40695 30250 40704
rect 30196 40656 30248 40662
rect 30196 40598 30248 40604
rect 30104 40044 30156 40050
rect 30104 39986 30156 39992
rect 30012 39840 30064 39846
rect 30012 39782 30064 39788
rect 30024 39284 30052 39782
rect 30116 39642 30144 39986
rect 30208 39914 30236 40598
rect 30196 39908 30248 39914
rect 30196 39850 30248 39856
rect 30104 39636 30156 39642
rect 30104 39578 30156 39584
rect 30944 39545 30972 41142
rect 31668 40996 31720 41002
rect 31668 40938 31720 40944
rect 31484 40928 31536 40934
rect 31484 40870 31536 40876
rect 31024 40520 31076 40526
rect 31024 40462 31076 40468
rect 31036 40186 31064 40462
rect 31024 40180 31076 40186
rect 31024 40122 31076 40128
rect 30930 39536 30986 39545
rect 30930 39471 30932 39480
rect 30984 39471 30986 39480
rect 30932 39442 30984 39448
rect 30104 39296 30156 39302
rect 30024 39256 30104 39284
rect 30104 39238 30156 39244
rect 30748 39296 30800 39302
rect 30748 39238 30800 39244
rect 30012 38888 30064 38894
rect 30012 38830 30064 38836
rect 29920 38344 29972 38350
rect 29920 38286 29972 38292
rect 29932 38010 29960 38286
rect 29552 38004 29604 38010
rect 29552 37946 29604 37952
rect 29920 38004 29972 38010
rect 29920 37946 29972 37952
rect 29090 37904 29146 37913
rect 29090 37839 29146 37848
rect 30024 37788 30052 38830
rect 30116 38486 30144 39238
rect 30656 39092 30708 39098
rect 30656 39034 30708 39040
rect 30668 38826 30696 39034
rect 30760 38894 30788 39238
rect 30748 38888 30800 38894
rect 30748 38830 30800 38836
rect 30656 38820 30708 38826
rect 30656 38762 30708 38768
rect 30288 38548 30340 38554
rect 30288 38490 30340 38496
rect 30104 38480 30156 38486
rect 30104 38422 30156 38428
rect 30194 37904 30250 37913
rect 30194 37839 30250 37848
rect 30104 37800 30156 37806
rect 30024 37760 30104 37788
rect 29736 37732 29788 37738
rect 29736 37674 29788 37680
rect 29000 37460 29052 37466
rect 29000 37402 29052 37408
rect 29644 37460 29696 37466
rect 29644 37402 29696 37408
rect 28632 37392 28684 37398
rect 28632 37334 28684 37340
rect 28540 37256 28592 37262
rect 28446 37224 28502 37233
rect 28540 37198 28592 37204
rect 28446 37159 28502 37168
rect 28356 36236 28408 36242
rect 28356 36178 28408 36184
rect 28448 36236 28500 36242
rect 28448 36178 28500 36184
rect 28368 36106 28396 36178
rect 28356 36100 28408 36106
rect 28356 36042 28408 36048
rect 28368 35698 28396 36042
rect 28460 35834 28488 36178
rect 28552 36174 28580 37198
rect 28644 36854 28672 37334
rect 28816 37256 28868 37262
rect 28816 37198 28868 37204
rect 28632 36848 28684 36854
rect 28632 36790 28684 36796
rect 28540 36168 28592 36174
rect 28540 36110 28592 36116
rect 28448 35828 28500 35834
rect 28448 35770 28500 35776
rect 28828 35766 28856 37198
rect 29656 36650 29684 37402
rect 29644 36644 29696 36650
rect 29644 36586 29696 36592
rect 29000 36576 29052 36582
rect 29000 36518 29052 36524
rect 29012 36310 29040 36518
rect 29656 36310 29684 36586
rect 29000 36304 29052 36310
rect 29000 36246 29052 36252
rect 29644 36304 29696 36310
rect 29644 36246 29696 36252
rect 29460 36236 29512 36242
rect 29460 36178 29512 36184
rect 28816 35760 28868 35766
rect 28816 35702 28868 35708
rect 28172 35692 28224 35698
rect 28172 35634 28224 35640
rect 28356 35692 28408 35698
rect 28356 35634 28408 35640
rect 28724 35692 28776 35698
rect 28724 35634 28776 35640
rect 28184 34950 28212 35634
rect 28736 35601 28764 35634
rect 28722 35592 28778 35601
rect 28722 35527 28778 35536
rect 28724 35488 28776 35494
rect 28724 35430 28776 35436
rect 28736 35086 28764 35430
rect 29472 35154 29500 36178
rect 29552 36168 29604 36174
rect 29552 36110 29604 36116
rect 29564 35834 29592 36110
rect 29656 35834 29684 36246
rect 29552 35828 29604 35834
rect 29552 35770 29604 35776
rect 29644 35828 29696 35834
rect 29644 35770 29696 35776
rect 29564 35222 29592 35770
rect 29552 35216 29604 35222
rect 29552 35158 29604 35164
rect 29000 35148 29052 35154
rect 29000 35090 29052 35096
rect 29460 35148 29512 35154
rect 29460 35090 29512 35096
rect 28724 35080 28776 35086
rect 28724 35022 28776 35028
rect 28172 34944 28224 34950
rect 28172 34886 28224 34892
rect 28184 34746 28212 34886
rect 28172 34740 28224 34746
rect 28172 34682 28224 34688
rect 29012 34678 29040 35090
rect 28356 34672 28408 34678
rect 28356 34614 28408 34620
rect 29000 34672 29052 34678
rect 29000 34614 29052 34620
rect 27712 33924 27764 33930
rect 27712 33866 27764 33872
rect 27804 33924 27856 33930
rect 27804 33866 27856 33872
rect 27620 33652 27672 33658
rect 27620 33594 27672 33600
rect 27816 33590 27844 33866
rect 27804 33584 27856 33590
rect 27804 33526 27856 33532
rect 27528 33448 27580 33454
rect 27528 33390 27580 33396
rect 28264 33448 28316 33454
rect 28264 33390 28316 33396
rect 28276 32978 28304 33390
rect 28080 32972 28132 32978
rect 28080 32914 28132 32920
rect 28264 32972 28316 32978
rect 28264 32914 28316 32920
rect 27436 32836 27488 32842
rect 27436 32778 27488 32784
rect 27988 32768 28040 32774
rect 27988 32710 28040 32716
rect 28000 32570 28028 32710
rect 27988 32564 28040 32570
rect 27988 32506 28040 32512
rect 27436 32428 27488 32434
rect 27436 32370 27488 32376
rect 26608 32292 26660 32298
rect 26608 32234 26660 32240
rect 26620 31958 26648 32234
rect 27448 32230 27476 32370
rect 27528 32292 27580 32298
rect 27528 32234 27580 32240
rect 26700 32224 26752 32230
rect 26700 32166 26752 32172
rect 27436 32224 27488 32230
rect 27436 32166 27488 32172
rect 26608 31952 26660 31958
rect 26608 31894 26660 31900
rect 26712 31822 26740 32166
rect 26700 31816 26752 31822
rect 26700 31758 26752 31764
rect 27160 31816 27212 31822
rect 27160 31758 27212 31764
rect 27068 30592 27120 30598
rect 27068 30534 27120 30540
rect 26608 29708 26660 29714
rect 26528 29668 26608 29696
rect 26608 29650 26660 29656
rect 26620 29034 26648 29650
rect 27080 29578 27108 30534
rect 27068 29572 27120 29578
rect 27068 29514 27120 29520
rect 26608 29028 26660 29034
rect 26608 28970 26660 28976
rect 26620 28937 26648 28970
rect 26606 28928 26662 28937
rect 26606 28863 26662 28872
rect 26700 28688 26752 28694
rect 26700 28630 26752 28636
rect 26608 28552 26660 28558
rect 26608 28494 26660 28500
rect 26620 28218 26648 28494
rect 26608 28212 26660 28218
rect 26608 28154 26660 28160
rect 26620 27674 26648 28154
rect 26712 28150 26740 28630
rect 26700 28144 26752 28150
rect 26700 28086 26752 28092
rect 26608 27668 26660 27674
rect 26608 27610 26660 27616
rect 27172 27334 27200 31758
rect 27448 31414 27476 32166
rect 27540 31890 27568 32234
rect 27804 32224 27856 32230
rect 27804 32166 27856 32172
rect 27528 31884 27580 31890
rect 27528 31826 27580 31832
rect 27436 31408 27488 31414
rect 27436 31350 27488 31356
rect 27448 30734 27476 31350
rect 27540 30802 27568 31826
rect 27816 31822 27844 32166
rect 27804 31816 27856 31822
rect 27724 31776 27804 31804
rect 27620 31204 27672 31210
rect 27620 31146 27672 31152
rect 27528 30796 27580 30802
rect 27528 30738 27580 30744
rect 27436 30728 27488 30734
rect 27436 30670 27488 30676
rect 27448 30054 27476 30670
rect 27436 30048 27488 30054
rect 27436 29990 27488 29996
rect 27342 28248 27398 28257
rect 27342 28183 27344 28192
rect 27396 28183 27398 28192
rect 27344 28154 27396 28160
rect 27356 28014 27384 28154
rect 27344 28008 27396 28014
rect 27344 27950 27396 27956
rect 27252 27532 27304 27538
rect 27252 27474 27304 27480
rect 27160 27328 27212 27334
rect 27160 27270 27212 27276
rect 26792 27056 26844 27062
rect 26792 26998 26844 27004
rect 26700 26988 26752 26994
rect 26700 26930 26752 26936
rect 26712 26586 26740 26930
rect 26700 26580 26752 26586
rect 26700 26522 26752 26528
rect 26516 26240 26568 26246
rect 26516 26182 26568 26188
rect 26528 25906 26556 26182
rect 26804 25906 26832 26998
rect 26976 26852 27028 26858
rect 26976 26794 27028 26800
rect 26516 25900 26568 25906
rect 26516 25842 26568 25848
rect 26792 25900 26844 25906
rect 26792 25842 26844 25848
rect 26516 25764 26568 25770
rect 26700 25764 26752 25770
rect 26568 25724 26700 25752
rect 26516 25706 26568 25712
rect 26424 25356 26476 25362
rect 26424 25298 26476 25304
rect 25412 25288 25464 25294
rect 25412 25230 25464 25236
rect 25424 24274 25452 25230
rect 26516 25152 26568 25158
rect 26516 25094 26568 25100
rect 25688 24744 25740 24750
rect 25688 24686 25740 24692
rect 25412 24268 25464 24274
rect 25412 24210 25464 24216
rect 25700 24070 25728 24686
rect 26424 24268 26476 24274
rect 26424 24210 26476 24216
rect 25688 24064 25740 24070
rect 25688 24006 25740 24012
rect 25700 23730 25728 24006
rect 26436 23866 26464 24210
rect 26424 23860 26476 23866
rect 26424 23802 26476 23808
rect 25688 23724 25740 23730
rect 25688 23666 25740 23672
rect 26332 23180 26384 23186
rect 26332 23122 26384 23128
rect 25320 23044 25372 23050
rect 25320 22986 25372 22992
rect 25228 22568 25280 22574
rect 25228 22510 25280 22516
rect 26148 22568 26200 22574
rect 26148 22510 26200 22516
rect 24676 22500 24728 22506
rect 24676 22442 24728 22448
rect 24688 22098 24716 22442
rect 25780 22432 25832 22438
rect 25780 22374 25832 22380
rect 24398 22063 24454 22072
rect 24492 22092 24544 22098
rect 24492 22034 24544 22040
rect 24676 22092 24728 22098
rect 24676 22034 24728 22040
rect 24124 22024 24176 22030
rect 24124 21966 24176 21972
rect 24136 21554 24164 21966
rect 24504 21690 24532 22034
rect 24688 21690 24716 22034
rect 24492 21684 24544 21690
rect 24492 21626 24544 21632
rect 24676 21684 24728 21690
rect 24676 21626 24728 21632
rect 24124 21548 24176 21554
rect 24124 21490 24176 21496
rect 24768 21072 24820 21078
rect 24768 21014 24820 21020
rect 24400 20936 24452 20942
rect 24400 20878 24452 20884
rect 23756 20800 23808 20806
rect 23756 20742 23808 20748
rect 23768 20330 23796 20742
rect 23756 20324 23808 20330
rect 23756 20266 23808 20272
rect 23768 19786 23796 20266
rect 23756 19780 23808 19786
rect 23756 19722 23808 19728
rect 24412 19718 24440 20878
rect 24780 20602 24808 21014
rect 24768 20596 24820 20602
rect 24768 20538 24820 20544
rect 25504 20596 25556 20602
rect 25504 20538 25556 20544
rect 25044 19848 25096 19854
rect 25044 19790 25096 19796
rect 24216 19712 24268 19718
rect 24216 19654 24268 19660
rect 24400 19712 24452 19718
rect 24400 19654 24452 19660
rect 24228 19378 24256 19654
rect 24216 19372 24268 19378
rect 24216 19314 24268 19320
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23572 18896 23624 18902
rect 23572 18838 23624 18844
rect 23478 18320 23534 18329
rect 23478 18255 23534 18264
rect 23124 17734 23244 17762
rect 23296 17808 23348 17814
rect 23296 17750 23348 17756
rect 22008 17536 22060 17542
rect 22008 17478 22060 17484
rect 21916 15972 21968 15978
rect 21916 15914 21968 15920
rect 21364 15904 21416 15910
rect 21364 15846 21416 15852
rect 21376 15706 21404 15846
rect 21272 15700 21324 15706
rect 21272 15642 21324 15648
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20916 15026 20944 15438
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20916 13938 20944 14962
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 21088 14952 21140 14958
rect 21088 14894 21140 14900
rect 21008 14618 21036 14894
rect 20996 14612 21048 14618
rect 20996 14554 21048 14560
rect 21100 14482 21128 14894
rect 21284 14890 21312 15642
rect 21272 14884 21324 14890
rect 21272 14826 21324 14832
rect 21088 14476 21140 14482
rect 21088 14418 21140 14424
rect 21100 14006 21128 14418
rect 21088 14000 21140 14006
rect 21088 13942 21140 13948
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 21008 12850 21036 13466
rect 21100 13394 21128 13942
rect 21088 13388 21140 13394
rect 21088 13330 21140 13336
rect 21180 13388 21232 13394
rect 21180 13330 21232 13336
rect 20996 12844 21048 12850
rect 20996 12786 21048 12792
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 20812 12096 20864 12102
rect 20812 12038 20864 12044
rect 21008 11762 21036 12174
rect 21088 12096 21140 12102
rect 21192 12084 21220 13330
rect 21284 12714 21312 14826
rect 21732 14476 21784 14482
rect 21732 14418 21784 14424
rect 21744 13734 21772 14418
rect 21732 13728 21784 13734
rect 21732 13670 21784 13676
rect 21272 12708 21324 12714
rect 21272 12650 21324 12656
rect 21284 12374 21312 12650
rect 21272 12368 21324 12374
rect 21272 12310 21324 12316
rect 21140 12056 21220 12084
rect 21088 12038 21140 12044
rect 21100 11830 21128 12038
rect 21284 11898 21312 12310
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 21088 11824 21140 11830
rect 21088 11766 21140 11772
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 20812 11688 20864 11694
rect 20812 11630 20864 11636
rect 20720 11280 20772 11286
rect 20720 11222 20772 11228
rect 20732 10810 20760 11222
rect 20824 11014 20852 11630
rect 20812 11008 20864 11014
rect 20812 10950 20864 10956
rect 20720 10804 20772 10810
rect 20456 8758 20576 8786
rect 20640 10764 20720 10792
rect 20456 8430 20484 8758
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20548 6186 20576 8570
rect 20536 6180 20588 6186
rect 20536 6122 20588 6128
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20272 5166 20300 5306
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20352 5160 20404 5166
rect 20352 5102 20404 5108
rect 20534 5128 20590 5137
rect 20364 4826 20392 5102
rect 20534 5063 20590 5072
rect 20352 4820 20404 4826
rect 20352 4762 20404 4768
rect 19984 4684 20036 4690
rect 19984 4626 20036 4632
rect 19892 4072 19944 4078
rect 19892 4014 19944 4020
rect 20548 4010 20576 5063
rect 20640 4622 20668 10764
rect 20720 10746 20772 10752
rect 20824 7449 20852 10950
rect 20904 10600 20956 10606
rect 20904 10542 20956 10548
rect 20916 9722 20944 10542
rect 20996 10532 21048 10538
rect 20996 10474 21048 10480
rect 21008 9994 21036 10474
rect 20996 9988 21048 9994
rect 20996 9930 21048 9936
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 20916 9518 20944 9658
rect 20904 9512 20956 9518
rect 20904 9454 20956 9460
rect 20916 8634 20944 9454
rect 21008 9382 21036 9930
rect 21100 9926 21128 11766
rect 21548 10532 21600 10538
rect 21548 10474 21600 10480
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 21088 9920 21140 9926
rect 21088 9862 21140 9868
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 20810 7440 20866 7449
rect 20810 7375 20866 7384
rect 20812 7336 20864 7342
rect 20812 7278 20864 7284
rect 20824 6866 20852 7278
rect 20812 6860 20864 6866
rect 20812 6802 20864 6808
rect 21008 6746 21036 9318
rect 21100 7954 21128 9862
rect 21468 9178 21496 10066
rect 21456 9172 21508 9178
rect 21456 9114 21508 9120
rect 21560 8974 21588 10474
rect 21744 9994 21772 13670
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21836 10130 21864 12582
rect 22020 12442 22048 17478
rect 23124 17202 23152 17734
rect 23204 17672 23256 17678
rect 23204 17614 23256 17620
rect 23112 17196 23164 17202
rect 23112 17138 23164 17144
rect 23216 16794 23244 17614
rect 23308 17338 23336 17750
rect 23296 17332 23348 17338
rect 23296 17274 23348 17280
rect 23584 16998 23612 18838
rect 23676 18358 23704 18906
rect 23848 18420 23900 18426
rect 23848 18362 23900 18368
rect 23664 18352 23716 18358
rect 23664 18294 23716 18300
rect 23860 18154 23888 18362
rect 24228 18290 24256 19314
rect 24412 19242 24440 19654
rect 24400 19236 24452 19242
rect 24400 19178 24452 19184
rect 24216 18284 24268 18290
rect 24216 18226 24268 18232
rect 23848 18148 23900 18154
rect 23848 18090 23900 18096
rect 24228 18086 24256 18226
rect 24216 18080 24268 18086
rect 24216 18022 24268 18028
rect 24412 17814 24440 19178
rect 24584 18828 24636 18834
rect 24584 18770 24636 18776
rect 24596 18426 24624 18770
rect 24860 18760 24912 18766
rect 24860 18702 24912 18708
rect 24584 18420 24636 18426
rect 24584 18362 24636 18368
rect 24872 17814 24900 18702
rect 25056 18630 25084 19790
rect 25516 19242 25544 20538
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 25608 19378 25636 19790
rect 25596 19372 25648 19378
rect 25596 19314 25648 19320
rect 25412 19236 25464 19242
rect 25412 19178 25464 19184
rect 25504 19236 25556 19242
rect 25504 19178 25556 19184
rect 25424 18970 25452 19178
rect 25412 18964 25464 18970
rect 25412 18906 25464 18912
rect 25044 18624 25096 18630
rect 25044 18566 25096 18572
rect 24952 18148 25004 18154
rect 24952 18090 25004 18096
rect 24400 17808 24452 17814
rect 24400 17750 24452 17756
rect 24860 17808 24912 17814
rect 24860 17750 24912 17756
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 23756 17060 23808 17066
rect 23756 17002 23808 17008
rect 23572 16992 23624 16998
rect 23572 16934 23624 16940
rect 23768 16794 23796 17002
rect 24780 16794 24808 17614
rect 24872 17338 24900 17750
rect 24860 17332 24912 17338
rect 24860 17274 24912 17280
rect 23204 16788 23256 16794
rect 23204 16730 23256 16736
rect 23756 16788 23808 16794
rect 23756 16730 23808 16736
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 22836 16720 22888 16726
rect 22888 16680 22968 16708
rect 22836 16662 22888 16668
rect 22284 16516 22336 16522
rect 22284 16458 22336 16464
rect 22100 16448 22152 16454
rect 22100 16390 22152 16396
rect 22112 16114 22140 16390
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 22296 15706 22324 16458
rect 22940 16182 22968 16680
rect 22928 16176 22980 16182
rect 22928 16118 22980 16124
rect 22744 15972 22796 15978
rect 22744 15914 22796 15920
rect 22284 15700 22336 15706
rect 22284 15642 22336 15648
rect 22560 15564 22612 15570
rect 22560 15506 22612 15512
rect 22572 14822 22600 15506
rect 22652 15360 22704 15366
rect 22652 15302 22704 15308
rect 22560 14816 22612 14822
rect 22560 14758 22612 14764
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22296 13734 22324 14350
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 22008 12436 22060 12442
rect 22008 12378 22060 12384
rect 22296 10266 22324 13670
rect 22572 12442 22600 14758
rect 22664 13530 22692 15302
rect 22756 14550 22784 15914
rect 22940 15910 22968 16118
rect 23216 16114 23244 16730
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 23204 16108 23256 16114
rect 23204 16050 23256 16056
rect 22928 15904 22980 15910
rect 22928 15846 22980 15852
rect 22744 14544 22796 14550
rect 22744 14486 22796 14492
rect 22756 14414 22784 14486
rect 22744 14408 22796 14414
rect 22744 14350 22796 14356
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 22652 13524 22704 13530
rect 22652 13466 22704 13472
rect 22664 12986 22692 13466
rect 22756 13190 22784 13806
rect 22836 13456 22888 13462
rect 22940 13444 22968 15846
rect 23308 14550 23336 16390
rect 23400 15910 23428 16594
rect 23768 16454 23796 16730
rect 23756 16448 23808 16454
rect 23756 16390 23808 16396
rect 24308 16448 24360 16454
rect 24308 16390 24360 16396
rect 24320 15978 24348 16390
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 24412 15978 24440 16186
rect 24308 15972 24360 15978
rect 24308 15914 24360 15920
rect 24400 15972 24452 15978
rect 24400 15914 24452 15920
rect 23388 15904 23440 15910
rect 23388 15846 23440 15852
rect 23400 15162 23428 15846
rect 24216 15496 24268 15502
rect 24216 15438 24268 15444
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 24228 15026 24256 15438
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 23388 14952 23440 14958
rect 23388 14894 23440 14900
rect 23756 14952 23808 14958
rect 23756 14894 23808 14900
rect 23296 14544 23348 14550
rect 23124 14504 23296 14532
rect 23020 13728 23072 13734
rect 23020 13670 23072 13676
rect 23032 13462 23060 13670
rect 22888 13416 22968 13444
rect 23020 13456 23072 13462
rect 22836 13398 22888 13404
rect 23020 13398 23072 13404
rect 22744 13184 22796 13190
rect 22744 13126 22796 13132
rect 22652 12980 22704 12986
rect 22652 12922 22704 12928
rect 22848 12918 22876 13398
rect 23124 13326 23152 14504
rect 23296 14486 23348 14492
rect 23400 14482 23428 14894
rect 23768 14618 23796 14894
rect 24228 14618 24256 14962
rect 23756 14612 23808 14618
rect 23756 14554 23808 14560
rect 24216 14612 24268 14618
rect 24216 14554 24268 14560
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 23204 14408 23256 14414
rect 23204 14350 23256 14356
rect 23216 13734 23244 14350
rect 23768 13814 23796 14554
rect 24320 14346 24348 15914
rect 24676 15632 24728 15638
rect 24676 15574 24728 15580
rect 24688 15162 24716 15574
rect 24676 15156 24728 15162
rect 24676 15098 24728 15104
rect 24308 14340 24360 14346
rect 24308 14282 24360 14288
rect 24780 13938 24808 16730
rect 24872 16250 24900 17274
rect 24964 16708 24992 18090
rect 25056 17678 25084 18566
rect 25424 18290 25452 18906
rect 25516 18834 25544 19178
rect 25504 18828 25556 18834
rect 25504 18770 25556 18776
rect 25412 18284 25464 18290
rect 25412 18226 25464 18232
rect 25044 17672 25096 17678
rect 25044 17614 25096 17620
rect 25056 17202 25084 17614
rect 25596 17536 25648 17542
rect 25596 17478 25648 17484
rect 25044 17196 25096 17202
rect 25044 17138 25096 17144
rect 25608 17066 25636 17478
rect 25688 17332 25740 17338
rect 25688 17274 25740 17280
rect 25700 17066 25728 17274
rect 25596 17060 25648 17066
rect 25596 17002 25648 17008
rect 25688 17060 25740 17066
rect 25688 17002 25740 17008
rect 25044 16720 25096 16726
rect 24964 16680 25044 16708
rect 25044 16662 25096 16668
rect 25056 16250 25084 16662
rect 25608 16590 25636 17002
rect 25596 16584 25648 16590
rect 25596 16526 25648 16532
rect 25412 16516 25464 16522
rect 25412 16458 25464 16464
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 25044 16244 25096 16250
rect 25044 16186 25096 16192
rect 24952 15972 25004 15978
rect 24952 15914 25004 15920
rect 24964 15434 24992 15914
rect 25424 15706 25452 16458
rect 25608 16114 25636 16526
rect 25596 16108 25648 16114
rect 25596 16050 25648 16056
rect 25412 15700 25464 15706
rect 25412 15642 25464 15648
rect 24952 15428 25004 15434
rect 24952 15370 25004 15376
rect 25136 14952 25188 14958
rect 25136 14894 25188 14900
rect 25148 14618 25176 14894
rect 25136 14612 25188 14618
rect 25136 14554 25188 14560
rect 24952 14476 25004 14482
rect 24952 14418 25004 14424
rect 25320 14476 25372 14482
rect 25320 14418 25372 14424
rect 24964 14074 24992 14418
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 25332 14006 25360 14418
rect 25320 14000 25372 14006
rect 25320 13942 25372 13948
rect 24768 13932 24820 13938
rect 24768 13874 24820 13880
rect 23676 13786 23796 13814
rect 24032 13796 24084 13802
rect 23204 13728 23256 13734
rect 23204 13670 23256 13676
rect 23112 13320 23164 13326
rect 23676 13297 23704 13786
rect 24032 13738 24084 13744
rect 24124 13796 24176 13802
rect 24124 13738 24176 13744
rect 23112 13262 23164 13268
rect 23662 13288 23718 13297
rect 23662 13223 23718 13232
rect 22928 13184 22980 13190
rect 22928 13126 22980 13132
rect 22836 12912 22888 12918
rect 22836 12854 22888 12860
rect 22560 12436 22612 12442
rect 22560 12378 22612 12384
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22560 11824 22612 11830
rect 22560 11766 22612 11772
rect 22468 11688 22520 11694
rect 22468 11630 22520 11636
rect 22480 11082 22508 11630
rect 22468 11076 22520 11082
rect 22468 11018 22520 11024
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 21824 10124 21876 10130
rect 21824 10066 21876 10072
rect 22100 10056 22152 10062
rect 22100 9998 22152 10004
rect 21732 9988 21784 9994
rect 21732 9930 21784 9936
rect 21916 9920 21968 9926
rect 21916 9862 21968 9868
rect 21732 9716 21784 9722
rect 21732 9658 21784 9664
rect 21744 9382 21772 9658
rect 21928 9586 21956 9862
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 22112 9450 22140 9998
rect 22480 9625 22508 11018
rect 22572 10266 22600 11766
rect 22756 11626 22784 12174
rect 22940 11898 22968 13126
rect 23388 12436 23440 12442
rect 23388 12378 23440 12384
rect 22928 11892 22980 11898
rect 22928 11834 22980 11840
rect 23400 11830 23428 12378
rect 23388 11824 23440 11830
rect 23388 11766 23440 11772
rect 23572 11756 23624 11762
rect 23572 11698 23624 11704
rect 23020 11688 23072 11694
rect 23020 11630 23072 11636
rect 22744 11620 22796 11626
rect 22744 11562 22796 11568
rect 22756 11354 22784 11562
rect 22744 11348 22796 11354
rect 22744 11290 22796 11296
rect 23032 11218 23060 11630
rect 23584 11286 23612 11698
rect 23572 11280 23624 11286
rect 23572 11222 23624 11228
rect 23676 11218 23704 13223
rect 24044 12986 24072 13738
rect 24136 13530 24164 13738
rect 24124 13524 24176 13530
rect 24124 13466 24176 13472
rect 24780 13326 24808 13874
rect 24584 13320 24636 13326
rect 24584 13262 24636 13268
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24596 12986 24624 13262
rect 24032 12980 24084 12986
rect 24032 12922 24084 12928
rect 24584 12980 24636 12986
rect 24584 12922 24636 12928
rect 23940 12776 23992 12782
rect 23940 12718 23992 12724
rect 25136 12776 25188 12782
rect 25136 12718 25188 12724
rect 23952 12442 23980 12718
rect 25148 12442 25176 12718
rect 23940 12436 23992 12442
rect 23940 12378 23992 12384
rect 25136 12436 25188 12442
rect 25136 12378 25188 12384
rect 24860 12300 24912 12306
rect 24860 12242 24912 12248
rect 25228 12300 25280 12306
rect 25228 12242 25280 12248
rect 24216 12096 24268 12102
rect 24216 12038 24268 12044
rect 24228 11762 24256 12038
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24872 11694 24900 12242
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24676 11620 24728 11626
rect 24676 11562 24728 11568
rect 24584 11348 24636 11354
rect 24584 11290 24636 11296
rect 23020 11212 23072 11218
rect 23020 11154 23072 11160
rect 23204 11212 23256 11218
rect 23204 11154 23256 11160
rect 23664 11212 23716 11218
rect 23664 11154 23716 11160
rect 24308 11212 24360 11218
rect 24308 11154 24360 11160
rect 22836 11008 22888 11014
rect 22836 10950 22888 10956
rect 22848 10606 22876 10950
rect 23032 10810 23060 11154
rect 23020 10804 23072 10810
rect 23020 10746 23072 10752
rect 22836 10600 22888 10606
rect 22836 10542 22888 10548
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 22572 9722 22600 10202
rect 22560 9716 22612 9722
rect 22560 9658 22612 9664
rect 22466 9616 22522 9625
rect 22466 9551 22522 9560
rect 22100 9444 22152 9450
rect 22100 9386 22152 9392
rect 21732 9376 21784 9382
rect 21732 9318 21784 9324
rect 21824 9376 21876 9382
rect 21824 9318 21876 9324
rect 21836 9178 21864 9318
rect 21824 9172 21876 9178
rect 21824 9114 21876 9120
rect 21548 8968 21600 8974
rect 21548 8910 21600 8916
rect 22112 8498 22140 9386
rect 22572 9110 22600 9658
rect 22848 9178 22876 10542
rect 23216 10470 23244 11154
rect 24320 10810 24348 11154
rect 24308 10804 24360 10810
rect 24308 10746 24360 10752
rect 23572 10600 23624 10606
rect 23572 10542 23624 10548
rect 23296 10532 23348 10538
rect 23296 10474 23348 10480
rect 22928 10464 22980 10470
rect 22928 10406 22980 10412
rect 23204 10464 23256 10470
rect 23204 10406 23256 10412
rect 22940 9994 22968 10406
rect 23216 10130 23244 10406
rect 23204 10124 23256 10130
rect 23204 10066 23256 10072
rect 22928 9988 22980 9994
rect 22928 9930 22980 9936
rect 23112 9512 23164 9518
rect 23112 9454 23164 9460
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22284 9104 22336 9110
rect 22284 9046 22336 9052
rect 22560 9104 22612 9110
rect 22560 9046 22612 9052
rect 22296 8634 22324 9046
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 22572 8634 22600 8910
rect 22284 8628 22336 8634
rect 22284 8570 22336 8576
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 21364 8492 21416 8498
rect 21364 8434 21416 8440
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 21272 8424 21324 8430
rect 21272 8366 21324 8372
rect 21088 7948 21140 7954
rect 21088 7890 21140 7896
rect 21100 7410 21128 7890
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 20824 6718 21036 6746
rect 20720 5092 20772 5098
rect 20720 5034 20772 5040
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 20640 4282 20668 4558
rect 20628 4276 20680 4282
rect 20628 4218 20680 4224
rect 20732 4010 20760 5034
rect 20824 4154 20852 6718
rect 21192 6254 21220 7482
rect 20904 6248 20956 6254
rect 20904 6190 20956 6196
rect 21180 6248 21232 6254
rect 21180 6190 21232 6196
rect 20916 5778 20944 6190
rect 20996 5908 21048 5914
rect 20996 5850 21048 5856
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 20916 5370 20944 5714
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 20824 4126 20944 4154
rect 21008 4146 21036 5850
rect 21192 5846 21220 6190
rect 21180 5840 21232 5846
rect 21180 5782 21232 5788
rect 21180 5092 21232 5098
rect 21180 5034 21232 5040
rect 20536 4004 20588 4010
rect 20536 3946 20588 3952
rect 20720 4004 20772 4010
rect 20720 3946 20772 3952
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 19892 3596 19944 3602
rect 19892 3538 19944 3544
rect 19904 3194 19932 3538
rect 19892 3188 19944 3194
rect 19892 3130 19944 3136
rect 20732 2922 20760 3946
rect 20916 3602 20944 4126
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 21008 3738 21036 4082
rect 20996 3732 21048 3738
rect 20996 3674 21048 3680
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 20916 3194 20944 3538
rect 21192 3466 21220 5034
rect 21284 4690 21312 8366
rect 21376 7954 21404 8434
rect 21456 8016 21508 8022
rect 21456 7958 21508 7964
rect 21364 7948 21416 7954
rect 21364 7890 21416 7896
rect 21376 7546 21404 7890
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 21376 6322 21404 6598
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 21468 5778 21496 7958
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 21836 7410 21864 7822
rect 22296 7546 22324 8570
rect 23020 8016 23072 8022
rect 23020 7958 23072 7964
rect 22836 7880 22888 7886
rect 22836 7822 22888 7828
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21824 7404 21876 7410
rect 21824 7346 21876 7352
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 21560 6254 21588 7142
rect 21548 6248 21600 6254
rect 21548 6190 21600 6196
rect 21456 5772 21508 5778
rect 21456 5714 21508 5720
rect 21468 5166 21496 5714
rect 21652 5166 21680 7346
rect 22296 7206 22324 7482
rect 22284 7200 22336 7206
rect 22284 7142 22336 7148
rect 22296 6934 22324 7142
rect 22848 7002 22876 7822
rect 23032 7546 23060 7958
rect 23124 7868 23152 9454
rect 23216 7970 23244 10066
rect 23308 8498 23336 10474
rect 23584 10266 23612 10542
rect 23572 10260 23624 10266
rect 23572 10202 23624 10208
rect 23480 10192 23532 10198
rect 23480 10134 23532 10140
rect 23388 9988 23440 9994
rect 23388 9930 23440 9936
rect 23400 9586 23428 9930
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23492 9382 23520 10134
rect 24320 10130 24348 10746
rect 24308 10124 24360 10130
rect 24308 10066 24360 10072
rect 24320 9722 24348 10066
rect 24308 9716 24360 9722
rect 24308 9658 24360 9664
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 24400 9376 24452 9382
rect 24400 9318 24452 9324
rect 23296 8492 23348 8498
rect 23296 8434 23348 8440
rect 23492 8430 23520 9318
rect 24308 9104 24360 9110
rect 24308 9046 24360 9052
rect 24216 8968 24268 8974
rect 24216 8910 24268 8916
rect 23940 8832 23992 8838
rect 23940 8774 23992 8780
rect 23952 8430 23980 8774
rect 24228 8634 24256 8910
rect 24216 8628 24268 8634
rect 24216 8570 24268 8576
rect 24320 8566 24348 9046
rect 24308 8560 24360 8566
rect 24308 8502 24360 8508
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 23480 8424 23532 8430
rect 23480 8366 23532 8372
rect 23940 8424 23992 8430
rect 23940 8366 23992 8372
rect 23216 7942 23612 7970
rect 23388 7880 23440 7886
rect 23124 7840 23244 7868
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 22836 6996 22888 7002
rect 22888 6956 22968 6984
rect 22836 6938 22888 6944
rect 22284 6928 22336 6934
rect 22284 6870 22336 6876
rect 22296 6458 22324 6870
rect 22284 6452 22336 6458
rect 22284 6394 22336 6400
rect 22192 6180 22244 6186
rect 22192 6122 22244 6128
rect 22204 5914 22232 6122
rect 22468 6112 22520 6118
rect 22468 6054 22520 6060
rect 22192 5908 22244 5914
rect 22192 5850 22244 5856
rect 21456 5160 21508 5166
rect 21456 5102 21508 5108
rect 21640 5160 21692 5166
rect 21640 5102 21692 5108
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 21284 4282 21312 4626
rect 21272 4276 21324 4282
rect 21272 4218 21324 4224
rect 21468 4154 21496 5102
rect 22480 4758 22508 6054
rect 22836 5840 22888 5846
rect 22836 5782 22888 5788
rect 22848 5370 22876 5782
rect 22940 5778 22968 6956
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 22940 5370 22968 5714
rect 23112 5704 23164 5710
rect 23112 5646 23164 5652
rect 22836 5364 22888 5370
rect 22836 5306 22888 5312
rect 22928 5364 22980 5370
rect 22928 5306 22980 5312
rect 22560 5228 22612 5234
rect 22560 5170 22612 5176
rect 22572 4826 22600 5170
rect 22836 5160 22888 5166
rect 22836 5102 22888 5108
rect 22560 4820 22612 4826
rect 22560 4762 22612 4768
rect 22468 4752 22520 4758
rect 22468 4694 22520 4700
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 21376 4126 21496 4154
rect 21376 3602 21404 4126
rect 21732 3936 21784 3942
rect 21732 3878 21784 3884
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21180 3460 21232 3466
rect 21180 3402 21232 3408
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 21192 3058 21220 3402
rect 21376 3126 21404 3538
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21364 3120 21416 3126
rect 21364 3062 21416 3068
rect 21180 3052 21232 3058
rect 21180 2994 21232 3000
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 20996 2916 21048 2922
rect 20996 2858 21048 2864
rect 19444 2650 19472 2858
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 21008 2650 21036 2858
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 20996 2644 21048 2650
rect 20996 2586 21048 2592
rect 21468 2514 21496 3470
rect 21456 2508 21508 2514
rect 21456 2450 21508 2456
rect 21744 1737 21772 3878
rect 22204 3602 22232 4558
rect 22572 4282 22600 4762
rect 22560 4276 22612 4282
rect 22560 4218 22612 4224
rect 22652 3664 22704 3670
rect 22652 3606 22704 3612
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 22204 3194 22232 3538
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22664 3126 22692 3606
rect 22652 3120 22704 3126
rect 22652 3062 22704 3068
rect 22664 2922 22692 3062
rect 22652 2916 22704 2922
rect 22652 2858 22704 2864
rect 22100 2848 22152 2854
rect 22100 2790 22152 2796
rect 22112 2145 22140 2790
rect 22848 2650 22876 5102
rect 23124 4690 23152 5646
rect 23112 4684 23164 4690
rect 23112 4626 23164 4632
rect 22928 4480 22980 4486
rect 22928 4422 22980 4428
rect 22940 4078 22968 4422
rect 22928 4072 22980 4078
rect 22928 4014 22980 4020
rect 23124 3194 23152 4626
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 22836 2644 22888 2650
rect 22836 2586 22888 2592
rect 22098 2136 22154 2145
rect 22098 2071 22154 2080
rect 21730 1728 21786 1737
rect 21730 1663 21786 1672
rect 19522 82 19578 480
rect 19352 54 19578 82
rect 5262 0 5318 54
rect 8850 0 8906 54
rect 12438 0 12494 54
rect 16026 0 16082 54
rect 19522 0 19578 54
rect 23110 82 23166 480
rect 23216 82 23244 7840
rect 23388 7822 23440 7828
rect 23400 5370 23428 7822
rect 23478 7440 23534 7449
rect 23478 7375 23534 7384
rect 23492 6866 23520 7375
rect 23480 6860 23532 6866
rect 23480 6802 23532 6808
rect 23492 6458 23520 6802
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23492 5846 23520 6394
rect 23584 6390 23612 7942
rect 23664 7744 23716 7750
rect 23664 7686 23716 7692
rect 23676 7410 23704 7686
rect 23756 7472 23808 7478
rect 23756 7414 23808 7420
rect 23664 7404 23716 7410
rect 23664 7346 23716 7352
rect 23676 7002 23704 7346
rect 23768 7274 23796 7414
rect 23756 7268 23808 7274
rect 23756 7210 23808 7216
rect 23664 6996 23716 7002
rect 23664 6938 23716 6944
rect 23952 6866 23980 8366
rect 24044 8090 24072 8434
rect 24320 8362 24348 8502
rect 24308 8356 24360 8362
rect 24308 8298 24360 8304
rect 24032 8084 24084 8090
rect 24032 8026 24084 8032
rect 24412 8022 24440 9318
rect 24400 8016 24452 8022
rect 24400 7958 24452 7964
rect 24308 7880 24360 7886
rect 24308 7822 24360 7828
rect 24320 7546 24348 7822
rect 24412 7546 24440 7958
rect 24308 7540 24360 7546
rect 24308 7482 24360 7488
rect 24400 7540 24452 7546
rect 24400 7482 24452 7488
rect 24320 7002 24348 7482
rect 24492 7336 24544 7342
rect 24492 7278 24544 7284
rect 24308 6996 24360 7002
rect 24308 6938 24360 6944
rect 24504 6866 24532 7278
rect 23940 6860 23992 6866
rect 23940 6802 23992 6808
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 23572 6384 23624 6390
rect 23572 6326 23624 6332
rect 23952 6322 23980 6802
rect 23940 6316 23992 6322
rect 23940 6258 23992 6264
rect 23952 5914 23980 6258
rect 23940 5908 23992 5914
rect 23940 5850 23992 5856
rect 23480 5840 23532 5846
rect 23480 5782 23532 5788
rect 24124 5704 24176 5710
rect 24124 5646 24176 5652
rect 24136 5370 24164 5646
rect 23388 5364 23440 5370
rect 23388 5306 23440 5312
rect 24124 5364 24176 5370
rect 24124 5306 24176 5312
rect 23664 5092 23716 5098
rect 23664 5034 23716 5040
rect 23676 4078 23704 5034
rect 24136 4154 24164 5306
rect 24596 5166 24624 11290
rect 24688 10538 24716 11562
rect 25240 11558 25268 12242
rect 25228 11552 25280 11558
rect 25228 11494 25280 11500
rect 25044 11212 25096 11218
rect 25044 11154 25096 11160
rect 24860 10600 24912 10606
rect 24860 10542 24912 10548
rect 24676 10532 24728 10538
rect 24676 10474 24728 10480
rect 24872 10198 24900 10542
rect 24860 10192 24912 10198
rect 24860 10134 24912 10140
rect 24860 9444 24912 9450
rect 24860 9386 24912 9392
rect 24872 8362 24900 9386
rect 24952 8968 25004 8974
rect 24952 8910 25004 8916
rect 24860 8356 24912 8362
rect 24860 8298 24912 8304
rect 24872 8265 24900 8298
rect 24858 8256 24914 8265
rect 24858 8191 24914 8200
rect 24964 8129 24992 8910
rect 24950 8120 25006 8129
rect 24950 8055 25006 8064
rect 24964 8022 24992 8055
rect 24952 8016 25004 8022
rect 24952 7958 25004 7964
rect 25056 7818 25084 11154
rect 25240 10985 25268 11494
rect 25332 11218 25360 13942
rect 25412 13864 25464 13870
rect 25464 13824 25636 13852
rect 25412 13806 25464 13812
rect 25608 13190 25636 13824
rect 25792 13814 25820 22374
rect 26160 21622 26188 22510
rect 26344 22506 26372 23122
rect 26424 23112 26476 23118
rect 26528 23100 26556 25094
rect 26620 24954 26648 25724
rect 26700 25706 26752 25712
rect 26804 25498 26832 25842
rect 26884 25696 26936 25702
rect 26884 25638 26936 25644
rect 26792 25492 26844 25498
rect 26792 25434 26844 25440
rect 26608 24948 26660 24954
rect 26608 24890 26660 24896
rect 26476 23072 26556 23100
rect 26424 23054 26476 23060
rect 26332 22500 26384 22506
rect 26332 22442 26384 22448
rect 26148 21616 26200 21622
rect 26148 21558 26200 21564
rect 26148 21480 26200 21486
rect 26148 21422 26200 21428
rect 26160 21146 26188 21422
rect 26240 21412 26292 21418
rect 26240 21354 26292 21360
rect 26148 21140 26200 21146
rect 26148 21082 26200 21088
rect 26148 20256 26200 20262
rect 26148 20198 26200 20204
rect 26160 20058 26188 20198
rect 26148 20052 26200 20058
rect 26148 19994 26200 20000
rect 26252 19990 26280 21354
rect 26344 21010 26372 22442
rect 26424 22432 26476 22438
rect 26424 22374 26476 22380
rect 26436 22166 26464 22374
rect 26424 22160 26476 22166
rect 26424 22102 26476 22108
rect 26332 21004 26384 21010
rect 26332 20946 26384 20952
rect 26344 20058 26372 20946
rect 26528 20466 26556 23072
rect 26700 22976 26752 22982
rect 26700 22918 26752 22924
rect 26516 20460 26568 20466
rect 26516 20402 26568 20408
rect 26712 20398 26740 22918
rect 26896 22080 26924 25638
rect 26988 23186 27016 26794
rect 27172 26246 27200 27270
rect 27264 26790 27292 27474
rect 27448 27452 27476 29990
rect 27540 29850 27568 30738
rect 27632 30598 27660 31146
rect 27724 31142 27752 31776
rect 27804 31758 27856 31764
rect 28000 31686 28028 32506
rect 28092 31958 28120 32914
rect 28264 32768 28316 32774
rect 28264 32710 28316 32716
rect 28276 32366 28304 32710
rect 28264 32360 28316 32366
rect 28264 32302 28316 32308
rect 28080 31952 28132 31958
rect 28080 31894 28132 31900
rect 28172 31748 28224 31754
rect 28172 31690 28224 31696
rect 27988 31680 28040 31686
rect 27988 31622 28040 31628
rect 28000 31346 28028 31622
rect 27988 31340 28040 31346
rect 27988 31282 28040 31288
rect 28184 31278 28212 31690
rect 28172 31272 28224 31278
rect 28172 31214 28224 31220
rect 27712 31136 27764 31142
rect 27712 31078 27764 31084
rect 27620 30592 27672 30598
rect 27620 30534 27672 30540
rect 27632 30054 27660 30534
rect 27620 30048 27672 30054
rect 27620 29990 27672 29996
rect 27528 29844 27580 29850
rect 27528 29786 27580 29792
rect 27632 29170 27660 29990
rect 27620 29164 27672 29170
rect 27620 29106 27672 29112
rect 27528 27464 27580 27470
rect 27448 27424 27528 27452
rect 27528 27406 27580 27412
rect 27540 26790 27568 27406
rect 27632 27334 27660 29106
rect 27724 28422 27752 31078
rect 28276 30938 28304 32302
rect 28264 30932 28316 30938
rect 28264 30874 28316 30880
rect 28368 29714 28396 34614
rect 29472 34610 29500 35090
rect 28540 34604 28592 34610
rect 28540 34546 28592 34552
rect 29460 34604 29512 34610
rect 29460 34546 29512 34552
rect 28448 32768 28500 32774
rect 28552 32756 28580 34546
rect 29656 34134 29684 35770
rect 29748 35630 29776 37674
rect 30024 37466 30052 37760
rect 30104 37742 30156 37748
rect 30208 37652 30236 37839
rect 30116 37624 30236 37652
rect 30012 37460 30064 37466
rect 30012 37402 30064 37408
rect 30024 36242 30052 37402
rect 30012 36236 30064 36242
rect 30012 36178 30064 36184
rect 29736 35624 29788 35630
rect 29736 35566 29788 35572
rect 29828 34400 29880 34406
rect 29828 34342 29880 34348
rect 29644 34128 29696 34134
rect 29644 34070 29696 34076
rect 29460 33992 29512 33998
rect 29460 33934 29512 33940
rect 28814 33824 28870 33833
rect 28814 33759 28870 33768
rect 28632 33448 28684 33454
rect 28632 33390 28684 33396
rect 28644 33017 28672 33390
rect 28828 33046 28856 33759
rect 29472 33318 29500 33934
rect 29656 33658 29684 34070
rect 29644 33652 29696 33658
rect 29644 33594 29696 33600
rect 29460 33312 29512 33318
rect 29460 33254 29512 33260
rect 29840 33046 29868 34342
rect 28816 33040 28868 33046
rect 28630 33008 28686 33017
rect 28816 32982 28868 32988
rect 29828 33040 29880 33046
rect 29828 32982 29880 32988
rect 28630 32943 28686 32952
rect 28632 32904 28684 32910
rect 28632 32846 28684 32852
rect 28500 32728 28580 32756
rect 28448 32710 28500 32716
rect 28460 31958 28488 32710
rect 28644 32230 28672 32846
rect 30012 32768 30064 32774
rect 30012 32710 30064 32716
rect 30024 32298 30052 32710
rect 29920 32292 29972 32298
rect 29920 32234 29972 32240
rect 30012 32292 30064 32298
rect 30012 32234 30064 32240
rect 28632 32224 28684 32230
rect 28632 32166 28684 32172
rect 28448 31952 28500 31958
rect 28448 31894 28500 31900
rect 29552 31816 29604 31822
rect 29552 31758 29604 31764
rect 29276 31680 29328 31686
rect 29276 31622 29328 31628
rect 29288 31346 29316 31622
rect 29276 31340 29328 31346
rect 29276 31282 29328 31288
rect 28632 31272 28684 31278
rect 28632 31214 28684 31220
rect 28722 31240 28778 31249
rect 28644 30734 28672 31214
rect 28722 31175 28778 31184
rect 28736 31142 28764 31175
rect 28724 31136 28776 31142
rect 28724 31078 28776 31084
rect 29000 31136 29052 31142
rect 29000 31078 29052 31084
rect 28632 30728 28684 30734
rect 28632 30670 28684 30676
rect 28538 30288 28594 30297
rect 28538 30223 28594 30232
rect 28356 29708 28408 29714
rect 28356 29650 28408 29656
rect 28368 29306 28396 29650
rect 28448 29572 28500 29578
rect 28448 29514 28500 29520
rect 28356 29300 28408 29306
rect 28356 29242 28408 29248
rect 27804 29096 27856 29102
rect 27804 29038 27856 29044
rect 27712 28416 27764 28422
rect 27712 28358 27764 28364
rect 27620 27328 27672 27334
rect 27620 27270 27672 27276
rect 27632 27130 27660 27270
rect 27620 27124 27672 27130
rect 27620 27066 27672 27072
rect 27252 26784 27304 26790
rect 27252 26726 27304 26732
rect 27528 26784 27580 26790
rect 27528 26726 27580 26732
rect 27264 26450 27292 26726
rect 27252 26444 27304 26450
rect 27252 26386 27304 26392
rect 27160 26240 27212 26246
rect 27160 26182 27212 26188
rect 27068 25356 27120 25362
rect 27068 25298 27120 25304
rect 27080 24954 27108 25298
rect 27068 24948 27120 24954
rect 27068 24890 27120 24896
rect 26976 23180 27028 23186
rect 26976 23122 27028 23128
rect 26976 22092 27028 22098
rect 26896 22052 26976 22080
rect 26976 22034 27028 22040
rect 26988 21350 27016 22034
rect 27080 22030 27108 24890
rect 27068 22024 27120 22030
rect 27068 21966 27120 21972
rect 27172 21690 27200 26182
rect 27264 25158 27292 26386
rect 27252 25152 27304 25158
rect 27252 25094 27304 25100
rect 27436 24744 27488 24750
rect 27436 24686 27488 24692
rect 27448 24313 27476 24686
rect 27434 24304 27490 24313
rect 27434 24239 27490 24248
rect 27448 24206 27476 24239
rect 27436 24200 27488 24206
rect 27436 24142 27488 24148
rect 27344 24064 27396 24070
rect 27344 24006 27396 24012
rect 27160 21684 27212 21690
rect 27160 21626 27212 21632
rect 26976 21344 27028 21350
rect 26976 21286 27028 21292
rect 26988 20942 27016 21286
rect 27172 21146 27200 21626
rect 27160 21140 27212 21146
rect 27160 21082 27212 21088
rect 26884 20936 26936 20942
rect 26884 20878 26936 20884
rect 26976 20936 27028 20942
rect 26976 20878 27028 20884
rect 26700 20392 26752 20398
rect 26700 20334 26752 20340
rect 26332 20052 26384 20058
rect 26332 19994 26384 20000
rect 26240 19984 26292 19990
rect 26240 19926 26292 19932
rect 26252 19514 26280 19926
rect 26896 19854 26924 20878
rect 27356 19922 27384 24006
rect 27448 20874 27476 24142
rect 27540 22030 27568 26726
rect 27620 26376 27672 26382
rect 27724 26364 27752 28358
rect 27672 26336 27752 26364
rect 27620 26318 27672 26324
rect 27632 25702 27660 26318
rect 27816 26246 27844 29038
rect 27896 28620 27948 28626
rect 27896 28562 27948 28568
rect 27908 27878 27936 28562
rect 27896 27872 27948 27878
rect 27896 27814 27948 27820
rect 28264 27872 28316 27878
rect 28264 27814 28316 27820
rect 27908 26761 27936 27814
rect 27894 26752 27950 26761
rect 27894 26687 27950 26696
rect 27804 26240 27856 26246
rect 27804 26182 27856 26188
rect 27816 25702 27844 26182
rect 27620 25696 27672 25702
rect 27620 25638 27672 25644
rect 27804 25696 27856 25702
rect 27804 25638 27856 25644
rect 27620 23860 27672 23866
rect 27620 23802 27672 23808
rect 27632 23662 27660 23802
rect 27620 23656 27672 23662
rect 27620 23598 27672 23604
rect 27712 23112 27764 23118
rect 27712 23054 27764 23060
rect 27724 22642 27752 23054
rect 27620 22636 27672 22642
rect 27620 22578 27672 22584
rect 27712 22636 27764 22642
rect 27712 22578 27764 22584
rect 27632 22545 27660 22578
rect 27618 22536 27674 22545
rect 27618 22471 27674 22480
rect 27528 22024 27580 22030
rect 27528 21966 27580 21972
rect 27712 22024 27764 22030
rect 27712 21966 27764 21972
rect 27620 21956 27672 21962
rect 27620 21898 27672 21904
rect 27528 21616 27580 21622
rect 27528 21558 27580 21564
rect 27540 21350 27568 21558
rect 27632 21486 27660 21898
rect 27724 21554 27752 21966
rect 27816 21604 27844 25638
rect 27908 24886 27936 26687
rect 27988 26512 28040 26518
rect 27988 26454 28040 26460
rect 27896 24880 27948 24886
rect 27896 24822 27948 24828
rect 27908 23866 27936 24822
rect 28000 24750 28028 26454
rect 28172 25288 28224 25294
rect 28172 25230 28224 25236
rect 27988 24744 28040 24750
rect 27988 24686 28040 24692
rect 28000 24410 28028 24686
rect 28184 24682 28212 25230
rect 28276 24721 28304 27814
rect 28356 26920 28408 26926
rect 28460 26908 28488 29514
rect 28408 26880 28488 26908
rect 28356 26862 28408 26868
rect 28368 26586 28396 26862
rect 28356 26580 28408 26586
rect 28356 26522 28408 26528
rect 28552 26042 28580 30223
rect 28644 29696 28672 30670
rect 28816 30048 28868 30054
rect 28816 29990 28868 29996
rect 28724 29708 28776 29714
rect 28644 29668 28724 29696
rect 28724 29650 28776 29656
rect 28736 29306 28764 29650
rect 28724 29300 28776 29306
rect 28724 29242 28776 29248
rect 28736 28626 28764 29242
rect 28724 28620 28776 28626
rect 28724 28562 28776 28568
rect 28632 28212 28684 28218
rect 28632 28154 28684 28160
rect 28540 26036 28592 26042
rect 28540 25978 28592 25984
rect 28356 25900 28408 25906
rect 28356 25842 28408 25848
rect 28368 25498 28396 25842
rect 28552 25838 28580 25978
rect 28540 25832 28592 25838
rect 28540 25774 28592 25780
rect 28540 25696 28592 25702
rect 28540 25638 28592 25644
rect 28356 25492 28408 25498
rect 28356 25434 28408 25440
rect 28262 24712 28318 24721
rect 28172 24676 28224 24682
rect 28262 24647 28318 24656
rect 28172 24618 28224 24624
rect 28184 24410 28212 24618
rect 28264 24608 28316 24614
rect 28368 24596 28396 25434
rect 28552 25294 28580 25638
rect 28540 25288 28592 25294
rect 28540 25230 28592 25236
rect 28316 24568 28396 24596
rect 28264 24550 28316 24556
rect 27988 24404 28040 24410
rect 27988 24346 28040 24352
rect 28172 24404 28224 24410
rect 28172 24346 28224 24352
rect 27896 23860 27948 23866
rect 27896 23802 27948 23808
rect 28000 23662 28028 24346
rect 27988 23656 28040 23662
rect 27988 23598 28040 23604
rect 27896 23316 27948 23322
rect 28000 23304 28028 23598
rect 28080 23588 28132 23594
rect 28080 23530 28132 23536
rect 27948 23276 28028 23304
rect 27896 23258 27948 23264
rect 28000 22574 28028 23276
rect 27988 22568 28040 22574
rect 27988 22510 28040 22516
rect 28092 22030 28120 23530
rect 28276 23254 28304 24550
rect 28264 23248 28316 23254
rect 28264 23190 28316 23196
rect 28276 22778 28304 23190
rect 28644 23066 28672 28154
rect 28724 27532 28776 27538
rect 28724 27474 28776 27480
rect 28736 27402 28764 27474
rect 28724 27396 28776 27402
rect 28724 27338 28776 27344
rect 28736 27130 28764 27338
rect 28724 27124 28776 27130
rect 28724 27066 28776 27072
rect 28736 27033 28764 27066
rect 28722 27024 28778 27033
rect 28722 26959 28778 26968
rect 28736 24274 28764 26959
rect 28828 25838 28856 29990
rect 28908 29096 28960 29102
rect 28908 29038 28960 29044
rect 28920 28694 28948 29038
rect 29012 28966 29040 31078
rect 29092 30796 29144 30802
rect 29092 30738 29144 30744
rect 29104 30258 29132 30738
rect 29564 30666 29592 31758
rect 29932 30977 29960 32234
rect 30024 31958 30052 32234
rect 30012 31952 30064 31958
rect 30012 31894 30064 31900
rect 30024 31482 30052 31894
rect 30012 31476 30064 31482
rect 30012 31418 30064 31424
rect 29918 30968 29974 30977
rect 30024 30938 30052 31418
rect 29918 30903 29974 30912
rect 30012 30932 30064 30938
rect 30012 30874 30064 30880
rect 30116 30818 30144 37624
rect 30300 33134 30328 38490
rect 30760 37874 30788 38830
rect 30944 38554 30972 39442
rect 31496 38654 31524 40870
rect 31680 39030 31708 40938
rect 31760 39840 31812 39846
rect 31760 39782 31812 39788
rect 31668 39024 31720 39030
rect 31668 38966 31720 38972
rect 31496 38626 31616 38654
rect 30932 38548 30984 38554
rect 30932 38490 30984 38496
rect 31588 38486 31616 38626
rect 31576 38480 31628 38486
rect 31576 38422 31628 38428
rect 30748 37868 30800 37874
rect 30748 37810 30800 37816
rect 31588 37466 31616 38422
rect 31680 37942 31708 38966
rect 31772 38758 31800 39782
rect 31760 38752 31812 38758
rect 31760 38694 31812 38700
rect 31772 38010 31800 38694
rect 31852 38344 31904 38350
rect 31852 38286 31904 38292
rect 32036 38344 32088 38350
rect 32036 38286 32088 38292
rect 31760 38004 31812 38010
rect 31760 37946 31812 37952
rect 31668 37936 31720 37942
rect 31668 37878 31720 37884
rect 31576 37460 31628 37466
rect 31576 37402 31628 37408
rect 31392 37392 31444 37398
rect 31392 37334 31444 37340
rect 30748 37324 30800 37330
rect 30748 37266 30800 37272
rect 30840 37324 30892 37330
rect 30840 37266 30892 37272
rect 30760 36650 30788 37266
rect 30852 36922 30880 37266
rect 30840 36916 30892 36922
rect 30840 36858 30892 36864
rect 31404 36786 31432 37334
rect 31576 37188 31628 37194
rect 31576 37130 31628 37136
rect 31392 36780 31444 36786
rect 31392 36722 31444 36728
rect 30748 36644 30800 36650
rect 30748 36586 30800 36592
rect 30472 36576 30524 36582
rect 30472 36518 30524 36524
rect 30484 36378 30512 36518
rect 30472 36372 30524 36378
rect 30472 36314 30524 36320
rect 30748 36372 30800 36378
rect 30748 36314 30800 36320
rect 30760 35562 30788 36314
rect 31404 36106 31432 36722
rect 31484 36644 31536 36650
rect 31484 36586 31536 36592
rect 31496 36242 31524 36586
rect 31588 36582 31616 37130
rect 31668 36780 31720 36786
rect 31668 36722 31720 36728
rect 31576 36576 31628 36582
rect 31576 36518 31628 36524
rect 31484 36236 31536 36242
rect 31484 36178 31536 36184
rect 31392 36100 31444 36106
rect 31392 36042 31444 36048
rect 31300 35692 31352 35698
rect 31300 35634 31352 35640
rect 30748 35556 30800 35562
rect 30748 35498 30800 35504
rect 30472 35148 30524 35154
rect 30472 35090 30524 35096
rect 30484 34474 30512 35090
rect 30564 35080 30616 35086
rect 30564 35022 30616 35028
rect 31208 35080 31260 35086
rect 31208 35022 31260 35028
rect 30472 34468 30524 34474
rect 30472 34410 30524 34416
rect 30484 34377 30512 34410
rect 30470 34368 30526 34377
rect 30470 34303 30526 34312
rect 30576 34134 30604 35022
rect 30748 34468 30800 34474
rect 30748 34410 30800 34416
rect 30760 34202 30788 34410
rect 30748 34196 30800 34202
rect 30748 34138 30800 34144
rect 30564 34128 30616 34134
rect 30564 34070 30616 34076
rect 30380 33652 30432 33658
rect 30380 33594 30432 33600
rect 30024 30790 30144 30818
rect 30208 33106 30328 33134
rect 29552 30660 29604 30666
rect 29552 30602 29604 30608
rect 29564 30394 29592 30602
rect 29644 30592 29696 30598
rect 29644 30534 29696 30540
rect 29552 30388 29604 30394
rect 29552 30330 29604 30336
rect 29656 30326 29684 30534
rect 29644 30320 29696 30326
rect 29550 30288 29606 30297
rect 29092 30252 29144 30258
rect 29644 30262 29696 30268
rect 29550 30223 29606 30232
rect 29092 30194 29144 30200
rect 29000 28960 29052 28966
rect 29000 28902 29052 28908
rect 28908 28688 28960 28694
rect 28908 28630 28960 28636
rect 29012 27878 29040 28902
rect 29104 28218 29132 30194
rect 29564 30190 29592 30223
rect 30024 30190 30052 30790
rect 30104 30728 30156 30734
rect 30104 30670 30156 30676
rect 30116 30394 30144 30670
rect 30104 30388 30156 30394
rect 30104 30330 30156 30336
rect 29552 30184 29604 30190
rect 29552 30126 29604 30132
rect 30012 30184 30064 30190
rect 30012 30126 30064 30132
rect 30116 29850 30144 30330
rect 30208 30258 30236 33106
rect 30288 31748 30340 31754
rect 30288 31690 30340 31696
rect 30196 30252 30248 30258
rect 30196 30194 30248 30200
rect 30104 29844 30156 29850
rect 30104 29786 30156 29792
rect 30300 29646 30328 31690
rect 30392 31142 30420 33594
rect 30576 33454 30604 34070
rect 31220 34066 31248 35022
rect 31312 34610 31340 35634
rect 31300 34604 31352 34610
rect 31300 34546 31352 34552
rect 31298 34368 31354 34377
rect 31298 34303 31354 34312
rect 31208 34060 31260 34066
rect 31208 34002 31260 34008
rect 30564 33448 30616 33454
rect 30564 33390 30616 33396
rect 31116 33448 31168 33454
rect 31116 33390 31168 33396
rect 30576 33134 30604 33390
rect 30576 33106 30788 33134
rect 30760 32978 30788 33106
rect 31128 32978 31156 33390
rect 30472 32972 30524 32978
rect 30472 32914 30524 32920
rect 30748 32972 30800 32978
rect 30748 32914 30800 32920
rect 31116 32972 31168 32978
rect 31116 32914 31168 32920
rect 30484 32230 30512 32914
rect 30564 32292 30616 32298
rect 30564 32234 30616 32240
rect 30472 32224 30524 32230
rect 30472 32166 30524 32172
rect 30484 31385 30512 32166
rect 30470 31376 30526 31385
rect 30470 31311 30526 31320
rect 30380 31136 30432 31142
rect 30380 31078 30432 31084
rect 30472 30864 30524 30870
rect 30472 30806 30524 30812
rect 30484 30394 30512 30806
rect 30576 30666 30604 32234
rect 30760 32026 30788 32914
rect 31312 32366 31340 34303
rect 31588 33134 31616 36518
rect 31680 35698 31708 36722
rect 31864 36666 31892 38286
rect 31944 38208 31996 38214
rect 32048 38185 32076 38286
rect 31944 38150 31996 38156
rect 32034 38176 32090 38185
rect 31956 37874 31984 38150
rect 32034 38111 32090 38120
rect 31944 37868 31996 37874
rect 31944 37810 31996 37816
rect 31772 36638 31892 36666
rect 31668 35692 31720 35698
rect 31668 35634 31720 35640
rect 31772 34610 31800 36638
rect 31852 36576 31904 36582
rect 31852 36518 31904 36524
rect 31864 36310 31892 36518
rect 31852 36304 31904 36310
rect 31852 36246 31904 36252
rect 31760 34604 31812 34610
rect 31760 34546 31812 34552
rect 31772 33930 31800 34546
rect 31760 33924 31812 33930
rect 31760 33866 31812 33872
rect 31496 33106 31616 33134
rect 31956 33134 31984 37810
rect 32036 37664 32088 37670
rect 32036 37606 32088 37612
rect 32048 36310 32076 37606
rect 32140 37233 32168 41142
rect 32588 40928 32640 40934
rect 32588 40870 32640 40876
rect 32496 40520 32548 40526
rect 32496 40462 32548 40468
rect 32404 40452 32456 40458
rect 32404 40394 32456 40400
rect 32220 40112 32272 40118
rect 32220 40054 32272 40060
rect 32126 37224 32182 37233
rect 32126 37159 32182 37168
rect 32232 36854 32260 40054
rect 32416 39370 32444 40394
rect 32508 39642 32536 40462
rect 32600 40050 32628 40870
rect 32680 40656 32732 40662
rect 32680 40598 32732 40604
rect 32588 40044 32640 40050
rect 32588 39986 32640 39992
rect 32588 39908 32640 39914
rect 32692 39896 32720 40598
rect 32640 39868 32720 39896
rect 32588 39850 32640 39856
rect 32496 39636 32548 39642
rect 32496 39578 32548 39584
rect 32404 39364 32456 39370
rect 32404 39306 32456 39312
rect 32416 39114 32444 39306
rect 32324 39086 32444 39114
rect 32324 37398 32352 39086
rect 32404 39024 32456 39030
rect 32404 38966 32456 38972
rect 32312 37392 32364 37398
rect 32312 37334 32364 37340
rect 32312 37256 32364 37262
rect 32312 37198 32364 37204
rect 32220 36848 32272 36854
rect 32220 36790 32272 36796
rect 32036 36304 32088 36310
rect 32036 36246 32088 36252
rect 32232 36145 32260 36790
rect 32324 36378 32352 37198
rect 32312 36372 32364 36378
rect 32312 36314 32364 36320
rect 32218 36136 32274 36145
rect 32218 36071 32274 36080
rect 32416 35766 32444 38966
rect 32600 38486 32628 39850
rect 32680 39568 32732 39574
rect 32680 39510 32732 39516
rect 32692 38758 32720 39510
rect 32680 38752 32732 38758
rect 32680 38694 32732 38700
rect 32588 38480 32640 38486
rect 32588 38422 32640 38428
rect 32600 38010 32628 38422
rect 32588 38004 32640 38010
rect 32588 37946 32640 37952
rect 32496 37460 32548 37466
rect 32496 37402 32548 37408
rect 32508 36582 32536 37402
rect 32692 37330 32720 38694
rect 32784 37874 32812 41414
rect 34940 41372 35236 41392
rect 34996 41370 35020 41372
rect 35076 41370 35100 41372
rect 35156 41370 35180 41372
rect 35018 41318 35020 41370
rect 35082 41318 35094 41370
rect 35156 41318 35158 41370
rect 34996 41316 35020 41318
rect 35076 41316 35100 41318
rect 35156 41316 35180 41318
rect 34940 41296 35236 41316
rect 35532 41132 35584 41138
rect 35532 41074 35584 41080
rect 32864 41064 32916 41070
rect 32864 41006 32916 41012
rect 32876 39681 32904 41006
rect 33048 40996 33100 41002
rect 33048 40938 33100 40944
rect 32956 40384 33008 40390
rect 32956 40326 33008 40332
rect 32862 39672 32918 39681
rect 32862 39607 32918 39616
rect 32864 39432 32916 39438
rect 32864 39374 32916 39380
rect 32876 39098 32904 39374
rect 32864 39092 32916 39098
rect 32864 39034 32916 39040
rect 32876 38486 32904 39034
rect 32864 38480 32916 38486
rect 32864 38422 32916 38428
rect 32864 38344 32916 38350
rect 32864 38286 32916 38292
rect 32876 38185 32904 38286
rect 32862 38176 32918 38185
rect 32862 38111 32918 38120
rect 32864 38004 32916 38010
rect 32864 37946 32916 37952
rect 32772 37868 32824 37874
rect 32772 37810 32824 37816
rect 32876 37738 32904 37946
rect 32864 37732 32916 37738
rect 32864 37674 32916 37680
rect 32680 37324 32732 37330
rect 32680 37266 32732 37272
rect 32692 36922 32720 37266
rect 32680 36916 32732 36922
rect 32680 36858 32732 36864
rect 32692 36650 32720 36858
rect 32968 36786 32996 40326
rect 33060 40186 33088 40938
rect 33784 40928 33836 40934
rect 33784 40870 33836 40876
rect 33232 40452 33284 40458
rect 33232 40394 33284 40400
rect 33048 40180 33100 40186
rect 33048 40122 33100 40128
rect 33140 39840 33192 39846
rect 33140 39782 33192 39788
rect 33048 39296 33100 39302
rect 33048 39238 33100 39244
rect 33060 38962 33088 39238
rect 33152 39030 33180 39782
rect 33140 39024 33192 39030
rect 33140 38966 33192 38972
rect 33048 38956 33100 38962
rect 33048 38898 33100 38904
rect 33060 38554 33088 38898
rect 33048 38548 33100 38554
rect 33048 38490 33100 38496
rect 33244 38400 33272 40394
rect 33152 38372 33272 38400
rect 32956 36780 33008 36786
rect 32956 36722 33008 36728
rect 32680 36644 32732 36650
rect 32680 36586 32732 36592
rect 32496 36576 32548 36582
rect 32496 36518 32548 36524
rect 33152 36394 33180 38372
rect 33232 37868 33284 37874
rect 33232 37810 33284 37816
rect 33244 37466 33272 37810
rect 33416 37732 33468 37738
rect 33416 37674 33468 37680
rect 33232 37460 33284 37466
rect 33232 37402 33284 37408
rect 33428 36854 33456 37674
rect 33796 37262 33824 40870
rect 33968 40588 34020 40594
rect 33968 40530 34020 40536
rect 35256 40588 35308 40594
rect 35256 40530 35308 40536
rect 33980 40118 34008 40530
rect 34940 40284 35236 40304
rect 34996 40282 35020 40284
rect 35076 40282 35100 40284
rect 35156 40282 35180 40284
rect 35018 40230 35020 40282
rect 35082 40230 35094 40282
rect 35156 40230 35158 40282
rect 34996 40228 35020 40230
rect 35076 40228 35100 40230
rect 35156 40228 35180 40230
rect 34940 40208 35236 40228
rect 35268 40186 35296 40530
rect 35256 40180 35308 40186
rect 35256 40122 35308 40128
rect 33968 40112 34020 40118
rect 33968 40054 34020 40060
rect 35544 39982 35572 41074
rect 35622 40760 35678 40769
rect 35622 40695 35678 40704
rect 35532 39976 35584 39982
rect 35532 39918 35584 39924
rect 34428 39500 34480 39506
rect 34428 39442 34480 39448
rect 34440 39001 34468 39442
rect 34940 39196 35236 39216
rect 34996 39194 35020 39196
rect 35076 39194 35100 39196
rect 35156 39194 35180 39196
rect 35018 39142 35020 39194
rect 35082 39142 35094 39194
rect 35156 39142 35158 39194
rect 34996 39140 35020 39142
rect 35076 39140 35100 39142
rect 35156 39140 35180 39142
rect 34940 39120 35236 39140
rect 35636 39098 35664 40695
rect 35716 39908 35768 39914
rect 35716 39850 35768 39856
rect 35624 39092 35676 39098
rect 35624 39034 35676 39040
rect 34426 38992 34482 39001
rect 34426 38927 34482 38936
rect 34440 38894 34468 38927
rect 35636 38894 35664 39034
rect 34428 38888 34480 38894
rect 34428 38830 34480 38836
rect 35624 38888 35676 38894
rect 35624 38830 35676 38836
rect 33968 38412 34020 38418
rect 33968 38354 34020 38360
rect 33980 38010 34008 38354
rect 34244 38344 34296 38350
rect 34244 38286 34296 38292
rect 35256 38344 35308 38350
rect 35256 38286 35308 38292
rect 33968 38004 34020 38010
rect 33968 37946 34020 37952
rect 34256 37262 34284 38286
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 35268 37466 35296 38286
rect 35728 38214 35756 39850
rect 35912 38758 35940 49558
rect 36082 49520 36138 49558
rect 41524 49558 41658 49586
rect 38198 40760 38254 40769
rect 38198 40695 38254 40704
rect 37464 40384 37516 40390
rect 37464 40326 37516 40332
rect 37476 39982 37504 40326
rect 37464 39976 37516 39982
rect 37464 39918 37516 39924
rect 36084 39840 36136 39846
rect 36084 39782 36136 39788
rect 36096 39642 36124 39782
rect 36084 39636 36136 39642
rect 36084 39578 36136 39584
rect 36452 39568 36504 39574
rect 36452 39510 36504 39516
rect 36464 38826 36492 39510
rect 36820 39432 36872 39438
rect 36820 39374 36872 39380
rect 36832 39030 36860 39374
rect 36820 39024 36872 39030
rect 36820 38966 36872 38972
rect 36452 38820 36504 38826
rect 36452 38762 36504 38768
rect 37004 38820 37056 38826
rect 37004 38762 37056 38768
rect 35900 38752 35952 38758
rect 35900 38694 35952 38700
rect 35808 38480 35860 38486
rect 35808 38422 35860 38428
rect 35716 38208 35768 38214
rect 35716 38150 35768 38156
rect 35820 37942 35848 38422
rect 35912 38418 35940 38694
rect 35900 38412 35952 38418
rect 35900 38354 35952 38360
rect 36464 38214 36492 38762
rect 36452 38208 36504 38214
rect 36452 38150 36504 38156
rect 36544 38208 36596 38214
rect 36544 38150 36596 38156
rect 35808 37936 35860 37942
rect 35808 37878 35860 37884
rect 35990 37904 36046 37913
rect 35990 37839 36046 37848
rect 36004 37806 36032 37839
rect 35992 37800 36044 37806
rect 36044 37760 36124 37788
rect 35992 37742 36044 37748
rect 35256 37460 35308 37466
rect 35256 37402 35308 37408
rect 35716 37324 35768 37330
rect 35716 37266 35768 37272
rect 35900 37324 35952 37330
rect 35900 37266 35952 37272
rect 33784 37256 33836 37262
rect 33784 37198 33836 37204
rect 34244 37256 34296 37262
rect 34244 37198 34296 37204
rect 33692 37120 33744 37126
rect 33692 37062 33744 37068
rect 33416 36848 33468 36854
rect 33416 36790 33468 36796
rect 33232 36576 33284 36582
rect 33232 36518 33284 36524
rect 33060 36366 33180 36394
rect 32864 36304 32916 36310
rect 32864 36246 32916 36252
rect 32496 35828 32548 35834
rect 32496 35770 32548 35776
rect 32404 35760 32456 35766
rect 32404 35702 32456 35708
rect 32404 35012 32456 35018
rect 32404 34954 32456 34960
rect 32416 34610 32444 34954
rect 32404 34604 32456 34610
rect 32404 34546 32456 34552
rect 32128 34400 32180 34406
rect 32128 34342 32180 34348
rect 32140 33658 32168 34342
rect 32312 34128 32364 34134
rect 32312 34070 32364 34076
rect 32128 33652 32180 33658
rect 32128 33594 32180 33600
rect 32324 33386 32352 34070
rect 32312 33380 32364 33386
rect 32312 33322 32364 33328
rect 32508 33134 32536 35770
rect 32876 35290 32904 36246
rect 33060 35698 33088 36366
rect 33140 36304 33192 36310
rect 33140 36246 33192 36252
rect 33048 35692 33100 35698
rect 33048 35634 33100 35640
rect 33152 35562 33180 36246
rect 33140 35556 33192 35562
rect 33140 35498 33192 35504
rect 32864 35284 32916 35290
rect 32864 35226 32916 35232
rect 33152 35222 33180 35498
rect 33140 35216 33192 35222
rect 33140 35158 33192 35164
rect 33048 35080 33100 35086
rect 33048 35022 33100 35028
rect 33060 34746 33088 35022
rect 32588 34740 32640 34746
rect 32588 34682 32640 34688
rect 33048 34740 33100 34746
rect 33048 34682 33100 34688
rect 32600 34474 32628 34682
rect 32588 34468 32640 34474
rect 32588 34410 32640 34416
rect 33060 34202 33088 34682
rect 33152 34406 33180 35158
rect 33140 34400 33192 34406
rect 33140 34342 33192 34348
rect 33048 34196 33100 34202
rect 33048 34138 33100 34144
rect 33152 34082 33180 34342
rect 33060 34054 33180 34082
rect 33060 33862 33088 34054
rect 33048 33856 33100 33862
rect 33048 33798 33100 33804
rect 33060 33658 33088 33798
rect 33048 33652 33100 33658
rect 33048 33594 33100 33600
rect 33244 33504 33272 36518
rect 33428 35086 33456 36790
rect 33704 36786 33732 37062
rect 33796 36922 33824 37198
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 33784 36916 33836 36922
rect 33784 36858 33836 36864
rect 33692 36780 33744 36786
rect 33692 36722 33744 36728
rect 35728 36718 35756 37266
rect 35912 36786 35940 37266
rect 35900 36780 35952 36786
rect 35900 36722 35952 36728
rect 34704 36712 34756 36718
rect 34704 36654 34756 36660
rect 35440 36712 35492 36718
rect 35440 36654 35492 36660
rect 35716 36712 35768 36718
rect 35716 36654 35768 36660
rect 34336 36236 34388 36242
rect 34336 36178 34388 36184
rect 34348 35834 34376 36178
rect 34336 35828 34388 35834
rect 34336 35770 34388 35776
rect 34716 35601 34744 36654
rect 35452 36038 35480 36654
rect 35624 36644 35676 36650
rect 35624 36586 35676 36592
rect 35636 36378 35664 36586
rect 35624 36372 35676 36378
rect 35624 36314 35676 36320
rect 34796 36032 34848 36038
rect 34796 35974 34848 35980
rect 35440 36032 35492 36038
rect 35440 35974 35492 35980
rect 34242 35592 34298 35601
rect 34242 35527 34298 35536
rect 34702 35592 34758 35601
rect 34702 35527 34758 35536
rect 33416 35080 33468 35086
rect 33416 35022 33468 35028
rect 33876 34060 33928 34066
rect 33876 34002 33928 34008
rect 33324 33924 33376 33930
rect 33324 33866 33376 33872
rect 33336 33522 33364 33866
rect 33888 33658 33916 34002
rect 33876 33652 33928 33658
rect 33876 33594 33928 33600
rect 33106 33476 33272 33504
rect 33106 33436 33134 33476
rect 32876 33408 33134 33436
rect 32772 33380 32824 33386
rect 32876 33368 32904 33408
rect 32824 33340 32904 33368
rect 32772 33322 32824 33328
rect 31956 33106 32168 33134
rect 31300 32360 31352 32366
rect 31300 32302 31352 32308
rect 30748 32020 30800 32026
rect 30748 31962 30800 31968
rect 30930 31376 30986 31385
rect 30930 31311 30986 31320
rect 30944 31278 30972 31311
rect 30932 31272 30984 31278
rect 30932 31214 30984 31220
rect 30840 30728 30892 30734
rect 30840 30670 30892 30676
rect 30564 30660 30616 30666
rect 30564 30602 30616 30608
rect 30472 30388 30524 30394
rect 30472 30330 30524 30336
rect 30380 29776 30432 29782
rect 30380 29718 30432 29724
rect 29184 29640 29236 29646
rect 29184 29582 29236 29588
rect 30288 29640 30340 29646
rect 30288 29582 30340 29588
rect 29196 28762 29224 29582
rect 29276 29504 29328 29510
rect 29276 29446 29328 29452
rect 29288 29102 29316 29446
rect 29276 29096 29328 29102
rect 29276 29038 29328 29044
rect 30196 28960 30248 28966
rect 30196 28902 30248 28908
rect 29184 28756 29236 28762
rect 29184 28698 29236 28704
rect 30104 28756 30156 28762
rect 30104 28698 30156 28704
rect 29092 28212 29144 28218
rect 29092 28154 29144 28160
rect 29196 28082 29224 28698
rect 29368 28620 29420 28626
rect 29368 28562 29420 28568
rect 29184 28076 29236 28082
rect 29184 28018 29236 28024
rect 29000 27872 29052 27878
rect 29000 27814 29052 27820
rect 28908 26512 28960 26518
rect 28908 26454 28960 26460
rect 28816 25832 28868 25838
rect 28816 25774 28868 25780
rect 28920 25702 28948 26454
rect 29012 25906 29040 27814
rect 29380 27538 29408 28562
rect 29736 28552 29788 28558
rect 29736 28494 29788 28500
rect 29748 27946 29776 28494
rect 29736 27940 29788 27946
rect 29736 27882 29788 27888
rect 29748 27538 29776 27882
rect 30116 27878 30144 28698
rect 30208 28218 30236 28902
rect 30300 28626 30328 29582
rect 30392 28966 30420 29718
rect 30576 29170 30604 30602
rect 30852 30258 30880 30670
rect 30932 30592 30984 30598
rect 30932 30534 30984 30540
rect 30840 30252 30892 30258
rect 30840 30194 30892 30200
rect 30944 30122 30972 30534
rect 31300 30252 31352 30258
rect 31300 30194 31352 30200
rect 30932 30116 30984 30122
rect 30932 30058 30984 30064
rect 30564 29164 30616 29170
rect 30564 29106 30616 29112
rect 30380 28960 30432 28966
rect 30380 28902 30432 28908
rect 30944 28762 30972 30058
rect 31312 29578 31340 30194
rect 31392 30048 31444 30054
rect 31392 29990 31444 29996
rect 31404 29646 31432 29990
rect 31496 29714 31524 33106
rect 32140 32978 32168 33106
rect 32220 33108 32272 33114
rect 32220 33050 32272 33056
rect 32416 33106 32536 33134
rect 33244 33114 33272 33476
rect 33324 33516 33376 33522
rect 33324 33458 33376 33464
rect 33232 33108 33284 33114
rect 32128 32972 32180 32978
rect 32128 32914 32180 32920
rect 31576 32768 31628 32774
rect 31576 32710 31628 32716
rect 31588 32434 31616 32710
rect 31576 32428 31628 32434
rect 31576 32370 31628 32376
rect 31588 31482 31616 32370
rect 31944 32360 31996 32366
rect 31944 32302 31996 32308
rect 31956 32026 31984 32302
rect 32128 32292 32180 32298
rect 32128 32234 32180 32240
rect 31944 32020 31996 32026
rect 31944 31962 31996 31968
rect 31576 31476 31628 31482
rect 31576 31418 31628 31424
rect 31956 29782 31984 31962
rect 32140 31822 32168 32234
rect 32128 31816 32180 31822
rect 32128 31758 32180 31764
rect 32232 31346 32260 33050
rect 32312 32904 32364 32910
rect 32312 32846 32364 32852
rect 32324 32230 32352 32846
rect 32416 32842 32444 33106
rect 33232 33050 33284 33056
rect 32496 32972 32548 32978
rect 32680 32972 32732 32978
rect 32548 32932 32628 32960
rect 32496 32914 32548 32920
rect 32404 32836 32456 32842
rect 32404 32778 32456 32784
rect 32312 32224 32364 32230
rect 32312 32166 32364 32172
rect 32220 31340 32272 31346
rect 32220 31282 32272 31288
rect 32232 30938 32260 31282
rect 32220 30932 32272 30938
rect 32220 30874 32272 30880
rect 31944 29776 31996 29782
rect 31944 29718 31996 29724
rect 31484 29708 31536 29714
rect 31484 29650 31536 29656
rect 32128 29708 32180 29714
rect 32128 29650 32180 29656
rect 31392 29640 31444 29646
rect 31392 29582 31444 29588
rect 31300 29572 31352 29578
rect 31300 29514 31352 29520
rect 31404 29170 31432 29582
rect 31300 29164 31352 29170
rect 31300 29106 31352 29112
rect 31392 29164 31444 29170
rect 31392 29106 31444 29112
rect 31944 29164 31996 29170
rect 31944 29106 31996 29112
rect 31312 28762 31340 29106
rect 31956 28762 31984 29106
rect 32140 28966 32168 29650
rect 32128 28960 32180 28966
rect 32128 28902 32180 28908
rect 30932 28756 30984 28762
rect 30932 28698 30984 28704
rect 31300 28756 31352 28762
rect 31300 28698 31352 28704
rect 31944 28756 31996 28762
rect 31944 28698 31996 28704
rect 30288 28620 30340 28626
rect 30288 28562 30340 28568
rect 30196 28212 30248 28218
rect 30196 28154 30248 28160
rect 30104 27872 30156 27878
rect 30104 27814 30156 27820
rect 31668 27872 31720 27878
rect 31668 27814 31720 27820
rect 30380 27600 30432 27606
rect 30380 27542 30432 27548
rect 29368 27532 29420 27538
rect 29368 27474 29420 27480
rect 29736 27532 29788 27538
rect 29736 27474 29788 27480
rect 29380 27130 29408 27474
rect 30392 27441 30420 27542
rect 31208 27464 31260 27470
rect 30378 27432 30434 27441
rect 31208 27406 31260 27412
rect 30378 27367 30434 27376
rect 30196 27328 30248 27334
rect 30196 27270 30248 27276
rect 29368 27124 29420 27130
rect 29368 27066 29420 27072
rect 30208 26926 30236 27270
rect 29092 26920 29144 26926
rect 29092 26862 29144 26868
rect 30196 26920 30248 26926
rect 30196 26862 30248 26868
rect 29104 26450 29132 26862
rect 30208 26586 30236 26862
rect 30840 26852 30892 26858
rect 30840 26794 30892 26800
rect 30852 26586 30880 26794
rect 31220 26790 31248 27406
rect 31680 26926 31708 27814
rect 32140 27062 32168 28902
rect 32220 28416 32272 28422
rect 32220 28358 32272 28364
rect 32232 28014 32260 28358
rect 32220 28008 32272 28014
rect 32220 27950 32272 27956
rect 32232 27674 32260 27950
rect 32220 27668 32272 27674
rect 32220 27610 32272 27616
rect 32324 27538 32352 32166
rect 32312 27532 32364 27538
rect 32312 27474 32364 27480
rect 32416 27112 32444 32778
rect 32600 32230 32628 32932
rect 32680 32914 32732 32920
rect 32692 32570 32720 32914
rect 32680 32564 32732 32570
rect 32680 32506 32732 32512
rect 34060 32564 34112 32570
rect 34060 32506 34112 32512
rect 32692 32366 32720 32506
rect 32772 32428 32824 32434
rect 32772 32370 32824 32376
rect 32680 32360 32732 32366
rect 32680 32302 32732 32308
rect 32588 32224 32640 32230
rect 32588 32166 32640 32172
rect 32496 32020 32548 32026
rect 32496 31962 32548 31968
rect 32508 31210 32536 31962
rect 32496 31204 32548 31210
rect 32496 31146 32548 31152
rect 32600 30716 32628 32166
rect 32680 31816 32732 31822
rect 32680 31758 32732 31764
rect 32692 30938 32720 31758
rect 32680 30932 32732 30938
rect 32680 30874 32732 30880
rect 32600 30688 32720 30716
rect 32496 29776 32548 29782
rect 32496 29718 32548 29724
rect 32508 28694 32536 29718
rect 32588 29708 32640 29714
rect 32588 29650 32640 29656
rect 32600 29306 32628 29650
rect 32588 29300 32640 29306
rect 32588 29242 32640 29248
rect 32496 28688 32548 28694
rect 32496 28630 32548 28636
rect 32508 28218 32536 28630
rect 32496 28212 32548 28218
rect 32496 28154 32548 28160
rect 32600 27538 32628 29242
rect 32588 27532 32640 27538
rect 32588 27474 32640 27480
rect 32600 27130 32628 27474
rect 32588 27124 32640 27130
rect 32416 27084 32536 27112
rect 32128 27056 32180 27062
rect 32128 26998 32180 27004
rect 32404 26988 32456 26994
rect 32404 26930 32456 26936
rect 31668 26920 31720 26926
rect 32416 26897 32444 26930
rect 31668 26862 31720 26868
rect 32402 26888 32458 26897
rect 32402 26823 32458 26832
rect 31208 26784 31260 26790
rect 31208 26726 31260 26732
rect 32220 26784 32272 26790
rect 32220 26726 32272 26732
rect 30196 26580 30248 26586
rect 30196 26522 30248 26528
rect 30840 26580 30892 26586
rect 30840 26522 30892 26528
rect 29092 26444 29144 26450
rect 29092 26386 29144 26392
rect 29276 26376 29328 26382
rect 29276 26318 29328 26324
rect 30012 26376 30064 26382
rect 30012 26318 30064 26324
rect 29288 26042 29316 26318
rect 29276 26036 29328 26042
rect 29276 25978 29328 25984
rect 29000 25900 29052 25906
rect 29000 25842 29052 25848
rect 28908 25696 28960 25702
rect 28908 25638 28960 25644
rect 28920 25158 28948 25638
rect 29920 25424 29972 25430
rect 29920 25366 29972 25372
rect 29368 25220 29420 25226
rect 29368 25162 29420 25168
rect 28908 25152 28960 25158
rect 28908 25094 28960 25100
rect 28920 24682 28948 25094
rect 29380 24818 29408 25162
rect 29368 24812 29420 24818
rect 29368 24754 29420 24760
rect 29828 24812 29880 24818
rect 29828 24754 29880 24760
rect 29366 24712 29422 24721
rect 28908 24676 28960 24682
rect 29366 24647 29422 24656
rect 28908 24618 28960 24624
rect 28816 24404 28868 24410
rect 28816 24346 28868 24352
rect 28724 24268 28776 24274
rect 28724 24210 28776 24216
rect 28736 23866 28764 24210
rect 28724 23860 28776 23866
rect 28724 23802 28776 23808
rect 28828 23118 28856 24346
rect 29000 23588 29052 23594
rect 29000 23530 29052 23536
rect 28816 23112 28868 23118
rect 28644 23038 28764 23066
rect 28816 23054 28868 23060
rect 28632 22976 28684 22982
rect 28632 22918 28684 22924
rect 28264 22772 28316 22778
rect 28264 22714 28316 22720
rect 28276 22438 28304 22714
rect 28644 22506 28672 22918
rect 28736 22710 28764 23038
rect 28828 22778 28856 23054
rect 28816 22772 28868 22778
rect 28816 22714 28868 22720
rect 28724 22704 28776 22710
rect 28724 22646 28776 22652
rect 28632 22500 28684 22506
rect 28632 22442 28684 22448
rect 28264 22432 28316 22438
rect 28264 22374 28316 22380
rect 28276 22166 28304 22374
rect 29012 22234 29040 23530
rect 29380 23474 29408 24647
rect 29460 24268 29512 24274
rect 29460 24210 29512 24216
rect 29472 23866 29500 24210
rect 29736 24064 29788 24070
rect 29736 24006 29788 24012
rect 29460 23860 29512 23866
rect 29460 23802 29512 23808
rect 29748 23526 29776 24006
rect 29840 23730 29868 24754
rect 29932 24614 29960 25366
rect 29920 24608 29972 24614
rect 29920 24550 29972 24556
rect 29828 23724 29880 23730
rect 29828 23666 29880 23672
rect 29736 23520 29788 23526
rect 29380 23446 29500 23474
rect 29736 23462 29788 23468
rect 29000 22228 29052 22234
rect 29000 22170 29052 22176
rect 28264 22160 28316 22166
rect 28264 22102 28316 22108
rect 28080 22024 28132 22030
rect 28080 21966 28132 21972
rect 28276 21690 28304 22102
rect 28816 22024 28868 22030
rect 28816 21966 28868 21972
rect 28264 21684 28316 21690
rect 28264 21626 28316 21632
rect 27896 21616 27948 21622
rect 27816 21576 27896 21604
rect 27896 21558 27948 21564
rect 27712 21548 27764 21554
rect 27712 21490 27764 21496
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 27528 21344 27580 21350
rect 27528 21286 27580 21292
rect 27436 20868 27488 20874
rect 27436 20810 27488 20816
rect 27436 20528 27488 20534
rect 27540 20516 27568 21286
rect 27632 21010 27660 21422
rect 27620 21004 27672 21010
rect 27620 20946 27672 20952
rect 27488 20488 27568 20516
rect 27436 20470 27488 20476
rect 27448 20262 27476 20470
rect 27436 20256 27488 20262
rect 27436 20198 27488 20204
rect 27344 19916 27396 19922
rect 27344 19858 27396 19864
rect 26700 19848 26752 19854
rect 26700 19790 26752 19796
rect 26884 19848 26936 19854
rect 26884 19790 26936 19796
rect 26240 19508 26292 19514
rect 26240 19450 26292 19456
rect 26712 18630 26740 19790
rect 26884 19712 26936 19718
rect 26884 19654 26936 19660
rect 26896 19174 26924 19654
rect 26884 19168 26936 19174
rect 26884 19110 26936 19116
rect 27068 18828 27120 18834
rect 27068 18770 27120 18776
rect 26700 18624 26752 18630
rect 26700 18566 26752 18572
rect 25872 18284 25924 18290
rect 25872 18226 25924 18232
rect 25884 17202 25912 18226
rect 25872 17196 25924 17202
rect 25872 17138 25924 17144
rect 26424 16652 26476 16658
rect 26424 16594 26476 16600
rect 25872 15972 25924 15978
rect 25872 15914 25924 15920
rect 26332 15972 26384 15978
rect 26332 15914 26384 15920
rect 25884 15366 25912 15914
rect 25872 15360 25924 15366
rect 25872 15302 25924 15308
rect 26344 14532 26372 15914
rect 26436 15910 26464 16594
rect 26424 15904 26476 15910
rect 26424 15846 26476 15852
rect 26436 15570 26464 15846
rect 26424 15564 26476 15570
rect 26424 15506 26476 15512
rect 26608 15496 26660 15502
rect 26608 15438 26660 15444
rect 26620 15162 26648 15438
rect 26712 15434 26740 18566
rect 27080 18426 27108 18770
rect 27068 18420 27120 18426
rect 27068 18362 27120 18368
rect 26792 18148 26844 18154
rect 26792 18090 26844 18096
rect 26804 16998 26832 18090
rect 27080 17882 27108 18362
rect 27068 17876 27120 17882
rect 27068 17818 27120 17824
rect 27356 17746 27384 19858
rect 27448 19718 27476 20198
rect 27632 20058 27660 20946
rect 27724 20806 27752 21490
rect 28828 21146 28856 21966
rect 28816 21140 28868 21146
rect 28816 21082 28868 21088
rect 28264 21004 28316 21010
rect 28264 20946 28316 20952
rect 29092 21004 29144 21010
rect 29092 20946 29144 20952
rect 27712 20800 27764 20806
rect 27712 20742 27764 20748
rect 28080 20800 28132 20806
rect 28080 20742 28132 20748
rect 27724 20330 27752 20742
rect 28092 20534 28120 20742
rect 28276 20602 28304 20946
rect 28632 20936 28684 20942
rect 28632 20878 28684 20884
rect 28644 20602 28672 20878
rect 29104 20602 29132 20946
rect 28264 20596 28316 20602
rect 28264 20538 28316 20544
rect 28632 20596 28684 20602
rect 28632 20538 28684 20544
rect 29092 20596 29144 20602
rect 29092 20538 29144 20544
rect 28080 20528 28132 20534
rect 28080 20470 28132 20476
rect 27712 20324 27764 20330
rect 27712 20266 27764 20272
rect 27620 20052 27672 20058
rect 27620 19994 27672 20000
rect 27436 19712 27488 19718
rect 27436 19654 27488 19660
rect 27896 19712 27948 19718
rect 27896 19654 27948 19660
rect 27908 19310 27936 19654
rect 28276 19514 28304 20538
rect 29472 19922 29500 23446
rect 30024 22642 30052 26318
rect 30852 25906 30880 26522
rect 30932 26444 30984 26450
rect 30932 26386 30984 26392
rect 30944 25974 30972 26386
rect 31220 25974 31248 26726
rect 31852 26376 31904 26382
rect 31852 26318 31904 26324
rect 30932 25968 30984 25974
rect 30932 25910 30984 25916
rect 31208 25968 31260 25974
rect 31208 25910 31260 25916
rect 30656 25900 30708 25906
rect 30656 25842 30708 25848
rect 30840 25900 30892 25906
rect 30840 25842 30892 25848
rect 30668 25770 30696 25842
rect 30656 25764 30708 25770
rect 30656 25706 30708 25712
rect 30104 25288 30156 25294
rect 30104 25230 30156 25236
rect 30116 24410 30144 25230
rect 30380 25220 30432 25226
rect 30380 25162 30432 25168
rect 30104 24404 30156 24410
rect 30104 24346 30156 24352
rect 30392 24206 30420 25162
rect 30944 25158 30972 25910
rect 30932 25152 30984 25158
rect 30932 25094 30984 25100
rect 30472 24336 30524 24342
rect 30472 24278 30524 24284
rect 30380 24200 30432 24206
rect 30380 24142 30432 24148
rect 30104 23724 30156 23730
rect 30104 23666 30156 23672
rect 30116 23322 30144 23666
rect 30104 23316 30156 23322
rect 30104 23258 30156 23264
rect 30392 23186 30420 24142
rect 30484 23866 30512 24278
rect 31024 24200 31076 24206
rect 31024 24142 31076 24148
rect 30472 23860 30524 23866
rect 30472 23802 30524 23808
rect 30484 23322 30512 23802
rect 31036 23798 31064 24142
rect 31024 23792 31076 23798
rect 31024 23734 31076 23740
rect 31036 23474 31064 23734
rect 30944 23446 31064 23474
rect 30472 23316 30524 23322
rect 30472 23258 30524 23264
rect 30380 23180 30432 23186
rect 30380 23122 30432 23128
rect 30104 22704 30156 22710
rect 30104 22646 30156 22652
rect 30012 22636 30064 22642
rect 30012 22578 30064 22584
rect 29828 22500 29880 22506
rect 29828 22442 29880 22448
rect 29644 22432 29696 22438
rect 29644 22374 29696 22380
rect 29552 21956 29604 21962
rect 29552 21898 29604 21904
rect 29564 21486 29592 21898
rect 29552 21480 29604 21486
rect 29552 21422 29604 21428
rect 28632 19916 28684 19922
rect 28632 19858 28684 19864
rect 29460 19916 29512 19922
rect 29460 19858 29512 19864
rect 28644 19514 28672 19858
rect 29472 19718 29500 19858
rect 29460 19712 29512 19718
rect 29460 19654 29512 19660
rect 29472 19514 29500 19654
rect 28264 19508 28316 19514
rect 28264 19450 28316 19456
rect 28632 19508 28684 19514
rect 28632 19450 28684 19456
rect 29460 19508 29512 19514
rect 29460 19450 29512 19456
rect 27896 19304 27948 19310
rect 27896 19246 27948 19252
rect 27436 19168 27488 19174
rect 27436 19110 27488 19116
rect 27448 18086 27476 19110
rect 29182 19000 29238 19009
rect 29182 18935 29238 18944
rect 29196 18834 29224 18935
rect 29184 18828 29236 18834
rect 29184 18770 29236 18776
rect 28540 18760 28592 18766
rect 28540 18702 28592 18708
rect 27712 18148 27764 18154
rect 27712 18090 27764 18096
rect 27436 18080 27488 18086
rect 27436 18022 27488 18028
rect 27344 17740 27396 17746
rect 27344 17682 27396 17688
rect 27356 17202 27384 17682
rect 27344 17196 27396 17202
rect 27344 17138 27396 17144
rect 26792 16992 26844 16998
rect 26792 16934 26844 16940
rect 27160 16992 27212 16998
rect 27160 16934 27212 16940
rect 26804 15638 26832 16934
rect 27172 15910 27200 16934
rect 27448 16250 27476 18022
rect 27724 17542 27752 18090
rect 28552 17814 28580 18702
rect 29196 18426 29224 18770
rect 29184 18420 29236 18426
rect 29184 18362 29236 18368
rect 28724 18284 28776 18290
rect 28724 18226 28776 18232
rect 28736 17814 28764 18226
rect 28816 18216 28868 18222
rect 28816 18158 28868 18164
rect 28540 17808 28592 17814
rect 28724 17808 28776 17814
rect 28592 17768 28672 17796
rect 28540 17750 28592 17756
rect 27712 17536 27764 17542
rect 27712 17478 27764 17484
rect 27620 17128 27672 17134
rect 27620 17070 27672 17076
rect 27528 16448 27580 16454
rect 27632 16436 27660 17070
rect 28644 16998 28672 17768
rect 28724 17750 28776 17756
rect 27804 16992 27856 16998
rect 27804 16934 27856 16940
rect 28632 16992 28684 16998
rect 28632 16934 28684 16940
rect 27816 16658 27844 16934
rect 28540 16720 28592 16726
rect 28540 16662 28592 16668
rect 27804 16652 27856 16658
rect 27804 16594 27856 16600
rect 27580 16408 27660 16436
rect 27528 16390 27580 16396
rect 27436 16244 27488 16250
rect 27436 16186 27488 16192
rect 27160 15904 27212 15910
rect 27160 15846 27212 15852
rect 26792 15632 26844 15638
rect 26792 15574 26844 15580
rect 26700 15428 26752 15434
rect 26700 15370 26752 15376
rect 26608 15156 26660 15162
rect 26608 15098 26660 15104
rect 26804 15094 26832 15574
rect 26884 15496 26936 15502
rect 26884 15438 26936 15444
rect 26792 15088 26844 15094
rect 26792 15030 26844 15036
rect 26424 14544 26476 14550
rect 26344 14504 26424 14532
rect 26424 14486 26476 14492
rect 26436 14006 26464 14486
rect 26608 14408 26660 14414
rect 26608 14350 26660 14356
rect 26620 14074 26648 14350
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26424 14000 26476 14006
rect 26424 13942 26476 13948
rect 26436 13870 26464 13942
rect 26700 13932 26752 13938
rect 26700 13874 26752 13880
rect 25700 13786 25820 13814
rect 26424 13864 26476 13870
rect 26424 13806 26476 13812
rect 26712 13802 26740 13874
rect 26700 13796 26752 13802
rect 25596 13184 25648 13190
rect 25596 13126 25648 13132
rect 25608 12986 25636 13126
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 25320 11212 25372 11218
rect 25320 11154 25372 11160
rect 25226 10976 25282 10985
rect 25226 10911 25282 10920
rect 25240 9994 25268 10911
rect 25228 9988 25280 9994
rect 25228 9930 25280 9936
rect 25700 9738 25728 13786
rect 26700 13738 26752 13744
rect 26332 13728 26384 13734
rect 26332 13670 26384 13676
rect 26344 13530 26372 13670
rect 26332 13524 26384 13530
rect 26332 13466 26384 13472
rect 26516 13320 26568 13326
rect 26516 13262 26568 13268
rect 26528 12102 26556 13262
rect 26792 12300 26844 12306
rect 26792 12242 26844 12248
rect 26516 12096 26568 12102
rect 26516 12038 26568 12044
rect 26528 11762 26556 12038
rect 26516 11756 26568 11762
rect 26516 11698 26568 11704
rect 25872 11688 25924 11694
rect 25792 11648 25872 11676
rect 25792 11257 25820 11648
rect 25872 11630 25924 11636
rect 26804 11626 26832 12242
rect 26896 11665 26924 15438
rect 26976 13456 27028 13462
rect 26976 13398 27028 13404
rect 26988 12918 27016 13398
rect 26976 12912 27028 12918
rect 26976 12854 27028 12860
rect 27172 12782 27200 15846
rect 27344 15360 27396 15366
rect 27344 15302 27396 15308
rect 27356 15162 27384 15302
rect 27252 15156 27304 15162
rect 27252 15098 27304 15104
rect 27344 15156 27396 15162
rect 27344 15098 27396 15104
rect 27264 14550 27292 15098
rect 27448 14600 27476 16186
rect 27540 16017 27568 16390
rect 27526 16008 27582 16017
rect 27526 15943 27582 15952
rect 27816 15706 27844 16594
rect 28080 16040 28132 16046
rect 28080 15982 28132 15988
rect 28170 16008 28226 16017
rect 27804 15700 27856 15706
rect 27804 15642 27856 15648
rect 28092 15502 28120 15982
rect 28170 15943 28226 15952
rect 28264 15972 28316 15978
rect 28080 15496 28132 15502
rect 28080 15438 28132 15444
rect 27528 14612 27580 14618
rect 27448 14572 27528 14600
rect 27528 14554 27580 14560
rect 27252 14544 27304 14550
rect 27252 14486 27304 14492
rect 27264 13938 27292 14486
rect 27252 13932 27304 13938
rect 27252 13874 27304 13880
rect 27540 13802 27568 14554
rect 27528 13796 27580 13802
rect 27528 13738 27580 13744
rect 27804 13184 27856 13190
rect 27804 13126 27856 13132
rect 27816 12782 27844 13126
rect 27160 12776 27212 12782
rect 27160 12718 27212 12724
rect 27804 12776 27856 12782
rect 27804 12718 27856 12724
rect 27436 12640 27488 12646
rect 27436 12582 27488 12588
rect 27448 12306 27476 12582
rect 27436 12300 27488 12306
rect 27436 12242 27488 12248
rect 27712 12300 27764 12306
rect 27712 12242 27764 12248
rect 27724 11801 27752 12242
rect 27710 11792 27766 11801
rect 27710 11727 27766 11736
rect 26882 11656 26938 11665
rect 26792 11620 26844 11626
rect 26938 11614 27016 11642
rect 26882 11591 26938 11600
rect 26792 11562 26844 11568
rect 26608 11348 26660 11354
rect 26608 11290 26660 11296
rect 25778 11248 25834 11257
rect 25778 11183 25834 11192
rect 26056 11212 26108 11218
rect 25792 11150 25820 11183
rect 26056 11154 26108 11160
rect 25780 11144 25832 11150
rect 25780 11086 25832 11092
rect 26068 10470 26096 11154
rect 26620 10674 26648 11290
rect 26700 11212 26752 11218
rect 26700 11154 26752 11160
rect 26608 10668 26660 10674
rect 26608 10610 26660 10616
rect 26056 10464 26108 10470
rect 26056 10406 26108 10412
rect 25700 9710 25820 9738
rect 25136 8288 25188 8294
rect 25136 8230 25188 8236
rect 25688 8288 25740 8294
rect 25688 8230 25740 8236
rect 25148 8022 25176 8230
rect 25136 8016 25188 8022
rect 25136 7958 25188 7964
rect 25044 7812 25096 7818
rect 25044 7754 25096 7760
rect 25056 6254 25084 7754
rect 25700 7750 25728 8230
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25700 7002 25728 7686
rect 25688 6996 25740 7002
rect 25688 6938 25740 6944
rect 25504 6860 25556 6866
rect 25504 6802 25556 6808
rect 25516 6458 25544 6802
rect 25504 6452 25556 6458
rect 25504 6394 25556 6400
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 25044 6248 25096 6254
rect 25044 6190 25096 6196
rect 24780 5846 24808 6190
rect 24768 5840 24820 5846
rect 24768 5782 24820 5788
rect 25044 5840 25096 5846
rect 25044 5782 25096 5788
rect 24780 5574 24808 5782
rect 24768 5568 24820 5574
rect 24768 5510 24820 5516
rect 24584 5160 24636 5166
rect 24584 5102 24636 5108
rect 24492 5092 24544 5098
rect 24492 5034 24544 5040
rect 24504 4758 24532 5034
rect 24596 4826 24624 5102
rect 24584 4820 24636 4826
rect 24584 4762 24636 4768
rect 25056 4758 25084 5782
rect 25792 5681 25820 9710
rect 25962 9616 26018 9625
rect 25962 9551 26018 9560
rect 25976 9518 26004 9551
rect 25964 9512 26016 9518
rect 25964 9454 26016 9460
rect 25872 9376 25924 9382
rect 25872 9318 25924 9324
rect 25884 8634 25912 9318
rect 25872 8628 25924 8634
rect 25872 8570 25924 8576
rect 25884 8362 25912 8570
rect 25872 8356 25924 8362
rect 25872 8298 25924 8304
rect 25976 6458 26004 9454
rect 26068 8090 26096 10406
rect 26620 10266 26648 10610
rect 26608 10260 26660 10266
rect 26608 10202 26660 10208
rect 26712 10010 26740 11154
rect 26620 9982 26740 10010
rect 26620 9926 26648 9982
rect 26608 9920 26660 9926
rect 26608 9862 26660 9868
rect 26620 9518 26648 9862
rect 26608 9512 26660 9518
rect 26608 9454 26660 9460
rect 26620 8838 26648 9454
rect 26884 9444 26936 9450
rect 26884 9386 26936 9392
rect 26896 9042 26924 9386
rect 26988 9042 27016 11614
rect 27528 11620 27580 11626
rect 27528 11562 27580 11568
rect 27540 11529 27568 11562
rect 27526 11520 27582 11529
rect 27526 11455 27582 11464
rect 27252 11076 27304 11082
rect 27252 11018 27304 11024
rect 27264 10198 27292 11018
rect 27252 10192 27304 10198
rect 27252 10134 27304 10140
rect 27344 10192 27396 10198
rect 27344 10134 27396 10140
rect 27264 9178 27292 10134
rect 27356 9722 27384 10134
rect 27344 9716 27396 9722
rect 27344 9658 27396 9664
rect 27160 9172 27212 9178
rect 27160 9114 27212 9120
rect 27252 9172 27304 9178
rect 27252 9114 27304 9120
rect 26884 9036 26936 9042
rect 26884 8978 26936 8984
rect 26976 9036 27028 9042
rect 26976 8978 27028 8984
rect 26608 8832 26660 8838
rect 26608 8774 26660 8780
rect 26896 8090 26924 8978
rect 27172 8566 27200 9114
rect 27356 8634 27384 9658
rect 27344 8628 27396 8634
rect 27344 8570 27396 8576
rect 27160 8560 27212 8566
rect 27160 8502 27212 8508
rect 26056 8084 26108 8090
rect 26056 8026 26108 8032
rect 26884 8084 26936 8090
rect 26884 8026 26936 8032
rect 26424 8016 26476 8022
rect 26424 7958 26476 7964
rect 26436 7546 26464 7958
rect 26608 7880 26660 7886
rect 26608 7822 26660 7828
rect 26424 7540 26476 7546
rect 26424 7482 26476 7488
rect 26620 7478 26648 7822
rect 27172 7546 27200 8502
rect 27252 8356 27304 8362
rect 27252 8298 27304 8304
rect 27264 7886 27292 8298
rect 27356 8294 27384 8570
rect 27344 8288 27396 8294
rect 27344 8230 27396 8236
rect 27540 8022 27568 11455
rect 27724 11354 27752 11727
rect 27896 11620 27948 11626
rect 27896 11562 27948 11568
rect 27712 11348 27764 11354
rect 27712 11290 27764 11296
rect 27908 10305 27936 11562
rect 27988 11552 28040 11558
rect 27988 11494 28040 11500
rect 28000 11218 28028 11494
rect 27988 11212 28040 11218
rect 27988 11154 28040 11160
rect 28000 10742 28028 11154
rect 27988 10736 28040 10742
rect 27988 10678 28040 10684
rect 27894 10296 27950 10305
rect 27894 10231 27950 10240
rect 27908 10198 27936 10231
rect 27896 10192 27948 10198
rect 27896 10134 27948 10140
rect 27620 9376 27672 9382
rect 27620 9318 27672 9324
rect 27988 9376 28040 9382
rect 27988 9318 28040 9324
rect 27528 8016 27580 8022
rect 27528 7958 27580 7964
rect 27252 7880 27304 7886
rect 27252 7822 27304 7828
rect 27160 7540 27212 7546
rect 27160 7482 27212 7488
rect 26608 7472 26660 7478
rect 26608 7414 26660 7420
rect 26792 7336 26844 7342
rect 26792 7278 26844 7284
rect 26332 7200 26384 7206
rect 26332 7142 26384 7148
rect 26700 7200 26752 7206
rect 26700 7142 26752 7148
rect 25964 6452 26016 6458
rect 25964 6394 26016 6400
rect 25976 6254 26004 6394
rect 25964 6248 26016 6254
rect 25964 6190 26016 6196
rect 25778 5672 25834 5681
rect 25778 5607 25834 5616
rect 25504 5024 25556 5030
rect 25504 4966 25556 4972
rect 24492 4752 24544 4758
rect 24492 4694 24544 4700
rect 25044 4752 25096 4758
rect 25044 4694 25096 4700
rect 24044 4126 24164 4154
rect 23664 4072 23716 4078
rect 23664 4014 23716 4020
rect 23296 3936 23348 3942
rect 23296 3878 23348 3884
rect 23308 2650 23336 3878
rect 23676 3738 23704 4014
rect 23848 4004 23900 4010
rect 23848 3946 23900 3952
rect 23664 3732 23716 3738
rect 23664 3674 23716 3680
rect 23860 3670 23888 3946
rect 23848 3664 23900 3670
rect 23848 3606 23900 3612
rect 23480 3392 23532 3398
rect 23480 3334 23532 3340
rect 23492 2990 23520 3334
rect 24044 3194 24072 4126
rect 24504 4010 24532 4694
rect 24492 4004 24544 4010
rect 24492 3946 24544 3952
rect 25056 3942 25084 4694
rect 25228 4616 25280 4622
rect 25228 4558 25280 4564
rect 25240 3942 25268 4558
rect 25412 4276 25464 4282
rect 25412 4218 25464 4224
rect 24584 3936 24636 3942
rect 24584 3878 24636 3884
rect 25044 3936 25096 3942
rect 25044 3878 25096 3884
rect 25228 3936 25280 3942
rect 25228 3878 25280 3884
rect 24032 3188 24084 3194
rect 24032 3130 24084 3136
rect 23480 2984 23532 2990
rect 23480 2926 23532 2932
rect 23296 2644 23348 2650
rect 23296 2586 23348 2592
rect 24596 2553 24624 3878
rect 25056 3670 25084 3878
rect 25044 3664 25096 3670
rect 25044 3606 25096 3612
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24780 2922 24808 3334
rect 24768 2916 24820 2922
rect 24768 2858 24820 2864
rect 24780 2689 24808 2858
rect 25056 2854 25084 3606
rect 25044 2848 25096 2854
rect 25096 2808 25176 2836
rect 25044 2790 25096 2796
rect 24766 2680 24822 2689
rect 24766 2615 24822 2624
rect 25148 2582 25176 2808
rect 25136 2576 25188 2582
rect 24582 2544 24638 2553
rect 25136 2518 25188 2524
rect 24582 2479 24638 2488
rect 25148 2446 25176 2518
rect 25136 2440 25188 2446
rect 25136 2382 25188 2388
rect 25240 1873 25268 3878
rect 25424 3058 25452 4218
rect 25516 4078 25544 4966
rect 25596 4548 25648 4554
rect 25596 4490 25648 4496
rect 25504 4072 25556 4078
rect 25504 4014 25556 4020
rect 25516 3738 25544 4014
rect 25504 3732 25556 3738
rect 25504 3674 25556 3680
rect 25412 3052 25464 3058
rect 25412 2994 25464 3000
rect 25424 2446 25452 2994
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 25608 2378 25636 4490
rect 26056 3936 26108 3942
rect 26056 3878 26108 3884
rect 26068 3534 26096 3878
rect 26056 3528 26108 3534
rect 26056 3470 26108 3476
rect 26068 3194 26096 3470
rect 26056 3188 26108 3194
rect 26056 3130 26108 3136
rect 26240 2440 26292 2446
rect 26238 2408 26240 2417
rect 26292 2408 26294 2417
rect 25596 2372 25648 2378
rect 26238 2343 26294 2352
rect 25596 2314 25648 2320
rect 26252 2310 26280 2343
rect 26240 2304 26292 2310
rect 26240 2246 26292 2252
rect 25226 1864 25282 1873
rect 25226 1799 25282 1808
rect 23110 54 23244 82
rect 26344 82 26372 7142
rect 26712 6866 26740 7142
rect 26804 7002 26832 7278
rect 27172 7274 27200 7482
rect 27160 7268 27212 7274
rect 27160 7210 27212 7216
rect 26792 6996 26844 7002
rect 26792 6938 26844 6944
rect 26516 6860 26568 6866
rect 26516 6802 26568 6808
rect 26700 6860 26752 6866
rect 26700 6802 26752 6808
rect 26528 6390 26556 6802
rect 26516 6384 26568 6390
rect 26516 6326 26568 6332
rect 26516 6248 26568 6254
rect 26516 6190 26568 6196
rect 26528 5574 26556 6190
rect 26712 5914 26740 6802
rect 26792 6248 26844 6254
rect 26792 6190 26844 6196
rect 26700 5908 26752 5914
rect 26700 5850 26752 5856
rect 26516 5568 26568 5574
rect 26516 5510 26568 5516
rect 26700 5296 26752 5302
rect 26700 5238 26752 5244
rect 26712 5098 26740 5238
rect 26700 5092 26752 5098
rect 26700 5034 26752 5040
rect 26516 5024 26568 5030
rect 26516 4966 26568 4972
rect 26424 3596 26476 3602
rect 26528 3584 26556 4966
rect 26608 4616 26660 4622
rect 26608 4558 26660 4564
rect 26620 3738 26648 4558
rect 26712 4214 26740 5034
rect 26804 4826 26832 6190
rect 26976 6180 27028 6186
rect 26976 6122 27028 6128
rect 26988 5778 27016 6122
rect 27172 5846 27200 7210
rect 27264 6905 27292 7822
rect 27250 6896 27306 6905
rect 27250 6831 27306 6840
rect 27540 6458 27568 7958
rect 27632 7546 27660 9318
rect 27896 8832 27948 8838
rect 27896 8774 27948 8780
rect 27712 8356 27764 8362
rect 27712 8298 27764 8304
rect 27724 8090 27752 8298
rect 27712 8084 27764 8090
rect 27712 8026 27764 8032
rect 27908 7954 27936 8774
rect 27896 7948 27948 7954
rect 27896 7890 27948 7896
rect 27908 7546 27936 7890
rect 27620 7540 27672 7546
rect 27620 7482 27672 7488
rect 27896 7540 27948 7546
rect 27896 7482 27948 7488
rect 28000 7002 28028 9318
rect 28184 7936 28212 15943
rect 28264 15914 28316 15920
rect 28276 15502 28304 15914
rect 28552 15910 28580 16662
rect 28540 15904 28592 15910
rect 28540 15846 28592 15852
rect 28552 15706 28580 15846
rect 28540 15700 28592 15706
rect 28540 15642 28592 15648
rect 28264 15496 28316 15502
rect 28264 15438 28316 15444
rect 28276 15162 28304 15438
rect 28264 15156 28316 15162
rect 28264 15098 28316 15104
rect 28552 15026 28580 15642
rect 28540 15020 28592 15026
rect 28540 14962 28592 14968
rect 28356 14816 28408 14822
rect 28356 14758 28408 14764
rect 28368 14550 28396 14758
rect 28356 14544 28408 14550
rect 28356 14486 28408 14492
rect 28368 14074 28396 14486
rect 28356 14068 28408 14074
rect 28356 14010 28408 14016
rect 28644 13870 28672 16934
rect 28828 16794 28856 18158
rect 29000 18080 29052 18086
rect 29000 18022 29052 18028
rect 29012 17678 29040 18022
rect 29000 17672 29052 17678
rect 29000 17614 29052 17620
rect 29012 17338 29040 17614
rect 29092 17536 29144 17542
rect 29092 17478 29144 17484
rect 29104 17338 29132 17478
rect 29000 17332 29052 17338
rect 29000 17274 29052 17280
rect 29092 17332 29144 17338
rect 29092 17274 29144 17280
rect 29184 17128 29236 17134
rect 29184 17070 29236 17076
rect 28816 16788 28868 16794
rect 28816 16730 28868 16736
rect 29196 16454 29224 17070
rect 29656 16658 29684 22374
rect 29840 22234 29868 22442
rect 30024 22234 30052 22578
rect 30116 22506 30144 22646
rect 30944 22642 30972 23446
rect 31024 23044 31076 23050
rect 31024 22986 31076 22992
rect 31036 22778 31064 22986
rect 31024 22772 31076 22778
rect 31024 22714 31076 22720
rect 30932 22636 30984 22642
rect 30932 22578 30984 22584
rect 30104 22500 30156 22506
rect 30104 22442 30156 22448
rect 29828 22228 29880 22234
rect 29828 22170 29880 22176
rect 30012 22228 30064 22234
rect 30012 22170 30064 22176
rect 29736 21480 29788 21486
rect 29736 21422 29788 21428
rect 29748 21078 29776 21422
rect 30012 21412 30064 21418
rect 30012 21354 30064 21360
rect 29828 21344 29880 21350
rect 29828 21286 29880 21292
rect 29736 21072 29788 21078
rect 29736 21014 29788 21020
rect 29748 18834 29776 21014
rect 29840 20398 29868 21286
rect 30024 20466 30052 21354
rect 30116 21010 30144 22442
rect 30944 22098 30972 22578
rect 30932 22092 30984 22098
rect 30932 22034 30984 22040
rect 30944 21690 30972 22034
rect 31220 21690 31248 25910
rect 31484 25832 31536 25838
rect 31484 25774 31536 25780
rect 30932 21684 30984 21690
rect 30932 21626 30984 21632
rect 31208 21684 31260 21690
rect 31208 21626 31260 21632
rect 30656 21548 30708 21554
rect 30656 21490 30708 21496
rect 30668 21457 30696 21490
rect 31220 21486 31248 21626
rect 31496 21486 31524 25774
rect 31668 25696 31720 25702
rect 31668 25638 31720 25644
rect 31680 24614 31708 25638
rect 31864 25498 31892 26318
rect 32232 25906 32260 26726
rect 32508 26518 32536 27084
rect 32588 27066 32640 27072
rect 32312 26512 32364 26518
rect 32312 26454 32364 26460
rect 32496 26512 32548 26518
rect 32496 26454 32548 26460
rect 32220 25900 32272 25906
rect 32220 25842 32272 25848
rect 32324 25702 32352 26454
rect 32312 25696 32364 25702
rect 32312 25638 32364 25644
rect 31852 25492 31904 25498
rect 31852 25434 31904 25440
rect 32324 25430 32352 25638
rect 32312 25424 32364 25430
rect 32312 25366 32364 25372
rect 32588 25288 32640 25294
rect 32588 25230 32640 25236
rect 32600 24682 32628 25230
rect 31760 24676 31812 24682
rect 31760 24618 31812 24624
rect 32404 24676 32456 24682
rect 32404 24618 32456 24624
rect 32588 24676 32640 24682
rect 32588 24618 32640 24624
rect 31668 24608 31720 24614
rect 31668 24550 31720 24556
rect 31772 24410 31800 24618
rect 32416 24585 32444 24618
rect 32402 24576 32458 24585
rect 32402 24511 32458 24520
rect 32600 24410 32628 24618
rect 31760 24404 31812 24410
rect 31760 24346 31812 24352
rect 32588 24404 32640 24410
rect 32588 24346 32640 24352
rect 31760 24268 31812 24274
rect 31760 24210 31812 24216
rect 31772 23526 31800 24210
rect 32692 24206 32720 30688
rect 32784 29238 32812 32370
rect 33048 32224 33100 32230
rect 33048 32166 33100 32172
rect 32864 31680 32916 31686
rect 32864 31622 32916 31628
rect 32876 31482 32904 31622
rect 32864 31476 32916 31482
rect 32864 31418 32916 31424
rect 32876 30938 32904 31418
rect 32864 30932 32916 30938
rect 32864 30874 32916 30880
rect 32876 30394 32904 30874
rect 33060 30870 33088 32166
rect 33968 31816 34020 31822
rect 33968 31758 34020 31764
rect 33980 31142 34008 31758
rect 33416 31136 33468 31142
rect 33416 31078 33468 31084
rect 33968 31136 34020 31142
rect 33968 31078 34020 31084
rect 33324 30932 33376 30938
rect 33324 30874 33376 30880
rect 33048 30864 33100 30870
rect 33048 30806 33100 30812
rect 32956 30660 33008 30666
rect 32956 30602 33008 30608
rect 32864 30388 32916 30394
rect 32864 30330 32916 30336
rect 32772 29232 32824 29238
rect 32772 29174 32824 29180
rect 32968 29170 32996 30602
rect 33060 30394 33088 30806
rect 33232 30728 33284 30734
rect 33232 30670 33284 30676
rect 33048 30388 33100 30394
rect 33048 30330 33100 30336
rect 33048 29640 33100 29646
rect 33048 29582 33100 29588
rect 32956 29164 33008 29170
rect 32956 29106 33008 29112
rect 32956 29028 33008 29034
rect 32876 28988 32956 29016
rect 32876 28422 32904 28988
rect 32956 28970 33008 28976
rect 33060 28626 33088 29582
rect 33048 28620 33100 28626
rect 33048 28562 33100 28568
rect 32864 28416 32916 28422
rect 32864 28358 32916 28364
rect 32876 28150 32904 28358
rect 32864 28144 32916 28150
rect 32864 28086 32916 28092
rect 33244 27878 33272 30670
rect 33336 30122 33364 30874
rect 33428 30122 33456 31078
rect 33506 30832 33562 30841
rect 33506 30767 33562 30776
rect 33520 30734 33548 30767
rect 33508 30728 33560 30734
rect 33508 30670 33560 30676
rect 33692 30728 33744 30734
rect 33692 30670 33744 30676
rect 33704 30122 33732 30670
rect 33980 30326 34008 31078
rect 33968 30320 34020 30326
rect 33968 30262 34020 30268
rect 33324 30116 33376 30122
rect 33324 30058 33376 30064
rect 33416 30116 33468 30122
rect 33416 30058 33468 30064
rect 33692 30116 33744 30122
rect 33692 30058 33744 30064
rect 33336 29850 33364 30058
rect 33324 29844 33376 29850
rect 33324 29786 33376 29792
rect 33428 29714 33456 30058
rect 33416 29708 33468 29714
rect 33416 29650 33468 29656
rect 33508 29232 33560 29238
rect 33508 29174 33560 29180
rect 33416 28756 33468 28762
rect 33416 28698 33468 28704
rect 33428 28150 33456 28698
rect 33416 28144 33468 28150
rect 33416 28086 33468 28092
rect 33428 27946 33456 28086
rect 33416 27940 33468 27946
rect 33416 27882 33468 27888
rect 33232 27872 33284 27878
rect 33232 27814 33284 27820
rect 32864 27464 32916 27470
rect 32864 27406 32916 27412
rect 32876 26790 32904 27406
rect 33520 26994 33548 29174
rect 33598 28928 33654 28937
rect 33598 28863 33654 28872
rect 33508 26988 33560 26994
rect 33508 26930 33560 26936
rect 33324 26920 33376 26926
rect 33324 26862 33376 26868
rect 32864 26784 32916 26790
rect 32864 26726 32916 26732
rect 32680 24200 32732 24206
rect 32680 24142 32732 24148
rect 31760 23520 31812 23526
rect 31758 23488 31760 23497
rect 31812 23488 31814 23497
rect 32876 23474 32904 26726
rect 33336 26246 33364 26862
rect 33324 26240 33376 26246
rect 33324 26182 33376 26188
rect 33232 25832 33284 25838
rect 33232 25774 33284 25780
rect 33244 23730 33272 25774
rect 33232 23724 33284 23730
rect 33232 23666 33284 23672
rect 33336 23594 33364 26182
rect 33416 25696 33468 25702
rect 33416 25638 33468 25644
rect 33324 23588 33376 23594
rect 33324 23530 33376 23536
rect 31758 23423 31814 23432
rect 32784 23446 32904 23474
rect 32956 23520 33008 23526
rect 32956 23462 33008 23468
rect 31668 22568 31720 22574
rect 31668 22510 31720 22516
rect 31680 22234 31708 22510
rect 31668 22228 31720 22234
rect 31668 22170 31720 22176
rect 31576 22024 31628 22030
rect 31576 21966 31628 21972
rect 31208 21480 31260 21486
rect 30654 21448 30710 21457
rect 31208 21422 31260 21428
rect 31484 21480 31536 21486
rect 31484 21422 31536 21428
rect 30654 21383 30710 21392
rect 30104 21004 30156 21010
rect 30104 20946 30156 20952
rect 30932 21004 30984 21010
rect 30932 20946 30984 20952
rect 30944 20602 30972 20946
rect 31116 20868 31168 20874
rect 31116 20810 31168 20816
rect 30932 20596 30984 20602
rect 30932 20538 30984 20544
rect 31128 20534 31156 20810
rect 31484 20800 31536 20806
rect 31484 20742 31536 20748
rect 31116 20528 31168 20534
rect 31116 20470 31168 20476
rect 30012 20460 30064 20466
rect 30012 20402 30064 20408
rect 29828 20392 29880 20398
rect 29880 20352 29960 20380
rect 29828 20334 29880 20340
rect 29932 20262 29960 20352
rect 29920 20256 29972 20262
rect 29920 20198 29972 20204
rect 29828 19304 29880 19310
rect 29828 19246 29880 19252
rect 29840 18902 29868 19246
rect 29932 19174 29960 20198
rect 30024 20058 30052 20402
rect 30194 20360 30250 20369
rect 30104 20324 30156 20330
rect 30156 20304 30194 20312
rect 31128 20330 31156 20470
rect 30156 20295 30250 20304
rect 31116 20324 31168 20330
rect 30156 20284 30236 20295
rect 30104 20266 30156 20272
rect 31116 20266 31168 20272
rect 30656 20256 30708 20262
rect 30656 20198 30708 20204
rect 30012 20052 30064 20058
rect 30012 19994 30064 20000
rect 30668 19990 30696 20198
rect 30656 19984 30708 19990
rect 30656 19926 30708 19932
rect 30668 19446 30696 19926
rect 31392 19848 31444 19854
rect 31392 19790 31444 19796
rect 31208 19780 31260 19786
rect 31208 19722 31260 19728
rect 30656 19440 30708 19446
rect 30656 19382 30708 19388
rect 29920 19168 29972 19174
rect 29920 19110 29972 19116
rect 30564 19168 30616 19174
rect 30564 19110 30616 19116
rect 30840 19168 30892 19174
rect 30840 19110 30892 19116
rect 29828 18896 29880 18902
rect 29828 18838 29880 18844
rect 29736 18828 29788 18834
rect 29736 18770 29788 18776
rect 29748 18426 29776 18770
rect 29736 18420 29788 18426
rect 29736 18362 29788 18368
rect 29748 17814 29776 18362
rect 30576 18086 30604 19110
rect 30852 18902 30880 19110
rect 31220 18902 31248 19722
rect 31404 19514 31432 19790
rect 31392 19508 31444 19514
rect 31392 19450 31444 19456
rect 30840 18896 30892 18902
rect 30840 18838 30892 18844
rect 31208 18896 31260 18902
rect 31260 18856 31340 18884
rect 31208 18838 31260 18844
rect 30656 18216 30708 18222
rect 30656 18158 30708 18164
rect 30564 18080 30616 18086
rect 30564 18022 30616 18028
rect 29736 17808 29788 17814
rect 29736 17750 29788 17756
rect 30288 17740 30340 17746
rect 30288 17682 30340 17688
rect 30472 17740 30524 17746
rect 30472 17682 30524 17688
rect 30300 17066 30328 17682
rect 30484 17338 30512 17682
rect 30472 17332 30524 17338
rect 30472 17274 30524 17280
rect 30288 17060 30340 17066
rect 30288 17002 30340 17008
rect 30484 16658 30512 17274
rect 29644 16652 29696 16658
rect 29644 16594 29696 16600
rect 29736 16652 29788 16658
rect 29736 16594 29788 16600
rect 30472 16652 30524 16658
rect 30472 16594 30524 16600
rect 29184 16448 29236 16454
rect 29184 16390 29236 16396
rect 29196 15706 29224 16390
rect 29656 16250 29684 16594
rect 29644 16244 29696 16250
rect 29644 16186 29696 16192
rect 29656 16017 29684 16186
rect 29642 16008 29698 16017
rect 29642 15943 29698 15952
rect 29748 15706 29776 16594
rect 30196 16584 30248 16590
rect 30196 16526 30248 16532
rect 30208 16114 30236 16526
rect 30196 16108 30248 16114
rect 30196 16050 30248 16056
rect 30208 15706 30236 16050
rect 30576 15978 30604 18022
rect 30668 17814 30696 18158
rect 30852 17882 30880 18838
rect 31116 18080 31168 18086
rect 31116 18022 31168 18028
rect 30840 17876 30892 17882
rect 30840 17818 30892 17824
rect 30656 17808 30708 17814
rect 30656 17750 30708 17756
rect 31128 17270 31156 18022
rect 31208 17672 31260 17678
rect 31208 17614 31260 17620
rect 31116 17264 31168 17270
rect 31116 17206 31168 17212
rect 31128 17048 31156 17206
rect 31220 17202 31248 17614
rect 31312 17202 31340 18856
rect 31496 18630 31524 20742
rect 31484 18624 31536 18630
rect 31484 18566 31536 18572
rect 31208 17196 31260 17202
rect 31208 17138 31260 17144
rect 31300 17196 31352 17202
rect 31300 17138 31352 17144
rect 31208 17060 31260 17066
rect 31128 17020 31208 17048
rect 31208 17002 31260 17008
rect 31220 16794 31248 17002
rect 31208 16788 31260 16794
rect 31208 16730 31260 16736
rect 31312 16114 31340 17138
rect 31300 16108 31352 16114
rect 31300 16050 31352 16056
rect 30564 15972 30616 15978
rect 30564 15914 30616 15920
rect 29184 15700 29236 15706
rect 29184 15642 29236 15648
rect 29736 15700 29788 15706
rect 29736 15642 29788 15648
rect 30196 15700 30248 15706
rect 30196 15642 30248 15648
rect 29748 15162 29776 15642
rect 31116 15564 31168 15570
rect 31116 15506 31168 15512
rect 30288 15428 30340 15434
rect 30288 15370 30340 15376
rect 30300 15162 30328 15370
rect 29736 15156 29788 15162
rect 29736 15098 29788 15104
rect 30288 15156 30340 15162
rect 30288 15098 30340 15104
rect 31128 14958 31156 15506
rect 29184 14952 29236 14958
rect 29184 14894 29236 14900
rect 31116 14952 31168 14958
rect 31116 14894 31168 14900
rect 28264 13864 28316 13870
rect 28264 13806 28316 13812
rect 28632 13864 28684 13870
rect 28632 13806 28684 13812
rect 29092 13864 29144 13870
rect 29092 13806 29144 13812
rect 28276 13530 28304 13806
rect 29104 13734 29132 13806
rect 29092 13728 29144 13734
rect 29092 13670 29144 13676
rect 28264 13524 28316 13530
rect 28264 13466 28316 13472
rect 28632 13524 28684 13530
rect 28632 13466 28684 13472
rect 28264 13320 28316 13326
rect 28264 13262 28316 13268
rect 28276 12374 28304 13262
rect 28644 12918 28672 13466
rect 29196 12986 29224 14894
rect 31128 14618 31156 14894
rect 31116 14612 31168 14618
rect 31116 14554 31168 14560
rect 30748 14476 30800 14482
rect 30748 14418 30800 14424
rect 29644 14408 29696 14414
rect 29644 14350 29696 14356
rect 29368 14272 29420 14278
rect 29368 14214 29420 14220
rect 29380 13802 29408 14214
rect 29656 13938 29684 14350
rect 30760 14006 30788 14418
rect 31128 14074 31156 14554
rect 31116 14068 31168 14074
rect 31116 14010 31168 14016
rect 30748 14000 30800 14006
rect 30748 13942 30800 13948
rect 29644 13932 29696 13938
rect 29644 13874 29696 13880
rect 29368 13796 29420 13802
rect 29368 13738 29420 13744
rect 29380 13530 29408 13738
rect 29368 13524 29420 13530
rect 29368 13466 29420 13472
rect 30760 13433 30788 13942
rect 31208 13864 31260 13870
rect 31208 13806 31260 13812
rect 30746 13424 30802 13433
rect 30472 13388 30524 13394
rect 30746 13359 30802 13368
rect 30472 13330 30524 13336
rect 29460 13184 29512 13190
rect 29460 13126 29512 13132
rect 29184 12980 29236 12986
rect 29184 12922 29236 12928
rect 28632 12912 28684 12918
rect 28632 12854 28684 12860
rect 28644 12714 28672 12854
rect 29472 12850 29500 13126
rect 30484 12986 30512 13330
rect 31024 13184 31076 13190
rect 31024 13126 31076 13132
rect 30472 12980 30524 12986
rect 30472 12922 30524 12928
rect 29460 12844 29512 12850
rect 29460 12786 29512 12792
rect 31036 12782 31064 13126
rect 28724 12776 28776 12782
rect 28724 12718 28776 12724
rect 30472 12776 30524 12782
rect 30472 12718 30524 12724
rect 31024 12776 31076 12782
rect 31024 12718 31076 12724
rect 28632 12708 28684 12714
rect 28632 12650 28684 12656
rect 28264 12368 28316 12374
rect 28264 12310 28316 12316
rect 28736 12306 28764 12718
rect 30484 12374 30512 12718
rect 30932 12708 30984 12714
rect 30932 12650 30984 12656
rect 30944 12374 30972 12650
rect 31220 12442 31248 13806
rect 31208 12436 31260 12442
rect 31208 12378 31260 12384
rect 30472 12368 30524 12374
rect 30472 12310 30524 12316
rect 30932 12368 30984 12374
rect 30932 12310 30984 12316
rect 28724 12300 28776 12306
rect 28724 12242 28776 12248
rect 28356 11756 28408 11762
rect 28356 11698 28408 11704
rect 28264 11620 28316 11626
rect 28264 11562 28316 11568
rect 28276 11354 28304 11562
rect 28264 11348 28316 11354
rect 28264 11290 28316 11296
rect 28264 11212 28316 11218
rect 28264 11154 28316 11160
rect 28276 10810 28304 11154
rect 28368 11014 28396 11698
rect 28736 11558 28764 12242
rect 30564 12232 30616 12238
rect 30564 12174 30616 12180
rect 30288 12096 30340 12102
rect 30288 12038 30340 12044
rect 30300 11694 30328 12038
rect 30288 11688 30340 11694
rect 30288 11630 30340 11636
rect 28724 11552 28776 11558
rect 28724 11494 28776 11500
rect 28736 11121 28764 11494
rect 30300 11286 30328 11630
rect 30576 11626 30604 12174
rect 30944 11898 30972 12310
rect 30932 11892 30984 11898
rect 30932 11834 30984 11840
rect 30380 11620 30432 11626
rect 30380 11562 30432 11568
rect 30564 11620 30616 11626
rect 30564 11562 30616 11568
rect 29184 11280 29236 11286
rect 29184 11222 29236 11228
rect 30288 11280 30340 11286
rect 30288 11222 30340 11228
rect 28722 11112 28778 11121
rect 28778 11070 28856 11098
rect 28722 11047 28778 11056
rect 28356 11008 28408 11014
rect 28356 10950 28408 10956
rect 28368 10810 28396 10950
rect 28264 10804 28316 10810
rect 28264 10746 28316 10752
rect 28356 10804 28408 10810
rect 28356 10746 28408 10752
rect 28724 9988 28776 9994
rect 28724 9930 28776 9936
rect 28736 9722 28764 9930
rect 28724 9716 28776 9722
rect 28724 9658 28776 9664
rect 28632 9036 28684 9042
rect 28632 8978 28684 8984
rect 28644 8634 28672 8978
rect 28736 8974 28764 9658
rect 28724 8968 28776 8974
rect 28724 8910 28776 8916
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 28356 8492 28408 8498
rect 28356 8434 28408 8440
rect 28368 8401 28396 8434
rect 28354 8392 28410 8401
rect 28354 8327 28410 8336
rect 28264 7948 28316 7954
rect 28184 7908 28264 7936
rect 28264 7890 28316 7896
rect 27988 6996 28040 7002
rect 27988 6938 28040 6944
rect 27528 6452 27580 6458
rect 27528 6394 27580 6400
rect 27540 6186 27568 6394
rect 28000 6322 28028 6938
rect 28368 6322 28396 8327
rect 27988 6316 28040 6322
rect 27988 6258 28040 6264
rect 28356 6316 28408 6322
rect 28356 6258 28408 6264
rect 27528 6180 27580 6186
rect 27528 6122 27580 6128
rect 28644 5914 28672 8570
rect 28828 7478 28856 11070
rect 29196 10742 29224 11222
rect 29736 11144 29788 11150
rect 29736 11086 29788 11092
rect 29276 11008 29328 11014
rect 29276 10950 29328 10956
rect 29184 10736 29236 10742
rect 29184 10678 29236 10684
rect 29196 10130 29224 10678
rect 29288 10606 29316 10950
rect 29748 10810 29776 11086
rect 29736 10804 29788 10810
rect 29736 10746 29788 10752
rect 29276 10600 29328 10606
rect 29276 10542 29328 10548
rect 29184 10124 29236 10130
rect 29184 10066 29236 10072
rect 29644 9512 29696 9518
rect 29644 9454 29696 9460
rect 29656 9110 29684 9454
rect 29644 9104 29696 9110
rect 29644 9046 29696 9052
rect 29000 9036 29052 9042
rect 29000 8978 29052 8984
rect 29012 8294 29040 8978
rect 29000 8288 29052 8294
rect 29000 8230 29052 8236
rect 29552 8288 29604 8294
rect 29552 8230 29604 8236
rect 29012 8022 29040 8230
rect 29564 8090 29592 8230
rect 29552 8084 29604 8090
rect 29552 8026 29604 8032
rect 29000 8016 29052 8022
rect 29000 7958 29052 7964
rect 28816 7472 28868 7478
rect 28816 7414 28868 7420
rect 29012 7206 29040 7958
rect 29460 7948 29512 7954
rect 29460 7890 29512 7896
rect 29472 7546 29500 7890
rect 29748 7546 29776 10746
rect 30288 9716 30340 9722
rect 30288 9658 30340 9664
rect 29920 8968 29972 8974
rect 29920 8910 29972 8916
rect 29932 8634 29960 8910
rect 30300 8634 30328 9658
rect 29920 8628 29972 8634
rect 29920 8570 29972 8576
rect 30288 8628 30340 8634
rect 30288 8570 30340 8576
rect 30300 8362 30328 8570
rect 30288 8356 30340 8362
rect 30288 8298 30340 8304
rect 29460 7540 29512 7546
rect 29460 7482 29512 7488
rect 29736 7540 29788 7546
rect 29736 7482 29788 7488
rect 29000 7200 29052 7206
rect 29000 7142 29052 7148
rect 28908 6928 28960 6934
rect 28908 6870 28960 6876
rect 28724 6792 28776 6798
rect 28724 6734 28776 6740
rect 28632 5908 28684 5914
rect 28632 5850 28684 5856
rect 27160 5840 27212 5846
rect 27160 5782 27212 5788
rect 27528 5840 27580 5846
rect 27528 5782 27580 5788
rect 26976 5772 27028 5778
rect 26976 5714 27028 5720
rect 26988 5370 27016 5714
rect 27160 5568 27212 5574
rect 27160 5510 27212 5516
rect 26976 5364 27028 5370
rect 26976 5306 27028 5312
rect 26792 4820 26844 4826
rect 26792 4762 26844 4768
rect 26700 4208 26752 4214
rect 26700 4150 26752 4156
rect 26712 4010 26740 4150
rect 26804 4146 26832 4762
rect 27068 4752 27120 4758
rect 27068 4694 27120 4700
rect 26792 4140 26844 4146
rect 26792 4082 26844 4088
rect 26700 4004 26752 4010
rect 26700 3946 26752 3952
rect 27080 3942 27108 4694
rect 27068 3936 27120 3942
rect 27068 3878 27120 3884
rect 26608 3732 26660 3738
rect 26608 3674 26660 3680
rect 26476 3556 26556 3584
rect 26424 3538 26476 3544
rect 26528 3194 26556 3556
rect 26976 3528 27028 3534
rect 26976 3470 27028 3476
rect 26988 3194 27016 3470
rect 26516 3188 26568 3194
rect 26516 3130 26568 3136
rect 26976 3188 27028 3194
rect 26976 3130 27028 3136
rect 27080 2922 27108 3878
rect 27172 3194 27200 5510
rect 27540 5302 27568 5782
rect 28736 5710 28764 6734
rect 28920 6118 28948 6870
rect 29472 6866 29500 7482
rect 30288 6996 30340 7002
rect 30288 6938 30340 6944
rect 29460 6860 29512 6866
rect 29460 6802 29512 6808
rect 30196 6860 30248 6866
rect 30196 6802 30248 6808
rect 30012 6792 30064 6798
rect 30012 6734 30064 6740
rect 29644 6656 29696 6662
rect 29644 6598 29696 6604
rect 29656 6322 29684 6598
rect 29644 6316 29696 6322
rect 29644 6258 29696 6264
rect 29460 6180 29512 6186
rect 29460 6122 29512 6128
rect 28908 6112 28960 6118
rect 28908 6054 28960 6060
rect 28724 5704 28776 5710
rect 28724 5646 28776 5652
rect 27528 5296 27580 5302
rect 27528 5238 27580 5244
rect 28816 5092 28868 5098
rect 28816 5034 28868 5040
rect 28448 5024 28500 5030
rect 28448 4966 28500 4972
rect 28172 4684 28224 4690
rect 28172 4626 28224 4632
rect 27344 4616 27396 4622
rect 27344 4558 27396 4564
rect 27356 4010 27384 4558
rect 28184 4214 28212 4626
rect 28172 4208 28224 4214
rect 28172 4150 28224 4156
rect 27344 4004 27396 4010
rect 27344 3946 27396 3952
rect 27356 3670 27384 3946
rect 28264 3936 28316 3942
rect 28264 3878 28316 3884
rect 27344 3664 27396 3670
rect 27344 3606 27396 3612
rect 28172 3664 28224 3670
rect 28172 3606 28224 3612
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 27160 3188 27212 3194
rect 27160 3130 27212 3136
rect 27172 2990 27200 3130
rect 27724 3058 27752 3334
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 27160 2984 27212 2990
rect 27160 2926 27212 2932
rect 27068 2916 27120 2922
rect 27068 2858 27120 2864
rect 27080 2582 27108 2858
rect 27724 2650 27752 2994
rect 28184 2854 28212 3606
rect 28172 2848 28224 2854
rect 28172 2790 28224 2796
rect 27712 2644 27764 2650
rect 27712 2586 27764 2592
rect 28276 2582 28304 3878
rect 28356 2916 28408 2922
rect 28356 2858 28408 2864
rect 28368 2582 28396 2858
rect 27068 2576 27120 2582
rect 27068 2518 27120 2524
rect 28264 2576 28316 2582
rect 28264 2518 28316 2524
rect 28356 2576 28408 2582
rect 28356 2518 28408 2524
rect 28460 2378 28488 4966
rect 28632 4480 28684 4486
rect 28632 4422 28684 4428
rect 28644 3738 28672 4422
rect 28632 3732 28684 3738
rect 28632 3674 28684 3680
rect 28828 3670 28856 5034
rect 28920 5030 28948 6054
rect 29368 5568 29420 5574
rect 29368 5510 29420 5516
rect 29092 5228 29144 5234
rect 29092 5170 29144 5176
rect 28908 5024 28960 5030
rect 28908 4966 28960 4972
rect 29104 4758 29132 5170
rect 29380 5098 29408 5510
rect 29368 5092 29420 5098
rect 29368 5034 29420 5040
rect 29092 4752 29144 4758
rect 29092 4694 29144 4700
rect 29104 4214 29132 4694
rect 29092 4208 29144 4214
rect 29092 4150 29144 4156
rect 29472 4010 29500 6122
rect 29552 5568 29604 5574
rect 29552 5510 29604 5516
rect 29564 4690 29592 5510
rect 29552 4684 29604 4690
rect 29552 4626 29604 4632
rect 29656 4554 29684 6258
rect 30024 6186 30052 6734
rect 30208 6458 30236 6802
rect 30196 6452 30248 6458
rect 30196 6394 30248 6400
rect 30012 6180 30064 6186
rect 30012 6122 30064 6128
rect 29828 5840 29880 5846
rect 29828 5782 29880 5788
rect 29840 5370 29868 5782
rect 30024 5642 30052 6122
rect 30300 5778 30328 6938
rect 30288 5772 30340 5778
rect 30288 5714 30340 5720
rect 30104 5704 30156 5710
rect 30104 5646 30156 5652
rect 30196 5704 30248 5710
rect 30196 5646 30248 5652
rect 30012 5636 30064 5642
rect 30012 5578 30064 5584
rect 29828 5364 29880 5370
rect 29828 5306 29880 5312
rect 29828 5228 29880 5234
rect 29828 5170 29880 5176
rect 29644 4548 29696 4554
rect 29644 4490 29696 4496
rect 29840 4146 29868 5170
rect 30012 4480 30064 4486
rect 30012 4422 30064 4428
rect 29828 4140 29880 4146
rect 29828 4082 29880 4088
rect 29460 4004 29512 4010
rect 29460 3946 29512 3952
rect 28816 3664 28868 3670
rect 28816 3606 28868 3612
rect 28828 3058 28856 3606
rect 29472 3602 29500 3946
rect 30024 3738 30052 4422
rect 30012 3732 30064 3738
rect 30012 3674 30064 3680
rect 29460 3596 29512 3602
rect 29460 3538 29512 3544
rect 29000 3528 29052 3534
rect 29000 3470 29052 3476
rect 29012 3194 29040 3470
rect 29000 3188 29052 3194
rect 29000 3130 29052 3136
rect 29920 3188 29972 3194
rect 29920 3130 29972 3136
rect 28816 3052 28868 3058
rect 28816 2994 28868 3000
rect 29932 2582 29960 3130
rect 30024 2990 30052 3674
rect 30012 2984 30064 2990
rect 30012 2926 30064 2932
rect 29920 2576 29972 2582
rect 29920 2518 29972 2524
rect 30116 2446 30144 5646
rect 30104 2440 30156 2446
rect 30104 2382 30156 2388
rect 28448 2372 28500 2378
rect 28448 2314 28500 2320
rect 26698 82 26754 480
rect 26344 54 26754 82
rect 30208 82 30236 5646
rect 30300 4826 30328 5714
rect 30392 5166 30420 11562
rect 30576 11354 30604 11562
rect 30564 11348 30616 11354
rect 30564 11290 30616 11296
rect 30564 11144 30616 11150
rect 30564 11086 30616 11092
rect 30576 10674 30604 11086
rect 30944 10810 30972 11834
rect 30932 10804 30984 10810
rect 30932 10746 30984 10752
rect 30564 10668 30616 10674
rect 30564 10610 30616 10616
rect 30944 10470 30972 10746
rect 30932 10464 30984 10470
rect 30932 10406 30984 10412
rect 31484 10464 31536 10470
rect 31484 10406 31536 10412
rect 30944 10130 30972 10406
rect 30932 10124 30984 10130
rect 30932 10066 30984 10072
rect 30944 9722 30972 10066
rect 31208 10056 31260 10062
rect 31208 9998 31260 10004
rect 31220 9722 31248 9998
rect 30932 9716 30984 9722
rect 30932 9658 30984 9664
rect 31208 9716 31260 9722
rect 31208 9658 31260 9664
rect 31496 9586 31524 10406
rect 31484 9580 31536 9586
rect 31484 9522 31536 9528
rect 30564 9376 30616 9382
rect 30564 9318 30616 9324
rect 30576 7954 30604 9318
rect 30656 9036 30708 9042
rect 30656 8978 30708 8984
rect 30564 7948 30616 7954
rect 30564 7890 30616 7896
rect 30564 7812 30616 7818
rect 30668 7800 30696 8978
rect 30932 8968 30984 8974
rect 30932 8910 30984 8916
rect 30616 7772 30696 7800
rect 30564 7754 30616 7760
rect 30576 7342 30604 7754
rect 30564 7336 30616 7342
rect 30564 7278 30616 7284
rect 30576 6866 30604 7278
rect 30840 7268 30892 7274
rect 30840 7210 30892 7216
rect 30852 6866 30880 7210
rect 30564 6860 30616 6866
rect 30564 6802 30616 6808
rect 30840 6860 30892 6866
rect 30840 6802 30892 6808
rect 30840 6452 30892 6458
rect 30840 6394 30892 6400
rect 30852 5370 30880 6394
rect 30944 5914 30972 8910
rect 31300 6996 31352 7002
rect 31300 6938 31352 6944
rect 31312 6322 31340 6938
rect 31300 6316 31352 6322
rect 31300 6258 31352 6264
rect 30932 5908 30984 5914
rect 30932 5850 30984 5856
rect 30840 5364 30892 5370
rect 30840 5306 30892 5312
rect 30380 5160 30432 5166
rect 30380 5102 30432 5108
rect 30852 5030 30880 5306
rect 30944 5234 30972 5850
rect 30932 5228 30984 5234
rect 30932 5170 30984 5176
rect 31024 5092 31076 5098
rect 31024 5034 31076 5040
rect 30840 5024 30892 5030
rect 30840 4966 30892 4972
rect 30288 4820 30340 4826
rect 30288 4762 30340 4768
rect 30852 4758 30880 4966
rect 30840 4752 30892 4758
rect 30840 4694 30892 4700
rect 30380 4684 30432 4690
rect 30380 4626 30432 4632
rect 30392 4282 30420 4626
rect 30932 4480 30984 4486
rect 30932 4422 30984 4428
rect 30380 4276 30432 4282
rect 30380 4218 30432 4224
rect 30944 4010 30972 4422
rect 31036 4282 31064 5034
rect 31024 4276 31076 4282
rect 31024 4218 31076 4224
rect 31036 4010 31064 4218
rect 30932 4004 30984 4010
rect 30932 3946 30984 3952
rect 31024 4004 31076 4010
rect 31024 3946 31076 3952
rect 30564 3664 30616 3670
rect 30748 3664 30800 3670
rect 30616 3624 30696 3652
rect 30564 3606 30616 3612
rect 30564 2916 30616 2922
rect 30564 2858 30616 2864
rect 30576 2650 30604 2858
rect 30564 2644 30616 2650
rect 30564 2586 30616 2592
rect 30668 2582 30696 3624
rect 30748 3606 30800 3612
rect 30760 3194 30788 3606
rect 31208 3528 31260 3534
rect 31208 3470 31260 3476
rect 30748 3188 30800 3194
rect 30748 3130 30800 3136
rect 31220 3058 31248 3470
rect 31208 3052 31260 3058
rect 31208 2994 31260 3000
rect 30656 2576 30708 2582
rect 30656 2518 30708 2524
rect 31588 2514 31616 21966
rect 31772 19310 31800 23423
rect 32588 23248 32640 23254
rect 32588 23190 32640 23196
rect 32128 23112 32180 23118
rect 32128 23054 32180 23060
rect 32140 22642 32168 23054
rect 32128 22636 32180 22642
rect 32128 22578 32180 22584
rect 32600 22438 32628 23190
rect 32784 23089 32812 23446
rect 32968 23322 32996 23462
rect 32956 23316 33008 23322
rect 32956 23258 33008 23264
rect 32770 23080 32826 23089
rect 32770 23015 32826 23024
rect 32680 22772 32732 22778
rect 32680 22714 32732 22720
rect 32588 22432 32640 22438
rect 32588 22374 32640 22380
rect 32404 22092 32456 22098
rect 32404 22034 32456 22040
rect 32416 22001 32444 22034
rect 32402 21992 32458 22001
rect 32402 21927 32458 21936
rect 32416 21554 32444 21927
rect 32496 21684 32548 21690
rect 32496 21626 32548 21632
rect 32404 21548 32456 21554
rect 32404 21490 32456 21496
rect 32128 21344 32180 21350
rect 32128 21286 32180 21292
rect 32036 20936 32088 20942
rect 32036 20878 32088 20884
rect 32048 20602 32076 20878
rect 32036 20596 32088 20602
rect 32036 20538 32088 20544
rect 32140 19854 32168 21286
rect 32404 21140 32456 21146
rect 32404 21082 32456 21088
rect 32416 20262 32444 21082
rect 32508 20602 32536 21626
rect 32600 21146 32628 22374
rect 32588 21140 32640 21146
rect 32588 21082 32640 21088
rect 32692 20602 32720 22714
rect 32784 22710 32812 23015
rect 32772 22704 32824 22710
rect 32772 22646 32824 22652
rect 33336 22574 33364 23530
rect 33324 22568 33376 22574
rect 33324 22510 33376 22516
rect 33428 22420 33456 25638
rect 33612 25362 33640 28863
rect 33692 28620 33744 28626
rect 33692 28562 33744 28568
rect 33704 28218 33732 28562
rect 33692 28212 33744 28218
rect 33692 28154 33744 28160
rect 34072 27538 34100 32506
rect 34256 31346 34284 35527
rect 34520 35148 34572 35154
rect 34520 35090 34572 35096
rect 34532 34474 34560 35090
rect 34520 34468 34572 34474
rect 34520 34410 34572 34416
rect 34520 33924 34572 33930
rect 34520 33866 34572 33872
rect 34532 33833 34560 33866
rect 34518 33824 34574 33833
rect 34518 33759 34574 33768
rect 34612 33380 34664 33386
rect 34612 33322 34664 33328
rect 34334 33144 34390 33153
rect 34334 33079 34390 33088
rect 34348 33046 34376 33079
rect 34336 33040 34388 33046
rect 34336 32982 34388 32988
rect 34348 32570 34376 32982
rect 34336 32564 34388 32570
rect 34336 32506 34388 32512
rect 34520 32224 34572 32230
rect 34520 32166 34572 32172
rect 34532 31958 34560 32166
rect 34520 31952 34572 31958
rect 34520 31894 34572 31900
rect 34532 31482 34560 31894
rect 34520 31476 34572 31482
rect 34520 31418 34572 31424
rect 34244 31340 34296 31346
rect 34244 31282 34296 31288
rect 34152 29776 34204 29782
rect 34152 29718 34204 29724
rect 34164 29306 34192 29718
rect 34152 29300 34204 29306
rect 34152 29242 34204 29248
rect 34164 28762 34192 29242
rect 34152 28756 34204 28762
rect 34152 28698 34204 28704
rect 34164 28218 34192 28698
rect 34152 28212 34204 28218
rect 34152 28154 34204 28160
rect 34060 27532 34112 27538
rect 34060 27474 34112 27480
rect 33876 26988 33928 26994
rect 33876 26930 33928 26936
rect 33600 25356 33652 25362
rect 33600 25298 33652 25304
rect 33612 24614 33640 25298
rect 33600 24608 33652 24614
rect 33600 24550 33652 24556
rect 33612 22710 33640 24550
rect 33784 24268 33836 24274
rect 33784 24210 33836 24216
rect 33796 23866 33824 24210
rect 33784 23860 33836 23866
rect 33784 23802 33836 23808
rect 33600 22704 33652 22710
rect 33600 22646 33652 22652
rect 33782 22672 33838 22681
rect 33782 22607 33838 22616
rect 33796 22574 33824 22607
rect 33784 22568 33836 22574
rect 33784 22510 33836 22516
rect 33428 22392 33548 22420
rect 33416 22160 33468 22166
rect 33416 22102 33468 22108
rect 33324 22024 33376 22030
rect 33324 21966 33376 21972
rect 32772 21888 32824 21894
rect 32772 21830 32824 21836
rect 33048 21888 33100 21894
rect 33048 21830 33100 21836
rect 32784 21554 32812 21830
rect 32772 21548 32824 21554
rect 32772 21490 32824 21496
rect 32784 21146 32812 21490
rect 32864 21480 32916 21486
rect 32864 21422 32916 21428
rect 32876 21185 32904 21422
rect 32956 21344 33008 21350
rect 33060 21332 33088 21830
rect 33336 21690 33364 21966
rect 33428 21690 33456 22102
rect 33324 21684 33376 21690
rect 33324 21626 33376 21632
rect 33416 21684 33468 21690
rect 33416 21626 33468 21632
rect 33008 21304 33088 21332
rect 32956 21286 33008 21292
rect 32862 21176 32918 21185
rect 32772 21140 32824 21146
rect 32862 21111 32918 21120
rect 32772 21082 32824 21088
rect 33060 21010 33088 21304
rect 33048 21004 33100 21010
rect 33100 20964 33180 20992
rect 33048 20946 33100 20952
rect 32496 20596 32548 20602
rect 32496 20538 32548 20544
rect 32680 20596 32732 20602
rect 32680 20538 32732 20544
rect 32692 20398 32720 20538
rect 32772 20528 32824 20534
rect 32772 20470 32824 20476
rect 32680 20392 32732 20398
rect 32680 20334 32732 20340
rect 32404 20256 32456 20262
rect 32404 20198 32456 20204
rect 32784 19922 32812 20470
rect 32954 20360 33010 20369
rect 32954 20295 33010 20304
rect 32772 19916 32824 19922
rect 32772 19858 32824 19864
rect 32864 19916 32916 19922
rect 32864 19858 32916 19864
rect 32128 19848 32180 19854
rect 32128 19790 32180 19796
rect 32784 19514 32812 19858
rect 32772 19508 32824 19514
rect 32772 19450 32824 19456
rect 32876 19446 32904 19858
rect 32864 19440 32916 19446
rect 32864 19382 32916 19388
rect 31760 19304 31812 19310
rect 31760 19246 31812 19252
rect 32864 19236 32916 19242
rect 32864 19178 32916 19184
rect 32876 18970 32904 19178
rect 32864 18964 32916 18970
rect 32864 18906 32916 18912
rect 32128 18828 32180 18834
rect 32180 18788 32260 18816
rect 32128 18770 32180 18776
rect 32232 18154 32260 18788
rect 32968 18737 32996 20295
rect 33152 20262 33180 20964
rect 33324 20324 33376 20330
rect 33324 20266 33376 20272
rect 33140 20256 33192 20262
rect 33140 20198 33192 20204
rect 33152 19990 33180 20198
rect 33140 19984 33192 19990
rect 33140 19926 33192 19932
rect 33336 19786 33364 20266
rect 33324 19780 33376 19786
rect 33324 19722 33376 19728
rect 33140 19440 33192 19446
rect 33140 19382 33192 19388
rect 33048 19372 33100 19378
rect 33048 19314 33100 19320
rect 32954 18728 33010 18737
rect 32954 18663 33010 18672
rect 32220 18148 32272 18154
rect 32220 18090 32272 18096
rect 32232 18057 32260 18090
rect 32218 18048 32274 18057
rect 32218 17983 32274 17992
rect 33060 17202 33088 19314
rect 33152 19310 33180 19382
rect 33140 19304 33192 19310
rect 33140 19246 33192 19252
rect 33520 18290 33548 22392
rect 33692 22024 33744 22030
rect 33692 21966 33744 21972
rect 33704 21554 33732 21966
rect 33692 21548 33744 21554
rect 33612 21508 33692 21536
rect 33612 19378 33640 21508
rect 33692 21490 33744 21496
rect 33692 20800 33744 20806
rect 33692 20742 33744 20748
rect 33704 20466 33732 20742
rect 33692 20460 33744 20466
rect 33692 20402 33744 20408
rect 33784 20460 33836 20466
rect 33784 20402 33836 20408
rect 33704 20058 33732 20402
rect 33692 20052 33744 20058
rect 33692 19994 33744 20000
rect 33796 19854 33824 20402
rect 33692 19848 33744 19854
rect 33692 19790 33744 19796
rect 33784 19848 33836 19854
rect 33784 19790 33836 19796
rect 33704 19514 33732 19790
rect 33692 19508 33744 19514
rect 33692 19450 33744 19456
rect 33600 19372 33652 19378
rect 33600 19314 33652 19320
rect 33692 19236 33744 19242
rect 33692 19178 33744 19184
rect 33704 18902 33732 19178
rect 33796 18970 33824 19790
rect 33784 18964 33836 18970
rect 33784 18906 33836 18912
rect 33692 18896 33744 18902
rect 33692 18838 33744 18844
rect 33600 18760 33652 18766
rect 33600 18702 33652 18708
rect 33612 18426 33640 18702
rect 33704 18426 33732 18838
rect 33600 18420 33652 18426
rect 33600 18362 33652 18368
rect 33692 18420 33744 18426
rect 33692 18362 33744 18368
rect 33508 18284 33560 18290
rect 33508 18226 33560 18232
rect 33508 18148 33560 18154
rect 33508 18090 33560 18096
rect 33232 18080 33284 18086
rect 33232 18022 33284 18028
rect 33140 17332 33192 17338
rect 33140 17274 33192 17280
rect 33048 17196 33100 17202
rect 33048 17138 33100 17144
rect 33152 17134 33180 17274
rect 33140 17128 33192 17134
rect 33140 17070 33192 17076
rect 32956 16652 33008 16658
rect 32956 16594 33008 16600
rect 32772 16176 32824 16182
rect 32772 16118 32824 16124
rect 31944 16108 31996 16114
rect 31944 16050 31996 16056
rect 31760 15972 31812 15978
rect 31760 15914 31812 15920
rect 31772 15638 31800 15914
rect 31956 15706 31984 16050
rect 31944 15700 31996 15706
rect 31944 15642 31996 15648
rect 32784 15638 32812 16118
rect 32968 15910 32996 16594
rect 32956 15904 33008 15910
rect 32956 15846 33008 15852
rect 31760 15632 31812 15638
rect 31760 15574 31812 15580
rect 32772 15632 32824 15638
rect 32772 15574 32824 15580
rect 31772 15162 31800 15574
rect 31760 15156 31812 15162
rect 31760 15098 31812 15104
rect 32496 14884 32548 14890
rect 32496 14826 32548 14832
rect 32508 14618 32536 14826
rect 32496 14612 32548 14618
rect 32496 14554 32548 14560
rect 31668 14408 31720 14414
rect 31668 14350 31720 14356
rect 31680 14074 31708 14350
rect 32508 14074 32536 14554
rect 32968 14521 32996 15846
rect 33244 15178 33272 18022
rect 33520 17814 33548 18090
rect 33704 17882 33732 18362
rect 33692 17876 33744 17882
rect 33692 17818 33744 17824
rect 33508 17808 33560 17814
rect 33508 17750 33560 17756
rect 33600 17808 33652 17814
rect 33600 17750 33652 17756
rect 33612 17270 33640 17750
rect 33796 17678 33824 18906
rect 33784 17672 33836 17678
rect 33784 17614 33836 17620
rect 33600 17264 33652 17270
rect 33600 17206 33652 17212
rect 33612 17066 33640 17206
rect 33324 17060 33376 17066
rect 33324 17002 33376 17008
rect 33600 17060 33652 17066
rect 33600 17002 33652 17008
rect 33336 16794 33364 17002
rect 33324 16788 33376 16794
rect 33324 16730 33376 16736
rect 33416 16720 33468 16726
rect 33416 16662 33468 16668
rect 33428 16250 33456 16662
rect 33416 16244 33468 16250
rect 33416 16186 33468 16192
rect 33152 15150 33272 15178
rect 33152 14890 33180 15150
rect 33140 14884 33192 14890
rect 33140 14826 33192 14832
rect 32954 14512 33010 14521
rect 32954 14447 33010 14456
rect 31668 14068 31720 14074
rect 31668 14010 31720 14016
rect 32496 14068 32548 14074
rect 32496 14010 32548 14016
rect 32508 13814 32536 14010
rect 32416 13786 32536 13814
rect 33152 13814 33180 14826
rect 33232 14816 33284 14822
rect 33232 14758 33284 14764
rect 33244 14550 33272 14758
rect 33232 14544 33284 14550
rect 33232 14486 33284 14492
rect 33796 14414 33824 17614
rect 33888 17338 33916 26930
rect 33968 26852 34020 26858
rect 33968 26794 34020 26800
rect 33980 26586 34008 26794
rect 34256 26761 34284 31282
rect 34336 30116 34388 30122
rect 34336 30058 34388 30064
rect 34348 29646 34376 30058
rect 34336 29640 34388 29646
rect 34336 29582 34388 29588
rect 34242 26752 34298 26761
rect 34242 26687 34298 26696
rect 33968 26580 34020 26586
rect 33968 26522 34020 26528
rect 33968 26444 34020 26450
rect 33968 26386 34020 26392
rect 33980 25702 34008 26386
rect 33968 25696 34020 25702
rect 33968 25638 34020 25644
rect 34428 25696 34480 25702
rect 34428 25638 34480 25644
rect 34060 24268 34112 24274
rect 34060 24210 34112 24216
rect 34072 23594 34100 24210
rect 34336 24200 34388 24206
rect 34336 24142 34388 24148
rect 34244 23860 34296 23866
rect 34244 23802 34296 23808
rect 34060 23588 34112 23594
rect 34060 23530 34112 23536
rect 34256 23497 34284 23802
rect 34242 23488 34298 23497
rect 34242 23423 34298 23432
rect 33968 22704 34020 22710
rect 33968 22646 34020 22652
rect 33980 18086 34008 22646
rect 34256 21962 34284 23423
rect 34348 23100 34376 24142
rect 34440 23254 34468 25638
rect 34520 25492 34572 25498
rect 34520 25434 34572 25440
rect 34532 24954 34560 25434
rect 34520 24948 34572 24954
rect 34520 24890 34572 24896
rect 34532 24682 34560 24890
rect 34520 24676 34572 24682
rect 34520 24618 34572 24624
rect 34624 23474 34652 33322
rect 34808 33114 34836 35974
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 35452 35154 35480 35974
rect 35636 35698 35664 36314
rect 35808 36168 35860 36174
rect 35808 36110 35860 36116
rect 35820 35698 35848 36110
rect 35624 35692 35676 35698
rect 35624 35634 35676 35640
rect 35808 35692 35860 35698
rect 35808 35634 35860 35640
rect 35820 35222 35848 35634
rect 35808 35216 35860 35222
rect 35808 35158 35860 35164
rect 35440 35148 35492 35154
rect 35440 35090 35492 35096
rect 35992 35148 36044 35154
rect 35992 35090 36044 35096
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 35452 34542 35480 35090
rect 35532 34604 35584 34610
rect 35532 34546 35584 34552
rect 35440 34536 35492 34542
rect 35440 34478 35492 34484
rect 35452 33930 35480 34478
rect 35544 33998 35572 34546
rect 35900 34468 35952 34474
rect 35900 34410 35952 34416
rect 35624 34060 35676 34066
rect 35624 34002 35676 34008
rect 35532 33992 35584 33998
rect 35532 33934 35584 33940
rect 35440 33924 35492 33930
rect 35440 33866 35492 33872
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 35544 33658 35572 33934
rect 35532 33652 35584 33658
rect 35532 33594 35584 33600
rect 34796 33108 34848 33114
rect 34796 33050 34848 33056
rect 34808 32434 34836 33050
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 34796 32428 34848 32434
rect 34796 32370 34848 32376
rect 35440 32428 35492 32434
rect 35440 32370 35492 32376
rect 35256 31816 35308 31822
rect 35256 31758 35308 31764
rect 34796 31680 34848 31686
rect 34796 31622 34848 31628
rect 34808 31210 34836 31622
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 35164 31340 35216 31346
rect 35164 31282 35216 31288
rect 35176 31210 35204 31282
rect 34704 31204 34756 31210
rect 34704 31146 34756 31152
rect 34796 31204 34848 31210
rect 34796 31146 34848 31152
rect 35164 31204 35216 31210
rect 35164 31146 35216 31152
rect 34716 30870 34744 31146
rect 34704 30864 34756 30870
rect 34704 30806 34756 30812
rect 34808 27606 34836 31146
rect 35268 30870 35296 31758
rect 35348 31748 35400 31754
rect 35348 31690 35400 31696
rect 35256 30864 35308 30870
rect 35254 30832 35256 30841
rect 35308 30832 35310 30841
rect 35254 30767 35310 30776
rect 35256 30592 35308 30598
rect 35256 30534 35308 30540
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 35268 30258 35296 30534
rect 35360 30258 35388 31690
rect 35452 31346 35480 32370
rect 35636 31385 35664 34002
rect 35912 31482 35940 34410
rect 36004 34406 36032 35090
rect 35992 34400 36044 34406
rect 35992 34342 36044 34348
rect 36004 32910 36032 34342
rect 36096 33522 36124 37760
rect 36464 37738 36492 38150
rect 36556 37874 36584 38150
rect 36544 37868 36596 37874
rect 36544 37810 36596 37816
rect 36452 37732 36504 37738
rect 36452 37674 36504 37680
rect 36464 37466 36492 37674
rect 36452 37460 36504 37466
rect 36452 37402 36504 37408
rect 36358 37224 36414 37233
rect 36358 37159 36414 37168
rect 36268 36712 36320 36718
rect 36268 36654 36320 36660
rect 36176 36372 36228 36378
rect 36176 36314 36228 36320
rect 36188 35562 36216 36314
rect 36176 35556 36228 35562
rect 36176 35498 36228 35504
rect 36188 35222 36216 35498
rect 36176 35216 36228 35222
rect 36176 35158 36228 35164
rect 36084 33516 36136 33522
rect 36084 33458 36136 33464
rect 36280 32978 36308 36654
rect 36268 32972 36320 32978
rect 36268 32914 36320 32920
rect 35992 32904 36044 32910
rect 35992 32846 36044 32852
rect 36084 32768 36136 32774
rect 36084 32710 36136 32716
rect 36096 31958 36124 32710
rect 36280 32230 36308 32914
rect 36268 32224 36320 32230
rect 36268 32166 36320 32172
rect 36084 31952 36136 31958
rect 36084 31894 36136 31900
rect 36176 31952 36228 31958
rect 36176 31894 36228 31900
rect 35900 31476 35952 31482
rect 35900 31418 35952 31424
rect 35622 31376 35678 31385
rect 35440 31340 35492 31346
rect 35622 31311 35678 31320
rect 35440 31282 35492 31288
rect 35256 30252 35308 30258
rect 35256 30194 35308 30200
rect 35348 30252 35400 30258
rect 35348 30194 35400 30200
rect 35360 30138 35388 30194
rect 35268 30110 35388 30138
rect 34980 30048 35032 30054
rect 34980 29990 35032 29996
rect 34992 29850 35020 29990
rect 34980 29844 35032 29850
rect 34980 29786 35032 29792
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 35072 29028 35124 29034
rect 35072 28970 35124 28976
rect 35084 28762 35112 28970
rect 35072 28756 35124 28762
rect 35072 28698 35124 28704
rect 35268 28694 35296 30110
rect 35452 29578 35480 31282
rect 35532 31136 35584 31142
rect 35532 31078 35584 31084
rect 35544 29714 35572 31078
rect 35532 29708 35584 29714
rect 35532 29650 35584 29656
rect 35440 29572 35492 29578
rect 35440 29514 35492 29520
rect 35348 29504 35400 29510
rect 35348 29446 35400 29452
rect 35360 29170 35388 29446
rect 35452 29170 35480 29514
rect 35348 29164 35400 29170
rect 35348 29106 35400 29112
rect 35440 29164 35492 29170
rect 35440 29106 35492 29112
rect 35256 28688 35308 28694
rect 35256 28630 35308 28636
rect 35256 28552 35308 28558
rect 35256 28494 35308 28500
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 35268 27674 35296 28494
rect 35256 27668 35308 27674
rect 35256 27610 35308 27616
rect 34796 27600 34848 27606
rect 34796 27542 34848 27548
rect 34704 27532 34756 27538
rect 34704 27474 34756 27480
rect 34716 27130 34744 27474
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 34704 27124 34756 27130
rect 34704 27066 34756 27072
rect 34888 26784 34940 26790
rect 34888 26726 34940 26732
rect 34796 26580 34848 26586
rect 34796 26522 34848 26528
rect 34704 26240 34756 26246
rect 34704 26182 34756 26188
rect 34716 25430 34744 26182
rect 34808 25906 34836 26522
rect 34900 26382 34928 26726
rect 35360 26586 35388 29106
rect 35440 29028 35492 29034
rect 35440 28970 35492 28976
rect 35348 26580 35400 26586
rect 35348 26522 35400 26528
rect 34888 26376 34940 26382
rect 34888 26318 34940 26324
rect 35256 26308 35308 26314
rect 35256 26250 35308 26256
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 34796 25900 34848 25906
rect 34796 25842 34848 25848
rect 34704 25424 34756 25430
rect 34756 25384 34836 25412
rect 34704 25366 34756 25372
rect 34704 25152 34756 25158
rect 34704 25094 34756 25100
rect 34716 24818 34744 25094
rect 34808 24954 34836 25384
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 34796 24948 34848 24954
rect 34796 24890 34848 24896
rect 35268 24818 35296 26250
rect 35348 25900 35400 25906
rect 35348 25842 35400 25848
rect 35360 24886 35388 25842
rect 35452 25226 35480 28970
rect 35544 28966 35572 29650
rect 35532 28960 35584 28966
rect 35532 28902 35584 28908
rect 35636 28626 35664 31311
rect 35992 30864 36044 30870
rect 36096 30852 36124 31894
rect 36188 31414 36216 31894
rect 36176 31408 36228 31414
rect 36176 31350 36228 31356
rect 36280 31249 36308 32166
rect 36266 31240 36322 31249
rect 36266 31175 36322 31184
rect 36044 30824 36124 30852
rect 35992 30806 36044 30812
rect 35900 29504 35952 29510
rect 35900 29446 35952 29452
rect 35992 29504 36044 29510
rect 35992 29446 36044 29452
rect 35624 28620 35676 28626
rect 35624 28562 35676 28568
rect 35912 28218 35940 29446
rect 36004 28558 36032 29446
rect 35992 28552 36044 28558
rect 35992 28494 36044 28500
rect 35900 28212 35952 28218
rect 35900 28154 35952 28160
rect 36176 27532 36228 27538
rect 36280 27520 36308 31175
rect 36372 30802 36400 37159
rect 36820 37120 36872 37126
rect 36820 37062 36872 37068
rect 36832 36650 36860 37062
rect 37016 36854 37044 38762
rect 37188 37732 37240 37738
rect 37188 37674 37240 37680
rect 37004 36848 37056 36854
rect 37004 36790 37056 36796
rect 36912 36780 36964 36786
rect 36912 36722 36964 36728
rect 36820 36644 36872 36650
rect 36820 36586 36872 36592
rect 36832 35834 36860 36586
rect 36924 36106 36952 36722
rect 36912 36100 36964 36106
rect 36912 36042 36964 36048
rect 36820 35828 36872 35834
rect 36820 35770 36872 35776
rect 36636 34672 36688 34678
rect 36636 34614 36688 34620
rect 36452 34604 36504 34610
rect 36452 34546 36504 34552
rect 36464 33454 36492 34546
rect 36544 34128 36596 34134
rect 36544 34070 36596 34076
rect 36452 33448 36504 33454
rect 36452 33390 36504 33396
rect 36556 33318 36584 34070
rect 36544 33312 36596 33318
rect 36544 33254 36596 33260
rect 36556 33114 36584 33254
rect 36544 33108 36596 33114
rect 36544 33050 36596 33056
rect 36544 32972 36596 32978
rect 36544 32914 36596 32920
rect 36556 32230 36584 32914
rect 36544 32224 36596 32230
rect 36544 32166 36596 32172
rect 36360 30796 36412 30802
rect 36360 30738 36412 30744
rect 36372 30394 36400 30738
rect 36360 30388 36412 30394
rect 36360 30330 36412 30336
rect 36228 27492 36308 27520
rect 36176 27474 36228 27480
rect 35716 27464 35768 27470
rect 35714 27432 35716 27441
rect 35768 27432 35770 27441
rect 35714 27367 35770 27376
rect 35728 27130 35756 27367
rect 35716 27124 35768 27130
rect 35716 27066 35768 27072
rect 36188 26790 36216 27474
rect 36176 26784 36228 26790
rect 36176 26726 36228 26732
rect 35808 26512 35860 26518
rect 35808 26454 35860 26460
rect 35624 26308 35676 26314
rect 35624 26250 35676 26256
rect 35636 25838 35664 26250
rect 35624 25832 35676 25838
rect 35624 25774 35676 25780
rect 35440 25220 35492 25226
rect 35440 25162 35492 25168
rect 35348 24880 35400 24886
rect 35348 24822 35400 24828
rect 34704 24812 34756 24818
rect 34704 24754 34756 24760
rect 35256 24812 35308 24818
rect 35256 24754 35308 24760
rect 35072 24676 35124 24682
rect 35072 24618 35124 24624
rect 35084 24410 35112 24618
rect 35072 24404 35124 24410
rect 35072 24346 35124 24352
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 34624 23446 34836 23474
rect 34428 23248 34480 23254
rect 34428 23190 34480 23196
rect 34704 23248 34756 23254
rect 34704 23190 34756 23196
rect 34520 23112 34572 23118
rect 34348 23072 34520 23100
rect 34520 23054 34572 23060
rect 34532 22234 34560 23054
rect 34716 22438 34744 23190
rect 34704 22432 34756 22438
rect 34704 22374 34756 22380
rect 34520 22228 34572 22234
rect 34520 22170 34572 22176
rect 34244 21956 34296 21962
rect 34244 21898 34296 21904
rect 34428 21956 34480 21962
rect 34428 21898 34480 21904
rect 34060 21684 34112 21690
rect 34060 21626 34112 21632
rect 34072 21078 34100 21626
rect 34060 21072 34112 21078
rect 34060 21014 34112 21020
rect 34244 21072 34296 21078
rect 34244 21014 34296 21020
rect 34072 20602 34100 21014
rect 34060 20596 34112 20602
rect 34060 20538 34112 20544
rect 34072 19990 34100 20538
rect 34060 19984 34112 19990
rect 34060 19926 34112 19932
rect 34072 19446 34100 19926
rect 34060 19440 34112 19446
rect 34060 19382 34112 19388
rect 34256 18902 34284 21014
rect 34244 18896 34296 18902
rect 34244 18838 34296 18844
rect 33968 18080 34020 18086
rect 33968 18022 34020 18028
rect 34256 17610 34284 18838
rect 34336 17808 34388 17814
rect 34336 17750 34388 17756
rect 34244 17604 34296 17610
rect 34164 17564 34244 17592
rect 33876 17332 33928 17338
rect 33928 17292 34100 17320
rect 33876 17274 33928 17280
rect 33968 17196 34020 17202
rect 33968 17138 34020 17144
rect 33876 16584 33928 16590
rect 33876 16526 33928 16532
rect 33888 16114 33916 16526
rect 33876 16108 33928 16114
rect 33876 16050 33928 16056
rect 33980 15638 34008 17138
rect 34072 16522 34100 17292
rect 34164 16794 34192 17564
rect 34244 17546 34296 17552
rect 34348 17338 34376 17750
rect 34336 17332 34388 17338
rect 34336 17274 34388 17280
rect 34440 17134 34468 21898
rect 34612 20936 34664 20942
rect 34612 20878 34664 20884
rect 34624 20602 34652 20878
rect 34612 20596 34664 20602
rect 34612 20538 34664 20544
rect 34716 20466 34744 22374
rect 34704 20460 34756 20466
rect 34704 20402 34756 20408
rect 34704 19168 34756 19174
rect 34704 19110 34756 19116
rect 34612 18896 34664 18902
rect 34612 18838 34664 18844
rect 34518 18728 34574 18737
rect 34518 18663 34574 18672
rect 34428 17128 34480 17134
rect 34428 17070 34480 17076
rect 34532 16794 34560 18663
rect 34624 18086 34652 18838
rect 34716 18766 34744 19110
rect 34704 18760 34756 18766
rect 34704 18702 34756 18708
rect 34704 18216 34756 18222
rect 34704 18158 34756 18164
rect 34612 18080 34664 18086
rect 34612 18022 34664 18028
rect 34152 16788 34204 16794
rect 34152 16730 34204 16736
rect 34520 16788 34572 16794
rect 34520 16730 34572 16736
rect 34244 16720 34296 16726
rect 34244 16662 34296 16668
rect 34060 16516 34112 16522
rect 34060 16458 34112 16464
rect 33968 15632 34020 15638
rect 33968 15574 34020 15580
rect 33876 15496 33928 15502
rect 33876 15438 33928 15444
rect 33888 15162 33916 15438
rect 34072 15162 34100 16458
rect 34256 15910 34284 16662
rect 34624 16250 34652 18022
rect 34716 17678 34744 18158
rect 34704 17672 34756 17678
rect 34704 17614 34756 17620
rect 34612 16244 34664 16250
rect 34612 16186 34664 16192
rect 34702 16144 34758 16153
rect 34520 16108 34572 16114
rect 34702 16079 34758 16088
rect 34520 16050 34572 16056
rect 34244 15904 34296 15910
rect 34244 15846 34296 15852
rect 34256 15706 34284 15846
rect 34244 15700 34296 15706
rect 34244 15642 34296 15648
rect 34336 15632 34388 15638
rect 34336 15574 34388 15580
rect 33876 15156 33928 15162
rect 33876 15098 33928 15104
rect 34060 15156 34112 15162
rect 34060 15098 34112 15104
rect 34244 14816 34296 14822
rect 34348 14804 34376 15574
rect 34532 15502 34560 16050
rect 34716 16046 34744 16079
rect 34704 16040 34756 16046
rect 34704 15982 34756 15988
rect 34520 15496 34572 15502
rect 34520 15438 34572 15444
rect 34296 14776 34376 14804
rect 34244 14758 34296 14764
rect 34256 14618 34284 14758
rect 34244 14612 34296 14618
rect 34244 14554 34296 14560
rect 34152 14544 34204 14550
rect 34152 14486 34204 14492
rect 33600 14408 33652 14414
rect 33600 14350 33652 14356
rect 33784 14408 33836 14414
rect 33784 14350 33836 14356
rect 33612 14074 33640 14350
rect 34164 14074 34192 14486
rect 34532 14346 34560 15438
rect 34520 14340 34572 14346
rect 34520 14282 34572 14288
rect 34532 14074 34560 14282
rect 33600 14068 33652 14074
rect 33600 14010 33652 14016
rect 34152 14068 34204 14074
rect 34152 14010 34204 14016
rect 34520 14068 34572 14074
rect 34520 14010 34572 14016
rect 34532 13870 34560 14010
rect 34520 13864 34572 13870
rect 33152 13786 33272 13814
rect 34520 13806 34572 13812
rect 32416 12714 32444 13786
rect 32680 13728 32732 13734
rect 32680 13670 32732 13676
rect 32588 13184 32640 13190
rect 32588 13126 32640 13132
rect 32600 12986 32628 13126
rect 32588 12980 32640 12986
rect 32588 12922 32640 12928
rect 32600 12782 32628 12922
rect 32588 12776 32640 12782
rect 32588 12718 32640 12724
rect 32404 12708 32456 12714
rect 32404 12650 32456 12656
rect 31944 12640 31996 12646
rect 31944 12582 31996 12588
rect 31956 11898 31984 12582
rect 32588 12368 32640 12374
rect 32588 12310 32640 12316
rect 32404 12300 32456 12306
rect 32404 12242 32456 12248
rect 32416 11898 32444 12242
rect 31944 11892 31996 11898
rect 31944 11834 31996 11840
rect 32404 11892 32456 11898
rect 32404 11834 32456 11840
rect 32600 11529 32628 12310
rect 32692 11762 32720 13670
rect 33140 13388 33192 13394
rect 33140 13330 33192 13336
rect 33152 12918 33180 13330
rect 33140 12912 33192 12918
rect 33140 12854 33192 12860
rect 32772 12708 32824 12714
rect 32772 12650 32824 12656
rect 32680 11756 32732 11762
rect 32680 11698 32732 11704
rect 32586 11520 32642 11529
rect 32586 11455 32642 11464
rect 31852 11212 31904 11218
rect 31852 11154 31904 11160
rect 31864 10470 31892 11154
rect 32496 11008 32548 11014
rect 32496 10950 32548 10956
rect 31852 10464 31904 10470
rect 31852 10406 31904 10412
rect 31864 10266 31892 10406
rect 31852 10260 31904 10266
rect 31852 10202 31904 10208
rect 32508 10198 32536 10950
rect 32600 10538 32628 11455
rect 32692 11354 32720 11698
rect 32784 11626 32812 12650
rect 32772 11620 32824 11626
rect 32772 11562 32824 11568
rect 32680 11348 32732 11354
rect 32680 11290 32732 11296
rect 32588 10532 32640 10538
rect 32588 10474 32640 10480
rect 32496 10192 32548 10198
rect 32496 10134 32548 10140
rect 32508 9654 32536 10134
rect 32496 9648 32548 9654
rect 32496 9590 32548 9596
rect 32128 9444 32180 9450
rect 32128 9386 32180 9392
rect 31760 8968 31812 8974
rect 31760 8910 31812 8916
rect 31772 8634 31800 8910
rect 31760 8628 31812 8634
rect 31760 8570 31812 8576
rect 31668 8356 31720 8362
rect 31668 8298 31720 8304
rect 31680 7478 31708 8298
rect 31772 8090 31800 8570
rect 32140 8498 32168 9386
rect 32600 9110 32628 10474
rect 32784 10198 32812 11562
rect 33140 10532 33192 10538
rect 33140 10474 33192 10480
rect 33152 10198 33180 10474
rect 32772 10192 32824 10198
rect 32772 10134 32824 10140
rect 33140 10192 33192 10198
rect 33140 10134 33192 10140
rect 32784 9450 32812 10134
rect 32772 9444 32824 9450
rect 32772 9386 32824 9392
rect 32956 9444 33008 9450
rect 32956 9386 33008 9392
rect 32968 9110 32996 9386
rect 32588 9104 32640 9110
rect 32588 9046 32640 9052
rect 32956 9104 33008 9110
rect 32956 9046 33008 9052
rect 32600 8634 32628 9046
rect 32588 8628 32640 8634
rect 32588 8570 32640 8576
rect 32128 8492 32180 8498
rect 32128 8434 32180 8440
rect 33140 8492 33192 8498
rect 33140 8434 33192 8440
rect 33152 8129 33180 8434
rect 33138 8120 33194 8129
rect 31760 8084 31812 8090
rect 31760 8026 31812 8032
rect 32220 8084 32272 8090
rect 33138 8055 33194 8064
rect 32220 8026 32272 8032
rect 32128 7948 32180 7954
rect 32128 7890 32180 7896
rect 32140 7546 32168 7890
rect 32128 7540 32180 7546
rect 32128 7482 32180 7488
rect 31668 7472 31720 7478
rect 31668 7414 31720 7420
rect 31680 7274 31708 7414
rect 31852 7336 31904 7342
rect 31852 7278 31904 7284
rect 31668 7268 31720 7274
rect 31668 7210 31720 7216
rect 31680 6458 31708 7210
rect 31864 6662 31892 7278
rect 32232 7002 32260 8026
rect 33152 8022 33180 8055
rect 33140 8016 33192 8022
rect 33140 7958 33192 7964
rect 33140 7880 33192 7886
rect 33140 7822 33192 7828
rect 33152 7546 33180 7822
rect 33140 7540 33192 7546
rect 33140 7482 33192 7488
rect 32496 7268 32548 7274
rect 32496 7210 32548 7216
rect 32508 7002 32536 7210
rect 32220 6996 32272 7002
rect 32220 6938 32272 6944
rect 32496 6996 32548 7002
rect 32496 6938 32548 6944
rect 31944 6860 31996 6866
rect 31944 6802 31996 6808
rect 31852 6656 31904 6662
rect 31852 6598 31904 6604
rect 31668 6452 31720 6458
rect 31668 6394 31720 6400
rect 31852 6112 31904 6118
rect 31852 6054 31904 6060
rect 31864 4690 31892 6054
rect 31956 5914 31984 6802
rect 32772 6656 32824 6662
rect 32772 6598 32824 6604
rect 31944 5908 31996 5914
rect 31944 5850 31996 5856
rect 32036 5908 32088 5914
rect 32036 5850 32088 5856
rect 31852 4684 31904 4690
rect 31852 4626 31904 4632
rect 32048 4622 32076 5850
rect 32128 5772 32180 5778
rect 32128 5714 32180 5720
rect 32140 5370 32168 5714
rect 32128 5364 32180 5370
rect 32128 5306 32180 5312
rect 32784 5030 32812 6598
rect 33140 6112 33192 6118
rect 33140 6054 33192 6060
rect 33152 5846 33180 6054
rect 33140 5840 33192 5846
rect 33140 5782 33192 5788
rect 32772 5024 32824 5030
rect 32772 4966 32824 4972
rect 33152 4758 33180 5782
rect 32220 4752 32272 4758
rect 32220 4694 32272 4700
rect 33140 4752 33192 4758
rect 33140 4694 33192 4700
rect 32036 4616 32088 4622
rect 32036 4558 32088 4564
rect 32232 4214 32260 4694
rect 33048 4548 33100 4554
rect 33048 4490 33100 4496
rect 32496 4480 32548 4486
rect 32496 4422 32548 4428
rect 32220 4208 32272 4214
rect 32220 4150 32272 4156
rect 31944 3936 31996 3942
rect 31944 3878 31996 3884
rect 31760 2984 31812 2990
rect 31760 2926 31812 2932
rect 31772 2650 31800 2926
rect 31956 2922 31984 3878
rect 32036 3732 32088 3738
rect 32036 3674 32088 3680
rect 32048 3194 32076 3674
rect 32232 3670 32260 4150
rect 32508 4146 32536 4422
rect 33060 4214 33088 4490
rect 33048 4208 33100 4214
rect 33048 4150 33100 4156
rect 32496 4140 32548 4146
rect 32496 4082 32548 4088
rect 32312 4004 32364 4010
rect 32312 3946 32364 3952
rect 32220 3664 32272 3670
rect 32220 3606 32272 3612
rect 32324 3534 32352 3946
rect 32508 3738 32536 4082
rect 32496 3732 32548 3738
rect 32496 3674 32548 3680
rect 33060 3670 33088 4150
rect 33048 3664 33100 3670
rect 33048 3606 33100 3612
rect 32220 3528 32272 3534
rect 32220 3470 32272 3476
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 32232 3194 32260 3470
rect 32036 3188 32088 3194
rect 32036 3130 32088 3136
rect 32220 3188 32272 3194
rect 32220 3130 32272 3136
rect 31944 2916 31996 2922
rect 31944 2858 31996 2864
rect 31760 2644 31812 2650
rect 31760 2586 31812 2592
rect 31576 2508 31628 2514
rect 31576 2450 31628 2456
rect 30286 82 30342 480
rect 33244 134 33272 13786
rect 33600 13728 33652 13734
rect 33600 13670 33652 13676
rect 33324 13184 33376 13190
rect 33324 13126 33376 13132
rect 33336 12306 33364 13126
rect 33324 12300 33376 12306
rect 33324 12242 33376 12248
rect 33508 10668 33560 10674
rect 33508 10610 33560 10616
rect 33520 10470 33548 10610
rect 33508 10464 33560 10470
rect 33508 10406 33560 10412
rect 33520 9722 33548 10406
rect 33508 9716 33560 9722
rect 33508 9658 33560 9664
rect 33612 7546 33640 13670
rect 34704 13388 34756 13394
rect 34704 13330 34756 13336
rect 34716 12646 34744 13330
rect 34704 12640 34756 12646
rect 34704 12582 34756 12588
rect 33784 12368 33836 12374
rect 34716 12345 34744 12582
rect 33784 12310 33836 12316
rect 34702 12336 34758 12345
rect 33796 11830 33824 12310
rect 34808 12306 34836 23446
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 35268 22642 35296 24754
rect 35636 24342 35664 25774
rect 35820 25702 35848 26454
rect 36084 26376 36136 26382
rect 36084 26318 36136 26324
rect 36096 26042 36124 26318
rect 36084 26036 36136 26042
rect 36084 25978 36136 25984
rect 35808 25696 35860 25702
rect 35808 25638 35860 25644
rect 35820 25430 35848 25638
rect 35808 25424 35860 25430
rect 35808 25366 35860 25372
rect 35808 25288 35860 25294
rect 35808 25230 35860 25236
rect 35348 24336 35400 24342
rect 35348 24278 35400 24284
rect 35624 24336 35676 24342
rect 35624 24278 35676 24284
rect 35360 23594 35388 24278
rect 35820 23798 35848 25230
rect 35992 25220 36044 25226
rect 35992 25162 36044 25168
rect 35808 23792 35860 23798
rect 35808 23734 35860 23740
rect 35348 23588 35400 23594
rect 35348 23530 35400 23536
rect 35360 22982 35388 23530
rect 35348 22976 35400 22982
rect 35348 22918 35400 22924
rect 35808 22976 35860 22982
rect 35808 22918 35860 22924
rect 35256 22636 35308 22642
rect 35256 22578 35308 22584
rect 35360 22506 35388 22918
rect 35438 22672 35494 22681
rect 35438 22607 35494 22616
rect 34888 22500 34940 22506
rect 34888 22442 34940 22448
rect 35348 22500 35400 22506
rect 35348 22442 35400 22448
rect 34900 22234 34928 22442
rect 34888 22228 34940 22234
rect 34888 22170 34940 22176
rect 35360 22166 35388 22442
rect 35348 22160 35400 22166
rect 35348 22102 35400 22108
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 34980 21548 35032 21554
rect 34980 21490 35032 21496
rect 35256 21548 35308 21554
rect 35256 21490 35308 21496
rect 34992 21146 35020 21490
rect 34980 21140 35032 21146
rect 34980 21082 35032 21088
rect 35268 21078 35296 21490
rect 35256 21072 35308 21078
rect 35256 21014 35308 21020
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 35452 20602 35480 22607
rect 35716 22432 35768 22438
rect 35716 22374 35768 22380
rect 35728 21010 35756 22374
rect 35820 22234 35848 22918
rect 35808 22228 35860 22234
rect 35808 22170 35860 22176
rect 35820 21146 35848 22170
rect 35900 22160 35952 22166
rect 35900 22102 35952 22108
rect 35912 21690 35940 22102
rect 35900 21684 35952 21690
rect 35900 21626 35952 21632
rect 35808 21140 35860 21146
rect 35808 21082 35860 21088
rect 35716 21004 35768 21010
rect 35716 20946 35768 20952
rect 35440 20596 35492 20602
rect 35440 20538 35492 20544
rect 35452 20398 35480 20538
rect 35440 20392 35492 20398
rect 35440 20334 35492 20340
rect 35728 19786 35756 20946
rect 36004 19990 36032 25162
rect 36188 22438 36216 26726
rect 36372 24750 36400 30330
rect 36648 29850 36676 34614
rect 36924 34610 36952 36042
rect 37016 36038 37044 36790
rect 37004 36032 37056 36038
rect 37004 35974 37056 35980
rect 37200 35018 37228 37674
rect 37476 36922 37504 39918
rect 37740 39908 37792 39914
rect 37740 39850 37792 39856
rect 37752 38418 37780 39850
rect 37832 39024 37884 39030
rect 37832 38966 37884 38972
rect 37740 38412 37792 38418
rect 37740 38354 37792 38360
rect 37752 38010 37780 38354
rect 37740 38004 37792 38010
rect 37740 37946 37792 37952
rect 37464 36916 37516 36922
rect 37464 36858 37516 36864
rect 37280 36780 37332 36786
rect 37280 36722 37332 36728
rect 37292 35766 37320 36722
rect 37740 36372 37792 36378
rect 37740 36314 37792 36320
rect 37752 35834 37780 36314
rect 37844 36310 37872 38966
rect 38108 38548 38160 38554
rect 38108 38490 38160 38496
rect 38120 37942 38148 38490
rect 38108 37936 38160 37942
rect 38108 37878 38160 37884
rect 38014 37224 38070 37233
rect 38014 37159 38070 37168
rect 38028 36718 38056 37159
rect 38016 36712 38068 36718
rect 38016 36654 38068 36660
rect 38028 36582 38056 36654
rect 38016 36576 38068 36582
rect 38016 36518 38068 36524
rect 37832 36304 37884 36310
rect 38016 36304 38068 36310
rect 37884 36264 38016 36292
rect 37832 36246 37884 36252
rect 38016 36246 38068 36252
rect 37740 35828 37792 35834
rect 37740 35770 37792 35776
rect 37280 35760 37332 35766
rect 37280 35702 37332 35708
rect 37844 35290 37872 36246
rect 37832 35284 37884 35290
rect 37832 35226 37884 35232
rect 37924 35216 37976 35222
rect 37924 35158 37976 35164
rect 37188 35012 37240 35018
rect 37188 34954 37240 34960
rect 36912 34604 36964 34610
rect 36912 34546 36964 34552
rect 36728 34468 36780 34474
rect 36728 34410 36780 34416
rect 36740 34202 36768 34410
rect 37200 34406 37228 34954
rect 37936 34610 37964 35158
rect 38108 35080 38160 35086
rect 38108 35022 38160 35028
rect 38120 34746 38148 35022
rect 38108 34740 38160 34746
rect 38108 34682 38160 34688
rect 37924 34604 37976 34610
rect 37924 34546 37976 34552
rect 37188 34400 37240 34406
rect 37188 34342 37240 34348
rect 36728 34196 36780 34202
rect 36728 34138 36780 34144
rect 37936 34134 37964 34546
rect 38212 34134 38240 40695
rect 38292 40588 38344 40594
rect 38292 40530 38344 40536
rect 38304 40118 38332 40530
rect 38752 40520 38804 40526
rect 38752 40462 38804 40468
rect 38568 40384 38620 40390
rect 38568 40326 38620 40332
rect 38292 40112 38344 40118
rect 38292 40054 38344 40060
rect 38580 39574 38608 40326
rect 38764 39914 38792 40462
rect 38844 40384 38896 40390
rect 38844 40326 38896 40332
rect 38856 39914 38884 40326
rect 39672 40180 39724 40186
rect 39672 40122 39724 40128
rect 39212 40112 39264 40118
rect 39212 40054 39264 40060
rect 38752 39908 38804 39914
rect 38752 39850 38804 39856
rect 38844 39908 38896 39914
rect 38844 39850 38896 39856
rect 38568 39568 38620 39574
rect 38568 39510 38620 39516
rect 38580 39098 38608 39510
rect 38568 39092 38620 39098
rect 38568 39034 38620 39040
rect 38568 38752 38620 38758
rect 38568 38694 38620 38700
rect 38476 36100 38528 36106
rect 38476 36042 38528 36048
rect 38384 35828 38436 35834
rect 38384 35770 38436 35776
rect 37924 34128 37976 34134
rect 37924 34070 37976 34076
rect 38200 34128 38252 34134
rect 38200 34070 38252 34076
rect 37924 33856 37976 33862
rect 37924 33798 37976 33804
rect 37464 33584 37516 33590
rect 37464 33526 37516 33532
rect 36728 32904 36780 32910
rect 36728 32846 36780 32852
rect 37188 32904 37240 32910
rect 37188 32846 37240 32852
rect 36636 29844 36688 29850
rect 36636 29786 36688 29792
rect 36452 29708 36504 29714
rect 36452 29650 36504 29656
rect 36464 29034 36492 29650
rect 36648 29102 36676 29786
rect 36740 29306 36768 32846
rect 37200 32570 37228 32846
rect 37188 32564 37240 32570
rect 37188 32506 37240 32512
rect 36820 32224 36872 32230
rect 36820 32166 36872 32172
rect 36832 31260 36860 32166
rect 37372 31340 37424 31346
rect 37372 31282 37424 31288
rect 36912 31272 36964 31278
rect 36832 31232 36912 31260
rect 36832 30977 36860 31232
rect 36912 31214 36964 31220
rect 36818 30968 36874 30977
rect 36818 30903 36874 30912
rect 36832 30870 36860 30903
rect 36820 30864 36872 30870
rect 36820 30806 36872 30812
rect 36728 29300 36780 29306
rect 36728 29242 36780 29248
rect 36832 29102 36860 30806
rect 37384 30258 37412 31282
rect 37476 30734 37504 33526
rect 37936 33522 37964 33798
rect 38212 33658 38240 34070
rect 38200 33652 38252 33658
rect 38200 33594 38252 33600
rect 37924 33516 37976 33522
rect 37924 33458 37976 33464
rect 38292 33516 38344 33522
rect 38292 33458 38344 33464
rect 37648 33448 37700 33454
rect 37648 33390 37700 33396
rect 37556 32768 37608 32774
rect 37556 32710 37608 32716
rect 37464 30728 37516 30734
rect 37464 30670 37516 30676
rect 37372 30252 37424 30258
rect 37372 30194 37424 30200
rect 37384 29850 37412 30194
rect 37372 29844 37424 29850
rect 37372 29786 37424 29792
rect 36636 29096 36688 29102
rect 36636 29038 36688 29044
rect 36820 29096 36872 29102
rect 36820 29038 36872 29044
rect 36452 29028 36504 29034
rect 36452 28970 36504 28976
rect 36648 27402 36676 29038
rect 36832 28762 36860 29038
rect 37568 28937 37596 32710
rect 37554 28928 37610 28937
rect 37554 28863 37610 28872
rect 36820 28756 36872 28762
rect 36820 28698 36872 28704
rect 36820 28620 36872 28626
rect 36820 28562 36872 28568
rect 37188 28620 37240 28626
rect 37188 28562 37240 28568
rect 36832 27878 36860 28562
rect 37200 28218 37228 28562
rect 37660 28558 37688 33390
rect 38108 33312 38160 33318
rect 38108 33254 38160 33260
rect 37832 33108 37884 33114
rect 37832 33050 37884 33056
rect 37844 32570 37872 33050
rect 38120 32842 38148 33254
rect 38108 32836 38160 32842
rect 38108 32778 38160 32784
rect 37832 32564 37884 32570
rect 37832 32506 37884 32512
rect 37740 32224 37792 32230
rect 37740 32166 37792 32172
rect 37752 31958 37780 32166
rect 37740 31952 37792 31958
rect 37740 31894 37792 31900
rect 37752 30938 37780 31894
rect 37740 30932 37792 30938
rect 37740 30874 37792 30880
rect 37844 30394 37872 32506
rect 38016 32224 38068 32230
rect 38016 32166 38068 32172
rect 37832 30388 37884 30394
rect 37832 30330 37884 30336
rect 37844 30122 37872 30330
rect 37832 30116 37884 30122
rect 37832 30058 37884 30064
rect 37844 29782 37872 30058
rect 37832 29776 37884 29782
rect 37832 29718 37884 29724
rect 37740 29640 37792 29646
rect 37740 29582 37792 29588
rect 37752 29170 37780 29582
rect 37844 29170 37872 29718
rect 37740 29164 37792 29170
rect 37740 29106 37792 29112
rect 37832 29164 37884 29170
rect 37884 29124 37964 29152
rect 37832 29106 37884 29112
rect 37752 28762 37780 29106
rect 37740 28756 37792 28762
rect 37740 28698 37792 28704
rect 37648 28552 37700 28558
rect 37648 28494 37700 28500
rect 37188 28212 37240 28218
rect 37188 28154 37240 28160
rect 36820 27872 36872 27878
rect 36820 27814 36872 27820
rect 36636 27396 36688 27402
rect 36636 27338 36688 27344
rect 36452 26852 36504 26858
rect 36452 26794 36504 26800
rect 36464 26761 36492 26794
rect 36450 26752 36506 26761
rect 36450 26687 36506 26696
rect 36544 26444 36596 26450
rect 36544 26386 36596 26392
rect 36556 25974 36584 26386
rect 36452 25968 36504 25974
rect 36452 25910 36504 25916
rect 36544 25968 36596 25974
rect 36544 25910 36596 25916
rect 36464 25362 36492 25910
rect 36452 25356 36504 25362
rect 36452 25298 36504 25304
rect 36464 24954 36492 25298
rect 36544 25152 36596 25158
rect 36544 25094 36596 25100
rect 36452 24948 36504 24954
rect 36452 24890 36504 24896
rect 36464 24857 36492 24890
rect 36450 24848 36506 24857
rect 36450 24783 36506 24792
rect 36360 24744 36412 24750
rect 36412 24704 36492 24732
rect 36360 24686 36412 24692
rect 36360 24608 36412 24614
rect 36360 24550 36412 24556
rect 36372 24206 36400 24550
rect 36464 24410 36492 24704
rect 36452 24404 36504 24410
rect 36452 24346 36504 24352
rect 36360 24200 36412 24206
rect 36360 24142 36412 24148
rect 36556 23866 36584 25094
rect 36648 23866 36676 27338
rect 36728 27328 36780 27334
rect 36728 27270 36780 27276
rect 36740 25906 36768 27270
rect 36728 25900 36780 25906
rect 36728 25842 36780 25848
rect 36740 25498 36768 25842
rect 36728 25492 36780 25498
rect 36728 25434 36780 25440
rect 36544 23860 36596 23866
rect 36544 23802 36596 23808
rect 36636 23860 36688 23866
rect 36636 23802 36688 23808
rect 36360 23656 36412 23662
rect 36360 23598 36412 23604
rect 36268 23180 36320 23186
rect 36268 23122 36320 23128
rect 36280 22778 36308 23122
rect 36268 22772 36320 22778
rect 36268 22714 36320 22720
rect 36176 22432 36228 22438
rect 36176 22374 36228 22380
rect 36176 21004 36228 21010
rect 36176 20946 36228 20952
rect 36188 20602 36216 20946
rect 36176 20596 36228 20602
rect 36176 20538 36228 20544
rect 36188 20369 36216 20538
rect 36174 20360 36230 20369
rect 36174 20295 36230 20304
rect 36268 20256 36320 20262
rect 36268 20198 36320 20204
rect 36280 19990 36308 20198
rect 35992 19984 36044 19990
rect 35992 19926 36044 19932
rect 36268 19984 36320 19990
rect 36268 19926 36320 19932
rect 35716 19780 35768 19786
rect 35716 19722 35768 19728
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 36004 19514 36032 19926
rect 36280 19514 36308 19926
rect 35992 19508 36044 19514
rect 35992 19450 36044 19456
rect 36268 19508 36320 19514
rect 36268 19450 36320 19456
rect 36082 19000 36138 19009
rect 36082 18935 36138 18944
rect 35256 18896 35308 18902
rect 35256 18838 35308 18844
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 35268 18426 35296 18838
rect 36096 18698 36124 18935
rect 36084 18692 36136 18698
rect 36084 18634 36136 18640
rect 35256 18420 35308 18426
rect 35256 18362 35308 18368
rect 35348 18216 35400 18222
rect 35348 18158 35400 18164
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 35360 17241 35388 18158
rect 35440 17672 35492 17678
rect 35440 17614 35492 17620
rect 35346 17232 35402 17241
rect 35346 17167 35402 17176
rect 35256 17128 35308 17134
rect 35256 17070 35308 17076
rect 35268 16794 35296 17070
rect 35256 16788 35308 16794
rect 35256 16730 35308 16736
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 35268 15502 35296 16730
rect 35360 16674 35388 17167
rect 35452 16794 35480 17614
rect 35992 17332 36044 17338
rect 35992 17274 36044 17280
rect 35808 17060 35860 17066
rect 35808 17002 35860 17008
rect 35440 16788 35492 16794
rect 35440 16730 35492 16736
rect 35360 16646 35480 16674
rect 35256 15496 35308 15502
rect 35256 15438 35308 15444
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 35268 14958 35296 15438
rect 35348 15428 35400 15434
rect 35348 15370 35400 15376
rect 35256 14952 35308 14958
rect 35256 14894 35308 14900
rect 35268 14618 35296 14894
rect 35256 14612 35308 14618
rect 35256 14554 35308 14560
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 35360 12782 35388 15370
rect 35348 12776 35400 12782
rect 35348 12718 35400 12724
rect 35360 12442 35388 12718
rect 35452 12714 35480 16646
rect 35820 16046 35848 17002
rect 36004 16726 36032 17274
rect 35992 16720 36044 16726
rect 35992 16662 36044 16668
rect 35900 16584 35952 16590
rect 35900 16526 35952 16532
rect 35912 16114 35940 16526
rect 36004 16182 36032 16662
rect 35992 16176 36044 16182
rect 35992 16118 36044 16124
rect 35900 16108 35952 16114
rect 35900 16050 35952 16056
rect 35808 16040 35860 16046
rect 35808 15982 35860 15988
rect 35716 15972 35768 15978
rect 35716 15914 35768 15920
rect 35624 14884 35676 14890
rect 35624 14826 35676 14832
rect 35532 14612 35584 14618
rect 35532 14554 35584 14560
rect 35544 13462 35572 14554
rect 35636 13938 35664 14826
rect 35728 14074 35756 15914
rect 35820 15638 35848 15982
rect 35912 15706 35940 16050
rect 35900 15700 35952 15706
rect 35900 15642 35952 15648
rect 35808 15632 35860 15638
rect 35808 15574 35860 15580
rect 36096 15570 36124 18634
rect 36372 17814 36400 23598
rect 36636 22092 36688 22098
rect 36636 22034 36688 22040
rect 36648 21350 36676 22034
rect 36832 22001 36860 27814
rect 37096 27532 37148 27538
rect 37096 27474 37148 27480
rect 37108 26926 37136 27474
rect 37464 27464 37516 27470
rect 37464 27406 37516 27412
rect 37096 26920 37148 26926
rect 37096 26862 37148 26868
rect 37108 26586 37136 26862
rect 37372 26852 37424 26858
rect 37372 26794 37424 26800
rect 37096 26580 37148 26586
rect 37096 26522 37148 26528
rect 36912 25900 36964 25906
rect 36912 25842 36964 25848
rect 36924 24585 36952 25842
rect 37004 25764 37056 25770
rect 37004 25706 37056 25712
rect 37016 25430 37044 25706
rect 37004 25424 37056 25430
rect 37004 25366 37056 25372
rect 37004 24948 37056 24954
rect 37004 24890 37056 24896
rect 36910 24576 36966 24585
rect 36910 24511 36966 24520
rect 36924 22030 36952 24511
rect 37016 22098 37044 24890
rect 37108 23644 37136 26522
rect 37384 26450 37412 26794
rect 37476 26586 37504 27406
rect 37464 26580 37516 26586
rect 37464 26522 37516 26528
rect 37372 26444 37424 26450
rect 37372 26386 37424 26392
rect 37384 26042 37412 26386
rect 37372 26036 37424 26042
rect 37372 25978 37424 25984
rect 37660 25362 37688 28494
rect 37832 28416 37884 28422
rect 37832 28358 37884 28364
rect 37648 25356 37700 25362
rect 37648 25298 37700 25304
rect 37660 24954 37688 25298
rect 37648 24948 37700 24954
rect 37648 24890 37700 24896
rect 37740 24812 37792 24818
rect 37740 24754 37792 24760
rect 37372 24404 37424 24410
rect 37372 24346 37424 24352
rect 37188 23656 37240 23662
rect 37108 23616 37188 23644
rect 37108 23322 37136 23616
rect 37188 23598 37240 23604
rect 37096 23316 37148 23322
rect 37096 23258 37148 23264
rect 37096 22568 37148 22574
rect 37096 22510 37148 22516
rect 37004 22092 37056 22098
rect 37004 22034 37056 22040
rect 36912 22024 36964 22030
rect 36818 21992 36874 22001
rect 36912 21966 36964 21972
rect 36818 21927 36874 21936
rect 37108 21894 37136 22510
rect 37004 21888 37056 21894
rect 37004 21830 37056 21836
rect 37096 21888 37148 21894
rect 37096 21830 37148 21836
rect 36912 21412 36964 21418
rect 36912 21354 36964 21360
rect 36452 21344 36504 21350
rect 36452 21286 36504 21292
rect 36636 21344 36688 21350
rect 36636 21286 36688 21292
rect 36820 21344 36872 21350
rect 36820 21286 36872 21292
rect 36464 21078 36492 21286
rect 36542 21176 36598 21185
rect 36542 21111 36598 21120
rect 36452 21072 36504 21078
rect 36452 21014 36504 21020
rect 36464 20466 36492 21014
rect 36452 20460 36504 20466
rect 36452 20402 36504 20408
rect 36360 17808 36412 17814
rect 36360 17750 36412 17756
rect 36084 15564 36136 15570
rect 36084 15506 36136 15512
rect 36096 15162 36124 15506
rect 36268 15496 36320 15502
rect 36268 15438 36320 15444
rect 36280 15162 36308 15438
rect 36084 15156 36136 15162
rect 36084 15098 36136 15104
rect 36268 15156 36320 15162
rect 36268 15098 36320 15104
rect 36372 15026 36400 17750
rect 36556 17746 36584 21111
rect 36648 20534 36676 21286
rect 36636 20528 36688 20534
rect 36636 20470 36688 20476
rect 36832 20330 36860 21286
rect 36924 20806 36952 21354
rect 37016 20942 37044 21830
rect 37108 21457 37136 21830
rect 37188 21548 37240 21554
rect 37188 21490 37240 21496
rect 37280 21548 37332 21554
rect 37280 21490 37332 21496
rect 37094 21448 37150 21457
rect 37094 21383 37150 21392
rect 37004 20936 37056 20942
rect 37004 20878 37056 20884
rect 36912 20800 36964 20806
rect 36912 20742 36964 20748
rect 36820 20324 36872 20330
rect 36820 20266 36872 20272
rect 36924 20262 36952 20742
rect 36912 20256 36964 20262
rect 36912 20198 36964 20204
rect 36820 19848 36872 19854
rect 36820 19790 36872 19796
rect 36728 19236 36780 19242
rect 36728 19178 36780 19184
rect 36740 18630 36768 19178
rect 36728 18624 36780 18630
rect 36728 18566 36780 18572
rect 36832 18358 36860 19790
rect 36912 19372 36964 19378
rect 36912 19314 36964 19320
rect 36924 18834 36952 19314
rect 37108 19242 37136 21383
rect 37200 20806 37228 21490
rect 37188 20800 37240 20806
rect 37188 20742 37240 20748
rect 37096 19236 37148 19242
rect 37096 19178 37148 19184
rect 36912 18828 36964 18834
rect 36912 18770 36964 18776
rect 36924 18426 36952 18770
rect 36912 18420 36964 18426
rect 36912 18362 36964 18368
rect 36820 18352 36872 18358
rect 36820 18294 36872 18300
rect 36544 17740 36596 17746
rect 36544 17682 36596 17688
rect 36556 17270 36584 17682
rect 36832 17270 36860 18294
rect 37096 18148 37148 18154
rect 37096 18090 37148 18096
rect 37108 17814 37136 18090
rect 37200 17882 37228 20742
rect 37292 19446 37320 21490
rect 37384 19718 37412 24346
rect 37752 23730 37780 24754
rect 37740 23724 37792 23730
rect 37740 23666 37792 23672
rect 37844 23610 37872 28358
rect 37936 27656 37964 29124
rect 38028 27878 38056 32166
rect 38120 31958 38148 32778
rect 38108 31952 38160 31958
rect 38108 31894 38160 31900
rect 38120 31482 38148 31894
rect 38108 31476 38160 31482
rect 38108 31418 38160 31424
rect 38304 29034 38332 33458
rect 38396 33153 38424 35770
rect 38488 35698 38516 36042
rect 38476 35692 38528 35698
rect 38476 35634 38528 35640
rect 38476 33992 38528 33998
rect 38476 33934 38528 33940
rect 38382 33144 38438 33153
rect 38382 33079 38438 33088
rect 38488 32434 38516 33934
rect 38580 33046 38608 38694
rect 38764 38554 38792 39850
rect 38856 39574 38884 39850
rect 38844 39568 38896 39574
rect 38844 39510 38896 39516
rect 38856 38826 38884 39510
rect 38844 38820 38896 38826
rect 38844 38762 38896 38768
rect 38752 38548 38804 38554
rect 38752 38490 38804 38496
rect 38856 38418 38884 38762
rect 38844 38412 38896 38418
rect 38844 38354 38896 38360
rect 38856 38010 38884 38354
rect 38936 38208 38988 38214
rect 38936 38150 38988 38156
rect 38844 38004 38896 38010
rect 38844 37946 38896 37952
rect 38856 37738 38884 37946
rect 38948 37874 38976 38150
rect 38936 37868 38988 37874
rect 38936 37810 38988 37816
rect 38844 37732 38896 37738
rect 38844 37674 38896 37680
rect 38844 37324 38896 37330
rect 38844 37266 38896 37272
rect 38856 36854 38884 37266
rect 38948 36922 38976 37810
rect 39028 37188 39080 37194
rect 39028 37130 39080 37136
rect 39040 36922 39068 37130
rect 38936 36916 38988 36922
rect 38936 36858 38988 36864
rect 39028 36916 39080 36922
rect 39028 36858 39080 36864
rect 38844 36848 38896 36854
rect 38844 36790 38896 36796
rect 38660 35488 38712 35494
rect 38660 35430 38712 35436
rect 38672 35290 38700 35430
rect 38660 35284 38712 35290
rect 38660 35226 38712 35232
rect 38660 34468 38712 34474
rect 38660 34410 38712 34416
rect 38672 34377 38700 34410
rect 38658 34368 38714 34377
rect 38658 34303 38714 34312
rect 38672 34134 38700 34303
rect 38660 34128 38712 34134
rect 38660 34070 38712 34076
rect 39040 34066 39068 36858
rect 39028 34060 39080 34066
rect 39028 34002 39080 34008
rect 39040 33658 39068 34002
rect 39028 33652 39080 33658
rect 39028 33594 39080 33600
rect 39224 33454 39252 40054
rect 39302 38992 39358 39001
rect 39302 38927 39358 38936
rect 39316 38894 39344 38927
rect 39304 38888 39356 38894
rect 39304 38830 39356 38836
rect 39580 38412 39632 38418
rect 39580 38354 39632 38360
rect 39592 37806 39620 38354
rect 39580 37800 39632 37806
rect 39580 37742 39632 37748
rect 39304 37732 39356 37738
rect 39304 37674 39356 37680
rect 39316 35766 39344 37674
rect 39684 36242 39712 40122
rect 41326 39536 41382 39545
rect 40776 39500 40828 39506
rect 41326 39471 41382 39480
rect 40776 39442 40828 39448
rect 39948 38888 40000 38894
rect 39948 38830 40000 38836
rect 39672 36236 39724 36242
rect 39672 36178 39724 36184
rect 39684 35834 39712 36178
rect 39672 35828 39724 35834
rect 39672 35770 39724 35776
rect 39304 35760 39356 35766
rect 39304 35702 39356 35708
rect 39580 35080 39632 35086
rect 39580 35022 39632 35028
rect 39592 34610 39620 35022
rect 39580 34604 39632 34610
rect 39580 34546 39632 34552
rect 39304 34536 39356 34542
rect 39304 34478 39356 34484
rect 39316 33930 39344 34478
rect 39396 34060 39448 34066
rect 39396 34002 39448 34008
rect 39304 33924 39356 33930
rect 39304 33866 39356 33872
rect 39212 33448 39264 33454
rect 39212 33390 39264 33396
rect 39408 33114 39436 34002
rect 39764 33992 39816 33998
rect 39764 33934 39816 33940
rect 39396 33108 39448 33114
rect 39396 33050 39448 33056
rect 38568 33040 38620 33046
rect 38568 32982 38620 32988
rect 38936 33040 38988 33046
rect 38936 32982 38988 32988
rect 38568 32836 38620 32842
rect 38568 32778 38620 32784
rect 38476 32428 38528 32434
rect 38476 32370 38528 32376
rect 38488 32026 38516 32370
rect 38580 32298 38608 32778
rect 38568 32292 38620 32298
rect 38568 32234 38620 32240
rect 38476 32020 38528 32026
rect 38476 31962 38528 31968
rect 38948 31890 38976 32982
rect 39408 32978 39436 33050
rect 39396 32972 39448 32978
rect 39396 32914 39448 32920
rect 39776 32910 39804 33934
rect 39856 33040 39908 33046
rect 39856 32982 39908 32988
rect 39764 32904 39816 32910
rect 39764 32846 39816 32852
rect 39776 32570 39804 32846
rect 39764 32564 39816 32570
rect 39764 32506 39816 32512
rect 39868 32502 39896 32982
rect 39856 32496 39908 32502
rect 39856 32438 39908 32444
rect 38936 31884 38988 31890
rect 38936 31826 38988 31832
rect 39856 31884 39908 31890
rect 39856 31826 39908 31832
rect 38384 31816 38436 31822
rect 38384 31758 38436 31764
rect 38396 30734 38424 31758
rect 39580 31204 39632 31210
rect 39580 31146 39632 31152
rect 38476 30864 38528 30870
rect 38476 30806 38528 30812
rect 38384 30728 38436 30734
rect 38384 30670 38436 30676
rect 38396 30326 38424 30670
rect 38488 30394 38516 30806
rect 38568 30728 38620 30734
rect 38568 30670 38620 30676
rect 38476 30388 38528 30394
rect 38476 30330 38528 30336
rect 38384 30320 38436 30326
rect 38384 30262 38436 30268
rect 38580 29170 38608 30670
rect 39028 30184 39080 30190
rect 39028 30126 39080 30132
rect 38660 29504 38712 29510
rect 38660 29446 38712 29452
rect 38568 29164 38620 29170
rect 38568 29106 38620 29112
rect 38292 29028 38344 29034
rect 38292 28970 38344 28976
rect 38304 28694 38332 28970
rect 38292 28688 38344 28694
rect 38292 28630 38344 28636
rect 38580 28626 38608 29106
rect 38672 29034 38700 29446
rect 38660 29028 38712 29034
rect 38660 28970 38712 28976
rect 38672 28762 38700 28970
rect 39040 28937 39068 30126
rect 39396 29776 39448 29782
rect 39396 29718 39448 29724
rect 39408 29170 39436 29718
rect 39592 29714 39620 31146
rect 39868 31142 39896 31826
rect 39960 31278 39988 38830
rect 40788 38826 40816 39442
rect 40960 39296 41012 39302
rect 40960 39238 41012 39244
rect 40776 38820 40828 38826
rect 40776 38762 40828 38768
rect 40868 38752 40920 38758
rect 40868 38694 40920 38700
rect 40880 38350 40908 38694
rect 40868 38344 40920 38350
rect 40868 38286 40920 38292
rect 40880 38010 40908 38286
rect 40868 38004 40920 38010
rect 40868 37946 40920 37952
rect 40040 37936 40092 37942
rect 40040 37878 40092 37884
rect 40052 37398 40080 37878
rect 40972 37874 41000 39238
rect 41340 38894 41368 39471
rect 41420 39432 41472 39438
rect 41420 39374 41472 39380
rect 41328 38888 41380 38894
rect 41328 38830 41380 38836
rect 41052 38480 41104 38486
rect 41052 38422 41104 38428
rect 40960 37868 41012 37874
rect 40960 37810 41012 37816
rect 40684 37800 40736 37806
rect 40684 37742 40736 37748
rect 40040 37392 40092 37398
rect 40040 37334 40092 37340
rect 40052 36582 40080 37334
rect 40132 37256 40184 37262
rect 40132 37198 40184 37204
rect 40040 36576 40092 36582
rect 40040 36518 40092 36524
rect 40052 35204 40080 36518
rect 40144 36378 40172 37198
rect 40314 36544 40370 36553
rect 40314 36479 40370 36488
rect 40132 36372 40184 36378
rect 40132 36314 40184 36320
rect 40052 35176 40172 35204
rect 40144 34406 40172 35176
rect 40132 34400 40184 34406
rect 40132 34342 40184 34348
rect 40040 33652 40092 33658
rect 40040 33594 40092 33600
rect 39948 31272 40000 31278
rect 39948 31214 40000 31220
rect 39856 31136 39908 31142
rect 39856 31078 39908 31084
rect 39580 29708 39632 29714
rect 39580 29650 39632 29656
rect 39396 29164 39448 29170
rect 39396 29106 39448 29112
rect 39026 28928 39082 28937
rect 39026 28863 39082 28872
rect 39592 28762 39620 29650
rect 39868 29646 39896 31078
rect 39856 29640 39908 29646
rect 39856 29582 39908 29588
rect 38660 28756 38712 28762
rect 38660 28698 38712 28704
rect 39580 28756 39632 28762
rect 39580 28698 39632 28704
rect 38568 28620 38620 28626
rect 38568 28562 38620 28568
rect 39304 28552 39356 28558
rect 39304 28494 39356 28500
rect 38936 28416 38988 28422
rect 38936 28358 38988 28364
rect 38568 28144 38620 28150
rect 38568 28086 38620 28092
rect 38016 27872 38068 27878
rect 38016 27814 38068 27820
rect 38108 27668 38160 27674
rect 37936 27628 38108 27656
rect 38108 27610 38160 27616
rect 38120 27130 38148 27610
rect 38108 27124 38160 27130
rect 38108 27066 38160 27072
rect 38120 26518 38148 27066
rect 38108 26512 38160 26518
rect 38108 26454 38160 26460
rect 38120 25702 38148 26454
rect 38108 25696 38160 25702
rect 38108 25638 38160 25644
rect 38016 24676 38068 24682
rect 38120 24664 38148 25638
rect 38200 25152 38252 25158
rect 38200 25094 38252 25100
rect 38212 24818 38240 25094
rect 38200 24812 38252 24818
rect 38200 24754 38252 24760
rect 38068 24636 38148 24664
rect 38016 24618 38068 24624
rect 38120 24342 38148 24636
rect 38108 24336 38160 24342
rect 38108 24278 38160 24284
rect 37924 24200 37976 24206
rect 37924 24142 37976 24148
rect 37752 23582 37872 23610
rect 37648 22500 37700 22506
rect 37648 22442 37700 22448
rect 37660 22098 37688 22442
rect 37648 22092 37700 22098
rect 37648 22034 37700 22040
rect 37660 21690 37688 22034
rect 37648 21684 37700 21690
rect 37648 21626 37700 21632
rect 37372 19712 37424 19718
rect 37370 19680 37372 19689
rect 37424 19680 37426 19689
rect 37370 19615 37426 19624
rect 37556 19508 37608 19514
rect 37556 19450 37608 19456
rect 37280 19440 37332 19446
rect 37280 19382 37332 19388
rect 37292 18154 37320 19382
rect 37372 18284 37424 18290
rect 37372 18226 37424 18232
rect 37280 18148 37332 18154
rect 37280 18090 37332 18096
rect 37188 17876 37240 17882
rect 37188 17818 37240 17824
rect 37096 17808 37148 17814
rect 37016 17768 37096 17796
rect 36544 17264 36596 17270
rect 36544 17206 36596 17212
rect 36820 17264 36872 17270
rect 36820 17206 36872 17212
rect 36360 15020 36412 15026
rect 36360 14962 36412 14968
rect 36176 14408 36228 14414
rect 36176 14350 36228 14356
rect 36188 14074 36216 14350
rect 35716 14068 35768 14074
rect 35716 14010 35768 14016
rect 35992 14068 36044 14074
rect 35992 14010 36044 14016
rect 36176 14068 36228 14074
rect 36176 14010 36228 14016
rect 35624 13932 35676 13938
rect 35624 13874 35676 13880
rect 35636 13530 35664 13874
rect 36004 13734 36032 14010
rect 36372 13814 36400 14962
rect 36832 14482 36860 17206
rect 37016 17066 37044 17768
rect 37096 17750 37148 17756
rect 37096 17196 37148 17202
rect 37096 17138 37148 17144
rect 37004 17060 37056 17066
rect 37004 17002 37056 17008
rect 37016 16794 37044 17002
rect 37004 16788 37056 16794
rect 37004 16730 37056 16736
rect 37108 16454 37136 17138
rect 37096 16448 37148 16454
rect 37096 16390 37148 16396
rect 37108 16250 37136 16390
rect 37096 16244 37148 16250
rect 37096 16186 37148 16192
rect 37004 15904 37056 15910
rect 37004 15846 37056 15852
rect 37016 15638 37044 15846
rect 37004 15632 37056 15638
rect 37004 15574 37056 15580
rect 37188 15360 37240 15366
rect 37188 15302 37240 15308
rect 37200 15162 37228 15302
rect 37188 15156 37240 15162
rect 37188 15098 37240 15104
rect 37292 14890 37320 18090
rect 37384 17882 37412 18226
rect 37372 17876 37424 17882
rect 37372 17818 37424 17824
rect 37384 16794 37412 17818
rect 37568 17218 37596 19450
rect 37648 18896 37700 18902
rect 37648 18838 37700 18844
rect 37660 18426 37688 18838
rect 37648 18420 37700 18426
rect 37648 18362 37700 18368
rect 37660 17814 37688 18362
rect 37648 17808 37700 17814
rect 37648 17750 37700 17756
rect 37568 17190 37688 17218
rect 37556 17128 37608 17134
rect 37556 17070 37608 17076
rect 37372 16788 37424 16794
rect 37372 16730 37424 16736
rect 37568 15434 37596 17070
rect 37660 16658 37688 17190
rect 37648 16652 37700 16658
rect 37648 16594 37700 16600
rect 37660 16250 37688 16594
rect 37648 16244 37700 16250
rect 37648 16186 37700 16192
rect 37556 15428 37608 15434
rect 37556 15370 37608 15376
rect 36912 14884 36964 14890
rect 36912 14826 36964 14832
rect 37280 14884 37332 14890
rect 37280 14826 37332 14832
rect 36924 14550 36952 14826
rect 36912 14544 36964 14550
rect 36912 14486 36964 14492
rect 36820 14476 36872 14482
rect 36820 14418 36872 14424
rect 36832 13814 36860 14418
rect 36912 14068 36964 14074
rect 36912 14010 36964 14016
rect 36280 13786 36400 13814
rect 36740 13786 36860 13814
rect 35992 13728 36044 13734
rect 35992 13670 36044 13676
rect 35624 13524 35676 13530
rect 35624 13466 35676 13472
rect 36004 13462 36032 13670
rect 35532 13456 35584 13462
rect 35532 13398 35584 13404
rect 35992 13456 36044 13462
rect 35992 13398 36044 13404
rect 35544 12782 35572 13398
rect 35808 13320 35860 13326
rect 35808 13262 35860 13268
rect 35820 12850 35848 13262
rect 35808 12844 35860 12850
rect 35808 12786 35860 12792
rect 35532 12776 35584 12782
rect 35532 12718 35584 12724
rect 35440 12708 35492 12714
rect 35440 12650 35492 12656
rect 35348 12436 35400 12442
rect 35348 12378 35400 12384
rect 34702 12271 34758 12280
rect 34796 12300 34848 12306
rect 34796 12242 34848 12248
rect 33968 12232 34020 12238
rect 33968 12174 34020 12180
rect 34244 12232 34296 12238
rect 34244 12174 34296 12180
rect 33980 11898 34008 12174
rect 33968 11892 34020 11898
rect 33968 11834 34020 11840
rect 33784 11824 33836 11830
rect 33784 11766 33836 11772
rect 34256 11762 34284 12174
rect 35256 12096 35308 12102
rect 35256 12038 35308 12044
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 34244 11756 34296 11762
rect 34244 11698 34296 11704
rect 34256 10198 34284 11698
rect 34336 11620 34388 11626
rect 34336 11562 34388 11568
rect 34348 10198 34376 11562
rect 35268 11218 35296 12038
rect 35256 11212 35308 11218
rect 35256 11154 35308 11160
rect 34704 11008 34756 11014
rect 34704 10950 34756 10956
rect 34716 10742 34744 10950
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 35268 10810 35296 11154
rect 35256 10804 35308 10810
rect 35256 10746 35308 10752
rect 34704 10736 34756 10742
rect 34704 10678 34756 10684
rect 34716 10470 34744 10678
rect 34980 10532 35032 10538
rect 34980 10474 35032 10480
rect 34704 10464 34756 10470
rect 34624 10424 34704 10452
rect 34244 10192 34296 10198
rect 34244 10134 34296 10140
rect 34336 10192 34388 10198
rect 34336 10134 34388 10140
rect 34256 10062 34284 10134
rect 34244 10056 34296 10062
rect 34244 9998 34296 10004
rect 34348 9722 34376 10134
rect 34336 9716 34388 9722
rect 34336 9658 34388 9664
rect 33784 9512 33836 9518
rect 33784 9454 33836 9460
rect 33796 9178 33824 9454
rect 34624 9178 34652 10424
rect 34704 10406 34756 10412
rect 34992 10266 35020 10474
rect 35162 10296 35218 10305
rect 34980 10260 35032 10266
rect 35162 10231 35218 10240
rect 34980 10202 35032 10208
rect 35176 10198 35204 10231
rect 35164 10192 35216 10198
rect 35216 10152 35296 10180
rect 35164 10134 35216 10140
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 35268 9586 35296 10152
rect 35256 9580 35308 9586
rect 35256 9522 35308 9528
rect 34704 9444 34756 9450
rect 34704 9386 34756 9392
rect 35072 9444 35124 9450
rect 35072 9386 35124 9392
rect 35164 9444 35216 9450
rect 35164 9386 35216 9392
rect 33784 9172 33836 9178
rect 33784 9114 33836 9120
rect 34244 9172 34296 9178
rect 34244 9114 34296 9120
rect 34612 9172 34664 9178
rect 34612 9114 34664 9120
rect 34060 8968 34112 8974
rect 34060 8910 34112 8916
rect 34072 8090 34100 8910
rect 34256 8634 34284 9114
rect 34716 8634 34744 9386
rect 35084 9110 35112 9386
rect 35072 9104 35124 9110
rect 35072 9046 35124 9052
rect 35176 9042 35204 9386
rect 35164 9036 35216 9042
rect 35164 8978 35216 8984
rect 34796 8832 34848 8838
rect 34796 8774 34848 8780
rect 34244 8628 34296 8634
rect 34244 8570 34296 8576
rect 34704 8628 34756 8634
rect 34704 8570 34756 8576
rect 34256 8362 34284 8570
rect 34716 8362 34744 8570
rect 34808 8480 34836 8774
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 34980 8492 35032 8498
rect 34808 8452 34980 8480
rect 34980 8434 35032 8440
rect 35256 8492 35308 8498
rect 35256 8434 35308 8440
rect 34992 8401 35020 8434
rect 34978 8392 35034 8401
rect 34244 8356 34296 8362
rect 34244 8298 34296 8304
rect 34704 8356 34756 8362
rect 34978 8327 35034 8336
rect 34704 8298 34756 8304
rect 34060 8084 34112 8090
rect 34060 8026 34112 8032
rect 34256 8022 34284 8298
rect 35268 8022 35296 8434
rect 34244 8016 34296 8022
rect 34244 7958 34296 7964
rect 35256 8016 35308 8022
rect 35256 7958 35308 7964
rect 34256 7546 34284 7958
rect 34520 7880 34572 7886
rect 34520 7822 34572 7828
rect 33416 7540 33468 7546
rect 33416 7482 33468 7488
rect 33600 7540 33652 7546
rect 33600 7482 33652 7488
rect 34244 7540 34296 7546
rect 34244 7482 34296 7488
rect 33324 6656 33376 6662
rect 33324 6598 33376 6604
rect 33336 6322 33364 6598
rect 33324 6316 33376 6322
rect 33324 6258 33376 6264
rect 33428 5914 33456 7482
rect 33612 7342 33640 7482
rect 33600 7336 33652 7342
rect 33600 7278 33652 7284
rect 34532 7206 34560 7822
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 33784 7200 33836 7206
rect 33784 7142 33836 7148
rect 34520 7200 34572 7206
rect 34520 7142 34572 7148
rect 34612 7200 34664 7206
rect 34612 7142 34664 7148
rect 33796 6458 33824 7142
rect 34336 6928 34388 6934
rect 34532 6905 34560 7142
rect 34336 6870 34388 6876
rect 34518 6896 34574 6905
rect 34060 6724 34112 6730
rect 34060 6666 34112 6672
rect 33784 6452 33836 6458
rect 33784 6394 33836 6400
rect 34072 6186 34100 6666
rect 34060 6180 34112 6186
rect 34060 6122 34112 6128
rect 33416 5908 33468 5914
rect 33416 5850 33468 5856
rect 33428 5778 33456 5850
rect 33416 5772 33468 5778
rect 33416 5714 33468 5720
rect 33428 5166 33456 5714
rect 33416 5160 33468 5166
rect 33416 5102 33468 5108
rect 34072 4622 34100 6122
rect 34348 6118 34376 6870
rect 34518 6831 34574 6840
rect 34336 6112 34388 6118
rect 34336 6054 34388 6060
rect 34152 5772 34204 5778
rect 34152 5714 34204 5720
rect 34164 5370 34192 5714
rect 34152 5364 34204 5370
rect 34152 5306 34204 5312
rect 34244 5024 34296 5030
rect 34244 4966 34296 4972
rect 34152 4752 34204 4758
rect 34152 4694 34204 4700
rect 33508 4616 33560 4622
rect 33508 4558 33560 4564
rect 34060 4616 34112 4622
rect 34060 4558 34112 4564
rect 33520 4282 33548 4558
rect 33324 4276 33376 4282
rect 33324 4218 33376 4224
rect 33508 4276 33560 4282
rect 33508 4218 33560 4224
rect 33336 3942 33364 4218
rect 34164 3942 34192 4694
rect 34256 4282 34284 4966
rect 34244 4276 34296 4282
rect 34244 4218 34296 4224
rect 34348 4010 34376 6054
rect 34624 5778 34652 7142
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 35256 6112 35308 6118
rect 35256 6054 35308 6060
rect 34612 5772 34664 5778
rect 34612 5714 34664 5720
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 35268 5137 35296 6054
rect 35452 5710 35480 12650
rect 35544 12220 35572 12718
rect 36176 12300 36228 12306
rect 36176 12242 36228 12248
rect 35624 12232 35676 12238
rect 35544 12192 35624 12220
rect 35544 11286 35572 12192
rect 35624 12174 35676 12180
rect 36188 11898 36216 12242
rect 36176 11892 36228 11898
rect 36176 11834 36228 11840
rect 36188 11354 36216 11834
rect 36176 11348 36228 11354
rect 36176 11290 36228 11296
rect 35532 11280 35584 11286
rect 35532 11222 35584 11228
rect 36280 11218 36308 13786
rect 36544 12640 36596 12646
rect 36544 12582 36596 12588
rect 36556 11626 36584 12582
rect 36636 12096 36688 12102
rect 36636 12038 36688 12044
rect 36648 11694 36676 12038
rect 36636 11688 36688 11694
rect 36636 11630 36688 11636
rect 36544 11620 36596 11626
rect 36544 11562 36596 11568
rect 36268 11212 36320 11218
rect 36268 11154 36320 11160
rect 36544 11212 36596 11218
rect 36544 11154 36596 11160
rect 36280 10810 36308 11154
rect 36556 10810 36584 11154
rect 36740 11150 36768 13786
rect 36924 12986 36952 14010
rect 37648 13456 37700 13462
rect 37648 13398 37700 13404
rect 37660 13190 37688 13398
rect 37648 13184 37700 13190
rect 37648 13126 37700 13132
rect 37660 12986 37688 13126
rect 36912 12980 36964 12986
rect 36912 12922 36964 12928
rect 37648 12980 37700 12986
rect 37648 12922 37700 12928
rect 36912 12096 36964 12102
rect 36912 12038 36964 12044
rect 36924 11762 36952 12038
rect 36912 11756 36964 11762
rect 36912 11698 36964 11704
rect 36924 11286 36952 11698
rect 37648 11552 37700 11558
rect 37648 11494 37700 11500
rect 37660 11286 37688 11494
rect 36912 11280 36964 11286
rect 36912 11222 36964 11228
rect 37648 11280 37700 11286
rect 37648 11222 37700 11228
rect 36728 11144 36780 11150
rect 36728 11086 36780 11092
rect 36740 10810 36768 11086
rect 37660 10810 37688 11222
rect 36268 10804 36320 10810
rect 36268 10746 36320 10752
rect 36544 10804 36596 10810
rect 36544 10746 36596 10752
rect 36728 10804 36780 10810
rect 36728 10746 36780 10752
rect 37648 10804 37700 10810
rect 37648 10746 37700 10752
rect 37752 10742 37780 23582
rect 37936 23322 37964 24142
rect 38120 23526 38148 24278
rect 38200 23656 38252 23662
rect 38580 23610 38608 28086
rect 38660 27940 38712 27946
rect 38660 27882 38712 27888
rect 38844 27940 38896 27946
rect 38844 27882 38896 27888
rect 38672 27674 38700 27882
rect 38752 27872 38804 27878
rect 38752 27814 38804 27820
rect 38660 27668 38712 27674
rect 38660 27610 38712 27616
rect 38672 26858 38700 27610
rect 38660 26852 38712 26858
rect 38660 26794 38712 26800
rect 38660 24608 38712 24614
rect 38660 24550 38712 24556
rect 38672 23866 38700 24550
rect 38764 24290 38792 27814
rect 38856 25294 38884 27882
rect 38948 27538 38976 28358
rect 39316 28218 39344 28494
rect 39580 28484 39632 28490
rect 39580 28426 39632 28432
rect 39304 28212 39356 28218
rect 39304 28154 39356 28160
rect 39488 27668 39540 27674
rect 39488 27610 39540 27616
rect 38936 27532 38988 27538
rect 38936 27474 38988 27480
rect 38948 26994 38976 27474
rect 39212 27396 39264 27402
rect 39212 27338 39264 27344
rect 38936 26988 38988 26994
rect 38936 26930 38988 26936
rect 39120 26852 39172 26858
rect 39120 26794 39172 26800
rect 38936 26240 38988 26246
rect 38936 26182 38988 26188
rect 38948 26042 38976 26182
rect 38936 26036 38988 26042
rect 38936 25978 38988 25984
rect 38948 25752 38976 25978
rect 39028 25764 39080 25770
rect 38948 25724 39028 25752
rect 39028 25706 39080 25712
rect 38936 25424 38988 25430
rect 38936 25366 38988 25372
rect 38844 25288 38896 25294
rect 38844 25230 38896 25236
rect 38856 24886 38884 25230
rect 38948 24954 38976 25366
rect 39028 25288 39080 25294
rect 39028 25230 39080 25236
rect 38936 24948 38988 24954
rect 38936 24890 38988 24896
rect 38844 24880 38896 24886
rect 38844 24822 38896 24828
rect 38948 24410 38976 24890
rect 38936 24404 38988 24410
rect 38936 24346 38988 24352
rect 38764 24262 38976 24290
rect 38660 23860 38712 23866
rect 38660 23802 38712 23808
rect 38200 23598 38252 23604
rect 38108 23520 38160 23526
rect 38108 23462 38160 23468
rect 37924 23316 37976 23322
rect 37924 23258 37976 23264
rect 37924 23180 37976 23186
rect 37924 23122 37976 23128
rect 37936 22545 37964 23122
rect 37922 22536 37978 22545
rect 37922 22471 37978 22480
rect 37936 22438 37964 22471
rect 37924 22432 37976 22438
rect 37924 22374 37976 22380
rect 38016 22432 38068 22438
rect 38016 22374 38068 22380
rect 37924 19984 37976 19990
rect 37924 19926 37976 19932
rect 37936 19174 37964 19926
rect 37924 19168 37976 19174
rect 37924 19110 37976 19116
rect 37936 18086 37964 19110
rect 37924 18080 37976 18086
rect 37924 18022 37976 18028
rect 37832 17740 37884 17746
rect 37832 17682 37884 17688
rect 37844 17270 37872 17682
rect 37832 17264 37884 17270
rect 37832 17206 37884 17212
rect 37936 15638 37964 18022
rect 37924 15632 37976 15638
rect 37924 15574 37976 15580
rect 37924 14884 37976 14890
rect 37924 14826 37976 14832
rect 37936 13326 37964 14826
rect 37924 13320 37976 13326
rect 37924 13262 37976 13268
rect 37832 13184 37884 13190
rect 37832 13126 37884 13132
rect 37844 12918 37872 13126
rect 37832 12912 37884 12918
rect 37832 12854 37884 12860
rect 37936 12442 37964 13262
rect 37924 12436 37976 12442
rect 37924 12378 37976 12384
rect 37740 10736 37792 10742
rect 37740 10678 37792 10684
rect 36176 10532 36228 10538
rect 36176 10474 36228 10480
rect 36188 10062 36216 10474
rect 37832 10464 37884 10470
rect 37832 10406 37884 10412
rect 36268 10192 36320 10198
rect 36268 10134 36320 10140
rect 36176 10056 36228 10062
rect 36176 9998 36228 10004
rect 36188 9722 36216 9998
rect 36176 9716 36228 9722
rect 36176 9658 36228 9664
rect 36280 9586 36308 10134
rect 37844 10130 37872 10406
rect 37832 10124 37884 10130
rect 37832 10066 37884 10072
rect 36820 10056 36872 10062
rect 36820 9998 36872 10004
rect 36268 9580 36320 9586
rect 36268 9522 36320 9528
rect 35808 8968 35860 8974
rect 35808 8910 35860 8916
rect 35532 8900 35584 8906
rect 35532 8842 35584 8848
rect 35544 8265 35572 8842
rect 35820 8566 35848 8910
rect 36280 8634 36308 9522
rect 36544 8832 36596 8838
rect 36544 8774 36596 8780
rect 36268 8628 36320 8634
rect 36268 8570 36320 8576
rect 35808 8560 35860 8566
rect 35808 8502 35860 8508
rect 35530 8256 35586 8265
rect 35530 8191 35586 8200
rect 35544 8090 35572 8191
rect 35532 8084 35584 8090
rect 35532 8026 35584 8032
rect 35820 7886 35848 8502
rect 36280 8362 36308 8570
rect 36556 8498 36584 8774
rect 36544 8492 36596 8498
rect 36544 8434 36596 8440
rect 36268 8356 36320 8362
rect 36268 8298 36320 8304
rect 36360 8288 36412 8294
rect 36280 8236 36360 8242
rect 36280 8230 36412 8236
rect 36280 8214 36400 8230
rect 36280 8022 36308 8214
rect 36360 8084 36412 8090
rect 36360 8026 36412 8032
rect 36268 8016 36320 8022
rect 36268 7958 36320 7964
rect 35808 7880 35860 7886
rect 35808 7822 35860 7828
rect 36176 7880 36228 7886
rect 36176 7822 36228 7828
rect 35808 7472 35860 7478
rect 35808 7414 35860 7420
rect 35820 6934 35848 7414
rect 36188 7002 36216 7822
rect 36280 7546 36308 7958
rect 36268 7540 36320 7546
rect 36268 7482 36320 7488
rect 36372 7410 36400 8026
rect 36832 8022 36860 9998
rect 37844 9722 37872 10066
rect 37832 9716 37884 9722
rect 37832 9658 37884 9664
rect 37832 9444 37884 9450
rect 37832 9386 37884 9392
rect 37844 8974 37872 9386
rect 37924 9376 37976 9382
rect 37924 9318 37976 9324
rect 37936 9110 37964 9318
rect 37924 9104 37976 9110
rect 37924 9046 37976 9052
rect 37832 8968 37884 8974
rect 37832 8910 37884 8916
rect 37844 8634 37872 8910
rect 37832 8628 37884 8634
rect 37832 8570 37884 8576
rect 37188 8492 37240 8498
rect 37188 8434 37240 8440
rect 37200 8090 37228 8434
rect 37936 8294 37964 9046
rect 38028 8430 38056 22374
rect 38120 22216 38148 23462
rect 38212 23168 38240 23598
rect 38396 23582 38608 23610
rect 38396 23497 38424 23582
rect 38382 23488 38438 23497
rect 38580 23474 38608 23582
rect 38672 23576 38700 23802
rect 38844 23588 38896 23594
rect 38672 23548 38844 23576
rect 38844 23530 38896 23536
rect 38750 23488 38806 23497
rect 38580 23446 38700 23474
rect 38382 23423 38438 23432
rect 38292 23180 38344 23186
rect 38212 23140 38292 23168
rect 38292 23122 38344 23128
rect 38304 22778 38332 23122
rect 38292 22772 38344 22778
rect 38292 22714 38344 22720
rect 38568 22704 38620 22710
rect 38568 22646 38620 22652
rect 38384 22500 38436 22506
rect 38384 22442 38436 22448
rect 38292 22228 38344 22234
rect 38120 22188 38292 22216
rect 38292 22170 38344 22176
rect 38304 21350 38332 22170
rect 38292 21344 38344 21350
rect 38292 21286 38344 21292
rect 38108 20460 38160 20466
rect 38108 20402 38160 20408
rect 38120 19718 38148 20402
rect 38108 19712 38160 19718
rect 38108 19654 38160 19660
rect 38120 19145 38148 19654
rect 38106 19136 38162 19145
rect 38106 19071 38162 19080
rect 38200 18148 38252 18154
rect 38120 18108 38200 18136
rect 38120 17882 38148 18108
rect 38200 18090 38252 18096
rect 38108 17876 38160 17882
rect 38108 17818 38160 17824
rect 38120 13258 38148 17818
rect 38396 17270 38424 22442
rect 38580 19446 38608 22646
rect 38672 22234 38700 23446
rect 38948 23474 38976 24262
rect 39040 23594 39068 25230
rect 39132 25208 39160 26794
rect 39224 26246 39252 27338
rect 39500 27130 39528 27610
rect 39592 27606 39620 28426
rect 39580 27600 39632 27606
rect 39580 27542 39632 27548
rect 39592 27130 39620 27542
rect 39488 27124 39540 27130
rect 39488 27066 39540 27072
rect 39580 27124 39632 27130
rect 39580 27066 39632 27072
rect 39764 27056 39816 27062
rect 39764 26998 39816 27004
rect 39776 26450 39804 26998
rect 39764 26444 39816 26450
rect 39764 26386 39816 26392
rect 39212 26240 39264 26246
rect 39212 26182 39264 26188
rect 39224 25906 39252 26182
rect 39776 26042 39804 26386
rect 39764 26036 39816 26042
rect 39684 25996 39764 26024
rect 39212 25900 39264 25906
rect 39212 25842 39264 25848
rect 39580 25764 39632 25770
rect 39580 25706 39632 25712
rect 39592 25294 39620 25706
rect 39580 25288 39632 25294
rect 39580 25230 39632 25236
rect 39212 25220 39264 25226
rect 39132 25180 39212 25208
rect 39132 23730 39160 25180
rect 39212 25162 39264 25168
rect 39488 24948 39540 24954
rect 39488 24890 39540 24896
rect 39120 23724 39172 23730
rect 39172 23684 39252 23712
rect 39120 23666 39172 23672
rect 39028 23588 39080 23594
rect 39028 23530 39080 23536
rect 38750 23423 38806 23432
rect 38856 23446 38976 23474
rect 38764 22710 38792 23423
rect 38752 22704 38804 22710
rect 38752 22646 38804 22652
rect 38752 22432 38804 22438
rect 38752 22374 38804 22380
rect 38660 22228 38712 22234
rect 38660 22170 38712 22176
rect 38660 19984 38712 19990
rect 38660 19926 38712 19932
rect 38672 19514 38700 19926
rect 38764 19854 38792 22374
rect 38856 21185 38884 23446
rect 39040 22574 39068 23530
rect 39224 23322 39252 23684
rect 39212 23316 39264 23322
rect 39212 23258 39264 23264
rect 39304 23180 39356 23186
rect 39304 23122 39356 23128
rect 39316 23089 39344 23122
rect 39302 23080 39358 23089
rect 39302 23015 39358 23024
rect 39316 22710 39344 23015
rect 39304 22704 39356 22710
rect 39304 22646 39356 22652
rect 39028 22568 39080 22574
rect 39028 22510 39080 22516
rect 39028 21888 39080 21894
rect 39028 21830 39080 21836
rect 39040 21418 39068 21830
rect 38936 21412 38988 21418
rect 38936 21354 38988 21360
rect 39028 21412 39080 21418
rect 39028 21354 39080 21360
rect 38842 21176 38898 21185
rect 38948 21146 38976 21354
rect 38842 21111 38898 21120
rect 38936 21140 38988 21146
rect 38856 21010 38884 21111
rect 38936 21082 38988 21088
rect 39040 21078 39068 21354
rect 39028 21072 39080 21078
rect 39028 21014 39080 21020
rect 38844 21004 38896 21010
rect 38844 20946 38896 20952
rect 38856 20602 38884 20946
rect 39040 20602 39068 21014
rect 38844 20596 38896 20602
rect 38844 20538 38896 20544
rect 39028 20596 39080 20602
rect 39028 20538 39080 20544
rect 39212 20324 39264 20330
rect 39212 20266 39264 20272
rect 39224 19854 39252 20266
rect 38752 19848 38804 19854
rect 38752 19790 38804 19796
rect 39212 19848 39264 19854
rect 39212 19790 39264 19796
rect 38660 19508 38712 19514
rect 38660 19450 38712 19456
rect 38568 19440 38620 19446
rect 38568 19382 38620 19388
rect 38580 19310 38608 19382
rect 38568 19304 38620 19310
rect 38568 19246 38620 19252
rect 38476 19236 38528 19242
rect 38476 19178 38528 19184
rect 38488 17746 38516 19178
rect 38580 18698 38608 19246
rect 38764 18970 38792 19790
rect 38752 18964 38804 18970
rect 38752 18906 38804 18912
rect 38844 18760 38896 18766
rect 38844 18702 38896 18708
rect 38568 18692 38620 18698
rect 38568 18634 38620 18640
rect 38568 18080 38620 18086
rect 38568 18022 38620 18028
rect 38580 17882 38608 18022
rect 38856 17882 38884 18702
rect 39224 18698 39252 19790
rect 39500 19378 39528 24890
rect 39684 23497 39712 25996
rect 39764 25978 39816 25984
rect 39764 25764 39816 25770
rect 39764 25706 39816 25712
rect 39670 23488 39726 23497
rect 39670 23423 39726 23432
rect 39776 23186 39804 25706
rect 39868 24750 39896 29582
rect 40052 25974 40080 33594
rect 40144 33046 40172 34342
rect 40328 34066 40356 36479
rect 40590 36136 40646 36145
rect 40590 36071 40646 36080
rect 40316 34060 40368 34066
rect 40316 34002 40368 34008
rect 40328 33658 40356 34002
rect 40316 33652 40368 33658
rect 40316 33594 40368 33600
rect 40500 33312 40552 33318
rect 40500 33254 40552 33260
rect 40132 33040 40184 33046
rect 40132 32982 40184 32988
rect 40316 31952 40368 31958
rect 40316 31894 40368 31900
rect 40328 31482 40356 31894
rect 40316 31476 40368 31482
rect 40316 31418 40368 31424
rect 40316 31272 40368 31278
rect 40316 31214 40368 31220
rect 40224 28552 40276 28558
rect 40224 28494 40276 28500
rect 40236 27878 40264 28494
rect 40224 27872 40276 27878
rect 40224 27814 40276 27820
rect 40236 27334 40264 27814
rect 40224 27328 40276 27334
rect 40224 27270 40276 27276
rect 40236 26994 40264 27270
rect 40224 26988 40276 26994
rect 40224 26930 40276 26936
rect 40236 26450 40264 26930
rect 40224 26444 40276 26450
rect 40224 26386 40276 26392
rect 40040 25968 40092 25974
rect 40040 25910 40092 25916
rect 39856 24744 39908 24750
rect 39856 24686 39908 24692
rect 40052 23474 40080 25910
rect 40236 25770 40264 26386
rect 40224 25764 40276 25770
rect 40224 25706 40276 25712
rect 40328 25362 40356 31214
rect 40408 30864 40460 30870
rect 40408 30806 40460 30812
rect 40420 30394 40448 30806
rect 40408 30388 40460 30394
rect 40408 30330 40460 30336
rect 40420 29850 40448 30330
rect 40408 29844 40460 29850
rect 40408 29786 40460 29792
rect 40512 27282 40540 33254
rect 40604 31414 40632 36071
rect 40592 31408 40644 31414
rect 40592 31350 40644 31356
rect 40696 30870 40724 37742
rect 40868 37664 40920 37670
rect 40868 37606 40920 37612
rect 40880 37466 40908 37606
rect 40972 37466 41000 37810
rect 41064 37738 41092 38422
rect 41432 38282 41460 39374
rect 41524 39098 41552 49558
rect 41602 49520 41658 49558
rect 46952 49558 47178 49586
rect 43074 43616 43130 43625
rect 43074 43551 43130 43560
rect 43088 40769 43116 43551
rect 43074 40760 43130 40769
rect 43074 40695 43130 40704
rect 42156 39908 42208 39914
rect 42156 39850 42208 39856
rect 41512 39092 41564 39098
rect 41512 39034 41564 39040
rect 41420 38276 41472 38282
rect 41420 38218 41472 38224
rect 41236 37868 41288 37874
rect 41236 37810 41288 37816
rect 41052 37732 41104 37738
rect 41052 37674 41104 37680
rect 40868 37460 40920 37466
rect 40868 37402 40920 37408
rect 40960 37460 41012 37466
rect 40960 37402 41012 37408
rect 41144 36712 41196 36718
rect 41144 36654 41196 36660
rect 40868 36304 40920 36310
rect 40868 36246 40920 36252
rect 40776 36032 40828 36038
rect 40776 35974 40828 35980
rect 40788 35698 40816 35974
rect 40776 35692 40828 35698
rect 40776 35634 40828 35640
rect 40788 35290 40816 35634
rect 40880 35562 40908 36246
rect 41156 36145 41184 36654
rect 41248 36378 41276 37810
rect 41236 36372 41288 36378
rect 41236 36314 41288 36320
rect 41142 36136 41198 36145
rect 41142 36071 41198 36080
rect 41432 36038 41460 38218
rect 42168 37942 42196 39850
rect 46952 38894 46980 49558
rect 47122 49520 47178 49558
rect 46940 38888 46992 38894
rect 46940 38830 46992 38836
rect 42524 38208 42576 38214
rect 42524 38150 42576 38156
rect 42156 37936 42208 37942
rect 42156 37878 42208 37884
rect 41604 37392 41656 37398
rect 41604 37334 41656 37340
rect 41616 36922 41644 37334
rect 41788 37256 41840 37262
rect 41788 37198 41840 37204
rect 41604 36916 41656 36922
rect 41604 36858 41656 36864
rect 41800 36854 41828 37198
rect 41788 36848 41840 36854
rect 41788 36790 41840 36796
rect 41696 36712 41748 36718
rect 41696 36654 41748 36660
rect 41708 36553 41736 36654
rect 41694 36544 41750 36553
rect 41694 36479 41750 36488
rect 41800 36378 41828 36790
rect 41788 36372 41840 36378
rect 41788 36314 41840 36320
rect 41696 36168 41748 36174
rect 41696 36110 41748 36116
rect 41420 36032 41472 36038
rect 41420 35974 41472 35980
rect 41432 35698 41460 35974
rect 41708 35834 41736 36110
rect 41696 35828 41748 35834
rect 41696 35770 41748 35776
rect 41420 35692 41472 35698
rect 41420 35634 41472 35640
rect 40868 35556 40920 35562
rect 40868 35498 40920 35504
rect 40776 35284 40828 35290
rect 40776 35226 40828 35232
rect 40880 35222 40908 35498
rect 40868 35216 40920 35222
rect 40868 35158 40920 35164
rect 41512 35216 41564 35222
rect 41512 35158 41564 35164
rect 41420 35080 41472 35086
rect 41420 35022 41472 35028
rect 41432 34202 41460 35022
rect 41524 34746 41552 35158
rect 41708 34746 41736 35770
rect 42064 35488 42116 35494
rect 42064 35430 42116 35436
rect 41512 34740 41564 34746
rect 41512 34682 41564 34688
rect 41696 34740 41748 34746
rect 41696 34682 41748 34688
rect 41972 34672 42024 34678
rect 41972 34614 42024 34620
rect 41420 34196 41472 34202
rect 41420 34138 41472 34144
rect 41696 34060 41748 34066
rect 41696 34002 41748 34008
rect 40776 33856 40828 33862
rect 40776 33798 40828 33804
rect 40788 33522 40816 33798
rect 41708 33658 41736 34002
rect 41512 33652 41564 33658
rect 41512 33594 41564 33600
rect 41696 33652 41748 33658
rect 41696 33594 41748 33600
rect 40776 33516 40828 33522
rect 40776 33458 40828 33464
rect 40868 33380 40920 33386
rect 40868 33322 40920 33328
rect 40880 33046 40908 33322
rect 40868 33040 40920 33046
rect 40868 32982 40920 32988
rect 40880 32774 40908 32982
rect 40868 32768 40920 32774
rect 40868 32710 40920 32716
rect 41052 32768 41104 32774
rect 41052 32710 41104 32716
rect 40880 32230 40908 32710
rect 41064 32298 41092 32710
rect 41144 32428 41196 32434
rect 41144 32370 41196 32376
rect 41052 32292 41104 32298
rect 41052 32234 41104 32240
rect 40868 32224 40920 32230
rect 40868 32166 40920 32172
rect 40880 31958 40908 32166
rect 40868 31952 40920 31958
rect 40868 31894 40920 31900
rect 40776 31816 40828 31822
rect 40776 31758 40828 31764
rect 40788 31210 40816 31758
rect 41064 31482 41092 32234
rect 41156 31822 41184 32370
rect 41144 31816 41196 31822
rect 41144 31758 41196 31764
rect 41156 31686 41184 31758
rect 41144 31680 41196 31686
rect 41144 31622 41196 31628
rect 41052 31476 41104 31482
rect 41052 31418 41104 31424
rect 40868 31408 40920 31414
rect 40868 31350 40920 31356
rect 40776 31204 40828 31210
rect 40776 31146 40828 31152
rect 40880 31142 40908 31350
rect 40868 31136 40920 31142
rect 40868 31078 40920 31084
rect 40684 30864 40736 30870
rect 40684 30806 40736 30812
rect 40776 30728 40828 30734
rect 40776 30670 40828 30676
rect 40788 29850 40816 30670
rect 40776 29844 40828 29850
rect 40776 29786 40828 29792
rect 40684 28688 40736 28694
rect 40684 28630 40736 28636
rect 40696 28218 40724 28630
rect 40684 28212 40736 28218
rect 40684 28154 40736 28160
rect 40420 27254 40540 27282
rect 40316 25356 40368 25362
rect 40316 25298 40368 25304
rect 40328 24954 40356 25298
rect 40316 24948 40368 24954
rect 40316 24890 40368 24896
rect 40052 23446 40264 23474
rect 40236 23186 40264 23446
rect 39764 23180 39816 23186
rect 39764 23122 39816 23128
rect 40224 23180 40276 23186
rect 40224 23122 40276 23128
rect 39776 22778 39804 23122
rect 39764 22772 39816 22778
rect 39764 22714 39816 22720
rect 40040 22160 40092 22166
rect 40040 22102 40092 22108
rect 39948 22024 40000 22030
rect 39948 21966 40000 21972
rect 39960 21690 39988 21966
rect 39948 21684 40000 21690
rect 39948 21626 40000 21632
rect 40052 21554 40080 22102
rect 40040 21548 40092 21554
rect 40040 21490 40092 21496
rect 39580 21412 39632 21418
rect 39580 21354 39632 21360
rect 39488 19372 39540 19378
rect 39488 19314 39540 19320
rect 39212 18692 39264 18698
rect 39212 18634 39264 18640
rect 38568 17876 38620 17882
rect 38568 17818 38620 17824
rect 38844 17876 38896 17882
rect 38844 17818 38896 17824
rect 38476 17740 38528 17746
rect 38476 17682 38528 17688
rect 38384 17264 38436 17270
rect 38384 17206 38436 17212
rect 38488 17116 38516 17682
rect 38568 17128 38620 17134
rect 38488 17088 38568 17116
rect 38568 17070 38620 17076
rect 38580 16794 38608 17070
rect 38568 16788 38620 16794
rect 38568 16730 38620 16736
rect 38292 16720 38344 16726
rect 38292 16662 38344 16668
rect 38304 15978 38332 16662
rect 39028 16448 39080 16454
rect 39028 16390 39080 16396
rect 39040 16114 39068 16390
rect 39028 16108 39080 16114
rect 39028 16050 39080 16056
rect 38292 15972 38344 15978
rect 38292 15914 38344 15920
rect 38844 15972 38896 15978
rect 38844 15914 38896 15920
rect 38304 15706 38332 15914
rect 38384 15904 38436 15910
rect 38384 15846 38436 15852
rect 38292 15700 38344 15706
rect 38292 15642 38344 15648
rect 38396 15586 38424 15846
rect 38304 15558 38424 15586
rect 38198 14512 38254 14521
rect 38198 14447 38254 14456
rect 38108 13252 38160 13258
rect 38108 13194 38160 13200
rect 38212 12986 38240 14447
rect 38304 14006 38332 15558
rect 38856 15502 38884 15914
rect 38476 15496 38528 15502
rect 38476 15438 38528 15444
rect 38844 15496 38896 15502
rect 38844 15438 38896 15444
rect 38488 15026 38516 15438
rect 38476 15020 38528 15026
rect 38476 14962 38528 14968
rect 38476 14544 38528 14550
rect 38396 14504 38476 14532
rect 38292 14000 38344 14006
rect 38292 13942 38344 13948
rect 38200 12980 38252 12986
rect 38200 12922 38252 12928
rect 38212 12782 38240 12922
rect 38200 12776 38252 12782
rect 38200 12718 38252 12724
rect 38304 11898 38332 13942
rect 38396 13734 38424 14504
rect 38476 14486 38528 14492
rect 38476 14408 38528 14414
rect 38476 14350 38528 14356
rect 38384 13728 38436 13734
rect 38384 13670 38436 13676
rect 38488 13716 38516 14350
rect 38856 13938 38884 15438
rect 39040 15162 39068 16050
rect 39120 15632 39172 15638
rect 39120 15574 39172 15580
rect 39028 15156 39080 15162
rect 39028 15098 39080 15104
rect 39132 15094 39160 15574
rect 39120 15088 39172 15094
rect 39120 15030 39172 15036
rect 39224 14414 39252 18634
rect 39592 18426 39620 21354
rect 40052 21078 40080 21490
rect 40040 21072 40092 21078
rect 40040 21014 40092 21020
rect 39672 20936 39724 20942
rect 39672 20878 39724 20884
rect 40040 20936 40092 20942
rect 40040 20878 40092 20884
rect 39684 20602 39712 20878
rect 39672 20596 39724 20602
rect 39672 20538 39724 20544
rect 40052 20466 40080 20878
rect 40040 20460 40092 20466
rect 40040 20402 40092 20408
rect 40132 19848 40184 19854
rect 40132 19790 40184 19796
rect 40144 19310 40172 19790
rect 40132 19304 40184 19310
rect 40132 19246 40184 19252
rect 40144 18970 40172 19246
rect 40132 18964 40184 18970
rect 40132 18906 40184 18912
rect 40236 18834 40264 23122
rect 40314 21992 40370 22001
rect 40314 21927 40370 21936
rect 40328 21486 40356 21927
rect 40316 21480 40368 21486
rect 40316 21422 40368 21428
rect 40224 18828 40276 18834
rect 40224 18770 40276 18776
rect 39580 18420 39632 18426
rect 39580 18362 39632 18368
rect 40236 18358 40264 18770
rect 40224 18352 40276 18358
rect 40224 18294 40276 18300
rect 39488 17808 39540 17814
rect 39488 17750 39540 17756
rect 39500 17338 39528 17750
rect 39856 17672 39908 17678
rect 39856 17614 39908 17620
rect 39868 17338 39896 17614
rect 39488 17332 39540 17338
rect 39488 17274 39540 17280
rect 39856 17332 39908 17338
rect 39856 17274 39908 17280
rect 39396 16652 39448 16658
rect 39396 16594 39448 16600
rect 39408 15910 39436 16594
rect 39500 16250 39528 17274
rect 39856 16652 39908 16658
rect 39856 16594 39908 16600
rect 39488 16244 39540 16250
rect 39488 16186 39540 16192
rect 39868 16182 39896 16594
rect 39856 16176 39908 16182
rect 40236 16153 40264 18294
rect 40316 17536 40368 17542
rect 40316 17478 40368 17484
rect 40328 17338 40356 17478
rect 40316 17332 40368 17338
rect 40316 17274 40368 17280
rect 40328 16998 40356 17274
rect 40316 16992 40368 16998
rect 40316 16934 40368 16940
rect 39856 16118 39908 16124
rect 40222 16144 40278 16153
rect 39396 15904 39448 15910
rect 39396 15846 39448 15852
rect 39868 15502 39896 16118
rect 40222 16079 40278 16088
rect 39856 15496 39908 15502
rect 39856 15438 39908 15444
rect 39868 15162 39896 15438
rect 39856 15156 39908 15162
rect 39856 15098 39908 15104
rect 39212 14408 39264 14414
rect 39212 14350 39264 14356
rect 38844 13932 38896 13938
rect 38844 13874 38896 13880
rect 38856 13814 38884 13874
rect 38856 13786 38976 13814
rect 38660 13728 38712 13734
rect 38488 13688 38660 13716
rect 38396 13530 38424 13670
rect 38384 13524 38436 13530
rect 38384 13466 38436 13472
rect 38384 13252 38436 13258
rect 38384 13194 38436 13200
rect 38396 12850 38424 13194
rect 38488 12918 38516 13688
rect 38660 13670 38712 13676
rect 38476 12912 38528 12918
rect 38476 12854 38528 12860
rect 38384 12844 38436 12850
rect 38384 12786 38436 12792
rect 38292 11892 38344 11898
rect 38292 11834 38344 11840
rect 38304 11694 38332 11834
rect 38292 11688 38344 11694
rect 38292 11630 38344 11636
rect 38292 11144 38344 11150
rect 38396 11132 38424 12786
rect 38948 12714 38976 13786
rect 39224 13326 39252 14350
rect 40236 13814 40264 16079
rect 40052 13786 40264 13814
rect 39580 13728 39632 13734
rect 39580 13670 39632 13676
rect 39488 13456 39540 13462
rect 39488 13398 39540 13404
rect 39212 13320 39264 13326
rect 39212 13262 39264 13268
rect 39500 12986 39528 13398
rect 39488 12980 39540 12986
rect 39488 12922 39540 12928
rect 38936 12708 38988 12714
rect 38936 12650 38988 12656
rect 38948 12442 38976 12650
rect 38936 12436 38988 12442
rect 38936 12378 38988 12384
rect 39396 12436 39448 12442
rect 39396 12378 39448 12384
rect 38844 12232 38896 12238
rect 38844 12174 38896 12180
rect 39028 12232 39080 12238
rect 39028 12174 39080 12180
rect 38856 11694 38884 12174
rect 39040 11762 39068 12174
rect 39408 11898 39436 12378
rect 39396 11892 39448 11898
rect 39396 11834 39448 11840
rect 39028 11756 39080 11762
rect 39028 11698 39080 11704
rect 38844 11688 38896 11694
rect 38896 11648 38976 11676
rect 38844 11630 38896 11636
rect 38344 11104 38424 11132
rect 38292 11086 38344 11092
rect 38108 8968 38160 8974
rect 38108 8910 38160 8916
rect 38120 8498 38148 8910
rect 38108 8492 38160 8498
rect 38108 8434 38160 8440
rect 38016 8424 38068 8430
rect 38016 8366 38068 8372
rect 37924 8288 37976 8294
rect 37924 8230 37976 8236
rect 38200 8288 38252 8294
rect 38200 8230 38252 8236
rect 37188 8084 37240 8090
rect 37188 8026 37240 8032
rect 36820 8016 36872 8022
rect 36820 7958 36872 7964
rect 37924 8016 37976 8022
rect 37924 7958 37976 7964
rect 37832 7880 37884 7886
rect 37832 7822 37884 7828
rect 37844 7546 37872 7822
rect 37832 7540 37884 7546
rect 37832 7482 37884 7488
rect 37280 7472 37332 7478
rect 37280 7414 37332 7420
rect 36360 7404 36412 7410
rect 36360 7346 36412 7352
rect 36360 7268 36412 7274
rect 36360 7210 36412 7216
rect 36176 6996 36228 7002
rect 36176 6938 36228 6944
rect 35808 6928 35860 6934
rect 35808 6870 35860 6876
rect 35900 6860 35952 6866
rect 35900 6802 35952 6808
rect 35912 6458 35940 6802
rect 36372 6798 36400 7210
rect 36912 6928 36964 6934
rect 36912 6870 36964 6876
rect 36360 6792 36412 6798
rect 36360 6734 36412 6740
rect 36924 6458 36952 6870
rect 37292 6458 37320 7414
rect 37936 7410 37964 7958
rect 38108 7880 38160 7886
rect 38108 7822 38160 7828
rect 38120 7478 38148 7822
rect 38108 7472 38160 7478
rect 38108 7414 38160 7420
rect 37924 7404 37976 7410
rect 37924 7346 37976 7352
rect 38212 7342 38240 8230
rect 38200 7336 38252 7342
rect 38200 7278 38252 7284
rect 35900 6452 35952 6458
rect 35900 6394 35952 6400
rect 36912 6452 36964 6458
rect 36912 6394 36964 6400
rect 37280 6452 37332 6458
rect 37280 6394 37332 6400
rect 36358 6352 36414 6361
rect 36358 6287 36414 6296
rect 36372 5846 36400 6287
rect 37292 6254 37320 6394
rect 38304 6254 38332 11086
rect 38948 10742 38976 11648
rect 39408 11626 39436 11834
rect 39396 11620 39448 11626
rect 39396 11562 39448 11568
rect 39396 11212 39448 11218
rect 39396 11154 39448 11160
rect 39408 10810 39436 11154
rect 39396 10804 39448 10810
rect 39396 10746 39448 10752
rect 38844 10736 38896 10742
rect 38844 10678 38896 10684
rect 38936 10736 38988 10742
rect 38936 10678 38988 10684
rect 38856 9518 38884 10678
rect 38844 9512 38896 9518
rect 38844 9454 38896 9460
rect 38476 8424 38528 8430
rect 38476 8366 38528 8372
rect 38488 7954 38516 8366
rect 38476 7948 38528 7954
rect 38476 7890 38528 7896
rect 39304 7948 39356 7954
rect 39304 7890 39356 7896
rect 38476 7744 38528 7750
rect 38476 7686 38528 7692
rect 38488 6866 38516 7686
rect 39316 7546 39344 7890
rect 39304 7540 39356 7546
rect 39304 7482 39356 7488
rect 38476 6860 38528 6866
rect 38476 6802 38528 6808
rect 38488 6458 38516 6802
rect 38476 6452 38528 6458
rect 38476 6394 38528 6400
rect 37280 6248 37332 6254
rect 37280 6190 37332 6196
rect 38292 6248 38344 6254
rect 38292 6190 38344 6196
rect 37832 6112 37884 6118
rect 37832 6054 37884 6060
rect 36084 5840 36136 5846
rect 36084 5782 36136 5788
rect 36360 5840 36412 5846
rect 36360 5782 36412 5788
rect 35440 5704 35492 5710
rect 35440 5646 35492 5652
rect 35254 5128 35310 5137
rect 35254 5063 35310 5072
rect 36096 5030 36124 5782
rect 36176 5636 36228 5642
rect 36228 5596 36308 5624
rect 36176 5578 36228 5584
rect 36084 5024 36136 5030
rect 36084 4966 36136 4972
rect 36096 4758 36124 4966
rect 36084 4752 36136 4758
rect 36084 4694 36136 4700
rect 35992 4684 36044 4690
rect 35992 4626 36044 4632
rect 34704 4616 34756 4622
rect 34704 4558 34756 4564
rect 34612 4548 34664 4554
rect 34612 4490 34664 4496
rect 34336 4004 34388 4010
rect 34336 3946 34388 3952
rect 33324 3936 33376 3942
rect 33324 3878 33376 3884
rect 34152 3936 34204 3942
rect 34152 3878 34204 3884
rect 33336 2446 33364 3878
rect 33508 3664 33560 3670
rect 33508 3606 33560 3612
rect 33876 3664 33928 3670
rect 33876 3606 33928 3612
rect 33520 3534 33548 3606
rect 33508 3528 33560 3534
rect 33508 3470 33560 3476
rect 33784 3528 33836 3534
rect 33784 3470 33836 3476
rect 33600 2848 33652 2854
rect 33600 2790 33652 2796
rect 33692 2848 33744 2854
rect 33692 2790 33744 2796
rect 33612 2553 33640 2790
rect 33704 2689 33732 2790
rect 33690 2680 33746 2689
rect 33690 2615 33746 2624
rect 33796 2582 33824 3470
rect 33888 3194 33916 3606
rect 34624 3466 34652 4490
rect 34716 3738 34744 4558
rect 34796 4480 34848 4486
rect 34796 4422 34848 4428
rect 35900 4480 35952 4486
rect 35900 4422 35952 4428
rect 34808 4146 34836 4422
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 35912 4146 35940 4422
rect 36004 4282 36032 4626
rect 35992 4276 36044 4282
rect 35992 4218 36044 4224
rect 36280 4146 36308 5596
rect 36372 4214 36400 5782
rect 37844 5778 37872 6054
rect 37832 5772 37884 5778
rect 37832 5714 37884 5720
rect 36912 5704 36964 5710
rect 36912 5646 36964 5652
rect 36544 5568 36596 5574
rect 36544 5510 36596 5516
rect 36556 5166 36584 5510
rect 36924 5370 36952 5646
rect 37844 5370 37872 5714
rect 36912 5364 36964 5370
rect 36912 5306 36964 5312
rect 37832 5364 37884 5370
rect 37832 5306 37884 5312
rect 36544 5160 36596 5166
rect 36544 5102 36596 5108
rect 36556 4826 36584 5102
rect 36636 5092 36688 5098
rect 36636 5034 36688 5040
rect 36544 4820 36596 4826
rect 36544 4762 36596 4768
rect 36648 4282 36676 5034
rect 36636 4276 36688 4282
rect 36636 4218 36688 4224
rect 36360 4208 36412 4214
rect 36360 4150 36412 4156
rect 36924 4154 36952 5306
rect 37844 5166 37872 5306
rect 37832 5160 37884 5166
rect 37832 5102 37884 5108
rect 37648 5024 37700 5030
rect 37648 4966 37700 4972
rect 37660 4690 37688 4966
rect 37648 4684 37700 4690
rect 37648 4626 37700 4632
rect 38108 4480 38160 4486
rect 38108 4422 38160 4428
rect 36832 4146 36952 4154
rect 38120 4146 38148 4422
rect 38200 4276 38252 4282
rect 38200 4218 38252 4224
rect 34796 4140 34848 4146
rect 34796 4082 34848 4088
rect 35900 4140 35952 4146
rect 35900 4082 35952 4088
rect 36268 4140 36320 4146
rect 36268 4082 36320 4088
rect 36820 4140 36952 4146
rect 36872 4126 36952 4140
rect 38108 4140 38160 4146
rect 36820 4082 36872 4088
rect 38108 4082 38160 4088
rect 35072 4004 35124 4010
rect 35072 3946 35124 3952
rect 34704 3732 34756 3738
rect 34704 3674 34756 3680
rect 35084 3670 35112 3946
rect 36280 3738 36308 4082
rect 36360 3936 36412 3942
rect 36360 3878 36412 3884
rect 36268 3732 36320 3738
rect 36268 3674 36320 3680
rect 35072 3664 35124 3670
rect 35072 3606 35124 3612
rect 35256 3664 35308 3670
rect 35256 3606 35308 3612
rect 34336 3460 34388 3466
rect 34336 3402 34388 3408
rect 34612 3460 34664 3466
rect 34612 3402 34664 3408
rect 33876 3188 33928 3194
rect 33876 3130 33928 3136
rect 33784 2576 33836 2582
rect 33598 2544 33654 2553
rect 33784 2518 33836 2524
rect 33598 2479 33654 2488
rect 34348 2446 34376 3402
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 35268 2650 35296 3606
rect 35440 3596 35492 3602
rect 35440 3538 35492 3544
rect 35452 2854 35480 3538
rect 36176 3392 36228 3398
rect 36176 3334 36228 3340
rect 36188 2990 36216 3334
rect 36372 3058 36400 3878
rect 36360 3052 36412 3058
rect 36360 2994 36412 3000
rect 36176 2984 36228 2990
rect 36176 2926 36228 2932
rect 35440 2848 35492 2854
rect 35440 2790 35492 2796
rect 35452 2650 35480 2790
rect 35256 2644 35308 2650
rect 35256 2586 35308 2592
rect 35440 2644 35492 2650
rect 35440 2586 35492 2592
rect 36832 2582 36860 4082
rect 37740 3596 37792 3602
rect 37740 3538 37792 3544
rect 37188 3528 37240 3534
rect 37188 3470 37240 3476
rect 37200 3058 37228 3470
rect 37752 3194 37780 3538
rect 37740 3188 37792 3194
rect 37740 3130 37792 3136
rect 37188 3052 37240 3058
rect 37188 2994 37240 3000
rect 37752 2650 37780 3130
rect 38120 3058 38148 4082
rect 38212 4010 38240 4218
rect 39592 4154 39620 13670
rect 39948 12980 40000 12986
rect 39948 12922 40000 12928
rect 39960 12442 39988 12922
rect 39948 12436 40000 12442
rect 39948 12378 40000 12384
rect 39764 11212 39816 11218
rect 39764 11154 39816 11160
rect 39776 10742 39804 11154
rect 39764 10736 39816 10742
rect 39764 10678 39816 10684
rect 39500 4126 39620 4154
rect 38200 4004 38252 4010
rect 38200 3946 38252 3952
rect 39500 3194 39528 4126
rect 39488 3188 39540 3194
rect 39488 3130 39540 3136
rect 38108 3052 38160 3058
rect 38108 2994 38160 3000
rect 37740 2644 37792 2650
rect 37740 2586 37792 2592
rect 36820 2576 36872 2582
rect 36820 2518 36872 2524
rect 33324 2440 33376 2446
rect 33324 2382 33376 2388
rect 34336 2440 34388 2446
rect 34336 2382 34388 2388
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 30208 54 30342 82
rect 33232 128 33284 134
rect 33232 70 33284 76
rect 33874 128 33930 480
rect 33874 76 33876 128
rect 33928 76 33930 128
rect 23110 0 23166 54
rect 26698 0 26754 54
rect 30286 0 30342 54
rect 33874 0 33930 76
rect 37370 0 37426 480
rect 40052 134 40080 13786
rect 40224 13320 40276 13326
rect 40224 13262 40276 13268
rect 40236 12986 40264 13262
rect 40420 13190 40448 27254
rect 40774 26888 40830 26897
rect 40880 26874 40908 31078
rect 41156 30734 41184 31622
rect 41236 31204 41288 31210
rect 41236 31146 41288 31152
rect 41248 30938 41276 31146
rect 41236 30932 41288 30938
rect 41236 30874 41288 30880
rect 41144 30728 41196 30734
rect 41144 30670 41196 30676
rect 41524 30326 41552 33594
rect 41984 33454 42012 34614
rect 42076 34610 42104 35430
rect 42168 35154 42196 37878
rect 42536 37738 42564 38150
rect 42524 37732 42576 37738
rect 42524 37674 42576 37680
rect 42536 36922 42564 37674
rect 42616 37256 42668 37262
rect 42616 37198 42668 37204
rect 42524 36916 42576 36922
rect 42524 36858 42576 36864
rect 42340 36644 42392 36650
rect 42340 36586 42392 36592
rect 42156 35148 42208 35154
rect 42156 35090 42208 35096
rect 42064 34604 42116 34610
rect 42064 34546 42116 34552
rect 42352 34524 42380 36586
rect 42432 36032 42484 36038
rect 42432 35974 42484 35980
rect 42444 35562 42472 35974
rect 42628 35698 42656 37198
rect 42616 35692 42668 35698
rect 42616 35634 42668 35640
rect 42432 35556 42484 35562
rect 42432 35498 42484 35504
rect 42444 35222 42472 35498
rect 42432 35216 42484 35222
rect 42432 35158 42484 35164
rect 42432 34536 42484 34542
rect 42352 34496 42432 34524
rect 42432 34478 42484 34484
rect 42248 34400 42300 34406
rect 42248 34342 42300 34348
rect 42340 34400 42392 34406
rect 42340 34342 42392 34348
rect 42156 34060 42208 34066
rect 42156 34002 42208 34008
rect 42168 33658 42196 34002
rect 42156 33652 42208 33658
rect 42076 33612 42156 33640
rect 41972 33448 42024 33454
rect 41972 33390 42024 33396
rect 42076 33114 42104 33612
rect 42156 33594 42208 33600
rect 42260 33134 42288 34342
rect 42352 34202 42380 34342
rect 42340 34196 42392 34202
rect 42340 34138 42392 34144
rect 42444 33134 42472 34478
rect 42616 33992 42668 33998
rect 42616 33934 42668 33940
rect 42064 33108 42116 33114
rect 42064 33050 42116 33056
rect 42168 33106 42288 33134
rect 42352 33106 42472 33134
rect 41604 32904 41656 32910
rect 41604 32846 41656 32852
rect 41616 32026 41644 32846
rect 42168 32842 42196 33106
rect 42156 32836 42208 32842
rect 42156 32778 42208 32784
rect 42168 32366 42196 32778
rect 42156 32360 42208 32366
rect 42156 32302 42208 32308
rect 41696 32292 41748 32298
rect 41696 32234 41748 32240
rect 41604 32020 41656 32026
rect 41604 31962 41656 31968
rect 41708 30938 41736 32234
rect 41696 30932 41748 30938
rect 41696 30874 41748 30880
rect 41708 30598 41736 30874
rect 41880 30660 41932 30666
rect 41880 30602 41932 30608
rect 41696 30592 41748 30598
rect 41696 30534 41748 30540
rect 41512 30320 41564 30326
rect 41512 30262 41564 30268
rect 41708 30258 41736 30534
rect 41696 30252 41748 30258
rect 41696 30194 41748 30200
rect 41892 30122 41920 30602
rect 41328 30116 41380 30122
rect 41328 30058 41380 30064
rect 41880 30116 41932 30122
rect 41880 30058 41932 30064
rect 41340 29850 41368 30058
rect 41328 29844 41380 29850
rect 41328 29786 41380 29792
rect 41144 29776 41196 29782
rect 41144 29718 41196 29724
rect 41052 29096 41104 29102
rect 41052 29038 41104 29044
rect 41064 28694 41092 29038
rect 41156 28966 41184 29718
rect 41236 29640 41288 29646
rect 41236 29582 41288 29588
rect 41248 29034 41276 29582
rect 41236 29028 41288 29034
rect 41236 28970 41288 28976
rect 41144 28960 41196 28966
rect 41144 28902 41196 28908
rect 41052 28688 41104 28694
rect 41052 28630 41104 28636
rect 41052 28552 41104 28558
rect 41052 28494 41104 28500
rect 41064 27538 41092 28494
rect 41156 28490 41184 28902
rect 41248 28762 41276 28970
rect 41236 28756 41288 28762
rect 41236 28698 41288 28704
rect 41144 28484 41196 28490
rect 41144 28426 41196 28432
rect 41156 28218 41184 28426
rect 41328 28416 41380 28422
rect 41328 28358 41380 28364
rect 41144 28212 41196 28218
rect 41144 28154 41196 28160
rect 41156 27946 41184 28154
rect 41340 28082 41368 28358
rect 41328 28076 41380 28082
rect 41328 28018 41380 28024
rect 41144 27940 41196 27946
rect 41144 27882 41196 27888
rect 41052 27532 41104 27538
rect 41052 27474 41104 27480
rect 40830 26846 40908 26874
rect 40774 26823 40830 26832
rect 40500 26376 40552 26382
rect 40500 26318 40552 26324
rect 40512 24274 40540 26318
rect 40500 24268 40552 24274
rect 40500 24210 40552 24216
rect 40512 23866 40540 24210
rect 40500 23860 40552 23866
rect 40500 23802 40552 23808
rect 40788 23662 40816 26823
rect 41064 26586 41092 27474
rect 41340 26994 41368 28018
rect 41880 28008 41932 28014
rect 41880 27950 41932 27956
rect 41512 27940 41564 27946
rect 41512 27882 41564 27888
rect 41524 27674 41552 27882
rect 41512 27668 41564 27674
rect 41512 27610 41564 27616
rect 41524 27130 41552 27610
rect 41512 27124 41564 27130
rect 41512 27066 41564 27072
rect 41328 26988 41380 26994
rect 41328 26930 41380 26936
rect 41052 26580 41104 26586
rect 41052 26522 41104 26528
rect 41892 26518 41920 27950
rect 42064 27328 42116 27334
rect 42064 27270 42116 27276
rect 42076 27130 42104 27270
rect 42064 27124 42116 27130
rect 42064 27066 42116 27072
rect 42076 26790 42104 27066
rect 42064 26784 42116 26790
rect 42064 26726 42116 26732
rect 42168 26518 42196 32302
rect 42248 31884 42300 31890
rect 42352 31872 42380 33106
rect 42628 32978 42656 33934
rect 43628 33856 43680 33862
rect 43628 33798 43680 33804
rect 43640 33522 43668 33798
rect 44180 33584 44232 33590
rect 44180 33526 44232 33532
rect 43628 33516 43680 33522
rect 43680 33476 43760 33504
rect 43628 33458 43680 33464
rect 43628 33108 43680 33114
rect 43628 33050 43680 33056
rect 42616 32972 42668 32978
rect 42616 32914 42668 32920
rect 42628 32570 42656 32914
rect 42984 32904 43036 32910
rect 42984 32846 43036 32852
rect 42616 32564 42668 32570
rect 42616 32506 42668 32512
rect 42300 31844 42380 31872
rect 42248 31826 42300 31832
rect 42352 31142 42380 31844
rect 42616 31816 42668 31822
rect 42616 31758 42668 31764
rect 42628 31482 42656 31758
rect 42616 31476 42668 31482
rect 42616 31418 42668 31424
rect 42996 31414 43024 32846
rect 43640 32570 43668 33050
rect 43628 32564 43680 32570
rect 43628 32506 43680 32512
rect 43628 32224 43680 32230
rect 43628 32166 43680 32172
rect 42984 31408 43036 31414
rect 42984 31350 43036 31356
rect 42340 31136 42392 31142
rect 42340 31078 42392 31084
rect 42248 30796 42300 30802
rect 42248 30738 42300 30744
rect 42260 30326 42288 30738
rect 42248 30320 42300 30326
rect 42248 30262 42300 30268
rect 42352 28626 42380 31078
rect 42996 30326 43024 31350
rect 43640 31346 43668 32166
rect 43732 32026 43760 33476
rect 44088 33380 44140 33386
rect 44088 33322 44140 33328
rect 44100 33114 44128 33322
rect 44088 33108 44140 33114
rect 44088 33050 44140 33056
rect 44100 32298 44128 33050
rect 44088 32292 44140 32298
rect 44088 32234 44140 32240
rect 43720 32020 43772 32026
rect 43720 31962 43772 31968
rect 43996 31952 44048 31958
rect 44100 31940 44128 32234
rect 44048 31912 44128 31940
rect 43996 31894 44048 31900
rect 44100 31754 44128 31912
rect 44192 31822 44220 33526
rect 44272 33380 44324 33386
rect 44272 33322 44324 33328
rect 44180 31816 44232 31822
rect 44180 31758 44232 31764
rect 44088 31748 44140 31754
rect 44088 31690 44140 31696
rect 44100 31482 44128 31690
rect 44284 31686 44312 33322
rect 45006 33144 45062 33153
rect 45006 33079 45062 33088
rect 44364 32496 44416 32502
rect 44364 32438 44416 32444
rect 44272 31680 44324 31686
rect 44272 31622 44324 31628
rect 43720 31476 43772 31482
rect 43720 31418 43772 31424
rect 44088 31476 44140 31482
rect 44088 31418 44140 31424
rect 43628 31340 43680 31346
rect 43628 31282 43680 31288
rect 43732 31210 43760 31418
rect 43720 31204 43772 31210
rect 43720 31146 43772 31152
rect 44284 30870 44312 31622
rect 43904 30864 43956 30870
rect 43904 30806 43956 30812
rect 44272 30864 44324 30870
rect 44272 30806 44324 30812
rect 43444 30728 43496 30734
rect 43444 30670 43496 30676
rect 43456 30394 43484 30670
rect 43444 30388 43496 30394
rect 43444 30330 43496 30336
rect 42984 30320 43036 30326
rect 42984 30262 43036 30268
rect 42800 30184 42852 30190
rect 42800 30126 42852 30132
rect 42432 29164 42484 29170
rect 42432 29106 42484 29112
rect 42708 29164 42760 29170
rect 42708 29106 42760 29112
rect 42444 28762 42472 29106
rect 42432 28756 42484 28762
rect 42432 28698 42484 28704
rect 42720 28694 42748 29106
rect 42708 28688 42760 28694
rect 42708 28630 42760 28636
rect 42340 28620 42392 28626
rect 42340 28562 42392 28568
rect 42812 28558 42840 30126
rect 42996 29238 43024 30262
rect 43456 29782 43484 30330
rect 43628 30252 43680 30258
rect 43628 30194 43680 30200
rect 43444 29776 43496 29782
rect 43444 29718 43496 29724
rect 43352 29640 43404 29646
rect 43352 29582 43404 29588
rect 42984 29232 43036 29238
rect 42984 29174 43036 29180
rect 43364 29170 43392 29582
rect 43352 29164 43404 29170
rect 43352 29106 43404 29112
rect 43352 28960 43404 28966
rect 43352 28902 43404 28908
rect 43260 28620 43312 28626
rect 43260 28562 43312 28568
rect 42524 28552 42576 28558
rect 42524 28494 42576 28500
rect 42800 28552 42852 28558
rect 42800 28494 42852 28500
rect 42248 28416 42300 28422
rect 42248 28358 42300 28364
rect 42260 27674 42288 28358
rect 42536 27878 42564 28494
rect 43272 28218 43300 28562
rect 43364 28490 43392 28902
rect 43640 28626 43668 30194
rect 43916 30122 43944 30806
rect 44272 30592 44324 30598
rect 44376 30580 44404 32438
rect 45020 31872 45048 33079
rect 45100 32904 45152 32910
rect 45100 32846 45152 32852
rect 45112 32570 45140 32846
rect 45100 32564 45152 32570
rect 45100 32506 45152 32512
rect 45100 31884 45152 31890
rect 45020 31844 45100 31872
rect 45100 31826 45152 31832
rect 45112 31385 45140 31826
rect 45284 31816 45336 31822
rect 45284 31758 45336 31764
rect 45098 31376 45154 31385
rect 45098 31311 45154 31320
rect 45112 31278 45140 31311
rect 44732 31272 44784 31278
rect 44732 31214 44784 31220
rect 45100 31272 45152 31278
rect 45100 31214 45152 31220
rect 44324 30552 44404 30580
rect 44272 30534 44324 30540
rect 44376 30326 44404 30552
rect 44456 30592 44508 30598
rect 44456 30534 44508 30540
rect 44468 30394 44496 30534
rect 44456 30388 44508 30394
rect 44456 30330 44508 30336
rect 44364 30320 44416 30326
rect 44364 30262 44416 30268
rect 44456 30184 44508 30190
rect 44456 30126 44508 30132
rect 43904 30116 43956 30122
rect 43904 30058 43956 30064
rect 43916 29850 43944 30058
rect 43904 29844 43956 29850
rect 43904 29786 43956 29792
rect 43916 29034 43944 29786
rect 43904 29028 43956 29034
rect 43904 28970 43956 28976
rect 43916 28762 43944 28970
rect 44364 28960 44416 28966
rect 44364 28902 44416 28908
rect 43904 28756 43956 28762
rect 43904 28698 43956 28704
rect 43628 28620 43680 28626
rect 43548 28580 43628 28608
rect 43352 28484 43404 28490
rect 43352 28426 43404 28432
rect 43260 28212 43312 28218
rect 43260 28154 43312 28160
rect 42524 27872 42576 27878
rect 42524 27814 42576 27820
rect 42248 27668 42300 27674
rect 42248 27610 42300 27616
rect 42260 26994 42288 27610
rect 42248 26988 42300 26994
rect 42248 26930 42300 26936
rect 42432 26988 42484 26994
rect 42432 26930 42484 26936
rect 41880 26512 41932 26518
rect 41880 26454 41932 26460
rect 42156 26512 42208 26518
rect 42156 26454 42208 26460
rect 41788 26376 41840 26382
rect 41788 26318 41840 26324
rect 41800 26042 41828 26318
rect 41788 26036 41840 26042
rect 41788 25978 41840 25984
rect 41892 25974 41920 26454
rect 42444 26382 42472 26930
rect 42064 26376 42116 26382
rect 42064 26318 42116 26324
rect 42432 26376 42484 26382
rect 42432 26318 42484 26324
rect 41880 25968 41932 25974
rect 41880 25910 41932 25916
rect 42076 25906 42104 26318
rect 42064 25900 42116 25906
rect 42064 25842 42116 25848
rect 41420 25764 41472 25770
rect 41420 25706 41472 25712
rect 41432 25498 41460 25706
rect 41696 25696 41748 25702
rect 41696 25638 41748 25644
rect 41420 25492 41472 25498
rect 41420 25434 41472 25440
rect 41708 25430 41736 25638
rect 41696 25424 41748 25430
rect 41696 25366 41748 25372
rect 41604 25288 41656 25294
rect 41604 25230 41656 25236
rect 40868 24744 40920 24750
rect 40868 24686 40920 24692
rect 40776 23656 40828 23662
rect 40776 23598 40828 23604
rect 40500 21616 40552 21622
rect 40500 21558 40552 21564
rect 40512 20058 40540 21558
rect 40500 20052 40552 20058
rect 40500 19994 40552 20000
rect 40512 19514 40540 19994
rect 40788 19854 40816 23598
rect 40880 19990 40908 24686
rect 41616 24410 41644 25230
rect 41708 24954 41736 25366
rect 41696 24948 41748 24954
rect 41696 24890 41748 24896
rect 41708 24614 41736 24890
rect 41696 24608 41748 24614
rect 41696 24550 41748 24556
rect 41604 24404 41656 24410
rect 41604 24346 41656 24352
rect 41708 24342 41736 24550
rect 41236 24336 41288 24342
rect 41236 24278 41288 24284
rect 41696 24336 41748 24342
rect 41696 24278 41748 24284
rect 41248 23866 41276 24278
rect 41236 23860 41288 23866
rect 41236 23802 41288 23808
rect 41248 23322 41276 23802
rect 42156 23724 42208 23730
rect 42156 23666 42208 23672
rect 41972 23588 42024 23594
rect 41972 23530 42024 23536
rect 41984 23322 42012 23530
rect 42168 23322 42196 23666
rect 41236 23316 41288 23322
rect 41236 23258 41288 23264
rect 41972 23316 42024 23322
rect 41972 23258 42024 23264
rect 42156 23316 42208 23322
rect 42156 23258 42208 23264
rect 41248 22778 41276 23258
rect 41696 23112 41748 23118
rect 41696 23054 41748 23060
rect 41708 22778 41736 23054
rect 41236 22772 41288 22778
rect 41236 22714 41288 22720
rect 41696 22772 41748 22778
rect 41696 22714 41748 22720
rect 41248 21622 41276 22714
rect 42536 22574 42564 27814
rect 43352 25832 43404 25838
rect 43352 25774 43404 25780
rect 43260 24336 43312 24342
rect 43260 24278 43312 24284
rect 42800 24268 42852 24274
rect 42800 24210 42852 24216
rect 42812 23526 42840 24210
rect 43272 23798 43300 24278
rect 43260 23792 43312 23798
rect 43260 23734 43312 23740
rect 42800 23520 42852 23526
rect 42800 23462 42852 23468
rect 42812 23186 42840 23462
rect 42800 23180 42852 23186
rect 42800 23122 42852 23128
rect 42524 22568 42576 22574
rect 42524 22510 42576 22516
rect 41420 22092 41472 22098
rect 41420 22034 41472 22040
rect 41432 21690 41460 22034
rect 41512 22024 41564 22030
rect 41512 21966 41564 21972
rect 42156 22024 42208 22030
rect 42156 21966 42208 21972
rect 41420 21684 41472 21690
rect 41420 21626 41472 21632
rect 41236 21616 41288 21622
rect 41236 21558 41288 21564
rect 41524 20942 41552 21966
rect 42168 21554 42196 21966
rect 42248 21956 42300 21962
rect 42248 21898 42300 21904
rect 43260 21956 43312 21962
rect 43260 21898 43312 21904
rect 42156 21548 42208 21554
rect 42156 21490 42208 21496
rect 42260 21146 42288 21898
rect 42984 21344 43036 21350
rect 42984 21286 43036 21292
rect 42248 21140 42300 21146
rect 42248 21082 42300 21088
rect 41604 21072 41656 21078
rect 41604 21014 41656 21020
rect 41144 20936 41196 20942
rect 41144 20878 41196 20884
rect 41512 20936 41564 20942
rect 41512 20878 41564 20884
rect 41156 20262 41184 20878
rect 41236 20868 41288 20874
rect 41236 20810 41288 20816
rect 41052 20256 41104 20262
rect 41052 20198 41104 20204
rect 41144 20256 41196 20262
rect 41144 20198 41196 20204
rect 40868 19984 40920 19990
rect 40868 19926 40920 19932
rect 41064 19922 41092 20198
rect 41052 19916 41104 19922
rect 41052 19858 41104 19864
rect 40776 19848 40828 19854
rect 40776 19790 40828 19796
rect 40500 19508 40552 19514
rect 40500 19450 40552 19456
rect 40592 18760 40644 18766
rect 40592 18702 40644 18708
rect 40604 18426 40632 18702
rect 40592 18420 40644 18426
rect 40592 18362 40644 18368
rect 40684 18148 40736 18154
rect 40684 18090 40736 18096
rect 40696 17746 40724 18090
rect 40788 18057 40816 19790
rect 40958 19680 41014 19689
rect 40958 19615 41014 19624
rect 40774 18048 40830 18057
rect 40774 17983 40830 17992
rect 40684 17740 40736 17746
rect 40684 17682 40736 17688
rect 40592 17604 40644 17610
rect 40592 17546 40644 17552
rect 40604 17066 40632 17546
rect 40592 17060 40644 17066
rect 40592 17002 40644 17008
rect 40604 16794 40632 17002
rect 40592 16788 40644 16794
rect 40592 16730 40644 16736
rect 40500 16584 40552 16590
rect 40500 16526 40552 16532
rect 40512 16114 40540 16526
rect 40500 16108 40552 16114
rect 40500 16050 40552 16056
rect 40498 16008 40554 16017
rect 40498 15943 40554 15952
rect 40512 15570 40540 15943
rect 40500 15564 40552 15570
rect 40500 15506 40552 15512
rect 40512 15162 40540 15506
rect 40500 15156 40552 15162
rect 40500 15098 40552 15104
rect 40408 13184 40460 13190
rect 40408 13126 40460 13132
rect 40224 12980 40276 12986
rect 40224 12922 40276 12928
rect 40512 11354 40540 15098
rect 40788 15094 40816 17983
rect 40972 15094 41000 19615
rect 41156 19514 41184 20198
rect 41144 19508 41196 19514
rect 41144 19450 41196 19456
rect 41248 18714 41276 20810
rect 41616 20330 41644 21014
rect 41972 20868 42024 20874
rect 41972 20810 42024 20816
rect 41984 20466 42012 20810
rect 41972 20460 42024 20466
rect 41972 20402 42024 20408
rect 41328 20324 41380 20330
rect 41328 20266 41380 20272
rect 41604 20324 41656 20330
rect 41604 20266 41656 20272
rect 41340 19718 41368 20266
rect 41616 19922 41644 20266
rect 41604 19916 41656 19922
rect 41604 19858 41656 19864
rect 41512 19780 41564 19786
rect 41512 19722 41564 19728
rect 41328 19712 41380 19718
rect 41328 19654 41380 19660
rect 41340 18970 41368 19654
rect 41328 18964 41380 18970
rect 41328 18906 41380 18912
rect 41524 18902 41552 19722
rect 41616 19174 41644 19858
rect 41788 19712 41840 19718
rect 41788 19654 41840 19660
rect 41800 19378 41828 19654
rect 41788 19372 41840 19378
rect 41788 19314 41840 19320
rect 41604 19168 41656 19174
rect 41604 19110 41656 19116
rect 41616 18902 41644 19110
rect 41512 18896 41564 18902
rect 41512 18838 41564 18844
rect 41604 18896 41656 18902
rect 41604 18838 41656 18844
rect 41156 18686 41276 18714
rect 41052 17672 41104 17678
rect 41052 17614 41104 17620
rect 41064 17202 41092 17614
rect 41052 17196 41104 17202
rect 41052 17138 41104 17144
rect 41156 16590 41184 18686
rect 41524 18426 41552 18838
rect 41512 18420 41564 18426
rect 41512 18362 41564 18368
rect 41616 18358 41644 18838
rect 41604 18352 41656 18358
rect 41604 18294 41656 18300
rect 41696 18352 41748 18358
rect 41696 18294 41748 18300
rect 41236 18148 41288 18154
rect 41236 18090 41288 18096
rect 41248 17270 41276 18090
rect 41512 17808 41564 17814
rect 41512 17750 41564 17756
rect 41524 17338 41552 17750
rect 41512 17332 41564 17338
rect 41512 17274 41564 17280
rect 41236 17264 41288 17270
rect 41288 17224 41368 17252
rect 41236 17206 41288 17212
rect 41236 16720 41288 16726
rect 41236 16662 41288 16668
rect 41144 16584 41196 16590
rect 41144 16526 41196 16532
rect 41052 16516 41104 16522
rect 41052 16458 41104 16464
rect 41064 16182 41092 16458
rect 41052 16176 41104 16182
rect 41052 16118 41104 16124
rect 41052 15972 41104 15978
rect 41052 15914 41104 15920
rect 40776 15088 40828 15094
rect 40776 15030 40828 15036
rect 40960 15088 41012 15094
rect 40960 15030 41012 15036
rect 41064 14550 41092 15914
rect 41156 15706 41184 16526
rect 41248 16250 41276 16662
rect 41340 16590 41368 17224
rect 41328 16584 41380 16590
rect 41328 16526 41380 16532
rect 41236 16244 41288 16250
rect 41236 16186 41288 16192
rect 41144 15700 41196 15706
rect 41144 15642 41196 15648
rect 41144 15496 41196 15502
rect 41144 15438 41196 15444
rect 41052 14544 41104 14550
rect 41052 14486 41104 14492
rect 41064 13938 41092 14486
rect 41156 14482 41184 15438
rect 41340 15094 41368 16526
rect 41328 15088 41380 15094
rect 41328 15030 41380 15036
rect 41236 14952 41288 14958
rect 41236 14894 41288 14900
rect 41144 14476 41196 14482
rect 41144 14418 41196 14424
rect 41156 14074 41184 14418
rect 41144 14068 41196 14074
rect 41144 14010 41196 14016
rect 41052 13932 41104 13938
rect 41052 13874 41104 13880
rect 41248 13814 41276 14894
rect 41340 14006 41368 15030
rect 41708 14890 41736 18294
rect 41984 17610 42012 20402
rect 42892 20392 42944 20398
rect 42892 20334 42944 20340
rect 42708 19916 42760 19922
rect 42708 19858 42760 19864
rect 42524 19848 42576 19854
rect 42524 19790 42576 19796
rect 42248 19780 42300 19786
rect 42248 19722 42300 19728
rect 42260 19689 42288 19722
rect 42246 19680 42302 19689
rect 42246 19615 42302 19624
rect 42536 19174 42564 19790
rect 42720 19514 42748 19858
rect 42708 19508 42760 19514
rect 42708 19450 42760 19456
rect 42524 19168 42576 19174
rect 42524 19110 42576 19116
rect 41972 17604 42024 17610
rect 41972 17546 42024 17552
rect 42432 17128 42484 17134
rect 42432 17070 42484 17076
rect 42444 16794 42472 17070
rect 42432 16788 42484 16794
rect 42432 16730 42484 16736
rect 42444 15910 42472 16730
rect 42708 16040 42760 16046
rect 42708 15982 42760 15988
rect 42432 15904 42484 15910
rect 42432 15846 42484 15852
rect 42720 15570 42748 15982
rect 42708 15564 42760 15570
rect 42708 15506 42760 15512
rect 41880 15360 41932 15366
rect 41880 15302 41932 15308
rect 41892 14890 41920 15302
rect 41696 14884 41748 14890
rect 41696 14826 41748 14832
rect 41880 14884 41932 14890
rect 41880 14826 41932 14832
rect 41892 14618 41920 14826
rect 41880 14612 41932 14618
rect 41880 14554 41932 14560
rect 41328 14000 41380 14006
rect 41328 13942 41380 13948
rect 41604 13932 41656 13938
rect 41604 13874 41656 13880
rect 41248 13786 41368 13814
rect 40868 12368 40920 12374
rect 40868 12310 40920 12316
rect 40880 11898 40908 12310
rect 41144 12232 41196 12238
rect 41144 12174 41196 12180
rect 40868 11892 40920 11898
rect 40868 11834 40920 11840
rect 41156 11558 41184 12174
rect 41144 11552 41196 11558
rect 41144 11494 41196 11500
rect 40500 11348 40552 11354
rect 40500 11290 40552 11296
rect 41156 11286 41184 11494
rect 41144 11280 41196 11286
rect 41144 11222 41196 11228
rect 40040 128 40092 134
rect 40040 70 40092 76
rect 40958 128 41014 480
rect 41340 134 41368 13786
rect 41616 12374 41644 13874
rect 41696 12640 41748 12646
rect 41696 12582 41748 12588
rect 41708 12442 41736 12582
rect 41696 12436 41748 12442
rect 41696 12378 41748 12384
rect 41604 12368 41656 12374
rect 42904 12345 42932 20334
rect 42996 20058 43024 21286
rect 43272 20942 43300 21898
rect 43260 20936 43312 20942
rect 43260 20878 43312 20884
rect 42984 20052 43036 20058
rect 42984 19994 43036 20000
rect 43260 19712 43312 19718
rect 43260 19654 43312 19660
rect 43272 19145 43300 19654
rect 43258 19136 43314 19145
rect 43258 19071 43314 19080
rect 43076 18624 43128 18630
rect 43076 18566 43128 18572
rect 43088 18290 43116 18566
rect 43258 18320 43314 18329
rect 43076 18284 43128 18290
rect 43258 18255 43314 18264
rect 43076 18226 43128 18232
rect 43272 17338 43300 18255
rect 43260 17332 43312 17338
rect 43260 17274 43312 17280
rect 43364 15570 43392 25774
rect 43548 24857 43576 28580
rect 43628 28562 43680 28568
rect 43720 28416 43772 28422
rect 43720 28358 43772 28364
rect 43732 28082 43760 28358
rect 43720 28076 43772 28082
rect 43720 28018 43772 28024
rect 43812 28076 43864 28082
rect 43812 28018 43864 28024
rect 43628 27872 43680 27878
rect 43628 27814 43680 27820
rect 43640 27606 43668 27814
rect 43628 27600 43680 27606
rect 43628 27542 43680 27548
rect 43640 27334 43668 27542
rect 43824 27402 43852 28018
rect 43904 27464 43956 27470
rect 43904 27406 43956 27412
rect 43812 27396 43864 27402
rect 43812 27338 43864 27344
rect 43628 27328 43680 27334
rect 43628 27270 43680 27276
rect 43640 26790 43668 27270
rect 43628 26784 43680 26790
rect 43628 26726 43680 26732
rect 43640 25430 43668 26726
rect 43720 26444 43772 26450
rect 43720 26386 43772 26392
rect 43732 26042 43760 26386
rect 43720 26036 43772 26042
rect 43720 25978 43772 25984
rect 43824 25922 43852 27338
rect 43916 26586 43944 27406
rect 44272 26988 44324 26994
rect 44272 26930 44324 26936
rect 44284 26858 44312 26930
rect 44180 26852 44232 26858
rect 44180 26794 44232 26800
rect 44272 26852 44324 26858
rect 44272 26794 44324 26800
rect 44192 26586 44220 26794
rect 43904 26580 43956 26586
rect 43904 26522 43956 26528
rect 44180 26580 44232 26586
rect 44180 26522 44232 26528
rect 44284 26518 44312 26794
rect 44272 26512 44324 26518
rect 44272 26454 44324 26460
rect 43732 25894 43852 25922
rect 43996 25900 44048 25906
rect 43628 25424 43680 25430
rect 43628 25366 43680 25372
rect 43640 24954 43668 25366
rect 43732 25294 43760 25894
rect 43996 25842 44048 25848
rect 44088 25900 44140 25906
rect 44088 25842 44140 25848
rect 43812 25696 43864 25702
rect 43812 25638 43864 25644
rect 43720 25288 43772 25294
rect 43720 25230 43772 25236
rect 43628 24948 43680 24954
rect 43628 24890 43680 24896
rect 43534 24848 43590 24857
rect 43534 24783 43590 24792
rect 43444 24200 43496 24206
rect 43444 24142 43496 24148
rect 43456 23866 43484 24142
rect 43444 23860 43496 23866
rect 43444 23802 43496 23808
rect 43444 22704 43496 22710
rect 43824 22681 43852 25638
rect 44008 24954 44036 25842
rect 44100 25226 44128 25842
rect 44284 25770 44312 26454
rect 44376 26450 44404 28902
rect 44364 26444 44416 26450
rect 44364 26386 44416 26392
rect 44272 25764 44324 25770
rect 44272 25706 44324 25712
rect 44376 25702 44404 26386
rect 44364 25696 44416 25702
rect 44364 25638 44416 25644
rect 44088 25220 44140 25226
rect 44088 25162 44140 25168
rect 43996 24948 44048 24954
rect 43996 24890 44048 24896
rect 43902 24848 43958 24857
rect 43902 24783 43958 24792
rect 43444 22646 43496 22652
rect 43810 22672 43866 22681
rect 43456 22030 43484 22646
rect 43810 22607 43866 22616
rect 43824 22574 43852 22607
rect 43812 22568 43864 22574
rect 43812 22510 43864 22516
rect 43720 22432 43772 22438
rect 43720 22374 43772 22380
rect 43628 22160 43680 22166
rect 43628 22102 43680 22108
rect 43444 22024 43496 22030
rect 43444 21966 43496 21972
rect 43456 21690 43484 21966
rect 43444 21684 43496 21690
rect 43444 21626 43496 21632
rect 43640 21350 43668 22102
rect 43732 21554 43760 22374
rect 43720 21548 43772 21554
rect 43720 21490 43772 21496
rect 43628 21344 43680 21350
rect 43628 21286 43680 21292
rect 43640 21078 43668 21286
rect 43732 21146 43760 21490
rect 43720 21140 43772 21146
rect 43720 21082 43772 21088
rect 43628 21072 43680 21078
rect 43628 21014 43680 21020
rect 43444 20936 43496 20942
rect 43444 20878 43496 20884
rect 43456 20602 43484 20878
rect 43444 20596 43496 20602
rect 43444 20538 43496 20544
rect 43444 20324 43496 20330
rect 43444 20266 43496 20272
rect 43456 19990 43484 20266
rect 43640 20262 43668 21014
rect 43916 20534 43944 24783
rect 44100 24206 44128 25162
rect 44468 24954 44496 30126
rect 44640 28620 44692 28626
rect 44640 28562 44692 28568
rect 44652 28218 44680 28562
rect 44640 28212 44692 28218
rect 44640 28154 44692 28160
rect 44744 26042 44772 31214
rect 45008 30864 45060 30870
rect 45008 30806 45060 30812
rect 45100 30864 45152 30870
rect 45100 30806 45152 30812
rect 45020 30326 45048 30806
rect 45008 30320 45060 30326
rect 45008 30262 45060 30268
rect 45112 30258 45140 30806
rect 45296 30734 45324 31758
rect 45284 30728 45336 30734
rect 45284 30670 45336 30676
rect 46572 30388 46624 30394
rect 46572 30330 46624 30336
rect 45100 30252 45152 30258
rect 45100 30194 45152 30200
rect 45112 29850 45140 30194
rect 46584 30190 46612 30330
rect 46572 30184 46624 30190
rect 46572 30126 46624 30132
rect 45100 29844 45152 29850
rect 45100 29786 45152 29792
rect 45100 29708 45152 29714
rect 45100 29650 45152 29656
rect 44824 29504 44876 29510
rect 44824 29446 44876 29452
rect 44836 29306 44864 29446
rect 44824 29300 44876 29306
rect 44824 29242 44876 29248
rect 45112 28966 45140 29650
rect 45100 28960 45152 28966
rect 45100 28902 45152 28908
rect 45468 28416 45520 28422
rect 45468 28358 45520 28364
rect 45480 27606 45508 28358
rect 45468 27600 45520 27606
rect 45468 27542 45520 27548
rect 45560 27600 45612 27606
rect 45560 27542 45612 27548
rect 44824 27464 44876 27470
rect 44824 27406 44876 27412
rect 44836 26858 44864 27406
rect 45480 27130 45508 27542
rect 45468 27124 45520 27130
rect 45468 27066 45520 27072
rect 45572 26994 45600 27542
rect 45560 26988 45612 26994
rect 45560 26930 45612 26936
rect 44824 26852 44876 26858
rect 44824 26794 44876 26800
rect 44732 26036 44784 26042
rect 44732 25978 44784 25984
rect 44640 25288 44692 25294
rect 44640 25230 44692 25236
rect 44652 24954 44680 25230
rect 44456 24948 44508 24954
rect 44456 24890 44508 24896
rect 44640 24948 44692 24954
rect 44640 24890 44692 24896
rect 44836 24886 44864 26794
rect 44824 24880 44876 24886
rect 44824 24822 44876 24828
rect 44272 24744 44324 24750
rect 44272 24686 44324 24692
rect 44088 24200 44140 24206
rect 44088 24142 44140 24148
rect 44100 23322 44128 24142
rect 44088 23316 44140 23322
rect 44088 23258 44140 23264
rect 44180 21548 44232 21554
rect 44180 21490 44232 21496
rect 43904 20528 43956 20534
rect 43904 20470 43956 20476
rect 43812 20392 43864 20398
rect 43812 20334 43864 20340
rect 43628 20256 43680 20262
rect 43628 20198 43680 20204
rect 43640 19990 43668 20198
rect 43444 19984 43496 19990
rect 43444 19926 43496 19932
rect 43628 19984 43680 19990
rect 43628 19926 43680 19932
rect 43456 19514 43484 19926
rect 43720 19848 43772 19854
rect 43720 19790 43772 19796
rect 43444 19508 43496 19514
rect 43444 19450 43496 19456
rect 43732 19446 43760 19790
rect 43824 19786 43852 20334
rect 44088 19984 44140 19990
rect 44088 19926 44140 19932
rect 43812 19780 43864 19786
rect 43812 19722 43864 19728
rect 44100 19514 44128 19926
rect 44088 19508 44140 19514
rect 44088 19450 44140 19456
rect 43720 19440 43772 19446
rect 43720 19382 43772 19388
rect 43536 18148 43588 18154
rect 43536 18090 43588 18096
rect 43548 17814 43576 18090
rect 43536 17808 43588 17814
rect 43536 17750 43588 17756
rect 43548 17338 43576 17750
rect 43536 17332 43588 17338
rect 43536 17274 43588 17280
rect 43548 16726 43576 17274
rect 43732 17202 43760 19382
rect 43996 18828 44048 18834
rect 43996 18770 44048 18776
rect 44008 18426 44036 18770
rect 44192 18766 44220 21490
rect 44284 20602 44312 24686
rect 44272 20596 44324 20602
rect 44272 20538 44324 20544
rect 44284 20398 44312 20538
rect 44272 20392 44324 20398
rect 44272 20334 44324 20340
rect 44916 19916 44968 19922
rect 44916 19858 44968 19864
rect 44928 19514 44956 19858
rect 44916 19508 44968 19514
rect 44916 19450 44968 19456
rect 44180 18760 44232 18766
rect 44180 18702 44232 18708
rect 43996 18420 44048 18426
rect 43996 18362 44048 18368
rect 44192 18290 44220 18702
rect 44180 18284 44232 18290
rect 44180 18226 44232 18232
rect 45192 17740 45244 17746
rect 45192 17682 45244 17688
rect 45204 17338 45232 17682
rect 44364 17332 44416 17338
rect 44364 17274 44416 17280
rect 45192 17332 45244 17338
rect 45192 17274 45244 17280
rect 43720 17196 43772 17202
rect 43720 17138 43772 17144
rect 43536 16720 43588 16726
rect 43536 16662 43588 16668
rect 43444 16584 43496 16590
rect 43444 16526 43496 16532
rect 43456 15978 43484 16526
rect 43548 16250 43576 16662
rect 43536 16244 43588 16250
rect 43536 16186 43588 16192
rect 43444 15972 43496 15978
rect 43444 15914 43496 15920
rect 43456 15706 43484 15914
rect 43444 15700 43496 15706
rect 43444 15642 43496 15648
rect 43352 15564 43404 15570
rect 43352 15506 43404 15512
rect 43364 15162 43392 15506
rect 43352 15156 43404 15162
rect 43352 15098 43404 15104
rect 43364 14521 43392 15098
rect 43732 15094 43760 17138
rect 44376 17066 44404 17274
rect 45204 17241 45232 17274
rect 45190 17232 45246 17241
rect 45190 17167 45246 17176
rect 44364 17060 44416 17066
rect 44364 17002 44416 17008
rect 43812 16992 43864 16998
rect 43812 16934 43864 16940
rect 43824 16114 43852 16934
rect 43812 16108 43864 16114
rect 43812 16050 43864 16056
rect 43720 15088 43772 15094
rect 43720 15030 43772 15036
rect 43350 14512 43406 14521
rect 43350 14447 43406 14456
rect 41604 12310 41656 12316
rect 42890 12336 42946 12345
rect 42890 12271 42946 12280
rect 44178 12336 44234 12345
rect 44178 12271 44234 12280
rect 40958 76 40960 128
rect 41012 76 41014 128
rect 40958 0 41014 76
rect 41328 128 41380 134
rect 41328 70 41380 76
rect 44192 82 44220 12271
rect 44546 82 44602 480
rect 44192 54 44602 82
rect 44546 0 44602 54
rect 48134 128 48190 480
rect 48134 76 48136 128
rect 48188 76 48190 128
rect 48134 0 48190 76
<< via2 >>
rect 4220 46810 4276 46812
rect 4300 46810 4356 46812
rect 4380 46810 4436 46812
rect 4460 46810 4516 46812
rect 4220 46758 4246 46810
rect 4246 46758 4276 46810
rect 4300 46758 4310 46810
rect 4310 46758 4356 46810
rect 4380 46758 4426 46810
rect 4426 46758 4436 46810
rect 4460 46758 4490 46810
rect 4490 46758 4516 46810
rect 4220 46756 4276 46758
rect 4300 46756 4356 46758
rect 4380 46756 4436 46758
rect 4460 46756 4516 46758
rect 4220 45722 4276 45724
rect 4300 45722 4356 45724
rect 4380 45722 4436 45724
rect 4460 45722 4516 45724
rect 4220 45670 4246 45722
rect 4246 45670 4276 45722
rect 4300 45670 4310 45722
rect 4310 45670 4356 45722
rect 4380 45670 4426 45722
rect 4426 45670 4436 45722
rect 4460 45670 4490 45722
rect 4490 45670 4516 45722
rect 4220 45668 4276 45670
rect 4300 45668 4356 45670
rect 4380 45668 4436 45670
rect 4460 45668 4516 45670
rect 4220 44634 4276 44636
rect 4300 44634 4356 44636
rect 4380 44634 4436 44636
rect 4460 44634 4516 44636
rect 4220 44582 4246 44634
rect 4246 44582 4276 44634
rect 4300 44582 4310 44634
rect 4310 44582 4356 44634
rect 4380 44582 4426 44634
rect 4426 44582 4436 44634
rect 4460 44582 4490 44634
rect 4490 44582 4516 44634
rect 4220 44580 4276 44582
rect 4300 44580 4356 44582
rect 4380 44580 4436 44582
rect 4460 44580 4516 44582
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4246 43546
rect 4246 43494 4276 43546
rect 4300 43494 4310 43546
rect 4310 43494 4356 43546
rect 4380 43494 4426 43546
rect 4426 43494 4436 43546
rect 4460 43494 4490 43546
rect 4490 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4246 42458
rect 4246 42406 4276 42458
rect 4300 42406 4310 42458
rect 4310 42406 4356 42458
rect 4380 42406 4426 42458
rect 4426 42406 4436 42458
rect 4460 42406 4490 42458
rect 4490 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4246 41370
rect 4246 41318 4276 41370
rect 4300 41318 4310 41370
rect 4310 41318 4356 41370
rect 4380 41318 4426 41370
rect 4426 41318 4436 41370
rect 4460 41318 4490 41370
rect 4490 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4246 40282
rect 4246 40230 4276 40282
rect 4300 40230 4310 40282
rect 4310 40230 4356 40282
rect 4380 40230 4426 40282
rect 4426 40230 4436 40282
rect 4460 40230 4490 40282
rect 4490 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 11426 41520 11482 41576
rect 11426 39888 11482 39944
rect 9954 31456 10010 31512
rect 8298 30912 8354 30968
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 9862 27512 9918 27568
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 9402 25200 9458 25256
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 2778 23024 2834 23080
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 11334 38664 11390 38720
rect 11886 37304 11942 37360
rect 11242 36624 11298 36680
rect 10414 31184 10470 31240
rect 10506 31048 10562 31104
rect 11058 25744 11114 25800
rect 9402 18692 9458 18728
rect 9402 18672 9404 18692
rect 9404 18672 9456 18692
rect 9456 18672 9458 18692
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 10138 13640 10194 13696
rect 10322 11192 10378 11248
rect 9678 10920 9734 10976
rect 10506 22616 10562 22672
rect 13358 39888 13414 39944
rect 13634 39208 13690 39264
rect 13082 31456 13138 31512
rect 14278 39208 14334 39264
rect 14554 38664 14610 38720
rect 14094 34484 14096 34504
rect 14096 34484 14148 34504
rect 14148 34484 14150 34504
rect 14094 34448 14150 34484
rect 11886 25880 11942 25936
rect 9770 9968 9826 10024
rect 10414 9968 10470 10024
rect 10782 13640 10838 13696
rect 14738 37168 14794 37224
rect 14554 33260 14556 33280
rect 14556 33260 14608 33280
rect 14608 33260 14610 33280
rect 14554 33224 14610 33260
rect 16026 36080 16082 36136
rect 15566 33224 15622 33280
rect 14278 28192 14334 28248
rect 14186 22072 14242 22128
rect 13634 19216 13690 19272
rect 14094 19216 14150 19272
rect 12714 11736 12770 11792
rect 12898 11056 12954 11112
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 10506 4800 10562 4856
rect 12438 5208 12494 5264
rect 15382 27512 15438 27568
rect 19580 47354 19636 47356
rect 19660 47354 19716 47356
rect 19740 47354 19796 47356
rect 19820 47354 19876 47356
rect 19580 47302 19606 47354
rect 19606 47302 19636 47354
rect 19660 47302 19670 47354
rect 19670 47302 19716 47354
rect 19740 47302 19786 47354
rect 19786 47302 19796 47354
rect 19820 47302 19850 47354
rect 19850 47302 19876 47354
rect 19580 47300 19636 47302
rect 19660 47300 19716 47302
rect 19740 47300 19796 47302
rect 19820 47300 19876 47302
rect 19580 46266 19636 46268
rect 19660 46266 19716 46268
rect 19740 46266 19796 46268
rect 19820 46266 19876 46268
rect 19580 46214 19606 46266
rect 19606 46214 19636 46266
rect 19660 46214 19670 46266
rect 19670 46214 19716 46266
rect 19740 46214 19786 46266
rect 19786 46214 19796 46266
rect 19820 46214 19850 46266
rect 19850 46214 19876 46266
rect 19580 46212 19636 46214
rect 19660 46212 19716 46214
rect 19740 46212 19796 46214
rect 19820 46212 19876 46214
rect 19580 45178 19636 45180
rect 19660 45178 19716 45180
rect 19740 45178 19796 45180
rect 19820 45178 19876 45180
rect 19580 45126 19606 45178
rect 19606 45126 19636 45178
rect 19660 45126 19670 45178
rect 19670 45126 19716 45178
rect 19740 45126 19786 45178
rect 19786 45126 19796 45178
rect 19820 45126 19850 45178
rect 19850 45126 19876 45178
rect 19580 45124 19636 45126
rect 19660 45124 19716 45126
rect 19740 45124 19796 45126
rect 19820 45124 19876 45126
rect 19580 44090 19636 44092
rect 19660 44090 19716 44092
rect 19740 44090 19796 44092
rect 19820 44090 19876 44092
rect 19580 44038 19606 44090
rect 19606 44038 19636 44090
rect 19660 44038 19670 44090
rect 19670 44038 19716 44090
rect 19740 44038 19786 44090
rect 19786 44038 19796 44090
rect 19820 44038 19850 44090
rect 19850 44038 19876 44090
rect 19580 44036 19636 44038
rect 19660 44036 19716 44038
rect 19740 44036 19796 44038
rect 19820 44036 19876 44038
rect 19580 43002 19636 43004
rect 19660 43002 19716 43004
rect 19740 43002 19796 43004
rect 19820 43002 19876 43004
rect 19580 42950 19606 43002
rect 19606 42950 19636 43002
rect 19660 42950 19670 43002
rect 19670 42950 19716 43002
rect 19740 42950 19786 43002
rect 19786 42950 19796 43002
rect 19820 42950 19850 43002
rect 19850 42950 19876 43002
rect 19580 42948 19636 42950
rect 19660 42948 19716 42950
rect 19740 42948 19796 42950
rect 19820 42948 19876 42950
rect 19580 41914 19636 41916
rect 19660 41914 19716 41916
rect 19740 41914 19796 41916
rect 19820 41914 19876 41916
rect 19580 41862 19606 41914
rect 19606 41862 19636 41914
rect 19660 41862 19670 41914
rect 19670 41862 19716 41914
rect 19740 41862 19786 41914
rect 19786 41862 19796 41914
rect 19820 41862 19850 41914
rect 19850 41862 19876 41914
rect 19580 41860 19636 41862
rect 19660 41860 19716 41862
rect 19740 41860 19796 41862
rect 19820 41860 19876 41862
rect 19062 41676 19118 41712
rect 19062 41656 19064 41676
rect 19064 41656 19116 41676
rect 19116 41656 19118 41676
rect 18786 41012 18788 41032
rect 18788 41012 18840 41032
rect 18840 41012 18842 41032
rect 17222 36080 17278 36136
rect 15750 28192 15806 28248
rect 16394 22616 16450 22672
rect 15106 18264 15162 18320
rect 18418 38412 18474 38448
rect 18418 38392 18420 38412
rect 18420 38392 18472 38412
rect 18472 38392 18474 38412
rect 18786 40976 18842 41012
rect 19580 40826 19636 40828
rect 19660 40826 19716 40828
rect 19740 40826 19796 40828
rect 19820 40826 19876 40828
rect 19580 40774 19606 40826
rect 19606 40774 19636 40826
rect 19660 40774 19670 40826
rect 19670 40774 19716 40826
rect 19740 40774 19786 40826
rect 19786 40774 19796 40826
rect 19820 40774 19850 40826
rect 19850 40774 19876 40826
rect 19580 40772 19636 40774
rect 19660 40772 19716 40774
rect 19740 40772 19796 40774
rect 19820 40772 19876 40774
rect 19580 39738 19636 39740
rect 19660 39738 19716 39740
rect 19740 39738 19796 39740
rect 19820 39738 19876 39740
rect 19580 39686 19606 39738
rect 19606 39686 19636 39738
rect 19660 39686 19670 39738
rect 19670 39686 19716 39738
rect 19740 39686 19786 39738
rect 19786 39686 19796 39738
rect 19820 39686 19850 39738
rect 19850 39686 19876 39738
rect 19580 39684 19636 39686
rect 19660 39684 19716 39686
rect 19740 39684 19796 39686
rect 19820 39684 19876 39686
rect 18786 39480 18842 39536
rect 19246 37168 19302 37224
rect 19338 37032 19394 37088
rect 17406 26016 17462 26072
rect 17774 24656 17830 24712
rect 18050 24248 18106 24304
rect 17314 22072 17370 22128
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 11426 2080 11482 2136
rect 11886 1808 11942 1864
rect 11058 1672 11114 1728
rect 14186 4140 14242 4176
rect 14186 4120 14188 4140
rect 14188 4120 14240 4140
rect 14240 4120 14242 4140
rect 15106 4120 15162 4176
rect 17774 18672 17830 18728
rect 18694 30912 18750 30968
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 19706 37304 19762 37360
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 19062 31048 19118 31104
rect 22650 39208 22706 39264
rect 21730 36236 21786 36272
rect 21730 36216 21732 36236
rect 21732 36216 21784 36236
rect 21784 36216 21786 36236
rect 21086 34448 21142 34504
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19982 30912 20038 30968
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 18602 28620 18658 28656
rect 18602 28600 18604 28620
rect 18604 28600 18656 28620
rect 18656 28600 18658 28620
rect 18418 23704 18474 23760
rect 18142 22888 18198 22944
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 18786 22480 18842 22536
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19246 22752 19302 22808
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 20810 31456 20866 31512
rect 20626 31184 20682 31240
rect 22282 32272 22338 32328
rect 21362 30232 21418 30288
rect 20902 29164 20958 29200
rect 20902 29144 20904 29164
rect 20904 29144 20956 29164
rect 20956 29144 20958 29164
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 17222 5208 17278 5264
rect 18050 11600 18106 11656
rect 18234 13232 18290 13288
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 18694 13388 18750 13424
rect 18694 13368 18696 13388
rect 18696 13368 18748 13388
rect 18748 13368 18750 13388
rect 18142 8880 18198 8936
rect 19338 18808 19394 18864
rect 19246 15952 19302 16008
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 19522 18808 19578 18864
rect 20626 23704 20682 23760
rect 20534 22888 20590 22944
rect 20258 22752 20314 22808
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 21086 25880 21142 25936
rect 34940 46810 34996 46812
rect 35020 46810 35076 46812
rect 35100 46810 35156 46812
rect 35180 46810 35236 46812
rect 34940 46758 34966 46810
rect 34966 46758 34996 46810
rect 35020 46758 35030 46810
rect 35030 46758 35076 46810
rect 35100 46758 35146 46810
rect 35146 46758 35156 46810
rect 35180 46758 35210 46810
rect 35210 46758 35236 46810
rect 34940 46756 34996 46758
rect 35020 46756 35076 46758
rect 35100 46756 35156 46758
rect 35180 46756 35236 46758
rect 34940 45722 34996 45724
rect 35020 45722 35076 45724
rect 35100 45722 35156 45724
rect 35180 45722 35236 45724
rect 34940 45670 34966 45722
rect 34966 45670 34996 45722
rect 35020 45670 35030 45722
rect 35030 45670 35076 45722
rect 35100 45670 35146 45722
rect 35146 45670 35156 45722
rect 35180 45670 35210 45722
rect 35210 45670 35236 45722
rect 34940 45668 34996 45670
rect 35020 45668 35076 45670
rect 35100 45668 35156 45670
rect 35180 45668 35236 45670
rect 34940 44634 34996 44636
rect 35020 44634 35076 44636
rect 35100 44634 35156 44636
rect 35180 44634 35236 44636
rect 34940 44582 34966 44634
rect 34966 44582 34996 44634
rect 35020 44582 35030 44634
rect 35030 44582 35076 44634
rect 35100 44582 35146 44634
rect 35146 44582 35156 44634
rect 35180 44582 35210 44634
rect 35210 44582 35236 44634
rect 34940 44580 34996 44582
rect 35020 44580 35076 44582
rect 35100 44580 35156 44582
rect 35180 44580 35236 44582
rect 34940 43546 34996 43548
rect 35020 43546 35076 43548
rect 35100 43546 35156 43548
rect 35180 43546 35236 43548
rect 34940 43494 34966 43546
rect 34966 43494 34996 43546
rect 35020 43494 35030 43546
rect 35030 43494 35076 43546
rect 35100 43494 35146 43546
rect 35146 43494 35156 43546
rect 35180 43494 35210 43546
rect 35210 43494 35236 43546
rect 34940 43492 34996 43494
rect 35020 43492 35076 43494
rect 35100 43492 35156 43494
rect 35180 43492 35236 43494
rect 34940 42458 34996 42460
rect 35020 42458 35076 42460
rect 35100 42458 35156 42460
rect 35180 42458 35236 42460
rect 34940 42406 34966 42458
rect 34966 42406 34996 42458
rect 35020 42406 35030 42458
rect 35030 42406 35076 42458
rect 35100 42406 35146 42458
rect 35146 42406 35156 42458
rect 35180 42406 35210 42458
rect 35210 42406 35236 42458
rect 34940 42404 34996 42406
rect 35020 42404 35076 42406
rect 35100 42404 35156 42406
rect 35180 42404 35236 42406
rect 24858 41656 24914 41712
rect 23202 39888 23258 39944
rect 25962 40996 26018 41032
rect 25962 40976 25964 40996
rect 25964 40976 26016 40996
rect 26016 40976 26018 40996
rect 24214 39480 24270 39536
rect 23478 38392 23534 38448
rect 22742 36080 22798 36136
rect 22926 34448 22982 34504
rect 24030 37032 24086 37088
rect 24306 36660 24308 36680
rect 24308 36660 24360 36680
rect 24360 36660 24362 36680
rect 24306 36624 24362 36660
rect 26882 36488 26938 36544
rect 26514 36216 26570 36272
rect 25686 34312 25742 34368
rect 25226 33088 25282 33144
rect 23018 29144 23074 29200
rect 21546 24248 21602 24304
rect 20534 13812 20536 13832
rect 20536 13812 20588 13832
rect 20588 13812 20590 13832
rect 20534 13776 20590 13812
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 19430 9968 19486 10024
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 17866 4800 17922 4856
rect 16394 2352 16450 2408
rect 19154 4120 19210 4176
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 20166 6296 20222 6352
rect 26422 33088 26478 33144
rect 24950 31320 25006 31376
rect 24950 30912 25006 30968
rect 23754 28600 23810 28656
rect 23938 26016 23994 26072
rect 24398 25744 24454 25800
rect 23938 22480 23994 22536
rect 24490 23432 24546 23488
rect 24490 23024 24546 23080
rect 24398 22072 24454 22128
rect 26882 33088 26938 33144
rect 30194 40704 30250 40760
rect 30930 39500 30986 39536
rect 30930 39480 30932 39500
rect 30932 39480 30984 39500
rect 30984 39480 30986 39500
rect 29090 37848 29146 37904
rect 30194 37848 30250 37904
rect 28446 37168 28502 37224
rect 28722 35536 28778 35592
rect 26606 28872 26662 28928
rect 27342 28212 27398 28248
rect 27342 28192 27344 28212
rect 27344 28192 27396 28212
rect 27396 28192 27398 28212
rect 23478 18264 23534 18320
rect 20534 5072 20590 5128
rect 20810 7384 20866 7440
rect 23662 13232 23718 13288
rect 22466 9560 22522 9616
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 22098 2080 22154 2136
rect 21730 1672 21786 1728
rect 23478 7384 23534 7440
rect 24858 8200 24914 8256
rect 24950 8064 25006 8120
rect 28814 33768 28870 33824
rect 28630 32952 28686 33008
rect 28722 31184 28778 31240
rect 28538 30232 28594 30288
rect 27434 24248 27490 24304
rect 27894 26696 27950 26752
rect 27618 22480 27674 22536
rect 28262 24656 28318 24712
rect 28722 26968 28778 27024
rect 29918 30912 29974 30968
rect 30470 34312 30526 34368
rect 29550 30232 29606 30288
rect 31298 34312 31354 34368
rect 30470 31320 30526 31376
rect 32034 38120 32090 38176
rect 32126 37168 32182 37224
rect 32218 36080 32274 36136
rect 34940 41370 34996 41372
rect 35020 41370 35076 41372
rect 35100 41370 35156 41372
rect 35180 41370 35236 41372
rect 34940 41318 34966 41370
rect 34966 41318 34996 41370
rect 35020 41318 35030 41370
rect 35030 41318 35076 41370
rect 35100 41318 35146 41370
rect 35146 41318 35156 41370
rect 35180 41318 35210 41370
rect 35210 41318 35236 41370
rect 34940 41316 34996 41318
rect 35020 41316 35076 41318
rect 35100 41316 35156 41318
rect 35180 41316 35236 41318
rect 32862 39616 32918 39672
rect 32862 38120 32918 38176
rect 34940 40282 34996 40284
rect 35020 40282 35076 40284
rect 35100 40282 35156 40284
rect 35180 40282 35236 40284
rect 34940 40230 34966 40282
rect 34966 40230 34996 40282
rect 35020 40230 35030 40282
rect 35030 40230 35076 40282
rect 35100 40230 35146 40282
rect 35146 40230 35156 40282
rect 35180 40230 35210 40282
rect 35210 40230 35236 40282
rect 34940 40228 34996 40230
rect 35020 40228 35076 40230
rect 35100 40228 35156 40230
rect 35180 40228 35236 40230
rect 35622 40704 35678 40760
rect 34940 39194 34996 39196
rect 35020 39194 35076 39196
rect 35100 39194 35156 39196
rect 35180 39194 35236 39196
rect 34940 39142 34966 39194
rect 34966 39142 34996 39194
rect 35020 39142 35030 39194
rect 35030 39142 35076 39194
rect 35100 39142 35146 39194
rect 35146 39142 35156 39194
rect 35180 39142 35210 39194
rect 35210 39142 35236 39194
rect 34940 39140 34996 39142
rect 35020 39140 35076 39142
rect 35100 39140 35156 39142
rect 35180 39140 35236 39142
rect 34426 38936 34482 38992
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 38198 40704 38254 40760
rect 35990 37848 36046 37904
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 34242 35536 34298 35592
rect 34702 35536 34758 35592
rect 30930 31320 30986 31376
rect 30378 27376 30434 27432
rect 32402 26832 32458 26888
rect 29366 24656 29422 24712
rect 29182 18944 29238 19000
rect 25226 10920 25282 10976
rect 27526 15952 27582 16008
rect 28170 15952 28226 16008
rect 27710 11736 27766 11792
rect 26882 11600 26938 11656
rect 25778 11192 25834 11248
rect 25962 9560 26018 9616
rect 27526 11464 27582 11520
rect 27894 10240 27950 10296
rect 25778 5616 25834 5672
rect 24766 2624 24822 2680
rect 24582 2488 24638 2544
rect 26238 2388 26240 2408
rect 26240 2388 26292 2408
rect 26292 2388 26294 2408
rect 26238 2352 26294 2388
rect 25226 1808 25282 1864
rect 27250 6840 27306 6896
rect 32402 24520 32458 24576
rect 33506 30776 33562 30832
rect 33598 28872 33654 28928
rect 31758 23468 31760 23488
rect 31760 23468 31812 23488
rect 31812 23468 31814 23488
rect 31758 23432 31814 23468
rect 30654 21392 30710 21448
rect 30194 20304 30250 20360
rect 29642 15952 29698 16008
rect 30746 13368 30802 13424
rect 28722 11056 28778 11112
rect 28354 8336 28410 8392
rect 32770 23024 32826 23080
rect 32402 21936 32458 21992
rect 34518 33768 34574 33824
rect 34334 33088 34390 33144
rect 33782 22616 33838 22672
rect 32862 21120 32918 21176
rect 32954 20304 33010 20360
rect 32954 18672 33010 18728
rect 32218 17992 32274 18048
rect 32954 14456 33010 14512
rect 34242 26696 34298 26752
rect 34242 23432 34298 23488
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 35254 30812 35256 30832
rect 35256 30812 35308 30832
rect 35308 30812 35310 30832
rect 35254 30776 35310 30812
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 36358 37168 36414 37224
rect 35622 31320 35678 31376
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 36266 31184 36322 31240
rect 35714 27412 35716 27432
rect 35716 27412 35768 27432
rect 35768 27412 35770 27432
rect 35714 27376 35770 27412
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34518 18672 34574 18728
rect 34702 16088 34758 16144
rect 32586 11464 32642 11520
rect 33138 8064 33194 8120
rect 34702 12280 34758 12336
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 35438 22616 35494 22672
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 38014 37168 38070 37224
rect 36818 30912 36874 30968
rect 37554 28872 37610 28928
rect 36450 26696 36506 26752
rect 36450 24792 36506 24848
rect 36174 20304 36230 20360
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 36082 18944 36138 19000
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 35346 17176 35402 17232
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 36910 24520 36966 24576
rect 36818 21936 36874 21992
rect 36542 21120 36598 21176
rect 37094 21392 37150 21448
rect 38382 33088 38438 33144
rect 38658 34312 38714 34368
rect 39302 38936 39358 38992
rect 41326 39480 41382 39536
rect 40314 36488 40370 36544
rect 39026 28872 39082 28928
rect 37370 19660 37372 19680
rect 37372 19660 37424 19680
rect 37424 19660 37426 19680
rect 37370 19624 37426 19660
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 35162 10240 35218 10296
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 34978 8336 35034 8392
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 34518 6840 34574 6896
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 37922 22480 37978 22536
rect 35530 8200 35586 8256
rect 38382 23432 38438 23488
rect 38106 19080 38162 19136
rect 38750 23432 38806 23488
rect 39302 23024 39358 23080
rect 38842 21120 38898 21176
rect 39670 23432 39726 23488
rect 40590 36080 40646 36136
rect 43074 43560 43130 43616
rect 43074 40704 43130 40760
rect 41142 36080 41198 36136
rect 41694 36488 41750 36544
rect 38198 14456 38254 14512
rect 40314 21936 40370 21992
rect 40222 16088 40278 16144
rect 36358 6296 36414 6352
rect 35254 5072 35310 5128
rect 33690 2624 33746 2680
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 33598 2488 33654 2544
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 40774 26832 40830 26888
rect 45006 33088 45062 33144
rect 45098 31320 45154 31376
rect 40958 19624 41014 19680
rect 40774 17992 40830 18048
rect 40498 15952 40554 16008
rect 42246 19624 42302 19680
rect 43258 19080 43314 19136
rect 43258 18264 43314 18320
rect 43534 24792 43590 24848
rect 43902 24792 43958 24848
rect 43810 22616 43866 22672
rect 45190 17176 45246 17232
rect 43350 14456 43406 14512
rect 42890 12280 42946 12336
rect 44178 12280 44234 12336
<< metal3 >>
rect 19568 47360 19888 47361
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 47295 19888 47296
rect 4208 46816 4528 46817
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 46751 4528 46752
rect 34928 46816 35248 46817
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 46751 35248 46752
rect 19568 46272 19888 46273
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 46207 19888 46208
rect 4208 45728 4528 45729
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 45663 4528 45664
rect 34928 45728 35248 45729
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 45663 35248 45664
rect 19568 45184 19888 45185
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 45119 19888 45120
rect 4208 44640 4528 44641
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 44575 4528 44576
rect 34928 44640 35248 44641
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 44575 35248 44576
rect 19568 44096 19888 44097
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 44031 19888 44032
rect 49520 43800 50000 43920
rect 43069 43618 43135 43621
rect 49558 43618 49618 43800
rect 43069 43616 49618 43618
rect 43069 43560 43074 43616
rect 43130 43560 49618 43616
rect 43069 43558 49618 43560
rect 43069 43555 43135 43558
rect 4208 43552 4528 43553
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 34928 43552 35248 43553
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 43487 35248 43488
rect 19568 43008 19888 43009
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 42943 19888 42944
rect 4208 42464 4528 42465
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 34928 42464 35248 42465
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 42399 35248 42400
rect 19568 41920 19888 41921
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 41855 19888 41856
rect 0 41716 480 41744
rect 0 41652 60 41716
rect 124 41652 480 41716
rect 0 41624 480 41652
rect 19057 41714 19123 41717
rect 24853 41714 24919 41717
rect 19057 41712 24919 41714
rect 19057 41656 19062 41712
rect 19118 41656 24858 41712
rect 24914 41656 24919 41712
rect 19057 41654 24919 41656
rect 19057 41651 19123 41654
rect 24853 41651 24919 41654
rect 11421 41578 11487 41581
rect 614 41576 11487 41578
rect 614 41520 11426 41576
rect 11482 41520 11487 41576
rect 614 41518 11487 41520
rect 54 41380 60 41444
rect 124 41442 130 41444
rect 614 41442 674 41518
rect 11421 41515 11487 41518
rect 124 41382 674 41442
rect 124 41380 130 41382
rect 4208 41376 4528 41377
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 34928 41376 35248 41377
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 41311 35248 41312
rect 18781 41034 18847 41037
rect 25957 41034 26023 41037
rect 18781 41032 26023 41034
rect 18781 40976 18786 41032
rect 18842 40976 25962 41032
rect 26018 40976 26023 41032
rect 18781 40974 26023 40976
rect 18781 40971 18847 40974
rect 25957 40971 26023 40974
rect 19568 40832 19888 40833
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 40767 19888 40768
rect 30189 40762 30255 40765
rect 35617 40762 35683 40765
rect 38193 40762 38259 40765
rect 43069 40762 43135 40765
rect 30189 40760 43135 40762
rect 30189 40704 30194 40760
rect 30250 40704 35622 40760
rect 35678 40704 38198 40760
rect 38254 40704 43074 40760
rect 43130 40704 43135 40760
rect 30189 40702 43135 40704
rect 30189 40699 30255 40702
rect 35617 40699 35683 40702
rect 38193 40699 38259 40702
rect 43069 40699 43135 40702
rect 4208 40288 4528 40289
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 34928 40288 35248 40289
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 40223 35248 40224
rect 11421 39946 11487 39949
rect 13353 39946 13419 39949
rect 23197 39946 23263 39949
rect 11421 39944 23263 39946
rect 11421 39888 11426 39944
rect 11482 39888 13358 39944
rect 13414 39888 23202 39944
rect 23258 39888 23263 39944
rect 11421 39886 23263 39888
rect 11421 39883 11487 39886
rect 13353 39883 13419 39886
rect 23197 39883 23263 39886
rect 19568 39744 19888 39745
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 39679 19888 39680
rect 32857 39674 32923 39677
rect 32990 39674 32996 39676
rect 32857 39672 32996 39674
rect 32857 39616 32862 39672
rect 32918 39616 32996 39672
rect 32857 39614 32996 39616
rect 32857 39611 32923 39614
rect 32990 39612 32996 39614
rect 33060 39612 33066 39676
rect 18781 39538 18847 39541
rect 24209 39538 24275 39541
rect 18781 39536 24275 39538
rect 18781 39480 18786 39536
rect 18842 39480 24214 39536
rect 24270 39480 24275 39536
rect 18781 39478 24275 39480
rect 18781 39475 18847 39478
rect 24209 39475 24275 39478
rect 30925 39538 30991 39541
rect 41321 39538 41387 39541
rect 30925 39536 41387 39538
rect 30925 39480 30930 39536
rect 30986 39480 41326 39536
rect 41382 39480 41387 39536
rect 30925 39478 41387 39480
rect 30925 39475 30991 39478
rect 41321 39475 41387 39478
rect 13629 39266 13695 39269
rect 14273 39266 14339 39269
rect 22645 39266 22711 39269
rect 13629 39264 22711 39266
rect 13629 39208 13634 39264
rect 13690 39208 14278 39264
rect 14334 39208 22650 39264
rect 22706 39208 22711 39264
rect 13629 39206 22711 39208
rect 13629 39203 13695 39206
rect 14273 39203 14339 39206
rect 22645 39203 22711 39206
rect 4208 39200 4528 39201
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 34928 39200 35248 39201
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 39135 35248 39136
rect 34421 38994 34487 38997
rect 39297 38994 39363 38997
rect 34421 38992 39363 38994
rect 34421 38936 34426 38992
rect 34482 38936 39302 38992
rect 39358 38936 39363 38992
rect 34421 38934 39363 38936
rect 34421 38931 34487 38934
rect 39297 38931 39363 38934
rect 11329 38722 11395 38725
rect 14549 38722 14615 38725
rect 11329 38720 14615 38722
rect 11329 38664 11334 38720
rect 11390 38664 14554 38720
rect 14610 38664 14615 38720
rect 11329 38662 14615 38664
rect 11329 38659 11395 38662
rect 14549 38659 14615 38662
rect 19568 38656 19888 38657
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 38591 19888 38592
rect 18413 38450 18479 38453
rect 23473 38450 23539 38453
rect 18413 38448 23539 38450
rect 18413 38392 18418 38448
rect 18474 38392 23478 38448
rect 23534 38392 23539 38448
rect 18413 38390 23539 38392
rect 18413 38387 18479 38390
rect 23473 38387 23539 38390
rect 32029 38178 32095 38181
rect 32857 38178 32923 38181
rect 32029 38176 32923 38178
rect 32029 38120 32034 38176
rect 32090 38120 32862 38176
rect 32918 38120 32923 38176
rect 32029 38118 32923 38120
rect 32029 38115 32095 38118
rect 32857 38115 32923 38118
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 38047 35248 38048
rect 29085 37906 29151 37909
rect 30189 37906 30255 37909
rect 35985 37906 36051 37909
rect 29085 37904 36051 37906
rect 29085 37848 29090 37904
rect 29146 37848 30194 37904
rect 30250 37848 35990 37904
rect 36046 37848 36051 37904
rect 29085 37846 36051 37848
rect 29085 37843 29151 37846
rect 30189 37843 30255 37846
rect 35985 37843 36051 37846
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 11881 37362 11947 37365
rect 19701 37362 19767 37365
rect 11881 37360 19767 37362
rect 11881 37304 11886 37360
rect 11942 37304 19706 37360
rect 19762 37304 19767 37360
rect 11881 37302 19767 37304
rect 11881 37299 11947 37302
rect 19701 37299 19767 37302
rect 14733 37226 14799 37229
rect 19241 37226 19307 37229
rect 14733 37224 19307 37226
rect 14733 37168 14738 37224
rect 14794 37168 19246 37224
rect 19302 37168 19307 37224
rect 14733 37166 19307 37168
rect 14733 37163 14799 37166
rect 19241 37163 19307 37166
rect 28441 37226 28507 37229
rect 32121 37226 32187 37229
rect 36353 37226 36419 37229
rect 38009 37226 38075 37229
rect 28441 37224 38075 37226
rect 28441 37168 28446 37224
rect 28502 37168 32126 37224
rect 32182 37168 36358 37224
rect 36414 37168 38014 37224
rect 38070 37168 38075 37224
rect 28441 37166 38075 37168
rect 28441 37163 28507 37166
rect 32121 37163 32187 37166
rect 36353 37163 36419 37166
rect 38009 37163 38075 37166
rect 19333 37090 19399 37093
rect 24025 37090 24091 37093
rect 19333 37088 24091 37090
rect 19333 37032 19338 37088
rect 19394 37032 24030 37088
rect 24086 37032 24091 37088
rect 19333 37030 24091 37032
rect 19333 37027 19399 37030
rect 24025 37027 24091 37030
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 11237 36682 11303 36685
rect 24301 36682 24367 36685
rect 11237 36680 24367 36682
rect 11237 36624 11242 36680
rect 11298 36624 24306 36680
rect 24362 36624 24367 36680
rect 11237 36622 24367 36624
rect 11237 36619 11303 36622
rect 24301 36619 24367 36622
rect 26877 36546 26943 36549
rect 32990 36546 32996 36548
rect 26877 36544 32996 36546
rect 26877 36488 26882 36544
rect 26938 36488 32996 36544
rect 26877 36486 32996 36488
rect 26877 36483 26943 36486
rect 32990 36484 32996 36486
rect 33060 36546 33066 36548
rect 40309 36546 40375 36549
rect 41689 36546 41755 36549
rect 33060 36544 41755 36546
rect 33060 36488 40314 36544
rect 40370 36488 41694 36544
rect 41750 36488 41755 36544
rect 33060 36486 41755 36488
rect 33060 36484 33066 36486
rect 40309 36483 40375 36486
rect 41689 36483 41755 36486
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 21725 36274 21791 36277
rect 26509 36274 26575 36277
rect 21725 36272 26575 36274
rect 21725 36216 21730 36272
rect 21786 36216 26514 36272
rect 26570 36216 26575 36272
rect 21725 36214 26575 36216
rect 21725 36211 21791 36214
rect 26509 36211 26575 36214
rect 16021 36138 16087 36141
rect 17217 36138 17283 36141
rect 22737 36138 22803 36141
rect 16021 36136 22803 36138
rect 16021 36080 16026 36136
rect 16082 36080 17222 36136
rect 17278 36080 22742 36136
rect 22798 36080 22803 36136
rect 16021 36078 22803 36080
rect 16021 36075 16087 36078
rect 17217 36075 17283 36078
rect 22737 36075 22803 36078
rect 32213 36138 32279 36141
rect 40585 36138 40651 36141
rect 41137 36138 41203 36141
rect 32213 36136 41203 36138
rect 32213 36080 32218 36136
rect 32274 36080 40590 36136
rect 40646 36080 41142 36136
rect 41198 36080 41203 36136
rect 32213 36078 41203 36080
rect 32213 36075 32279 36078
rect 40585 36075 40651 36078
rect 41137 36075 41203 36078
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 28717 35594 28783 35597
rect 34237 35594 34303 35597
rect 34697 35594 34763 35597
rect 28717 35592 34763 35594
rect 28717 35536 28722 35592
rect 28778 35536 34242 35592
rect 34298 35536 34702 35592
rect 34758 35536 34763 35592
rect 28717 35534 34763 35536
rect 28717 35531 28783 35534
rect 34237 35531 34303 35534
rect 34697 35531 34763 35534
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 14089 34506 14155 34509
rect 21081 34506 21147 34509
rect 22921 34506 22987 34509
rect 14089 34504 22987 34506
rect 14089 34448 14094 34504
rect 14150 34448 21086 34504
rect 21142 34448 22926 34504
rect 22982 34448 22987 34504
rect 14089 34446 22987 34448
rect 14089 34443 14155 34446
rect 21081 34443 21147 34446
rect 22921 34443 22987 34446
rect 25681 34370 25747 34373
rect 30465 34370 30531 34373
rect 31293 34370 31359 34373
rect 38653 34370 38719 34373
rect 25681 34368 38719 34370
rect 25681 34312 25686 34368
rect 25742 34312 30470 34368
rect 30526 34312 31298 34368
rect 31354 34312 38658 34368
rect 38714 34312 38719 34368
rect 25681 34310 38719 34312
rect 25681 34307 25747 34310
rect 30465 34307 30531 34310
rect 31293 34307 31359 34310
rect 38653 34307 38719 34310
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 28809 33826 28875 33829
rect 34513 33826 34579 33829
rect 28809 33824 34579 33826
rect 28809 33768 28814 33824
rect 28870 33768 34518 33824
rect 34574 33768 34579 33824
rect 28809 33766 34579 33768
rect 28809 33763 28875 33766
rect 34513 33763 34579 33766
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 14549 33282 14615 33285
rect 15561 33282 15627 33285
rect 14549 33280 15627 33282
rect 14549 33224 14554 33280
rect 14610 33224 15566 33280
rect 15622 33224 15627 33280
rect 14549 33222 15627 33224
rect 14549 33219 14615 33222
rect 15561 33219 15627 33222
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 25221 33146 25287 33149
rect 26417 33146 26483 33149
rect 26877 33146 26943 33149
rect 25221 33144 26943 33146
rect 25221 33088 25226 33144
rect 25282 33088 26422 33144
rect 26478 33088 26882 33144
rect 26938 33088 26943 33144
rect 25221 33086 26943 33088
rect 25221 33083 25287 33086
rect 26417 33083 26483 33086
rect 26877 33083 26943 33086
rect 34329 33146 34395 33149
rect 38377 33146 38443 33149
rect 45001 33146 45067 33149
rect 34329 33144 45067 33146
rect 34329 33088 34334 33144
rect 34390 33088 38382 33144
rect 38438 33088 45006 33144
rect 45062 33088 45067 33144
rect 34329 33086 45067 33088
rect 34329 33083 34395 33086
rect 38377 33083 38443 33086
rect 45001 33083 45067 33086
rect 23422 32948 23428 33012
rect 23492 33010 23498 33012
rect 28625 33010 28691 33013
rect 23492 33008 28691 33010
rect 23492 32952 28630 33008
rect 28686 32952 28691 33008
rect 23492 32950 28691 32952
rect 23492 32948 23498 32950
rect 28625 32947 28691 32950
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 22277 32330 22343 32333
rect 23422 32330 23428 32332
rect 22277 32328 23428 32330
rect 22277 32272 22282 32328
rect 22338 32272 23428 32328
rect 22277 32270 23428 32272
rect 22277 32267 22343 32270
rect 23422 32268 23428 32270
rect 23492 32268 23498 32332
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 9949 31514 10015 31517
rect 13077 31514 13143 31517
rect 20805 31514 20871 31517
rect 9949 31512 20871 31514
rect 9949 31456 9954 31512
rect 10010 31456 13082 31512
rect 13138 31456 20810 31512
rect 20866 31456 20871 31512
rect 9949 31454 20871 31456
rect 9949 31451 10015 31454
rect 13077 31451 13143 31454
rect 20805 31451 20871 31454
rect 24945 31378 25011 31381
rect 30465 31378 30531 31381
rect 24945 31376 30531 31378
rect 24945 31320 24950 31376
rect 25006 31320 30470 31376
rect 30526 31320 30531 31376
rect 24945 31318 30531 31320
rect 24945 31315 25011 31318
rect 30465 31315 30531 31318
rect 30925 31378 30991 31381
rect 35617 31378 35683 31381
rect 30925 31376 35683 31378
rect 30925 31320 30930 31376
rect 30986 31320 35622 31376
rect 35678 31320 35683 31376
rect 30925 31318 35683 31320
rect 30925 31315 30991 31318
rect 35617 31315 35683 31318
rect 45093 31378 45159 31381
rect 49520 31378 50000 31408
rect 45093 31376 50000 31378
rect 45093 31320 45098 31376
rect 45154 31320 50000 31376
rect 45093 31318 50000 31320
rect 45093 31315 45159 31318
rect 49520 31288 50000 31318
rect 10409 31242 10475 31245
rect 20621 31242 20687 31245
rect 10409 31240 20687 31242
rect 10409 31184 10414 31240
rect 10470 31184 20626 31240
rect 20682 31184 20687 31240
rect 10409 31182 20687 31184
rect 10409 31179 10475 31182
rect 20621 31179 20687 31182
rect 28717 31242 28783 31245
rect 36261 31242 36327 31245
rect 28717 31240 36327 31242
rect 28717 31184 28722 31240
rect 28778 31184 36266 31240
rect 36322 31184 36327 31240
rect 28717 31182 36327 31184
rect 28717 31179 28783 31182
rect 36261 31179 36327 31182
rect 10501 31106 10567 31109
rect 19057 31106 19123 31109
rect 10501 31104 19123 31106
rect 10501 31048 10506 31104
rect 10562 31048 19062 31104
rect 19118 31048 19123 31104
rect 10501 31046 19123 31048
rect 10501 31043 10567 31046
rect 19057 31043 19123 31046
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 8293 30970 8359 30973
rect 18689 30970 18755 30973
rect 8293 30968 18755 30970
rect 8293 30912 8298 30968
rect 8354 30912 18694 30968
rect 18750 30912 18755 30968
rect 8293 30910 18755 30912
rect 8293 30907 8359 30910
rect 18689 30907 18755 30910
rect 19977 30970 20043 30973
rect 24945 30970 25011 30973
rect 19977 30968 25011 30970
rect 19977 30912 19982 30968
rect 20038 30912 24950 30968
rect 25006 30912 25011 30968
rect 19977 30910 25011 30912
rect 19977 30907 20043 30910
rect 24945 30907 25011 30910
rect 29913 30970 29979 30973
rect 36813 30970 36879 30973
rect 29913 30968 36879 30970
rect 29913 30912 29918 30968
rect 29974 30912 36818 30968
rect 36874 30912 36879 30968
rect 29913 30910 36879 30912
rect 29913 30907 29979 30910
rect 36813 30907 36879 30910
rect 33501 30834 33567 30837
rect 35249 30834 35315 30837
rect 33501 30832 35315 30834
rect 33501 30776 33506 30832
rect 33562 30776 35254 30832
rect 35310 30776 35315 30832
rect 33501 30774 35315 30776
rect 33501 30771 33567 30774
rect 35249 30771 35315 30774
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 21357 30290 21423 30293
rect 28533 30290 28599 30293
rect 29545 30290 29611 30293
rect 21357 30288 29611 30290
rect 21357 30232 21362 30288
rect 21418 30232 28538 30288
rect 28594 30232 29550 30288
rect 29606 30232 29611 30288
rect 21357 30230 29611 30232
rect 21357 30227 21423 30230
rect 28533 30227 28599 30230
rect 29545 30227 29611 30230
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 20897 29202 20963 29205
rect 23013 29202 23079 29205
rect 20897 29200 23079 29202
rect 20897 29144 20902 29200
rect 20958 29144 23018 29200
rect 23074 29144 23079 29200
rect 20897 29142 23079 29144
rect 20897 29139 20963 29142
rect 23013 29139 23079 29142
rect 26601 28930 26667 28933
rect 33593 28930 33659 28933
rect 37549 28930 37615 28933
rect 39021 28930 39087 28933
rect 26601 28928 39087 28930
rect 26601 28872 26606 28928
rect 26662 28872 33598 28928
rect 33654 28872 37554 28928
rect 37610 28872 39026 28928
rect 39082 28872 39087 28928
rect 26601 28870 39087 28872
rect 26601 28867 26667 28870
rect 33593 28867 33659 28870
rect 37549 28867 37615 28870
rect 39021 28867 39087 28870
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 18597 28658 18663 28661
rect 23749 28658 23815 28661
rect 18597 28656 23815 28658
rect 18597 28600 18602 28656
rect 18658 28600 23754 28656
rect 23810 28600 23815 28656
rect 18597 28598 23815 28600
rect 18597 28595 18663 28598
rect 23749 28595 23815 28598
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 14273 28250 14339 28253
rect 15745 28250 15811 28253
rect 27337 28250 27403 28253
rect 14273 28248 27403 28250
rect 14273 28192 14278 28248
rect 14334 28192 15750 28248
rect 15806 28192 27342 28248
rect 27398 28192 27403 28248
rect 14273 28190 27403 28192
rect 14273 28187 14339 28190
rect 15745 28187 15811 28190
rect 27337 28187 27403 28190
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 9857 27570 9923 27573
rect 15377 27570 15443 27573
rect 9857 27568 15443 27570
rect 9857 27512 9862 27568
rect 9918 27512 15382 27568
rect 15438 27512 15443 27568
rect 9857 27510 15443 27512
rect 9857 27507 9923 27510
rect 15377 27507 15443 27510
rect 30373 27434 30439 27437
rect 35709 27434 35775 27437
rect 30373 27432 35775 27434
rect 30373 27376 30378 27432
rect 30434 27376 35714 27432
rect 35770 27376 35775 27432
rect 30373 27374 35775 27376
rect 30373 27371 30439 27374
rect 35709 27371 35775 27374
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 27167 35248 27168
rect 23422 26964 23428 27028
rect 23492 27026 23498 27028
rect 28717 27026 28783 27029
rect 23492 27024 28783 27026
rect 23492 26968 28722 27024
rect 28778 26968 28783 27024
rect 23492 26966 28783 26968
rect 23492 26964 23498 26966
rect 28717 26963 28783 26966
rect 32397 26890 32463 26893
rect 40769 26890 40835 26893
rect 32397 26888 40835 26890
rect 32397 26832 32402 26888
rect 32458 26832 40774 26888
rect 40830 26832 40835 26888
rect 32397 26830 40835 26832
rect 32397 26827 32463 26830
rect 40769 26827 40835 26830
rect 27889 26754 27955 26757
rect 34237 26754 34303 26757
rect 36445 26754 36511 26757
rect 27889 26752 36511 26754
rect 27889 26696 27894 26752
rect 27950 26696 34242 26752
rect 34298 26696 36450 26752
rect 36506 26696 36511 26752
rect 27889 26694 36511 26696
rect 27889 26691 27955 26694
rect 34237 26691 34303 26694
rect 36445 26691 36511 26694
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 17401 26074 17467 26077
rect 23933 26074 23999 26077
rect 17401 26072 23999 26074
rect 17401 26016 17406 26072
rect 17462 26016 23938 26072
rect 23994 26016 23999 26072
rect 17401 26014 23999 26016
rect 17401 26011 17467 26014
rect 23933 26011 23999 26014
rect 11881 25938 11947 25941
rect 21081 25938 21147 25941
rect 11881 25936 21147 25938
rect 11881 25880 11886 25936
rect 11942 25880 21086 25936
rect 21142 25880 21147 25936
rect 11881 25878 21147 25880
rect 11881 25875 11947 25878
rect 21081 25875 21147 25878
rect 11053 25802 11119 25805
rect 24393 25802 24459 25805
rect 11053 25800 24459 25802
rect 11053 25744 11058 25800
rect 11114 25744 24398 25800
rect 24454 25744 24459 25800
rect 11053 25742 24459 25744
rect 11053 25739 11119 25742
rect 24393 25739 24459 25742
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 9397 25258 9463 25261
rect 62 25256 9463 25258
rect 62 25200 9402 25256
rect 9458 25200 9463 25256
rect 62 25198 9463 25200
rect 62 25016 122 25198
rect 9397 25195 9463 25198
rect 4208 25056 4528 25057
rect 0 24896 480 25016
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 36445 24850 36511 24853
rect 43529 24850 43595 24853
rect 43897 24850 43963 24853
rect 36445 24848 43963 24850
rect 36445 24792 36450 24848
rect 36506 24792 43534 24848
rect 43590 24792 43902 24848
rect 43958 24792 43963 24848
rect 36445 24790 43963 24792
rect 36445 24787 36511 24790
rect 43529 24787 43595 24790
rect 43897 24787 43963 24790
rect 17769 24714 17835 24717
rect 28257 24714 28323 24717
rect 29361 24714 29427 24717
rect 17769 24712 29427 24714
rect 17769 24656 17774 24712
rect 17830 24656 28262 24712
rect 28318 24656 29366 24712
rect 29422 24656 29427 24712
rect 17769 24654 29427 24656
rect 17769 24651 17835 24654
rect 28257 24651 28323 24654
rect 29361 24651 29427 24654
rect 32397 24578 32463 24581
rect 36905 24578 36971 24581
rect 32397 24576 36971 24578
rect 32397 24520 32402 24576
rect 32458 24520 36910 24576
rect 36966 24520 36971 24576
rect 32397 24518 36971 24520
rect 32397 24515 32463 24518
rect 36905 24515 36971 24518
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 18045 24306 18111 24309
rect 21541 24306 21607 24309
rect 27429 24306 27495 24309
rect 18045 24304 27495 24306
rect 18045 24248 18050 24304
rect 18106 24248 21546 24304
rect 21602 24248 27434 24304
rect 27490 24248 27495 24304
rect 18045 24246 27495 24248
rect 18045 24243 18111 24246
rect 21541 24243 21607 24246
rect 27429 24243 27495 24246
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 18413 23762 18479 23765
rect 20621 23762 20687 23765
rect 18413 23760 20687 23762
rect 18413 23704 18418 23760
rect 18474 23704 20626 23760
rect 20682 23704 20687 23760
rect 18413 23702 20687 23704
rect 18413 23699 18479 23702
rect 20621 23699 20687 23702
rect 24485 23490 24551 23493
rect 31753 23490 31819 23493
rect 24485 23488 31819 23490
rect 24485 23432 24490 23488
rect 24546 23432 31758 23488
rect 31814 23432 31819 23488
rect 24485 23430 31819 23432
rect 24485 23427 24551 23430
rect 31753 23427 31819 23430
rect 34237 23490 34303 23493
rect 38377 23490 38443 23493
rect 34237 23488 38443 23490
rect 34237 23432 34242 23488
rect 34298 23432 38382 23488
rect 38438 23432 38443 23488
rect 34237 23430 38443 23432
rect 34237 23427 34303 23430
rect 38377 23427 38443 23430
rect 38745 23490 38811 23493
rect 39665 23490 39731 23493
rect 38745 23488 39731 23490
rect 38745 23432 38750 23488
rect 38806 23432 39670 23488
rect 39726 23432 39731 23488
rect 38745 23430 39731 23432
rect 38745 23427 38811 23430
rect 39665 23427 39731 23430
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 2773 23082 2839 23085
rect 24485 23082 24551 23085
rect 2773 23080 24551 23082
rect 2773 23024 2778 23080
rect 2834 23024 24490 23080
rect 24546 23024 24551 23080
rect 2773 23022 24551 23024
rect 2773 23019 2839 23022
rect 24485 23019 24551 23022
rect 32765 23082 32831 23085
rect 39297 23082 39363 23085
rect 32765 23080 39363 23082
rect 32765 23024 32770 23080
rect 32826 23024 39302 23080
rect 39358 23024 39363 23080
rect 32765 23022 39363 23024
rect 32765 23019 32831 23022
rect 39297 23019 39363 23022
rect 18137 22946 18203 22949
rect 20529 22946 20595 22949
rect 18137 22944 20595 22946
rect 18137 22888 18142 22944
rect 18198 22888 20534 22944
rect 20590 22888 20595 22944
rect 18137 22886 20595 22888
rect 18137 22883 18203 22886
rect 20529 22883 20595 22886
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 19241 22810 19307 22813
rect 20253 22810 20319 22813
rect 19241 22808 20319 22810
rect 19241 22752 19246 22808
rect 19302 22752 20258 22808
rect 20314 22752 20319 22808
rect 19241 22750 20319 22752
rect 19241 22747 19307 22750
rect 20253 22747 20319 22750
rect 10501 22674 10567 22677
rect 16389 22674 16455 22677
rect 10501 22672 16455 22674
rect 10501 22616 10506 22672
rect 10562 22616 16394 22672
rect 16450 22616 16455 22672
rect 10501 22614 16455 22616
rect 10501 22611 10567 22614
rect 16389 22611 16455 22614
rect 33777 22674 33843 22677
rect 35433 22674 35499 22677
rect 43805 22674 43871 22677
rect 33777 22672 43871 22674
rect 33777 22616 33782 22672
rect 33838 22616 35438 22672
rect 35494 22616 43810 22672
rect 43866 22616 43871 22672
rect 33777 22614 43871 22616
rect 33777 22611 33843 22614
rect 35433 22611 35499 22614
rect 43805 22611 43871 22614
rect 18781 22538 18847 22541
rect 23933 22538 23999 22541
rect 18781 22536 23999 22538
rect 18781 22480 18786 22536
rect 18842 22480 23938 22536
rect 23994 22480 23999 22536
rect 18781 22478 23999 22480
rect 18781 22475 18847 22478
rect 23933 22475 23999 22478
rect 27613 22538 27679 22541
rect 37917 22538 37983 22541
rect 27613 22536 37983 22538
rect 27613 22480 27618 22536
rect 27674 22480 37922 22536
rect 37978 22480 37983 22536
rect 27613 22478 37983 22480
rect 27613 22475 27679 22478
rect 37917 22475 37983 22478
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 14181 22130 14247 22133
rect 17309 22130 17375 22133
rect 24393 22130 24459 22133
rect 14181 22128 24459 22130
rect 14181 22072 14186 22128
rect 14242 22072 17314 22128
rect 17370 22072 24398 22128
rect 24454 22072 24459 22128
rect 14181 22070 24459 22072
rect 14181 22067 14247 22070
rect 17309 22067 17375 22070
rect 24393 22067 24459 22070
rect 32397 21994 32463 21997
rect 36813 21994 36879 21997
rect 40309 21994 40375 21997
rect 32397 21992 40375 21994
rect 32397 21936 32402 21992
rect 32458 21936 36818 21992
rect 36874 21936 40314 21992
rect 40370 21936 40375 21992
rect 32397 21934 40375 21936
rect 32397 21931 32463 21934
rect 36813 21931 36879 21934
rect 40309 21931 40375 21934
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 30649 21450 30715 21453
rect 37089 21450 37155 21453
rect 30649 21448 37155 21450
rect 30649 21392 30654 21448
rect 30710 21392 37094 21448
rect 37150 21392 37155 21448
rect 30649 21390 37155 21392
rect 30649 21387 30715 21390
rect 37089 21387 37155 21390
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 32857 21178 32923 21181
rect 36537 21178 36603 21181
rect 38837 21178 38903 21181
rect 32857 21176 38903 21178
rect 32857 21120 32862 21176
rect 32918 21120 36542 21176
rect 36598 21120 38842 21176
rect 38898 21120 38903 21176
rect 32857 21118 38903 21120
rect 32857 21115 32923 21118
rect 36537 21115 36603 21118
rect 38837 21115 38903 21118
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 30189 20362 30255 20365
rect 32949 20362 33015 20365
rect 36169 20362 36235 20365
rect 30189 20360 36235 20362
rect 30189 20304 30194 20360
rect 30250 20304 32954 20360
rect 33010 20304 36174 20360
rect 36230 20304 36235 20360
rect 30189 20302 36235 20304
rect 30189 20299 30255 20302
rect 32949 20299 33015 20302
rect 36169 20299 36235 20302
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 37365 19682 37431 19685
rect 40953 19682 41019 19685
rect 42241 19682 42307 19685
rect 37365 19680 42307 19682
rect 37365 19624 37370 19680
rect 37426 19624 40958 19680
rect 41014 19624 42246 19680
rect 42302 19624 42307 19680
rect 37365 19622 42307 19624
rect 37365 19619 37431 19622
rect 40953 19619 41019 19622
rect 42241 19619 42307 19622
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 13629 19274 13695 19277
rect 14089 19274 14155 19277
rect 13629 19272 14155 19274
rect 13629 19216 13634 19272
rect 13690 19216 14094 19272
rect 14150 19216 14155 19272
rect 13629 19214 14155 19216
rect 13629 19211 13695 19214
rect 14089 19211 14155 19214
rect 38101 19138 38167 19141
rect 43253 19138 43319 19141
rect 38101 19136 43319 19138
rect 38101 19080 38106 19136
rect 38162 19080 43258 19136
rect 43314 19080 43319 19136
rect 38101 19078 43319 19080
rect 38101 19075 38167 19078
rect 43253 19075 43319 19078
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 29177 19002 29243 19005
rect 36077 19002 36143 19005
rect 29177 19000 36143 19002
rect 29177 18944 29182 19000
rect 29238 18944 36082 19000
rect 36138 18944 36143 19000
rect 29177 18942 36143 18944
rect 29177 18939 29243 18942
rect 36077 18939 36143 18942
rect 19333 18866 19399 18869
rect 19517 18866 19583 18869
rect 19333 18864 19583 18866
rect 19333 18808 19338 18864
rect 19394 18808 19522 18864
rect 19578 18808 19583 18864
rect 19333 18806 19583 18808
rect 19333 18803 19399 18806
rect 19517 18803 19583 18806
rect 49520 18776 50000 18896
rect 9397 18730 9463 18733
rect 17769 18730 17835 18733
rect 9397 18728 17835 18730
rect 9397 18672 9402 18728
rect 9458 18672 17774 18728
rect 17830 18672 17835 18728
rect 9397 18670 17835 18672
rect 9397 18667 9463 18670
rect 17769 18667 17835 18670
rect 32949 18730 33015 18733
rect 34513 18730 34579 18733
rect 32949 18728 34579 18730
rect 32949 18672 32954 18728
rect 33010 18672 34518 18728
rect 34574 18672 34579 18728
rect 32949 18670 34579 18672
rect 32949 18667 33015 18670
rect 34513 18667 34579 18670
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 15101 18322 15167 18325
rect 23473 18322 23539 18325
rect 15101 18320 23539 18322
rect 15101 18264 15106 18320
rect 15162 18264 23478 18320
rect 23534 18264 23539 18320
rect 15101 18262 23539 18264
rect 15101 18259 15167 18262
rect 23473 18259 23539 18262
rect 43253 18322 43319 18325
rect 49558 18322 49618 18776
rect 43253 18320 49618 18322
rect 43253 18264 43258 18320
rect 43314 18264 49618 18320
rect 43253 18262 49618 18264
rect 43253 18259 43319 18262
rect 32213 18050 32279 18053
rect 40769 18050 40835 18053
rect 32213 18048 40835 18050
rect 32213 17992 32218 18048
rect 32274 17992 40774 18048
rect 40830 17992 40835 18048
rect 32213 17990 40835 17992
rect 32213 17987 32279 17990
rect 40769 17987 40835 17990
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 35341 17234 35407 17237
rect 45185 17234 45251 17237
rect 35341 17232 45251 17234
rect 35341 17176 35346 17232
rect 35402 17176 45190 17232
rect 45246 17176 45251 17232
rect 35341 17174 45251 17176
rect 35341 17171 35407 17174
rect 45185 17171 45251 17174
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 34697 16146 34763 16149
rect 40217 16146 40283 16149
rect 34697 16144 40283 16146
rect 34697 16088 34702 16144
rect 34758 16088 40222 16144
rect 40278 16088 40283 16144
rect 34697 16086 40283 16088
rect 34697 16083 34763 16086
rect 40217 16083 40283 16086
rect 19241 16010 19307 16013
rect 27521 16010 27587 16013
rect 28165 16010 28231 16013
rect 19241 16008 28231 16010
rect 19241 15952 19246 16008
rect 19302 15952 27526 16008
rect 27582 15952 28170 16008
rect 28226 15952 28231 16008
rect 19241 15950 28231 15952
rect 19241 15947 19307 15950
rect 27521 15947 27587 15950
rect 28165 15947 28231 15950
rect 29637 16010 29703 16013
rect 40493 16010 40559 16013
rect 29637 16008 40559 16010
rect 29637 15952 29642 16008
rect 29698 15952 40498 16008
rect 40554 15952 40559 16008
rect 29637 15950 40559 15952
rect 29637 15947 29703 15950
rect 40493 15947 40559 15950
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 32949 14514 33015 14517
rect 38193 14514 38259 14517
rect 43345 14514 43411 14517
rect 32949 14512 43411 14514
rect 32949 14456 32954 14512
rect 33010 14456 38198 14512
rect 38254 14456 43350 14512
rect 43406 14456 43411 14512
rect 32949 14454 43411 14456
rect 32949 14451 33015 14454
rect 38193 14451 38259 14454
rect 43345 14451 43411 14454
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 20529 13834 20595 13837
rect 19290 13832 20595 13834
rect 19290 13776 20534 13832
rect 20590 13776 20595 13832
rect 19290 13774 20595 13776
rect 10133 13698 10199 13701
rect 10777 13698 10843 13701
rect 19290 13698 19350 13774
rect 20529 13771 20595 13774
rect 10133 13696 19350 13698
rect 10133 13640 10138 13696
rect 10194 13640 10782 13696
rect 10838 13640 19350 13696
rect 10133 13638 19350 13640
rect 10133 13635 10199 13638
rect 10777 13635 10843 13638
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 18689 13426 18755 13429
rect 30741 13426 30807 13429
rect 18689 13424 30807 13426
rect 18689 13368 18694 13424
rect 18750 13368 30746 13424
rect 30802 13368 30807 13424
rect 18689 13366 30807 13368
rect 18689 13363 18755 13366
rect 30741 13363 30807 13366
rect 18229 13290 18295 13293
rect 23657 13290 23723 13293
rect 18229 13288 23723 13290
rect 18229 13232 18234 13288
rect 18290 13232 23662 13288
rect 23718 13232 23723 13288
rect 18229 13230 23723 13232
rect 18229 13227 18295 13230
rect 23657 13227 23723 13230
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 13023 35248 13024
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 34697 12338 34763 12341
rect 42885 12338 42951 12341
rect 44173 12338 44239 12341
rect 34697 12336 44239 12338
rect 34697 12280 34702 12336
rect 34758 12280 42890 12336
rect 42946 12280 44178 12336
rect 44234 12280 44239 12336
rect 34697 12278 44239 12280
rect 34697 12275 34763 12278
rect 42885 12275 42951 12278
rect 44173 12275 44239 12278
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 12709 11794 12775 11797
rect 27705 11794 27771 11797
rect 12709 11792 27771 11794
rect 12709 11736 12714 11792
rect 12770 11736 27710 11792
rect 27766 11736 27771 11792
rect 12709 11734 27771 11736
rect 12709 11731 12775 11734
rect 27705 11731 27771 11734
rect 18045 11658 18111 11661
rect 26877 11658 26943 11661
rect 18045 11656 26943 11658
rect 18045 11600 18050 11656
rect 18106 11600 26882 11656
rect 26938 11600 26943 11656
rect 18045 11598 26943 11600
rect 18045 11595 18111 11598
rect 26877 11595 26943 11598
rect 27521 11522 27587 11525
rect 32581 11522 32647 11525
rect 27521 11520 32647 11522
rect 27521 11464 27526 11520
rect 27582 11464 32586 11520
rect 32642 11464 32647 11520
rect 27521 11462 32647 11464
rect 27521 11459 27587 11462
rect 32581 11459 32647 11462
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 10317 11250 10383 11253
rect 25773 11250 25839 11253
rect 10317 11248 25839 11250
rect 10317 11192 10322 11248
rect 10378 11192 25778 11248
rect 25834 11192 25839 11248
rect 10317 11190 25839 11192
rect 10317 11187 10383 11190
rect 25773 11187 25839 11190
rect 12893 11114 12959 11117
rect 28717 11114 28783 11117
rect 12893 11112 28783 11114
rect 12893 11056 12898 11112
rect 12954 11056 28722 11112
rect 28778 11056 28783 11112
rect 12893 11054 28783 11056
rect 12893 11051 12959 11054
rect 28717 11051 28783 11054
rect 9673 10978 9739 10981
rect 25221 10978 25287 10981
rect 9673 10976 25287 10978
rect 9673 10920 9678 10976
rect 9734 10920 25226 10976
rect 25282 10920 25287 10976
rect 9673 10918 25287 10920
rect 9673 10915 9739 10918
rect 25221 10915 25287 10918
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 27889 10298 27955 10301
rect 35157 10298 35223 10301
rect 27889 10296 35223 10298
rect 27889 10240 27894 10296
rect 27950 10240 35162 10296
rect 35218 10240 35223 10296
rect 27889 10238 35223 10240
rect 27889 10235 27955 10238
rect 35157 10235 35223 10238
rect 9765 10026 9831 10029
rect 10409 10026 10475 10029
rect 19425 10026 19491 10029
rect 9765 10024 19491 10026
rect 9765 9968 9770 10024
rect 9826 9968 10414 10024
rect 10470 9968 19430 10024
rect 19486 9968 19491 10024
rect 9765 9966 19491 9968
rect 9765 9963 9831 9966
rect 10409 9963 10475 9966
rect 19425 9963 19491 9966
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 22461 9618 22527 9621
rect 25957 9618 26023 9621
rect 22461 9616 26023 9618
rect 22461 9560 22466 9616
rect 22522 9560 25962 9616
rect 26018 9560 26023 9616
rect 22461 9558 26023 9560
rect 22461 9555 22527 9558
rect 25957 9555 26023 9558
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 18137 8938 18203 8941
rect 62 8936 18203 8938
rect 62 8880 18142 8936
rect 18198 8880 18203 8936
rect 62 8878 18203 8880
rect 62 8424 122 8878
rect 18137 8875 18203 8878
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 0 8304 480 8424
rect 28349 8394 28415 8397
rect 34973 8394 35039 8397
rect 28349 8392 35039 8394
rect 28349 8336 28354 8392
rect 28410 8336 34978 8392
rect 35034 8336 35039 8392
rect 28349 8334 35039 8336
rect 28349 8331 28415 8334
rect 34973 8331 35039 8334
rect 24853 8258 24919 8261
rect 35525 8258 35591 8261
rect 24853 8256 35591 8258
rect 24853 8200 24858 8256
rect 24914 8200 35530 8256
rect 35586 8200 35591 8256
rect 24853 8198 35591 8200
rect 24853 8195 24919 8198
rect 35525 8195 35591 8198
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 24945 8122 25011 8125
rect 33133 8122 33199 8125
rect 24945 8120 33199 8122
rect 24945 8064 24950 8120
rect 25006 8064 33138 8120
rect 33194 8064 33199 8120
rect 24945 8062 33199 8064
rect 24945 8059 25011 8062
rect 33133 8059 33199 8062
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 20805 7442 20871 7445
rect 23473 7442 23539 7445
rect 20805 7440 23539 7442
rect 20805 7384 20810 7440
rect 20866 7384 23478 7440
rect 23534 7384 23539 7440
rect 20805 7382 23539 7384
rect 20805 7379 20871 7382
rect 23473 7379 23539 7382
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 27245 6898 27311 6901
rect 34513 6898 34579 6901
rect 27245 6896 34579 6898
rect 27245 6840 27250 6896
rect 27306 6840 34518 6896
rect 34574 6840 34579 6896
rect 27245 6838 34579 6840
rect 27245 6835 27311 6838
rect 34513 6835 34579 6838
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 20161 6354 20227 6357
rect 36353 6354 36419 6357
rect 20161 6352 36419 6354
rect 20161 6296 20166 6352
rect 20222 6296 36358 6352
rect 36414 6296 36419 6352
rect 20161 6294 36419 6296
rect 20161 6291 20227 6294
rect 36353 6291 36419 6294
rect 49520 6264 50000 6384
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 25773 5674 25839 5677
rect 49558 5674 49618 6264
rect 25773 5672 49618 5674
rect 25773 5616 25778 5672
rect 25834 5616 49618 5672
rect 25773 5614 49618 5616
rect 25773 5611 25839 5614
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 12433 5266 12499 5269
rect 17217 5266 17283 5269
rect 12433 5264 17283 5266
rect 12433 5208 12438 5264
rect 12494 5208 17222 5264
rect 17278 5208 17283 5264
rect 12433 5206 17283 5208
rect 12433 5203 12499 5206
rect 17217 5203 17283 5206
rect 20529 5130 20595 5133
rect 35249 5130 35315 5133
rect 20529 5128 35315 5130
rect 20529 5072 20534 5128
rect 20590 5072 35254 5128
rect 35310 5072 35315 5128
rect 20529 5070 35315 5072
rect 20529 5067 20595 5070
rect 35249 5067 35315 5070
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 10501 4858 10567 4861
rect 17861 4858 17927 4861
rect 10501 4856 17927 4858
rect 10501 4800 10506 4856
rect 10562 4800 17866 4856
rect 17922 4800 17927 4856
rect 10501 4798 17927 4800
rect 10501 4795 10567 4798
rect 17861 4795 17927 4798
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 14181 4178 14247 4181
rect 15101 4178 15167 4181
rect 19149 4178 19215 4181
rect 14181 4176 19215 4178
rect 14181 4120 14186 4176
rect 14242 4120 15106 4176
rect 15162 4120 19154 4176
rect 19210 4120 19215 4176
rect 14181 4118 19215 4120
rect 14181 4115 14247 4118
rect 15101 4115 15167 4118
rect 19149 4115 19215 4118
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 24761 2682 24827 2685
rect 33685 2682 33751 2685
rect 24761 2680 33751 2682
rect 24761 2624 24766 2680
rect 24822 2624 33690 2680
rect 33746 2624 33751 2680
rect 24761 2622 33751 2624
rect 24761 2619 24827 2622
rect 33685 2619 33751 2622
rect 24577 2546 24643 2549
rect 33593 2546 33659 2549
rect 24577 2544 33659 2546
rect 24577 2488 24582 2544
rect 24638 2488 33598 2544
rect 33654 2488 33659 2544
rect 24577 2486 33659 2488
rect 24577 2483 24643 2486
rect 33593 2483 33659 2486
rect 16389 2410 16455 2413
rect 26233 2410 26299 2413
rect 16389 2408 26299 2410
rect 16389 2352 16394 2408
rect 16450 2352 26238 2408
rect 26294 2352 26299 2408
rect 16389 2350 26299 2352
rect 16389 2347 16455 2350
rect 26233 2347 26299 2350
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
rect 11421 2138 11487 2141
rect 22093 2138 22159 2141
rect 11421 2136 22159 2138
rect 11421 2080 11426 2136
rect 11482 2080 22098 2136
rect 22154 2080 22159 2136
rect 11421 2078 22159 2080
rect 11421 2075 11487 2078
rect 22093 2075 22159 2078
rect 11881 1866 11947 1869
rect 25221 1866 25287 1869
rect 11881 1864 25287 1866
rect 11881 1808 11886 1864
rect 11942 1808 25226 1864
rect 25282 1808 25287 1864
rect 11881 1806 25287 1808
rect 11881 1803 11947 1806
rect 25221 1803 25287 1806
rect 11053 1730 11119 1733
rect 21725 1730 21791 1733
rect 11053 1728 21791 1730
rect 11053 1672 11058 1728
rect 11114 1672 21730 1728
rect 21786 1672 21791 1728
rect 11053 1670 21791 1672
rect 11053 1667 11119 1670
rect 21725 1667 21791 1670
<< via3 >>
rect 19576 47356 19640 47360
rect 19576 47300 19580 47356
rect 19580 47300 19636 47356
rect 19636 47300 19640 47356
rect 19576 47296 19640 47300
rect 19656 47356 19720 47360
rect 19656 47300 19660 47356
rect 19660 47300 19716 47356
rect 19716 47300 19720 47356
rect 19656 47296 19720 47300
rect 19736 47356 19800 47360
rect 19736 47300 19740 47356
rect 19740 47300 19796 47356
rect 19796 47300 19800 47356
rect 19736 47296 19800 47300
rect 19816 47356 19880 47360
rect 19816 47300 19820 47356
rect 19820 47300 19876 47356
rect 19876 47300 19880 47356
rect 19816 47296 19880 47300
rect 4216 46812 4280 46816
rect 4216 46756 4220 46812
rect 4220 46756 4276 46812
rect 4276 46756 4280 46812
rect 4216 46752 4280 46756
rect 4296 46812 4360 46816
rect 4296 46756 4300 46812
rect 4300 46756 4356 46812
rect 4356 46756 4360 46812
rect 4296 46752 4360 46756
rect 4376 46812 4440 46816
rect 4376 46756 4380 46812
rect 4380 46756 4436 46812
rect 4436 46756 4440 46812
rect 4376 46752 4440 46756
rect 4456 46812 4520 46816
rect 4456 46756 4460 46812
rect 4460 46756 4516 46812
rect 4516 46756 4520 46812
rect 4456 46752 4520 46756
rect 34936 46812 35000 46816
rect 34936 46756 34940 46812
rect 34940 46756 34996 46812
rect 34996 46756 35000 46812
rect 34936 46752 35000 46756
rect 35016 46812 35080 46816
rect 35016 46756 35020 46812
rect 35020 46756 35076 46812
rect 35076 46756 35080 46812
rect 35016 46752 35080 46756
rect 35096 46812 35160 46816
rect 35096 46756 35100 46812
rect 35100 46756 35156 46812
rect 35156 46756 35160 46812
rect 35096 46752 35160 46756
rect 35176 46812 35240 46816
rect 35176 46756 35180 46812
rect 35180 46756 35236 46812
rect 35236 46756 35240 46812
rect 35176 46752 35240 46756
rect 19576 46268 19640 46272
rect 19576 46212 19580 46268
rect 19580 46212 19636 46268
rect 19636 46212 19640 46268
rect 19576 46208 19640 46212
rect 19656 46268 19720 46272
rect 19656 46212 19660 46268
rect 19660 46212 19716 46268
rect 19716 46212 19720 46268
rect 19656 46208 19720 46212
rect 19736 46268 19800 46272
rect 19736 46212 19740 46268
rect 19740 46212 19796 46268
rect 19796 46212 19800 46268
rect 19736 46208 19800 46212
rect 19816 46268 19880 46272
rect 19816 46212 19820 46268
rect 19820 46212 19876 46268
rect 19876 46212 19880 46268
rect 19816 46208 19880 46212
rect 4216 45724 4280 45728
rect 4216 45668 4220 45724
rect 4220 45668 4276 45724
rect 4276 45668 4280 45724
rect 4216 45664 4280 45668
rect 4296 45724 4360 45728
rect 4296 45668 4300 45724
rect 4300 45668 4356 45724
rect 4356 45668 4360 45724
rect 4296 45664 4360 45668
rect 4376 45724 4440 45728
rect 4376 45668 4380 45724
rect 4380 45668 4436 45724
rect 4436 45668 4440 45724
rect 4376 45664 4440 45668
rect 4456 45724 4520 45728
rect 4456 45668 4460 45724
rect 4460 45668 4516 45724
rect 4516 45668 4520 45724
rect 4456 45664 4520 45668
rect 34936 45724 35000 45728
rect 34936 45668 34940 45724
rect 34940 45668 34996 45724
rect 34996 45668 35000 45724
rect 34936 45664 35000 45668
rect 35016 45724 35080 45728
rect 35016 45668 35020 45724
rect 35020 45668 35076 45724
rect 35076 45668 35080 45724
rect 35016 45664 35080 45668
rect 35096 45724 35160 45728
rect 35096 45668 35100 45724
rect 35100 45668 35156 45724
rect 35156 45668 35160 45724
rect 35096 45664 35160 45668
rect 35176 45724 35240 45728
rect 35176 45668 35180 45724
rect 35180 45668 35236 45724
rect 35236 45668 35240 45724
rect 35176 45664 35240 45668
rect 19576 45180 19640 45184
rect 19576 45124 19580 45180
rect 19580 45124 19636 45180
rect 19636 45124 19640 45180
rect 19576 45120 19640 45124
rect 19656 45180 19720 45184
rect 19656 45124 19660 45180
rect 19660 45124 19716 45180
rect 19716 45124 19720 45180
rect 19656 45120 19720 45124
rect 19736 45180 19800 45184
rect 19736 45124 19740 45180
rect 19740 45124 19796 45180
rect 19796 45124 19800 45180
rect 19736 45120 19800 45124
rect 19816 45180 19880 45184
rect 19816 45124 19820 45180
rect 19820 45124 19876 45180
rect 19876 45124 19880 45180
rect 19816 45120 19880 45124
rect 4216 44636 4280 44640
rect 4216 44580 4220 44636
rect 4220 44580 4276 44636
rect 4276 44580 4280 44636
rect 4216 44576 4280 44580
rect 4296 44636 4360 44640
rect 4296 44580 4300 44636
rect 4300 44580 4356 44636
rect 4356 44580 4360 44636
rect 4296 44576 4360 44580
rect 4376 44636 4440 44640
rect 4376 44580 4380 44636
rect 4380 44580 4436 44636
rect 4436 44580 4440 44636
rect 4376 44576 4440 44580
rect 4456 44636 4520 44640
rect 4456 44580 4460 44636
rect 4460 44580 4516 44636
rect 4516 44580 4520 44636
rect 4456 44576 4520 44580
rect 34936 44636 35000 44640
rect 34936 44580 34940 44636
rect 34940 44580 34996 44636
rect 34996 44580 35000 44636
rect 34936 44576 35000 44580
rect 35016 44636 35080 44640
rect 35016 44580 35020 44636
rect 35020 44580 35076 44636
rect 35076 44580 35080 44636
rect 35016 44576 35080 44580
rect 35096 44636 35160 44640
rect 35096 44580 35100 44636
rect 35100 44580 35156 44636
rect 35156 44580 35160 44636
rect 35096 44576 35160 44580
rect 35176 44636 35240 44640
rect 35176 44580 35180 44636
rect 35180 44580 35236 44636
rect 35236 44580 35240 44636
rect 35176 44576 35240 44580
rect 19576 44092 19640 44096
rect 19576 44036 19580 44092
rect 19580 44036 19636 44092
rect 19636 44036 19640 44092
rect 19576 44032 19640 44036
rect 19656 44092 19720 44096
rect 19656 44036 19660 44092
rect 19660 44036 19716 44092
rect 19716 44036 19720 44092
rect 19656 44032 19720 44036
rect 19736 44092 19800 44096
rect 19736 44036 19740 44092
rect 19740 44036 19796 44092
rect 19796 44036 19800 44092
rect 19736 44032 19800 44036
rect 19816 44092 19880 44096
rect 19816 44036 19820 44092
rect 19820 44036 19876 44092
rect 19876 44036 19880 44092
rect 19816 44032 19880 44036
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 34936 43548 35000 43552
rect 34936 43492 34940 43548
rect 34940 43492 34996 43548
rect 34996 43492 35000 43548
rect 34936 43488 35000 43492
rect 35016 43548 35080 43552
rect 35016 43492 35020 43548
rect 35020 43492 35076 43548
rect 35076 43492 35080 43548
rect 35016 43488 35080 43492
rect 35096 43548 35160 43552
rect 35096 43492 35100 43548
rect 35100 43492 35156 43548
rect 35156 43492 35160 43548
rect 35096 43488 35160 43492
rect 35176 43548 35240 43552
rect 35176 43492 35180 43548
rect 35180 43492 35236 43548
rect 35236 43492 35240 43548
rect 35176 43488 35240 43492
rect 19576 43004 19640 43008
rect 19576 42948 19580 43004
rect 19580 42948 19636 43004
rect 19636 42948 19640 43004
rect 19576 42944 19640 42948
rect 19656 43004 19720 43008
rect 19656 42948 19660 43004
rect 19660 42948 19716 43004
rect 19716 42948 19720 43004
rect 19656 42944 19720 42948
rect 19736 43004 19800 43008
rect 19736 42948 19740 43004
rect 19740 42948 19796 43004
rect 19796 42948 19800 43004
rect 19736 42944 19800 42948
rect 19816 43004 19880 43008
rect 19816 42948 19820 43004
rect 19820 42948 19876 43004
rect 19876 42948 19880 43004
rect 19816 42944 19880 42948
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 34936 42460 35000 42464
rect 34936 42404 34940 42460
rect 34940 42404 34996 42460
rect 34996 42404 35000 42460
rect 34936 42400 35000 42404
rect 35016 42460 35080 42464
rect 35016 42404 35020 42460
rect 35020 42404 35076 42460
rect 35076 42404 35080 42460
rect 35016 42400 35080 42404
rect 35096 42460 35160 42464
rect 35096 42404 35100 42460
rect 35100 42404 35156 42460
rect 35156 42404 35160 42460
rect 35096 42400 35160 42404
rect 35176 42460 35240 42464
rect 35176 42404 35180 42460
rect 35180 42404 35236 42460
rect 35236 42404 35240 42460
rect 35176 42400 35240 42404
rect 19576 41916 19640 41920
rect 19576 41860 19580 41916
rect 19580 41860 19636 41916
rect 19636 41860 19640 41916
rect 19576 41856 19640 41860
rect 19656 41916 19720 41920
rect 19656 41860 19660 41916
rect 19660 41860 19716 41916
rect 19716 41860 19720 41916
rect 19656 41856 19720 41860
rect 19736 41916 19800 41920
rect 19736 41860 19740 41916
rect 19740 41860 19796 41916
rect 19796 41860 19800 41916
rect 19736 41856 19800 41860
rect 19816 41916 19880 41920
rect 19816 41860 19820 41916
rect 19820 41860 19876 41916
rect 19876 41860 19880 41916
rect 19816 41856 19880 41860
rect 60 41652 124 41716
rect 60 41380 124 41444
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 34936 41372 35000 41376
rect 34936 41316 34940 41372
rect 34940 41316 34996 41372
rect 34996 41316 35000 41372
rect 34936 41312 35000 41316
rect 35016 41372 35080 41376
rect 35016 41316 35020 41372
rect 35020 41316 35076 41372
rect 35076 41316 35080 41372
rect 35016 41312 35080 41316
rect 35096 41372 35160 41376
rect 35096 41316 35100 41372
rect 35100 41316 35156 41372
rect 35156 41316 35160 41372
rect 35096 41312 35160 41316
rect 35176 41372 35240 41376
rect 35176 41316 35180 41372
rect 35180 41316 35236 41372
rect 35236 41316 35240 41372
rect 35176 41312 35240 41316
rect 19576 40828 19640 40832
rect 19576 40772 19580 40828
rect 19580 40772 19636 40828
rect 19636 40772 19640 40828
rect 19576 40768 19640 40772
rect 19656 40828 19720 40832
rect 19656 40772 19660 40828
rect 19660 40772 19716 40828
rect 19716 40772 19720 40828
rect 19656 40768 19720 40772
rect 19736 40828 19800 40832
rect 19736 40772 19740 40828
rect 19740 40772 19796 40828
rect 19796 40772 19800 40828
rect 19736 40768 19800 40772
rect 19816 40828 19880 40832
rect 19816 40772 19820 40828
rect 19820 40772 19876 40828
rect 19876 40772 19880 40828
rect 19816 40768 19880 40772
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 34936 40284 35000 40288
rect 34936 40228 34940 40284
rect 34940 40228 34996 40284
rect 34996 40228 35000 40284
rect 34936 40224 35000 40228
rect 35016 40284 35080 40288
rect 35016 40228 35020 40284
rect 35020 40228 35076 40284
rect 35076 40228 35080 40284
rect 35016 40224 35080 40228
rect 35096 40284 35160 40288
rect 35096 40228 35100 40284
rect 35100 40228 35156 40284
rect 35156 40228 35160 40284
rect 35096 40224 35160 40228
rect 35176 40284 35240 40288
rect 35176 40228 35180 40284
rect 35180 40228 35236 40284
rect 35236 40228 35240 40284
rect 35176 40224 35240 40228
rect 19576 39740 19640 39744
rect 19576 39684 19580 39740
rect 19580 39684 19636 39740
rect 19636 39684 19640 39740
rect 19576 39680 19640 39684
rect 19656 39740 19720 39744
rect 19656 39684 19660 39740
rect 19660 39684 19716 39740
rect 19716 39684 19720 39740
rect 19656 39680 19720 39684
rect 19736 39740 19800 39744
rect 19736 39684 19740 39740
rect 19740 39684 19796 39740
rect 19796 39684 19800 39740
rect 19736 39680 19800 39684
rect 19816 39740 19880 39744
rect 19816 39684 19820 39740
rect 19820 39684 19876 39740
rect 19876 39684 19880 39740
rect 19816 39680 19880 39684
rect 32996 39612 33060 39676
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 34936 39196 35000 39200
rect 34936 39140 34940 39196
rect 34940 39140 34996 39196
rect 34996 39140 35000 39196
rect 34936 39136 35000 39140
rect 35016 39196 35080 39200
rect 35016 39140 35020 39196
rect 35020 39140 35076 39196
rect 35076 39140 35080 39196
rect 35016 39136 35080 39140
rect 35096 39196 35160 39200
rect 35096 39140 35100 39196
rect 35100 39140 35156 39196
rect 35156 39140 35160 39196
rect 35096 39136 35160 39140
rect 35176 39196 35240 39200
rect 35176 39140 35180 39196
rect 35180 39140 35236 39196
rect 35236 39140 35240 39196
rect 35176 39136 35240 39140
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 32996 36484 33060 36548
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 23428 32948 23492 33012
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 23428 32268 23492 32332
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 23428 26964 23492 27028
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
<< metal4 >>
rect 4208 46816 4528 47376
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 45728 4528 46752
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 44640 4528 45664
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 43552 4528 44576
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 42464 4528 43488
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 59 41716 125 41717
rect 59 41652 60 41716
rect 124 41652 125 41716
rect 59 41651 125 41652
rect 62 41445 122 41651
rect 59 41444 125 41445
rect 59 41380 60 41444
rect 124 41380 125 41444
rect 59 41379 125 41380
rect 4208 41376 4528 42400
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 47360 19888 47376
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 46272 19888 47296
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 45184 19888 46208
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 44096 19888 45120
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 43008 19888 44032
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 41920 19888 42944
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 40832 19888 41856
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 39744 19888 40768
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 38656 19888 39680
rect 34928 46816 35248 47376
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 45728 35248 46752
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 44640 35248 45664
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 43552 35248 44576
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 42464 35248 43488
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 41376 35248 42400
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 40288 35248 41312
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 32995 39676 33061 39677
rect 32995 39612 32996 39676
rect 33060 39612 33061 39676
rect 32995 39611 33061 39612
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 32998 36549 33058 39611
rect 34928 39200 35248 40224
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 38112 35248 39136
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 32995 36548 33061 36549
rect 32995 36484 32996 36548
rect 33060 36484 33061 36548
rect 32995 36483 33061 36484
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 23427 33012 23493 33013
rect 23427 32948 23428 33012
rect 23492 32948 23493 33012
rect 23427 32947 23493 32948
rect 23430 32333 23490 32947
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 23427 32332 23493 32333
rect 23427 32268 23428 32332
rect 23492 32268 23493 32332
rect 23427 32267 23493 32268
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 23430 27029 23490 32267
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 23427 27028 23493 27029
rect 23427 26964 23428 27028
rect 23492 26964 23493 27028
rect 23427 26963 23493 26964
rect 23430 26836 23490 26963
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2128 35248 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_84
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_90
timestamp 1586364061
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_87 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
timestamp 1586364061
transform 1 0 9200 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_105
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 314 592
use scs8hd_dfbbp_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 2430 592
use scs8hd_fill_2  FILLER_0_109
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_119
timestamp 1586364061
transform 1 0 12052 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
timestamp 1586364061
transform 1 0 12604 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_130
timestamp 1586364061
transform 1 0 13064 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12788 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_134
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_conb_1  _430_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_140
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_136
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14352 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_160
timestamp 1586364061
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15640 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_dfbbp_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 2430 592
use scs8hd_fill_2  FILLER_1_168
timestamp 1586364061
transform 1 0 16560 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_164
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 16008 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 2720
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 16192 0 -1 2720
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_175
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_179
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18216 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_188
timestamp 1586364061
transform 1 0 18400 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18676 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18492 0 -1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_206
timestamp 1586364061
transform 1 0 20056 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_202
timestamp 1586364061
transform 1 0 19688 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__409__B
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_214
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__409__A
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
timestamp 1586364061
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
timestamp 1586364061
transform 1 0 21344 0 -1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
timestamp 1586364061
transform 1 0 21160 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_239
timestamp 1586364061
transform 1 0 23092 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_235
timestamp 1586364061
transform 1 0 22724 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_229
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_231
timestamp 1586364061
transform 1 0 22356 0 -1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22908 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
timestamp 1586364061
transform 1 0 22540 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23276 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_248
timestamp 1586364061
transform 1 0 23920 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_243
timestamp 1586364061
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_247
timestamp 1586364061
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_243
timestamp 1586364061
transform 1 0 23460 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_252
timestamp 1586364061
transform 1 0 24288 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_255
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24380 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24748 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24656 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_265
timestamp 1586364061
transform 1 0 25484 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_268
timestamp 1586364061
transform 1 0 25760 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25668 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_273
timestamp 1586364061
transform 1 0 26220 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_272
timestamp 1586364061
transform 1 0 26128 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26036 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26404 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26588 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26588 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_284
timestamp 1586364061
transform 1 0 27232 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_280
timestamp 1586364061
transform 1 0 26864 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27048 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27416 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 1 2720
box -38 -48 866 592
use scs8hd_decap_6  FILLER_0_289
timestamp 1586364061
transform 1 0 27692 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28244 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_301
timestamp 1586364061
transform 1 0 28796 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_297
timestamp 1586364061
transform 1 0 28428 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_300
timestamp 1586364061
transform 1 0 28704 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28980 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28612 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28428 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_311
timestamp 1586364061
transform 1 0 29716 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_306
timestamp 1586364061
transform 1 0 29256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29900 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29440 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29440 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_315
timestamp 1586364061
transform 1 0 30084 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_320
timestamp 1586364061
transform 1 0 30544 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30268 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30452 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_328
timestamp 1586364061
transform 1 0 31280 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_328
timestamp 1586364061
transform 1 0 31280 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_324
timestamp 1586364061
transform 1 0 30912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31096 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31464 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_334
timestamp 1586364061
transform 1 0 31832 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_337
timestamp 1586364061
transform 1 0 32108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_333
timestamp 1586364061
transform 1 0 31740 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 32292 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 31648 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32016 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_8  _150_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 32200 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_347
timestamp 1586364061
transform 1 0 33028 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _149_
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_358
timestamp 1586364061
transform 1 0 34040 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_351
timestamp 1586364061
transform 1 0 33396 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_356
timestamp 1586364061
transform 1 0 33856 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_351
timestamp 1586364061
transform 1 0 33396 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33672 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33212 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33580 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33764 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_362
timestamp 1586364061
transform 1 0 34408 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_362
timestamp 1586364061
transform 1 0 34408 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 34592 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 34592 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 34132 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_371
timestamp 1586364061
transform 1 0 35236 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 35328 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35144 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _151_
timestamp 1586364061
transform 1 0 35512 0 1 2720
box -38 -48 866 592
use scs8hd_decap_6  FILLER_1_383
timestamp 1586364061
transform 1 0 36340 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_382
timestamp 1586364061
transform 1 0 36248 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36432 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_393
timestamp 1586364061
transform 1 0 37260 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_386
timestamp 1586364061
transform 1 0 36616 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37444 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36892 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36984 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_400
timestamp 1586364061
transform 1 0 37904 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 38088 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 40388 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_416
timestamp 1586364061
transform 1 0 39376 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_428
timestamp 1586364061
transform 1 0 40480 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_404
timestamp 1586364061
transform 1 0 38272 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_416
timestamp 1586364061
transform 1 0 39376 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  FILLER_1_424
timestamp 1586364061
transform 1 0 40112 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_428
timestamp 1586364061
transform 1 0 40480 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 41032 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_435
timestamp 1586364061
transform 1 0 41124 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_447
timestamp 1586364061
transform 1 0 42228 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_440
timestamp 1586364061
transform 1 0 41584 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_452
timestamp 1586364061
transform 1 0 42688 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 43884 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_459
timestamp 1586364061
transform 1 0 43332 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_466
timestamp 1586364061
transform 1 0 43976 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_478
timestamp 1586364061
transform 1 0 45080 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_464
timestamp 1586364061
transform 1 0 43792 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_476
timestamp 1586364061
transform 1 0 44896 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 46736 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 46000 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_490
timestamp 1586364061
transform 1 0 46184 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_497
timestamp 1586364061
transform 1 0 46828 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_509
timestamp 1586364061
transform 1 0 47932 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_489
timestamp 1586364061
transform 1 0 46092 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_501
timestamp 1586364061
transform 1 0 47196 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 48852 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 48852 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_515
timestamp 1586364061
transform 1 0 48484 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_513
timestamp 1586364061
transform 1 0 48300 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_90
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use scs8hd_dfbbp_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 2430 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_109
timestamp 1586364061
transform 1 0 11132 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_113
timestamp 1586364061
transform 1 0 11500 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_SETB
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_143
timestamp 1586364061
transform 1 0 14260 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_147
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_151
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16192 0 -1 3808
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17940 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16008 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_175
timestamp 1586364061
transform 1 0 17204 0 -1 3808
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19504 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_192
timestamp 1586364061
transform 1 0 18768 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_196
timestamp 1586364061
transform 1 0 19136 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_203
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_211
timestamp 1586364061
transform 1 0 20516 0 -1 3808
box -38 -48 130 592
use scs8hd_nor2_4  _409_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
timestamp 1586364061
transform 1 0 22540 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_224
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_228
timestamp 1586364061
transform 1 0 22080 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_232
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 23736 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24104 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_244
timestamp 1586364061
transform 1 0 23552 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_248
timestamp 1586364061
transform 1 0 23920 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_252
timestamp 1586364061
transform 1 0 24288 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_267
timestamp 1586364061
transform 1 0 25668 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_271
timestamp 1586364061
transform 1 0 26036 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25852 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_287
timestamp 1586364061
transform 1 0 27508 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_283
timestamp 1586364061
transform 1 0 27140 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_279
timestamp 1586364061
transform 1 0 26772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26956 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27600 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_290
timestamp 1586364061
transform 1 0 27784 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27968 0 -1 3808
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30452 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29256 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29624 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_301
timestamp 1586364061
transform 1 0 28796 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_305
timestamp 1586364061
transform 1 0 29164 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_308
timestamp 1586364061
transform 1 0 29440 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_312
timestamp 1586364061
transform 1 0 29808 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_318
timestamp 1586364061
transform 1 0 30360 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33120 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_328
timestamp 1586364061
transform 1 0 31280 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_346
timestamp 1586364061
transform 1 0 32936 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _152_
timestamp 1586364061
transform 1 0 35512 0 -1 3808
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33672 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34684 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_350
timestamp 1586364061
transform 1 0 33304 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_363
timestamp 1586364061
transform 1 0 34500 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_367
timestamp 1586364061
transform 1 0 34868 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_373
timestamp 1586364061
transform 1 0 35420 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36524 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37076 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_383
timestamp 1586364061
transform 1 0 36340 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_387
timestamp 1586364061
transform 1 0 36708 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_2_393
timestamp 1586364061
transform 1 0 37260 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_401
timestamp 1586364061
transform 1 0 37996 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_413
timestamp 1586364061
transform 1 0 39100 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_425
timestamp 1586364061
transform 1 0 40204 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_437
timestamp 1586364061
transform 1 0 41308 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_449
timestamp 1586364061
transform 1 0 42412 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 43240 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_457
timestamp 1586364061
transform 1 0 43148 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_459
timestamp 1586364061
transform 1 0 43332 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_471
timestamp 1586364061
transform 1 0 44436 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_483
timestamp 1586364061
transform 1 0 45540 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_495
timestamp 1586364061
transform 1 0 46644 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_507
timestamp 1586364061
transform 1 0 47748 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 48852 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_515
timestamp 1586364061
transform 1 0 48484 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__213__A
timestamp 1586364061
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__213__B
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_94
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_102
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 314 592
use scs8hd_or2_4  _177_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_130
timestamp 1586364061
transform 1 0 13064 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_134
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_dfbbp_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 2430 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_CLK
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_168
timestamp 1586364061
transform 1 0 16560 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_164
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__404__B
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__404__A
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_fill_2  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__211__A
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_204
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__211__B
timestamp 1586364061
transform 1 0 20056 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23092 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__408__A
timestamp 1586364061
transform 1 0 21988 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__408__B
timestamp 1586364061
transform 1 0 22356 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_225
timestamp 1586364061
transform 1 0 21804 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_229
timestamp 1586364061
transform 1 0 22172 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_236
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_241
timestamp 1586364061
transform 1 0 23276 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_256
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_260
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_264
timestamp 1586364061
transform 1 0 25392 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
timestamp 1586364061
transform 1 0 26772 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 26588 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26220 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_275
timestamp 1586364061
transform 1 0 26404 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_290
timestamp 1586364061
transform 1 0 27784 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_295
timestamp 1586364061
transform 1 0 28244 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30636 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30268 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28612 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_301
timestamp 1586364061
transform 1 0 28796 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_315
timestamp 1586364061
transform 1 0 30084 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_319
timestamp 1586364061
transform 1 0 30452 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32384 0 1 3808
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30820 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32200 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31832 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_332
timestamp 1586364061
transform 1 0 31648 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_336
timestamp 1586364061
transform 1 0 32016 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33948 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33396 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_349
timestamp 1586364061
transform 1 0 33212 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_353
timestamp 1586364061
transform 1 0 33580 0 1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_3_359
timestamp 1586364061
transform 1 0 34132 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_363
timestamp 1586364061
transform 1 0 34500 0 1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 3808
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37996 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36248 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37812 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 35880 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_376
timestamp 1586364061
transform 1 0 35696 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_380
timestamp 1586364061
transform 1 0 36064 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_393
timestamp 1586364061
transform 1 0 37260 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 40388 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_410
timestamp 1586364061
transform 1 0 38824 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_3_422
timestamp 1586364061
transform 1 0 39928 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_426
timestamp 1586364061
transform 1 0 40296 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_428
timestamp 1586364061
transform 1 0 40480 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_440
timestamp 1586364061
transform 1 0 41584 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_452
timestamp 1586364061
transform 1 0 42688 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_464
timestamp 1586364061
transform 1 0 43792 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_476
timestamp 1586364061
transform 1 0 44896 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 46000 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_489
timestamp 1586364061
transform 1 0 46092 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_501
timestamp 1586364061
transform 1 0 47196 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 48852 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_513
timestamp 1586364061
transform 1 0 48300 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_nor2_4  _213_
timestamp 1586364061
transform 1 0 10304 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_99
timestamp 1586364061
transform 1 0 10212 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_113
timestamp 1586364061
transform 1 0 11500 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_109
timestamp 1586364061
transform 1 0 11132 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11316 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_124
timestamp 1586364061
transform 1 0 12512 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_120
timestamp 1586364061
transform 1 0 12144 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_131
timestamp 1586364061
transform 1 0 13156 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_128
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__214__B
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 866 592
use scs8hd_fill_2  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_RESETB
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__ff_0.DFFSRQ_0_.dff_D
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__405__A
timestamp 1586364061
transform 1 0 15548 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_159
timestamp 1586364061
transform 1 0 15732 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__403__B
timestamp 1586364061
transform 1 0 15916 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _404_
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16100 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_174
timestamp 1586364061
transform 1 0 17112 0 -1 4896
box -38 -48 590 592
use scs8hd_or2_4  _211_
timestamp 1586364061
transform 1 0 19412 0 -1 4896
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__410__B
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_191
timestamp 1586364061
transform 1 0 18676 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_195
timestamp 1586364061
transform 1 0 19044 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_219
timestamp 1586364061
transform 1 0 21252 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__411__B
timestamp 1586364061
transform 1 0 21068 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _408_
timestamp 1586364061
transform 1 0 21436 0 -1 4896
box -38 -48 866 592
use scs8hd_fill_1  FILLER_4_238
timestamp 1586364061
transform 1 0 23000 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_234
timestamp 1586364061
transform 1 0 22632 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_230
timestamp 1586364061
transform 1 0 22264 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22816 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__423__B
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24288 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_250
timestamp 1586364061
transform 1 0 24104 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_254
timestamp 1586364061
transform 1 0 24472 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_267
timestamp 1586364061
transform 1 0 25668 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28060 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27508 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_285
timestamp 1586364061
transform 1 0 27324 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_289
timestamp 1586364061
transform 1 0 27692 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
timestamp 1586364061
transform 1 0 29072 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30268 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28888 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_296
timestamp 1586364061
transform 1 0 28336 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_2  FILLER_4_315
timestamp 1586364061
transform 1 0 30084 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_319
timestamp 1586364061
transform 1 0 30452 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31004 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32384 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30820 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_328
timestamp 1586364061
transform 1 0 31280 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_337
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33948 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34960 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_349
timestamp 1586364061
transform 1 0 33212 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_366
timestamp 1586364061
transform 1 0 34776 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_370
timestamp 1586364061
transform 1 0 35144 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_8  _153_
timestamp 1586364061
transform 1 0 36064 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 35880 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37996 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_389
timestamp 1586364061
transform 1 0 36892 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_403
timestamp 1586364061
transform 1 0 38180 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_415
timestamp 1586364061
transform 1 0 39284 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_427
timestamp 1586364061
transform 1 0 40388 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_439
timestamp 1586364061
transform 1 0 41492 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_4_451
timestamp 1586364061
transform 1 0 42596 0 -1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 43240 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_457
timestamp 1586364061
transform 1 0 43148 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_459
timestamp 1586364061
transform 1 0 43332 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_471
timestamp 1586364061
transform 1 0 44436 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_483
timestamp 1586364061
transform 1 0 45540 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_495
timestamp 1586364061
transform 1 0 46644 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_507
timestamp 1586364061
transform 1 0 47748 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 48852 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_515
timestamp 1586364061
transform 1 0 48484 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_conb_1  _428_
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 590 592
use scs8hd_fill_2  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_99
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13156 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__214__A
timestamp 1586364061
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _403_
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__403__A
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__405__B
timestamp 1586364061
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_142
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_146
timestamp 1586364061
transform 1 0 14536 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_150
timestamp 1586364061
transform 1 0 14904 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_153
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_166
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_172
timestamp 1586364061
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_176
timestamp 1586364061
transform 1 0 17296 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_180
timestamp 1586364061
transform 1 0 17664 0 1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _410_
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__410__A
timestamp 1586364061
transform 1 0 20056 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_195
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_199
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_205
timestamp 1586364061
transform 1 0 19964 0 1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _423_
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__411__A
timestamp 1586364061
transform 1 0 21252 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__422__A
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__423__A
timestamp 1586364061
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__422__B
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_217
timestamp 1586364061
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_221
timestamp 1586364061
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_234
timestamp 1586364061
transform 1 0 22632 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_238
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
timestamp 1586364061
transform 1 0 24564 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 24380 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24012 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_242
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_251
timestamp 1586364061
transform 1 0 24196 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_266
timestamp 1586364061
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28060 0 1 4896
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
timestamp 1586364061
transform 1 0 26312 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 26128 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 27508 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27876 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_270
timestamp 1586364061
transform 1 0 25944 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_285
timestamp 1586364061
transform 1 0 27324 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_289
timestamp 1586364061
transform 1 0 27692 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_300
timestamp 1586364061
transform 1 0 28704 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_296
timestamp 1586364061
transform 1 0 28336 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28520 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  FILLER_5_319
timestamp 1586364061
transform 1 0 30452 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_315
timestamp 1586364061
transform 1 0 30084 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 30268 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
timestamp 1586364061
transform 1 0 30728 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _413_
timestamp 1586364061
transform 1 0 32660 0 1 4896
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
timestamp 1586364061
transform 1 0 30912 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__413__A
timestamp 1586364061
transform 1 0 32476 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__418__A
timestamp 1586364061
transform 1 0 32108 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_335
timestamp 1586364061
transform 1 0 31924 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_339
timestamp 1586364061
transform 1 0 32292 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_352
timestamp 1586364061
transform 1 0 33488 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_356
timestamp 1586364061
transform 1 0 33856 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 34040 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__418__B
timestamp 1586364061
transform 1 0 33672 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_360
timestamp 1586364061
transform 1 0 34224 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34592 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_370
timestamp 1586364061
transform 1 0 35144 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_374
timestamp 1586364061
transform 1 0 35512 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35604 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _154_
timestamp 1586364061
transform 1 0 35880 0 1 4896
box -38 -48 866 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 37444 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 37904 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36892 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_377
timestamp 1586364061
transform 1 0 35788 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_387
timestamp 1586364061
transform 1 0 36708 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_391
timestamp 1586364061
transform 1 0 37076 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_398
timestamp 1586364061
transform 1 0 37720 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_402
timestamp 1586364061
transform 1 0 38088 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 40388 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38272 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_406
timestamp 1586364061
transform 1 0 38456 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_418
timestamp 1586364061
transform 1 0 39560 0 1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_5_426
timestamp 1586364061
transform 1 0 40296 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_428
timestamp 1586364061
transform 1 0 40480 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_440
timestamp 1586364061
transform 1 0 41584 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_452
timestamp 1586364061
transform 1 0 42688 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_464
timestamp 1586364061
transform 1 0 43792 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_476
timestamp 1586364061
transform 1 0 44896 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 46000 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_489
timestamp 1586364061
transform 1 0 46092 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_501
timestamp 1586364061
transform 1 0 47196 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 48852 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_513
timestamp 1586364061
transform 1 0 48300 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_90
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__381__B
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__212__B
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_94
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_100
timestamp 1586364061
transform 1 0 10304 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_97
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__212__A
timestamp 1586364061
transform 1 0 10120 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__381__A
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 1050 592
use scs8hd_nor2_4  _212_
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 866 592
use scs8hd_decap_8  FILLER_7_107
timestamp 1586364061
transform 1 0 10948 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_115
timestamp 1586364061
transform 1 0 11684 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_113
timestamp 1586364061
transform 1 0 11500 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_125
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_121
timestamp 1586364061
transform 1 0 12236 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__383__B
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__383__A
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use scs8hd_decap_6  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 590 592
use scs8hd_nor2_4  _214_
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_141
timestamp 1586364061
transform 1 0 14076 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_138
timestamp 1586364061
transform 1 0 13800 0 -1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _125_
timestamp 1586364061
transform 1 0 14444 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_158
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_154
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_150
timestamp 1586364061
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__425__B
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _405_
timestamp 1586364061
transform 1 0 15548 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__425__A
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 774 592
use scs8hd_nor2_4  _425_
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_187
timestamp 1586364061
transform 1 0 18308 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_183
timestamp 1586364061
transform 1 0 17940 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18124 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__426__A
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _426_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_200
timestamp 1586364061
transform 1 0 19504 0 -1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_204
timestamp 1586364061
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__389__B
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__389__A
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 314 592
use scs8hd_nor2_4  _389_
timestamp 1586364061
transform 1 0 20608 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_226
timestamp 1586364061
transform 1 0 21896 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_221
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
timestamp 1586364061
transform 1 0 21712 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _411_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_231
timestamp 1586364061
transform 1 0 22356 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_228
timestamp 1586364061
transform 1 0 22080 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__402__B
timestamp 1586364061
transform 1 0 22172 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__402__A
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _422_
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 866 592
use scs8hd_or2_4  _402_
timestamp 1586364061
transform 1 0 22172 0 1 5984
box -38 -48 682 592
use scs8hd_decap_12  FILLER_6_241
timestamp 1586364061
transform 1 0 23276 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_249
timestamp 1586364061
transform 1 0 24012 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__400__B
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__400__A
timestamp 1586364061
transform 1 0 23828 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_253
timestamp 1586364061
transform 1 0 24380 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__420__B
timestamp 1586364061
transform 1 0 24472 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__420__A
timestamp 1586364061
transform 1 0 24288 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24656 0 -1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _420_
timestamp 1586364061
transform 1 0 24472 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_267
timestamp 1586364061
transform 1 0 25668 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_263
timestamp 1586364061
transform 1 0 25300 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_265
timestamp 1586364061
transform 1 0 25484 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_280
timestamp 1586364061
transform 1 0 26864 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_280
timestamp 1586364061
transform 1 0 26864 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_273
timestamp 1586364061
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__421__B
timestamp 1586364061
transform 1 0 26036 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__398__B
timestamp 1586364061
transform 1 0 26680 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__421__A
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _421_
timestamp 1586364061
transform 1 0 26036 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_284
timestamp 1586364061
transform 1 0 27232 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__398__A
timestamp 1586364061
transform 1 0 27048 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27416 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
timestamp 1586364061
transform 1 0 27048 0 -1 5984
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_6_293
timestamp 1586364061
transform 1 0 28060 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28612 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28612 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_301
timestamp 1586364061
transform 1 0 28796 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_297
timestamp 1586364061
transform 1 0 28428 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_301
timestamp 1586364061
transform 1 0 28796 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29256 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_305
timestamp 1586364061
transform 1 0 29164 0 -1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_315
timestamp 1586364061
transform 1 0 30084 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__419__A
timestamp 1586364061
transform 1 0 30268 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
timestamp 1586364061
transform 1 0 29440 0 -1 5984
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_7_319
timestamp 1586364061
transform 1 0 30452 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_319
timestamp 1586364061
transform 1 0 30452 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__419__B
timestamp 1586364061
transform 1 0 30636 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
timestamp 1586364061
transform 1 0 30728 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_333
timestamp 1586364061
transform 1 0 31740 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_327
timestamp 1586364061
transform 1 0 31188 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_6_323
timestamp 1586364061
transform 1 0 30820 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31004 0 -1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
timestamp 1586364061
transform 1 0 30912 0 1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_345
timestamp 1586364061
transform 1 0 32844 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_339
timestamp 1586364061
transform 1 0 32292 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_335
timestamp 1586364061
transform 1 0 31924 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31832 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32660 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
timestamp 1586364061
transform 1 0 32108 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _418_
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_346
timestamp 1586364061
transform 1 0 32936 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__413__B
timestamp 1586364061
transform 1 0 33120 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33028 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_358
timestamp 1586364061
transform 1 0 34040 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_354
timestamp 1586364061
transform 1 0 33672 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_350
timestamp 1586364061
transform 1 0 33304 0 -1 5984
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 5984
box -38 -48 866 592
use scs8hd_inv_8  _148_
timestamp 1586364061
transform 1 0 33764 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_362
timestamp 1586364061
transform 1 0 34408 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_364
timestamp 1586364061
transform 1 0 34592 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 34592 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_inv_8  _147_
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 866 592
use scs8hd_decap_3  FILLER_6_372
timestamp 1586364061
transform 1 0 35328 0 -1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35604 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_387
timestamp 1586364061
transform 1 0 36708 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_380
timestamp 1586364061
transform 1 0 36064 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_376
timestamp 1586364061
transform 1 0 35696 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_384
timestamp 1586364061
transform 1 0 36432 0 -1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35880 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36432 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36892 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37260 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_391
timestamp 1586364061
transform 1 0 37076 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37444 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 37904 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_396
timestamp 1586364061
transform 1 0 37536 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_398
timestamp 1586364061
transform 1 0 37720 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_401
timestamp 1586364061
transform 1 0 37996 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_402
timestamp 1586364061
transform 1 0 38088 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 40388 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38272 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_413
timestamp 1586364061
transform 1 0 39100 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_425
timestamp 1586364061
transform 1 0 40204 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_406
timestamp 1586364061
transform 1 0 38456 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_418
timestamp 1586364061
transform 1 0 39560 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_426
timestamp 1586364061
transform 1 0 40296 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_428
timestamp 1586364061
transform 1 0 40480 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_437
timestamp 1586364061
transform 1 0 41308 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_449
timestamp 1586364061
transform 1 0 42412 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_440
timestamp 1586364061
transform 1 0 41584 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_452
timestamp 1586364061
transform 1 0 42688 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 43240 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_457
timestamp 1586364061
transform 1 0 43148 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_459
timestamp 1586364061
transform 1 0 43332 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_471
timestamp 1586364061
transform 1 0 44436 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_483
timestamp 1586364061
transform 1 0 45540 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_464
timestamp 1586364061
transform 1 0 43792 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_476
timestamp 1586364061
transform 1 0 44896 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 46000 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_495
timestamp 1586364061
transform 1 0 46644 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_507
timestamp 1586364061
transform 1 0 47748 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_489
timestamp 1586364061
transform 1 0 46092 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_501
timestamp 1586364061
transform 1 0 47196 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 48852 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 48852 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_515
timestamp 1586364061
transform 1 0 48484 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_513
timestamp 1586364061
transform 1 0 48300 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 774 592
use scs8hd_nor2_4  _381_
timestamp 1586364061
transform 1 0 9936 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _383_
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_109
timestamp 1586364061
transform 1 0 11132 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_120
timestamp 1586364061
transform 1 0 12144 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_132
timestamp 1586364061
transform 1 0 13248 0 -1 7072
box -38 -48 774 592
use scs8hd_conb_1  _429_
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_143
timestamp 1586364061
transform 1 0 14260 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_151
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_160
timestamp 1586364061
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16560 0 -1 7072
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__207__C
timestamp 1586364061
transform 1 0 16008 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__426__B
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_164
timestamp 1586364061
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_179
timestamp 1586364061
transform 1 0 17572 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_183
timestamp 1586364061
transform 1 0 17940 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__407__B
timestamp 1586364061
transform 1 0 19412 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_196
timestamp 1586364061
transform 1 0 19136 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_201
timestamp 1586364061
transform 1 0 19596 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_213
timestamp 1586364061
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__417__B
timestamp 1586364061
transform 1 0 22908 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21528 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_219
timestamp 1586364061
transform 1 0 21252 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_235
timestamp 1586364061
transform 1 0 22724 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 406 592
use scs8hd_nor2_4  _400_
timestamp 1586364061
transform 1 0 23460 0 -1 7072
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24472 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_252
timestamp 1586364061
transform 1 0 24288 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_256
timestamp 1586364061
transform 1 0 24656 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 774 592
use scs8hd_nor2_4  _398_
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27600 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_271
timestamp 1586364061
transform 1 0 26036 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_285
timestamp 1586364061
transform 1 0 27324 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_290
timestamp 1586364061
transform 1 0 27784 0 -1 7072
box -38 -48 774 592
use scs8hd_nor2_4  _419_
timestamp 1586364061
transform 1 0 30176 0 -1 7072
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28612 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29624 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_298
timestamp 1586364061
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_308
timestamp 1586364061
transform 1 0 29440 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_312
timestamp 1586364061
transform 1 0 29808 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31832 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31188 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_325
timestamp 1586364061
transform 1 0 31004 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_329
timestamp 1586364061
transform 1 0 31372 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_333
timestamp 1586364061
transform 1 0 31740 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_8_348
timestamp 1586364061
transform 1 0 33120 0 -1 7072
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35420 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33856 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33672 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_365
timestamp 1586364061
transform 1 0 34684 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_383
timestamp 1586364061
transform 1 0 36340 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_380
timestamp 1586364061
transform 1 0 36064 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_376
timestamp 1586364061
transform 1 0 35696 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36156 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36432 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_8_391
timestamp 1586364061
transform 1 0 37076 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_2  FILLER_8_387
timestamp 1586364061
transform 1 0 36708 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36892 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_8  _146_
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_12  FILLER_8_407
timestamp 1586364061
transform 1 0 38548 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_419
timestamp 1586364061
transform 1 0 39652 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_431
timestamp 1586364061
transform 1 0 40756 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_443
timestamp 1586364061
transform 1 0 41860 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_8_455
timestamp 1586364061
transform 1 0 42964 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 43240 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_459
timestamp 1586364061
transform 1 0 43332 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_471
timestamp 1586364061
transform 1 0 44436 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_483
timestamp 1586364061
transform 1 0 45540 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_495
timestamp 1586364061
transform 1 0 46644 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_507
timestamp 1586364061
transform 1 0 47748 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 48852 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_515
timestamp 1586364061
transform 1 0 48484 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_78
timestamp 1586364061
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use scs8hd_or2_4  _171_
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 682 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_88
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_92
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_107
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_111
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_115
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_134
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_142
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_138
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__B
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_150
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_146
timestamp 1586364061
transform 1 0 14536 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__D
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use scs8hd_or4_4  _205_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 866 592
use scs8hd_fill_2  FILLER_9_167
timestamp 1586364061
transform 1 0 16468 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_163
timestamp 1586364061
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__207__D
timestamp 1586364061
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__207__B
timestamp 1586364061
transform 1 0 16284 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__427__A
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__427__B
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_inv_8  _126_
timestamp 1586364061
transform 1 0 18952 0 1 7072
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20792 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__407__A
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 18768 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__401__B
timestamp 1586364061
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_203
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_207
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_211
timestamp 1586364061
transform 1 0 20516 0 1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21804 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__417__A
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__401__A
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_217
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_221
timestamp 1586364061
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_240
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_256
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_260
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_267
timestamp 1586364061
transform 1 0 25668 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
timestamp 1586364061
transform 1 0 26772 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 26588 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26220 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27968 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_271
timestamp 1586364061
transform 1 0 26036 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_275
timestamp 1586364061
transform 1 0 26404 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_290
timestamp 1586364061
transform 1 0 27784 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_294
timestamp 1586364061
transform 1 0 28152 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_302
timestamp 1586364061
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_298
timestamp 1586364061
transform 1 0 28520 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28336 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__397__B
timestamp 1586364061
transform 1 0 28980 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_310
timestamp 1586364061
transform 1 0 29624 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_306
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__397__A
timestamp 1586364061
transform 1 0 29440 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__412__A
timestamp 1586364061
transform 1 0 29900 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _412_
timestamp 1586364061
transform 1 0 30084 0 1 7072
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
timestamp 1586364061
transform 1 0 31832 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
timestamp 1586364061
transform 1 0 31648 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__414__A
timestamp 1586364061
transform 1 0 31280 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__414__B
timestamp 1586364061
transform 1 0 33028 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_324
timestamp 1586364061
transform 1 0 30912 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_330
timestamp 1586364061
transform 1 0 31464 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_345
timestamp 1586364061
transform 1 0 32844 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_349
timestamp 1586364061
transform 1 0 33212 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 33396 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 33580 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_356
timestamp 1586364061
transform 1 0 33856 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_361
timestamp 1586364061
transform 1 0 34316 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34500 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34132 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_365
timestamp 1586364061
transform 1 0 34684 0 1 7072
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_370
timestamp 1586364061
transform 1 0 35144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35328 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_374
timestamp 1586364061
transform 1 0 35512 0 1 7072
box -38 -48 406 592
use scs8hd_inv_8  _145_
timestamp 1586364061
transform 1 0 37720 0 1 7072
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36156 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35972 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37536 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 37168 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_378
timestamp 1586364061
transform 1 0 35880 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_390
timestamp 1586364061
transform 1 0 36984 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_394
timestamp 1586364061
transform 1 0 37352 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 40388 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39284 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38732 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_407
timestamp 1586364061
transform 1 0 38548 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_411
timestamp 1586364061
transform 1 0 38916 0 1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_9_417
timestamp 1586364061
transform 1 0 39468 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_425
timestamp 1586364061
transform 1 0 40204 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_428
timestamp 1586364061
transform 1 0 40480 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_440
timestamp 1586364061
transform 1 0 41584 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_452
timestamp 1586364061
transform 1 0 42688 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_464
timestamp 1586364061
transform 1 0 43792 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_476
timestamp 1586364061
transform 1 0 44896 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 46000 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_489
timestamp 1586364061
transform 1 0 46092 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_501
timestamp 1586364061
transform 1 0 47196 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 48852 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_513
timestamp 1586364061
transform 1 0 48300 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 130 592
use scs8hd_conb_1  _431_
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__382__A
timestamp 1586364061
transform 1 0 10028 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_4  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_99
timestamp 1586364061
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11960 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_110
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_4  FILLER_10_127
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_131
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_134
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _124_
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use scs8hd_or4_4  _207_
timestamp 1586364061
transform 1 0 15824 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__205__C
timestamp 1586364061
transform 1 0 15456 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_158
timestamp 1586364061
transform 1 0 15640 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _427_
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_1.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_169
timestamp 1586364061
transform 1 0 16652 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_174
timestamp 1586364061
transform 1 0 17112 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_6  FILLER_10_186
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 590 592
use scs8hd_or2_4  _407_
timestamp 1586364061
transform 1 0 19412 0 -1 8160
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__424__B
timestamp 1586364061
transform 1 0 18768 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_194
timestamp 1586364061
transform 1 0 18952 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_198
timestamp 1586364061
transform 1 0 19320 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 774 592
use scs8hd_nor2_4  _401_
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use scs8hd_nor2_4  _417_
timestamp 1586364061
transform 1 0 22632 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_228
timestamp 1586364061
transform 1 0 22080 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25668 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24012 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_243
timestamp 1586364061
transform 1 0 23460 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_247
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_260
timestamp 1586364061
transform 1 0 25024 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_266
timestamp 1586364061
transform 1 0 25576 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28060 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27600 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_269
timestamp 1586364061
transform 1 0 25852 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_3  FILLER_10_285
timestamp 1586364061
transform 1 0 27324 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_290
timestamp 1586364061
transform 1 0 27784 0 -1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _397_
timestamp 1586364061
transform 1 0 29256 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__415__B
timestamp 1586364061
transform 1 0 30268 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__412__B
timestamp 1586364061
transform 1 0 30636 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_296
timestamp 1586364061
transform 1 0 28336 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_304
timestamp 1586364061
transform 1 0 29072 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_315
timestamp 1586364061
transform 1 0 30084 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_319
timestamp 1586364061
transform 1 0 30452 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _414_
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30912 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31372 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_323
timestamp 1586364061
transform 1 0 30820 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_327
timestamp 1586364061
transform 1 0 31188 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_331
timestamp 1586364061
transform 1 0 31556 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_335
timestamp 1586364061
transform 1 0 31924 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_346
timestamp 1586364061
transform 1 0 32936 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34132 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33948 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33212 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35512 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_351
timestamp 1586364061
transform 1 0 33396 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_6  FILLER_10_368
timestamp 1586364061
transform 1 0 34960 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36064 0 -1 8160
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35880 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_376
timestamp 1586364061
transform 1 0 35696 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_389
timestamp 1586364061
transform 1 0 36892 0 -1 8160
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39284 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_407
timestamp 1586364061
transform 1 0 38548 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_12  FILLER_10_418
timestamp 1586364061
transform 1 0 39560 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_430
timestamp 1586364061
transform 1 0 40664 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_442
timestamp 1586364061
transform 1 0 41768 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_454
timestamp 1586364061
transform 1 0 42872 0 -1 8160
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 43240 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_459
timestamp 1586364061
transform 1 0 43332 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_471
timestamp 1586364061
transform 1 0 44436 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_483
timestamp 1586364061
transform 1 0 45540 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_495
timestamp 1586364061
transform 1 0 46644 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_507
timestamp 1586364061
transform 1 0 47748 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 48852 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_515
timestamp 1586364061
transform 1 0 48484 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_80
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _382_
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__382__B
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_83
timestamp 1586364061
transform 1 0 8740 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_89
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_93
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_106
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_11_115
timestamp 1586364061
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 11868 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_119
timestamp 1586364061
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_128
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__C
timestamp 1586364061
transform 1 0 13064 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _123_
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 866 592
use scs8hd_or3_4  _198_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__198__C
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__B
timestamp 1586364061
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_141
timestamp 1586364061
transform 1 0 14076 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_145
timestamp 1586364061
transform 1 0 14444 0 1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_11_153
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_157
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__198__B
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__380__A
timestamp 1586364061
transform 1 0 18216 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__380__B
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_170
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_178
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_188
timestamp 1586364061
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__424__A
timestamp 1586364061
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use scs8hd_or2_4  _424_
timestamp 1586364061
transform 1 0 18768 0 1 8160
box -38 -48 682 592
use scs8hd_fill_2  FILLER_11_203
timestamp 1586364061
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_199
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__385__A
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_211
timestamp 1586364061
transform 1 0 20516 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_207
timestamp 1586364061
transform 1 0 20148 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__385__B
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_214
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__386__B
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _386_
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__386__A
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_227
timestamp 1586364061
transform 1 0 21988 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_231
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_235
timestamp 1586364061
transform 1 0 22724 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_241
timestamp 1586364061
transform 1 0 23276 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 1 8160
box -38 -48 866 592
use scs8hd_fill_2  FILLER_11_259
timestamp 1586364061
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_263
timestamp 1586364061
transform 1 0 25300 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 26772 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27416 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_276
timestamp 1586364061
transform 1 0 26496 0 1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_11_281
timestamp 1586364061
transform 1 0 26956 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_285
timestamp 1586364061
transform 1 0 27324 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_306
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_301
timestamp 1586364061
transform 1 0 28796 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_297
timestamp 1586364061
transform 1 0 28428 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__396__B
timestamp 1586364061
transform 1 0 28980 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__396__A
timestamp 1586364061
transform 1 0 28612 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_315
timestamp 1586364061
transform 1 0 30084 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_311
timestamp 1586364061
transform 1 0 29716 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__415__A
timestamp 1586364061
transform 1 0 29900 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 30268 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
timestamp 1586364061
transform 1 0 30452 0 1 8160
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32200 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32660 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33028 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32016 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31648 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_330
timestamp 1586364061
transform 1 0 31464 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_334
timestamp 1586364061
transform 1 0 31832 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_341
timestamp 1586364061
transform 1 0 32476 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_345
timestamp 1586364061
transform 1 0 32844 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_358
timestamp 1586364061
transform 1 0 34040 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_362
timestamp 1586364061
transform 1 0 34408 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_380
timestamp 1586364061
transform 1 0 36064 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_376
timestamp 1586364061
transform 1 0 35696 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36248 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 8160
box -38 -48 866 592
use scs8hd_decap_4  FILLER_11_393
timestamp 1586364061
transform 1 0 37260 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_400
timestamp 1586364061
transform 1 0 37904 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_397
timestamp 1586364061
transform 1 0 37628 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37720 0 1 8160
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 37996 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 40388 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 38456 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38824 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_404
timestamp 1586364061
transform 1 0 38272 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_408
timestamp 1586364061
transform 1 0 38640 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_412
timestamp 1586364061
transform 1 0 39008 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_11_424
timestamp 1586364061
transform 1 0 40112 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_428
timestamp 1586364061
transform 1 0 40480 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_440
timestamp 1586364061
transform 1 0 41584 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_452
timestamp 1586364061
transform 1 0 42688 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_464
timestamp 1586364061
transform 1 0 43792 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_476
timestamp 1586364061
transform 1 0 44896 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 46000 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_489
timestamp 1586364061
transform 1 0 46092 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_501
timestamp 1586364061
transform 1 0 47196 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 48852 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_513
timestamp 1586364061
transform 1 0 48300 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mem_ble4_out_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_116
timestamp 1586364061
transform 1 0 11776 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_112
timestamp 1586364061
transform 1 0 11408 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_108
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__B
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use scs8hd_or2_4  _174_
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 682 592
use scs8hd_fill_2  FILLER_12_124
timestamp 1586364061
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__D
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_128
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 13064 0 -1 9248
box -38 -48 222 592
use scs8hd_or3_4  _195_
timestamp 1586364061
transform 1 0 13248 0 -1 9248
box -38 -48 866 592
use scs8hd_or3_4  _168_
timestamp 1586364061
transform 1 0 15640 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 15456 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 222 592
use scs8hd_or2_4  _380_
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 682 592
use scs8hd_decap_12  FILLER_12_167
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_179
timestamp 1586364061
transform 1 0 17572 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_183
timestamp 1586364061
transform 1 0 17940 0 -1 9248
box -38 -48 130 592
use scs8hd_or2_4  _385_
timestamp 1586364061
transform 1 0 19412 0 -1 9248
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__388__A
timestamp 1586364061
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__199__B
timestamp 1586364061
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_191
timestamp 1586364061
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_195
timestamp 1586364061
transform 1 0 19044 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
timestamp 1586364061
transform 1 0 21896 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_218
timestamp 1586364061
transform 1 0 21160 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_222
timestamp 1586364061
transform 1 0 21528 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_237
timestamp 1586364061
transform 1 0 22908 0 -1 9248
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_12_249
timestamp 1586364061
transform 1 0 24012 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_259
timestamp 1586364061
transform 1 0 24932 0 -1 9248
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
timestamp 1586364061
transform 1 0 26772 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__399__B
timestamp 1586364061
transform 1 0 26128 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27968 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_271
timestamp 1586364061
transform 1 0 26036 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_274
timestamp 1586364061
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_290
timestamp 1586364061
transform 1 0 27784 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_294
timestamp 1586364061
transform 1 0 28152 0 -1 9248
box -38 -48 406 592
use scs8hd_nor2_4  _396_
timestamp 1586364061
transform 1 0 28612 0 -1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _415_
timestamp 1586364061
transform 1 0 30176 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29624 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_298
timestamp 1586364061
transform 1 0 28520 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_308
timestamp 1586364061
transform 1 0 29440 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_312
timestamp 1586364061
transform 1 0 29808 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_325
timestamp 1586364061
transform 1 0 31004 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_333
timestamp 1586364061
transform 1 0 31740 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_346
timestamp 1586364061
transform 1 0 32936 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33948 0 -1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35512 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33764 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34960 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_354
timestamp 1586364061
transform 1 0 33672 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_366
timestamp 1586364061
transform 1 0 34776 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_370
timestamp 1586364061
transform 1 0 35144 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36524 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_383
timestamp 1586364061
transform 1 0 36340 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_387
timestamp 1586364061
transform 1 0 36708 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_395
timestamp 1586364061
transform 1 0 37444 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_407
timestamp 1586364061
transform 1 0 38548 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_419
timestamp 1586364061
transform 1 0 39652 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_431
timestamp 1586364061
transform 1 0 40756 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_443
timestamp 1586364061
transform 1 0 41860 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_12_455
timestamp 1586364061
transform 1 0 42964 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 43240 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_459
timestamp 1586364061
transform 1 0 43332 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_471
timestamp 1586364061
transform 1 0 44436 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_483
timestamp 1586364061
transform 1 0 45540 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_495
timestamp 1586364061
transform 1 0 46644 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_507
timestamp 1586364061
transform 1 0 47748 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 48852 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_515
timestamp 1586364061
transform 1 0 48484 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_286
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_80
timestamp 1586364061
transform 1 0 8464 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_13_84
timestamp 1586364061
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__190__B
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use scs8hd_or2_4  _190_
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 682 592
use scs8hd_decap_3  FILLER_14_99
timestamp 1586364061
transform 1 0 10212 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_99
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__370__A
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_287
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 866 592
use scs8hd_or2_4  _188_
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 682 592
use scs8hd_decap_4  FILLER_14_113
timestamp 1586364061
transform 1 0 11500 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_109
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_116
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_112
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use scs8hd_or2_4  _187_
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 682 592
use scs8hd_fill_2  FILLER_14_124
timestamp 1586364061
transform 1 0 12512 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_13_119
timestamp 1586364061
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__187__B
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__C
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_128
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_129
timestamp 1586364061
transform 1 0 12972 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__B
timestamp 1586364061
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__C
timestamp 1586364061
transform 1 0 13156 0 1 9248
box -38 -48 222 592
use scs8hd_or3_4  _184_
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 866 592
use scs8hd_or4_4  _172_
timestamp 1586364061
transform 1 0 13340 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_142
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_150
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_146
timestamp 1586364061
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_288
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_160
timestamp 1586364061
transform 1 0 15824 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_154
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 15640 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__D
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use scs8hd_or4_4  _175_
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_167
timestamp 1586364061
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__C
timestamp 1586364061
transform 1 0 16008 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use scs8hd_inv_8  _122_
timestamp 1586364061
transform 1 0 16192 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_173
timestamp 1586364061
transform 1 0 17020 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__203__B
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__C
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_181
timestamp 1586364061
transform 1 0 17756 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_or2_4  _203_
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 682 592
use scs8hd_or2_4  _199_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 682 592
use scs8hd_decap_6  FILLER_14_191
timestamp 1586364061
transform 1 0 18676 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_4  FILLER_13_195
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_191
timestamp 1586364061
transform 1 0 18676 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__363__B
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_206
timestamp 1586364061
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_201
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _388_
timestamp 1586364061
transform 1 0 19780 0 1 9248
box -38 -48 866 592
use scs8hd_or2_4  _209_
timestamp 1586364061
transform 1 0 19412 0 -1 10336
box -38 -48 682 592
use scs8hd_decap_4  FILLER_14_210
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_212
timestamp 1586364061
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__388__B
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__209__B
timestamp 1586364061
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_289
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_220
timestamp 1586364061
transform 1 0 21344 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_216
timestamp 1586364061
transform 1 0 20976 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__387__A
timestamp 1586364061
transform 1 0 21528 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
timestamp 1586364061
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21068 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_235
timestamp 1586364061
transform 1 0 22724 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_231
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22908 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
timestamp 1586364061
transform 1 0 22540 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
timestamp 1586364061
transform 1 0 22080 0 -1 10336
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 590 592
use scs8hd_decap_3  FILLER_13_239
timestamp 1586364061
transform 1 0 23092 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_247
timestamp 1586364061
transform 1 0 23828 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23644 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24104 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__394__B
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_261
timestamp 1586364061
transform 1 0 25116 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_259
timestamp 1586364061
transform 1 0 24932 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__394__A
timestamp 1586364061
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _394_
timestamp 1586364061
transform 1 0 24288 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_265
timestamp 1586364061
transform 1 0 25484 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_6  FILLER_13_263
timestamp 1586364061
transform 1 0 25300 0 1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__395__B
timestamp 1586364061
transform 1 0 26680 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__399__A
timestamp 1586364061
transform 1 0 25944 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_290
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_nor2_4  _399_
timestamp 1586364061
transform 1 0 26128 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_280
timestamp 1586364061
transform 1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_285
timestamp 1586364061
transform 1 0 27324 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_281
timestamp 1586364061
transform 1 0 26956 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27508 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27140 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27140 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_292
timestamp 1586364061
transform 1 0 27968 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_4  FILLER_13_292
timestamp 1586364061
transform 1 0 27968 0 1 9248
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27692 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_306
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_302
timestamp 1586364061
transform 1 0 28888 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_298
timestamp 1586364061
transform 1 0 28520 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__393__B
timestamp 1586364061
transform 1 0 28336 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__393__A
timestamp 1586364061
transform 1 0 28704 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_nor2_4  _393_
timestamp 1586364061
transform 1 0 28704 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_309
timestamp 1586364061
transform 1 0 29532 0 -1 10336
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 29440 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
timestamp 1586364061
transform 1 0 30268 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
timestamp 1586364061
transform 1 0 29624 0 1 9248
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_13_321
timestamp 1586364061
transform 1 0 30636 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_328
timestamp 1586364061
transform 1 0 31280 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_329
timestamp 1586364061
transform 1 0 31372 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_325
timestamp 1586364061
transform 1 0 31004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31188 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
timestamp 1586364061
transform 1 0 30820 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_334
timestamp 1586364061
transform 1 0 31832 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31648 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32016 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_291
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32384 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32200 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_347
timestamp 1586364061
transform 1 0 33028 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_349
timestamp 1586364061
transform 1 0 33212 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_358
timestamp 1586364061
transform 1 0 34040 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_351
timestamp 1586364061
transform 1 0 33396 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33948 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33580 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33212 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33764 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_368
timestamp 1586364061
transform 1 0 34960 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_362
timestamp 1586364061
transform 1 0 34408 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34132 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_372
timestamp 1586364061
transform 1 0 35328 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35512 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35144 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_376
timestamp 1586364061
transform 1 0 35696 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_382
timestamp 1586364061
transform 1 0 36248 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_376
timestamp 1586364061
transform 1 0 35696 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36432 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36064 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36064 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_389
timestamp 1586364061
transform 1 0 36892 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_13_390
timestamp 1586364061
transform 1 0 36984 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_386
timestamp 1586364061
transform 1 0 36616 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 37076 0 1 9248
box -38 -48 222 592
use scs8hd_inv_8  _143_
timestamp 1586364061
transform 1 0 37260 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_402
timestamp 1586364061
transform 1 0 38088 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_292
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_8  _144_
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_12  FILLER_14_407
timestamp 1586364061
transform 1 0 38548 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_13_413
timestamp 1586364061
transform 1 0 39100 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_406
timestamp 1586364061
transform 1 0 38456 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 38272 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 39284 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 38824 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_419
timestamp 1586364061
transform 1 0 39652 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_428
timestamp 1586364061
transform 1 0 40480 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_13_425
timestamp 1586364061
transform 1 0 40204 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_417
timestamp 1586364061
transform 1 0 39468 0 1 9248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 40388 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_440
timestamp 1586364061
transform 1 0 41584 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_452
timestamp 1586364061
transform 1 0 42688 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_431
timestamp 1586364061
transform 1 0 40756 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_443
timestamp 1586364061
transform 1 0 41860 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_14_455
timestamp 1586364061
transform 1 0 42964 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_293
timestamp 1586364061
transform 1 0 43240 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_464
timestamp 1586364061
transform 1 0 43792 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_476
timestamp 1586364061
transform 1 0 44896 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_459
timestamp 1586364061
transform 1 0 43332 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_471
timestamp 1586364061
transform 1 0 44436 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_483
timestamp 1586364061
transform 1 0 45540 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 46000 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_489
timestamp 1586364061
transform 1 0 46092 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_501
timestamp 1586364061
transform 1 0 47196 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_495
timestamp 1586364061
transform 1 0 46644 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_507
timestamp 1586364061
transform 1 0 47748 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 48852 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 48852 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_513
timestamp 1586364061
transform 1 0 48300 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_515
timestamp 1586364061
transform 1 0 48484 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_294
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 774 592
use scs8hd_or2_4  _169_
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 682 592
use scs8hd_or2_4  _191_
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__191__B
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_82
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_94
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_113
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_109
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__B
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_295
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_or2_4  _185_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 682 592
use scs8hd_fill_2  FILLER_15_130
timestamp 1586364061
transform 1 0 13064 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_134
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_139
timestamp 1586364061
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__B
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 13708 0 1 10336
box -38 -48 222 592
use scs8hd_or2_4  _179_
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 682 592
use scs8hd_fill_2  FILLER_15_154
timestamp 1586364061
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_150
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__B
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_158
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_or3_4  _181_
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__378__B
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__378__A
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__376__B
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__376__A
timestamp 1586364061
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_296
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_188
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__B
timestamp 1586364061
transform 1 0 18584 0 1 10336
box -38 -48 222 592
use scs8hd_or2_4  _201_
timestamp 1586364061
transform 1 0 18768 0 1 10336
box -38 -48 682 592
use scs8hd_decap_4  FILLER_15_207
timestamp 1586364061
transform 1 0 20148 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_203
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_199
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__363__A
timestamp 1586364061
transform 1 0 19964 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_211
timestamp 1586364061
transform 1 0 20516 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _387_
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__387__B
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_223
timestamp 1586364061
transform 1 0 21620 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_227
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_231
timestamp 1586364061
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
timestamp 1586364061
transform 1 0 24840 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_297
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 24656 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__416__A
timestamp 1586364061
transform 1 0 24288 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__B
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_248
timestamp 1586364061
transform 1 0 23920 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_254
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
timestamp 1586364061
transform 1 0 26588 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 26404 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__395__A
timestamp 1586364061
transform 1 0 26036 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28060 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_273
timestamp 1586364061
transform 1 0 26220 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_288
timestamp 1586364061
transform 1 0 27600 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_292
timestamp 1586364061
transform 1 0 27968 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_295
timestamp 1586364061
transform 1 0 28244 0 1 10336
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
timestamp 1586364061
transform 1 0 30544 0 1 10336
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_298
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
timestamp 1586364061
transform 1 0 30360 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__392__A
timestamp 1586364061
transform 1 0 29716 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__392__B
timestamp 1586364061
transform 1 0 28980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_309
timestamp 1586364061
transform 1 0 29532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_313
timestamp 1586364061
transform 1 0 29900 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_317
timestamp 1586364061
transform 1 0 30268 0 1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32384 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32200 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31832 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_331
timestamp 1586364061
transform 1 0 31556 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_336
timestamp 1586364061
transform 1 0 32016 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_299
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 34224 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33396 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_349
timestamp 1586364061
transform 1 0 33212 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_353
timestamp 1586364061
transform 1 0 33580 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_359
timestamp 1586364061
transform 1 0 34132 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_362
timestamp 1586364061
transform 1 0 34408 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_382
timestamp 1586364061
transform 1 0 36248 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_376
timestamp 1586364061
transform 1 0 35696 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__294__A
timestamp 1586364061
transform 1 0 36064 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_386
timestamp 1586364061
transform 1 0 36616 0 1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__294__B
timestamp 1586364061
transform 1 0 36432 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_392
timestamp 1586364061
transform 1 0 37168 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37260 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37444 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_402
timestamp 1586364061
transform 1 0 38088 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_398
timestamp 1586364061
transform 1 0 37720 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37904 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_300
timestamp 1586364061
transform 1 0 40388 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__291__A
timestamp 1586364061
transform 1 0 39284 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__291__B
timestamp 1586364061
transform 1 0 39652 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38272 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_406
timestamp 1586364061
transform 1 0 38456 0 1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_15_414
timestamp 1586364061
transform 1 0 39192 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_417
timestamp 1586364061
transform 1 0 39468 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_421
timestamp 1586364061
transform 1 0 39836 0 1 10336
box -38 -48 590 592
use scs8hd_decap_12  FILLER_15_428
timestamp 1586364061
transform 1 0 40480 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_440
timestamp 1586364061
transform 1 0 41584 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_452
timestamp 1586364061
transform 1 0 42688 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_464
timestamp 1586364061
transform 1 0 43792 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_476
timestamp 1586364061
transform 1 0 44896 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_301
timestamp 1586364061
transform 1 0 46000 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_489
timestamp 1586364061
transform 1 0 46092 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_501
timestamp 1586364061
transform 1 0 47196 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 48852 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_513
timestamp 1586364061
transform 1 0 48300 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_302
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_nor2_4  _370_
timestamp 1586364061
transform 1 0 10028 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_303
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__370__B
timestamp 1586364061
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_106
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 222 592
use scs8hd_or2_4  _182_
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__185__B
timestamp 1586364061
transform 1 0 13156 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11040 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_110
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_133
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 406 592
use scs8hd_or2_4  _178_
timestamp 1586364061
transform 1 0 13708 0 -1 11424
box -38 -48 682 592
use scs8hd_nor2_4  _378_
timestamp 1586364061
transform 1 0 15916 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_304
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_144
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_152
timestamp 1586364061
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_160
timestamp 1586364061
transform 1 0 15824 0 -1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _376_
timestamp 1586364061
transform 1 0 17848 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_170
timestamp 1586364061
transform 1 0 16744 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 222 592
use scs8hd_or2_4  _363_
timestamp 1586364061
transform 1 0 19412 0 -1 11424
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_305
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__208__B
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__379__B
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_191
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_195
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_4  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_212
timestamp 1586364061
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use scs8hd_or2_4  _167_
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 682 592
use scs8hd_nor2_4  _204_
timestamp 1586364061
transform 1 0 22816 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__206__B
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22540 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_222
timestamp 1586364061
transform 1 0 21528 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_226
timestamp 1586364061
transform 1 0 21896 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_229
timestamp 1586364061
transform 1 0 22172 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_235
timestamp 1586364061
transform 1 0 22724 0 -1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _416_
timestamp 1586364061
transform 1 0 24380 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__189__B
timestamp 1586364061
transform 1 0 25760 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__416__B
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23828 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_245
timestamp 1586364061
transform 1 0 23644 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_249
timestamp 1586364061
transform 1 0 24012 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_262
timestamp 1586364061
transform 1 0 25208 0 -1 11424
box -38 -48 590 592
use scs8hd_nor2_4  _395_
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28060 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_306
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__186__B
timestamp 1586364061
transform 1 0 27508 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27876 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_270
timestamp 1586364061
transform 1 0 25944 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_285
timestamp 1586364061
transform 1 0 27324 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_289
timestamp 1586364061
transform 1 0 27692 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _392_
timestamp 1586364061
transform 1 0 29532 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29256 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30544 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_296
timestamp 1586364061
transform 1 0 28336 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_304
timestamp 1586364061
transform 1 0 29072 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_308
timestamp 1586364061
transform 1 0 29440 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_318
timestamp 1586364061
transform 1 0 30360 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_322
timestamp 1586364061
transform 1 0 30728 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_307
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32568 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30912 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_326
timestamp 1586364061
transform 1 0 31096 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_334
timestamp 1586364061
transform 1 0 31832 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_340
timestamp 1586364061
transform 1 0 32384 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_344
timestamp 1586364061
transform 1 0 32752 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_8  _142_
timestamp 1586364061
transform 1 0 34500 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35512 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_356
timestamp 1586364061
transform 1 0 33856 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_362
timestamp 1586364061
transform 1 0 34408 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_372
timestamp 1586364061
transform 1 0 35328 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _294_
timestamp 1586364061
transform 1 0 36064 0 -1 11424
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_308
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_376
timestamp 1586364061
transform 1 0 35696 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_389
timestamp 1586364061
transform 1 0 36892 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _291_
timestamp 1586364061
transform 1 0 39284 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_8  FILLER_16_407
timestamp 1586364061
transform 1 0 38548 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_16_424
timestamp 1586364061
transform 1 0 40112 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_436
timestamp 1586364061
transform 1 0 41216 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_448
timestamp 1586364061
transform 1 0 42320 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_456
timestamp 1586364061
transform 1 0 43056 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_309
timestamp 1586364061
transform 1 0 43240 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_459
timestamp 1586364061
transform 1 0 43332 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_471
timestamp 1586364061
transform 1 0 44436 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_483
timestamp 1586364061
transform 1 0 45540 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_495
timestamp 1586364061
transform 1 0 46644 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_507
timestamp 1586364061
transform 1 0 47748 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 48852 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_515
timestamp 1586364061
transform 1 0 48484 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_310
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_92
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_96
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _369_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_311
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__369__A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__369__B
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_111
timestamp 1586364061
transform 1 0 11316 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_115
timestamp 1586364061
transform 1 0 11684 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
timestamp 1586364061
transform 1 0 14904 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_161
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_165
timestamp 1586364061
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_172
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_180
timestamp 1586364061
transform 1 0 17664 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_176
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 406 592
use scs8hd_decap_4  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_312
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _208_
timestamp 1586364061
transform 1 0 20424 0 1 11424
box -38 -48 866 592
use scs8hd_nor2_4  _379_
timestamp 1586364061
transform 1 0 18584 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__379__A
timestamp 1586364061
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_199
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  FILLER_17_205
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _206_
timestamp 1586364061
transform 1 0 21988 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 21804 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_219
timestamp 1586364061
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_223
timestamp 1586364061
transform 1 0 21620 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_236
timestamp 1586364061
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_313
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_17_264
timestamp 1586364061
transform 1 0 25392 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_260
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_256
timestamp 1586364061
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__B
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _189_
timestamp 1586364061
transform 1 0 25760 0 1 11424
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27324 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27140 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 26772 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_277
timestamp 1586364061
transform 1 0 26588 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_281
timestamp 1586364061
transform 1 0 26956 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_294
timestamp 1586364061
transform 1 0 28152 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _391_
timestamp 1586364061
transform 1 0 29808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_314
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__390__A
timestamp 1586364061
transform 1 0 28704 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__391__A
timestamp 1586364061
transform 1 0 29624 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__390__B
timestamp 1586364061
transform 1 0 28336 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_298
timestamp 1586364061
transform 1 0 28520 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_302
timestamp 1586364061
transform 1 0 28888 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_306
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_321
timestamp 1586364061
transform 1 0 30636 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31556 0 1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32568 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
timestamp 1586364061
transform 1 0 30820 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32384 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 32016 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31372 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_325
timestamp 1586364061
transform 1 0 31004 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_334
timestamp 1586364061
transform 1 0 31832 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_338
timestamp 1586364061
transform 1 0 32200 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _141_
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_315
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33856 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 34592 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34224 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_351
timestamp 1586364061
transform 1 0 33396 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_355
timestamp 1586364061
transform 1 0 33764 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_358
timestamp 1586364061
transform 1 0 34040 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_362
timestamp 1586364061
transform 1 0 34408 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 36708 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 36524 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 36156 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_376
timestamp 1586364061
transform 1 0 35696 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_380
timestamp 1586364061
transform 1 0 36064 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_383
timestamp 1586364061
transform 1 0 36340 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_398
timestamp 1586364061
transform 1 0 37720 0 1 11424
box -38 -48 590 592
use scs8hd_nor2_4  _292_
timestamp 1586364061
transform 1 0 38456 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_316
timestamp 1586364061
transform 1 0 40388 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 39468 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__292__A
timestamp 1586364061
transform 1 0 38272 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39836 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_415
timestamp 1586364061
transform 1 0 39284 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_419
timestamp 1586364061
transform 1 0 39652 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_423
timestamp 1586364061
transform 1 0 40020 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  FILLER_17_428
timestamp 1586364061
transform 1 0 40480 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 40756 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 41124 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_433
timestamp 1586364061
transform 1 0 40940 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_437
timestamp 1586364061
transform 1 0 41308 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_449
timestamp 1586364061
transform 1 0 42412 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_461
timestamp 1586364061
transform 1 0 43516 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_473
timestamp 1586364061
transform 1 0 44620 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_317
timestamp 1586364061
transform 1 0 46000 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_485
timestamp 1586364061
transform 1 0 45724 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_489
timestamp 1586364061
transform 1 0 46092 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_501
timestamp 1586364061
transform 1 0 47196 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 48852 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_513
timestamp 1586364061
transform 1 0 48300 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_318
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
timestamp 1586364061
transform 1 0 10212 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_319
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__365__B
timestamp 1586364061
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_97
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_18_110
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_18_122
timestamp 1586364061
transform 1 0 12328 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_139
timestamp 1586364061
transform 1 0 13892 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_135
timestamp 1586364061
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13708 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_147
timestamp 1586364061
transform 1 0 14628 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__377__B
timestamp 1586364061
transform 1 0 14904 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_158
timestamp 1586364061
transform 1 0 15640 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_152
timestamp 1586364061
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_320
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16008 0 -1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch
timestamp 1586364061
transform 1 0 17756 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_18_173
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_321
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__196__B
timestamp 1586364061
transform 1 0 18952 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_192
timestamp 1586364061
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_196
timestamp 1586364061
transform 1 0 19136 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21252 0 -1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_2_.latch
timestamp 1586364061
transform 1 0 23000 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__210__B
timestamp 1586364061
transform 1 0 21068 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_230
timestamp 1586364061
transform 1 0 22264 0 -1 12512
box -38 -48 774 592
use scs8hd_nor2_4  _192_
timestamp 1586364061
transform 1 0 24840 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_249
timestamp 1586364061
transform 1 0 24012 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_253
timestamp 1586364061
transform 1 0 24380 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_257
timestamp 1586364061
transform 1 0 24748 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_267
timestamp 1586364061
transform 1 0 25668 0 -1 12512
box -38 -48 774 592
use scs8hd_nor2_4  _186_
timestamp 1586364061
transform 1 0 27140 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_322
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28244 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26680 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_280
timestamp 1586364061
transform 1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_292
timestamp 1586364061
transform 1 0 27968 0 -1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _390_
timestamp 1586364061
transform 1 0 28704 0 -1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
timestamp 1586364061
transform 1 0 30268 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__391__B
timestamp 1586364061
transform 1 0 29808 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_297
timestamp 1586364061
transform 1 0 28428 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_309
timestamp 1586364061
transform 1 0 29532 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_314
timestamp 1586364061
transform 1 0 29992 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_8  _139_
timestamp 1586364061
transform 1 0 32292 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_323
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_328
timestamp 1586364061
transform 1 0 31280 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_337
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_348
timestamp 1586364061
transform 1 0 33120 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35420 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33856 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__293__A
timestamp 1586364061
transform 1 0 35052 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_365
timestamp 1586364061
transform 1 0 34684 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_371
timestamp 1586364061
transform 1 0 35236 0 -1 12512
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 36432 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_324
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36892 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37904 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_376
timestamp 1586364061
transform 1 0 35696 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_387
timestamp 1586364061
transform 1 0 36708 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_391
timestamp 1586364061
transform 1 0 37076 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_402
timestamp 1586364061
transform 1 0 38088 0 -1 12512
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_6_.latch
timestamp 1586364061
transform 1 0 39008 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__292__B
timestamp 1586364061
transform 1 0 38456 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38824 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_408
timestamp 1586364061
transform 1 0 38640 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_423
timestamp 1586364061
transform 1 0 40020 0 -1 12512
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_7_.latch
timestamp 1586364061
transform 1 0 40756 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_18_442
timestamp 1586364061
transform 1 0 41768 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_454
timestamp 1586364061
transform 1 0 42872 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_325
timestamp 1586364061
transform 1 0 43240 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_459
timestamp 1586364061
transform 1 0 43332 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_471
timestamp 1586364061
transform 1 0 44436 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_483
timestamp 1586364061
transform 1 0 45540 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_495
timestamp 1586364061
transform 1 0 46644 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_507
timestamp 1586364061
transform 1 0 47748 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 48852 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_515
timestamp 1586364061
transform 1 0 48484 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_334
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8096 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_326
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_79
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_19_90
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_83
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_96
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__365__A
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_335
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _371_
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _365_
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_107
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_103
timestamp 1586364061
transform 1 0 10580 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_107
timestamp 1586364061
transform 1 0 10948 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__371__A
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_111
timestamp 1586364061
transform 1 0 11316 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_118
timestamp 1586364061
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_114
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_111
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__371__B
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_327
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__368__A
timestamp 1586364061
transform 1 0 12604 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
timestamp 1586364061
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_127
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _368_
timestamp 1586364061
transform 1 0 13156 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
timestamp 1586364061
transform 1 0 13156 0 -1 13600
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_20_121
timestamp 1586364061
transform 1 0 12236 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_6  FILLER_20_142
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_4  FILLER_19_144
timestamp 1586364061
transform 1 0 14352 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_140
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__368__B
timestamp 1586364061
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_150
timestamp 1586364061
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14720 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__377__A
timestamp 1586364061
transform 1 0 14720 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_336
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _377_
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 866 592
use scs8hd_decap_6  FILLER_20_161
timestamp 1586364061
transform 1 0 15916 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_157
timestamp 1586364061
transform 1 0 15548 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_167
timestamp 1586364061
transform 1 0 16468 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_164
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__B
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16744 0 -1 13600
box -38 -48 866 592
use scs8hd_or2_4  _193_
timestamp 1586364061
transform 1 0 16560 0 1 12512
box -38 -48 682 592
use scs8hd_fill_2  FILLER_20_179
timestamp 1586364061
transform 1 0 17572 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_183
timestamp 1586364061
transform 1 0 17940 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18216 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_328
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_192
timestamp 1586364061
transform 1 0 18768 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_189
timestamp 1586364061
transform 1 0 18492 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_199
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__373__A
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18400 0 1 12512
box -38 -48 1050 592
use scs8hd_or2_4  _196_
timestamp 1586364061
transform 1 0 18860 0 -1 13600
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19964 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_203
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__210__A
timestamp 1586364061
transform 1 0 20332 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 20332 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_207
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_211
timestamp 1586364061
transform 1 0 20516 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_208
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_200
timestamp 1586364061
transform 1 0 19504 0 -1 13600
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20700 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_337
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_8  FILLER_19_226
timestamp 1586364061
transform 1 0 21896 0 1 12512
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 1050 592
use scs8hd_nor2_4  _210_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22632 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_240
timestamp 1586364061
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_329
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_243
timestamp 1586364061
transform 1 0 23460 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_247
timestamp 1586364061
transform 1 0 23828 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24196 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_248
timestamp 1586364061
transform 1 0 23920 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_253
timestamp 1586364061
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_250
timestamp 1586364061
transform 1 0 24104 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_1  FILLER_20_264
timestamp 1586364061
transform 1 0 25392 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_260
timestamp 1586364061
transform 1 0 25024 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_262
timestamp 1586364061
transform 1 0 25208 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25024 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch_D
timestamp 1586364061
transform 1 0 25392 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_267
timestamp 1586364061
transform 1 0 25668 0 -1 13600
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_8_.latch
timestamp 1586364061
transform 1 0 25576 0 1 12512
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_19_277
timestamp 1586364061
transform 1 0 26588 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch_D
timestamp 1586364061
transform 1 0 26772 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_338
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_9_.latch
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_20_291
timestamp 1586364061
transform 1 0 27876 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_287
timestamp 1586364061
transform 1 0 27508 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_285
timestamp 1586364061
transform 1 0 27324 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_281
timestamp 1586364061
transform 1 0 26956 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__183__B
timestamp 1586364061
transform 1 0 27692 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 27416 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _183_
timestamp 1586364061
transform 1 0 27600 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28060 0 -1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch
timestamp 1586364061
transform 1 0 28244 0 -1 13600
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_20_306
timestamp 1586364061
transform 1 0 29256 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_301
timestamp 1586364061
transform 1 0 28796 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_297
timestamp 1586364061
transform 1 0 28428 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_10_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_330
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_20_317
timestamp 1586364061
transform 1 0 30268 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_4  FILLER_20_310
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_317
timestamp 1586364061
transform 1 0 30268 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29440 0 -1 13600
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29992 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_321
timestamp 1586364061
transform 1 0 30636 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30452 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_327
timestamp 1586364061
transform 1 0 31188 0 -1 13600
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31004 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch_D
timestamp 1586364061
transform 1 0 30820 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_11_.latch
timestamp 1586364061
transform 1 0 31004 0 1 12512
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_20_340
timestamp 1586364061
transform 1 0 32384 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_335
timestamp 1586364061
transform 1 0 31924 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_340
timestamp 1586364061
transform 1 0 32384 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_336
timestamp 1586364061
transform 1 0 32016 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 32568 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32200 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_339
timestamp 1586364061
transform 1 0 32016 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32108 0 -1 13600
box -38 -48 314 592
use scs8hd_inv_8  _140_
timestamp 1586364061
transform 1 0 32752 0 1 12512
box -38 -48 866 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 33120 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_351
timestamp 1586364061
transform 1 0 33396 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_19_357
timestamp 1586364061
transform 1 0 33948 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_353
timestamp 1586364061
transform 1 0 33580 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 33764 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34776 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_331
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34592 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_363
timestamp 1586364061
transform 1 0 34500 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_367
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_363
timestamp 1586364061
transform 1 0 34500 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__293__B
timestamp 1586364061
transform 1 0 35236 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_369
timestamp 1586364061
transform 1 0 35052 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_373
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _293_
timestamp 1586364061
transform 1 0 35052 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35604 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_382
timestamp 1586364061
transform 1 0 36248 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_378
timestamp 1586364061
transform 1 0 35880 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36432 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 36064 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36616 0 1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 35788 0 -1 13600
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_20_396
timestamp 1586364061
transform 1 0 37536 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_388
timestamp 1586364061
transform 1 0 36800 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_4  FILLER_19_393
timestamp 1586364061
transform 1 0 37260 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_389
timestamp 1586364061
transform 1 0 36892 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37628 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37076 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_340
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37720 0 -1 13600
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37812 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_402
timestamp 1586364061
transform 1 0 38088 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_411
timestamp 1586364061
transform 1 0 38916 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_407
timestamp 1586364061
transform 1 0 38548 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_406
timestamp 1586364061
transform 1 0 38456 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38640 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38732 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38272 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38824 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 39284 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_12  FILLER_20_424
timestamp 1586364061
transform 1 0 40112 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_428
timestamp 1586364061
transform 1 0 40480 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_19_423
timestamp 1586364061
transform 1 0 40020 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_419
timestamp 1586364061
transform 1 0 39652 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40204 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39836 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_332
timestamp 1586364061
transform 1 0 40388 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_440
timestamp 1586364061
transform 1 0 41584 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_452
timestamp 1586364061
transform 1 0 42688 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_436
timestamp 1586364061
transform 1 0 41216 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_448
timestamp 1586364061
transform 1 0 42320 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_456
timestamp 1586364061
transform 1 0 43056 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_341
timestamp 1586364061
transform 1 0 43240 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_464
timestamp 1586364061
transform 1 0 43792 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_476
timestamp 1586364061
transform 1 0 44896 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_459
timestamp 1586364061
transform 1 0 43332 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_471
timestamp 1586364061
transform 1 0 44436 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_483
timestamp 1586364061
transform 1 0 45540 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_333
timestamp 1586364061
transform 1 0 46000 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_489
timestamp 1586364061
transform 1 0 46092 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_501
timestamp 1586364061
transform 1 0 47196 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_495
timestamp 1586364061
transform 1 0 46644 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_507
timestamp 1586364061
transform 1 0 47748 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 48852 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 48852 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_513
timestamp 1586364061
transform 1 0 48300 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_515
timestamp 1586364061
transform 1 0 48484 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_342
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use scs8hd_nor2_4  _364_
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
timestamp 1586364061
transform 1 0 10764 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__364__A
timestamp 1586364061
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__364__B
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_90
timestamp 1586364061
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_103
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_107
timestamp 1586364061
transform 1 0 10948 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_127
timestamp 1586364061
transform 1 0 12788 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_343
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14720 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_140
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_144
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_157
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_161
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_344
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__372__A
timestamp 1586364061
transform 1 0 18308 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__373__B
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__372__B
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_174
timestamp 1586364061
transform 1 0 17112 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _170_
timestamp 1586364061
transform 1 0 20332 0 1 13600
box -38 -48 866 592
use scs8hd_nor2_4  _373_
timestamp 1586364061
transform 1 0 18584 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 20148 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_189
timestamp 1586364061
transform 1 0 18492 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_199
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_218
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_222
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 21712 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_226
timestamp 1586364061
transform 1 0 21896 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_230
timestamp 1586364061
transform 1 0 22264 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22356 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_345
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23920 0 1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_21_261
timestamp 1586364061
transform 1 0 25116 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 24932 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_268
timestamp 1586364061
transform 1 0 25760 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__B
timestamp 1586364061
transform 1 0 25300 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25484 0 1 13600
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28060 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26312 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25944 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27876 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27508 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_272
timestamp 1586364061
transform 1 0 26128 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_285
timestamp 1586364061
transform 1 0 27324 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_289
timestamp 1586364061
transform 1 0 27692 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_346
timestamp 1586364061
transform 1 0 29164 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28520 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__319__A
timestamp 1586364061
transform 1 0 30452 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_296
timestamp 1586364061
transform 1 0 28336 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_300
timestamp 1586364061
transform 1 0 28704 0 1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_21_315
timestamp 1586364061
transform 1 0 30084 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_321
timestamp 1586364061
transform 1 0 30636 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_325
timestamp 1586364061
transform 1 0 31004 0 1 13600
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__319__B
timestamp 1586364061
transform 1 0 30820 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_331
timestamp 1586364061
transform 1 0 31556 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31648 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31832 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_341
timestamp 1586364061
transform 1 0 32476 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_337
timestamp 1586364061
transform 1 0 32108 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 32292 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_345
timestamp 1586364061
transform 1 0 32844 0 1 13600
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_2.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32660 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_357
timestamp 1586364061
transform 1 0 33948 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_351
timestamp 1586364061
transform 1 0 33396 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33488 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34132 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33672 0 1 13600
box -38 -48 314 592
use scs8hd_decap_6  FILLER_21_367
timestamp 1586364061
transform 1 0 34868 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_365
timestamp 1586364061
transform 1 0 34684 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_361
timestamp 1586364061
transform 1 0 34316 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34500 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_347
timestamp 1586364061
transform 1 0 34776 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 35420 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 35604 0 1 13600
box -38 -48 1050 592
use scs8hd_conb_1  _439_
timestamp 1586364061
transform 1 0 37352 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37812 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36800 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37168 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_386
timestamp 1586364061
transform 1 0 36616 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_390
timestamp 1586364061
transform 1 0 36984 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_397
timestamp 1586364061
transform 1 0 37628 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_401
timestamp 1586364061
transform 1 0 37996 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38364 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_348
timestamp 1586364061
transform 1 0 40388 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38180 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40204 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39376 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_414
timestamp 1586364061
transform 1 0 39192 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_418
timestamp 1586364061
transform 1 0 39560 0 1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_21_424
timestamp 1586364061
transform 1 0 40112 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 41124 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 41492 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_431
timestamp 1586364061
transform 1 0 40756 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_437
timestamp 1586364061
transform 1 0 41308 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_441
timestamp 1586364061
transform 1 0 41676 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_453
timestamp 1586364061
transform 1 0 42780 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_465
timestamp 1586364061
transform 1 0 43884 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_477
timestamp 1586364061
transform 1 0 44988 0 1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_349
timestamp 1586364061
transform 1 0 46000 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_485
timestamp 1586364061
transform 1 0 45724 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_489
timestamp 1586364061
transform 1 0 46092 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_501
timestamp 1586364061
transform 1 0 47196 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 48852 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_513
timestamp 1586364061
transform 1 0 48300 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_350
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_351
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11776 0 -1 14688
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13156 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_108
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_6  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_352
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_142
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_146
timestamp 1586364061
transform 1 0 14536 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _372_
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17296 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18124 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_170
timestamp 1586364061
transform 1 0 16744 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_6  FILLER_22_179
timestamp 1586364061
transform 1 0 17572 0 -1 14688
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_353
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_196
timestamp 1586364061
transform 1 0 19136 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_22_208
timestamp 1586364061
transform 1 0 20240 0 -1 14688
box -38 -48 590 592
use scs8hd_nor2_4  _173_
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_4  FILLER_22_241
timestamp 1586364061
transform 1 0 23276 0 -1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _197_
timestamp 1586364061
transform 1 0 24840 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__194__B
timestamp 1586364061
transform 1 0 23644 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24104 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_247
timestamp 1586364061
transform 1 0 23828 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_22_252
timestamp 1586364061
transform 1 0 24288 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_8  FILLER_22_267
timestamp 1586364061
transform 1 0 25668 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_4_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28244 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_354
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_285
timestamp 1586364061
transform 1 0 27324 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_293
timestamp 1586364061
transform 1 0 28060 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _319_
timestamp 1586364061
transform 1 0 30452 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__320__B
timestamp 1586364061
transform 1 0 30268 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_5_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29256 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_304
timestamp 1586364061
transform 1 0 29072 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_308
timestamp 1586364061
transform 1 0 29440 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_316
timestamp 1586364061
transform 1 0 30176 0 -1 14688
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_355
timestamp 1586364061
transform 1 0 32016 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_328
timestamp 1586364061
transform 1 0 31280 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_8  FILLER_22_348
timestamp 1586364061
transform 1 0 33120 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33856 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__296__B
timestamp 1586364061
transform 1 0 34868 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_365
timestamp 1586364061
transform 1 0 34684 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_369
timestamp 1586364061
transform 1 0 35052 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36064 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_356
timestamp 1586364061
transform 1 0 37628 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37076 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_377
timestamp 1586364061
transform 1 0 35788 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_389
timestamp 1586364061
transform 1 0 36892 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_393
timestamp 1586364061
transform 1 0 37260 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_6  FILLER_22_398
timestamp 1586364061
transform 1 0 37720 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38364 0 -1 14688
box -38 -48 866 592
use scs8hd_fill_1  FILLER_22_404
timestamp 1586364061
transform 1 0 38272 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_414
timestamp 1586364061
transform 1 0 39192 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_426
timestamp 1586364061
transform 1 0 40296 0 -1 14688
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_7_.latch
timestamp 1586364061
transform 1 0 41124 0 -1 14688
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_22_434
timestamp 1586364061
transform 1 0 41032 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_446
timestamp 1586364061
transform 1 0 42136 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_357
timestamp 1586364061
transform 1 0 43240 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_459
timestamp 1586364061
transform 1 0 43332 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_471
timestamp 1586364061
transform 1 0 44436 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_483
timestamp 1586364061
transform 1 0 45540 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_495
timestamp 1586364061
transform 1 0 46644 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_507
timestamp 1586364061
transform 1 0 47748 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 48852 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_515
timestamp 1586364061
transform 1 0 48484 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_358
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
timestamp 1586364061
transform 1 0 9936 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_88
timestamp 1586364061
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_92
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_107
timestamp 1586364061
transform 1 0 10948 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_111
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_121
timestamp 1586364061
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_23_115
timestamp 1586364061
transform 1 0 11684 0 1 14688
box -38 -48 590 592
use scs8hd_fill_2  FILLER_23_127
timestamp 1586364061
transform 1 0 12788 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_359
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_131
timestamp 1586364061
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13340 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_136
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_140
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_144
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_156
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_160
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16192 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_167
timestamp 1586364061
transform 1 0 16468 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_360
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 18216 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
timestamp 1586364061
transform 1 0 18400 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_D
timestamp 1586364061
transform 1 0 20792 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_D
timestamp 1586364061
transform 1 0 20424 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20056 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_199
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_203
timestamp 1586364061
transform 1 0 19780 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_212
timestamp 1586364061
transform 1 0 20608 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_14_.latch
timestamp 1586364061
transform 1 0 20976 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22632 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22172 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_227
timestamp 1586364061
transform 1 0 21988 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_231
timestamp 1586364061
transform 1 0 22356 0 1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_23_236
timestamp 1586364061
transform 1 0 22816 0 1 14688
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_361
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _194_
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use scs8hd_fill_2  FILLER_23_262
timestamp 1586364061
transform 1 0 25208 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_258
timestamp 1586364061
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_254
timestamp 1586364061
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 25392 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_6_.latch
timestamp 1586364061
transform 1 0 25576 0 1 14688
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27324 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 28244 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26772 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27784 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27140 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_277
timestamp 1586364061
transform 1 0 26588 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_281
timestamp 1586364061
transform 1 0 26956 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_288
timestamp 1586364061
transform 1 0 27600 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_292
timestamp 1586364061
transform 1 0 27968 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_301
timestamp 1586364061
transform 1 0 28796 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_297
timestamp 1586364061
transform 1 0 28428 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28612 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28980 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_362
timestamp 1586364061
transform 1 0 29164 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_314
timestamp 1586364061
transform 1 0 29992 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_309
timestamp 1586364061
transform 1 0 29532 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__321__B
timestamp 1586364061
transform 1 0 29808 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_318
timestamp 1586364061
transform 1 0 30360 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__320__A
timestamp 1586364061
transform 1 0 30176 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__321__A
timestamp 1586364061
transform 1 0 30544 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _321_
timestamp 1586364061
transform 1 0 30728 0 1 14688
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 32292 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 32108 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 31740 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_331
timestamp 1586364061
transform 1 0 31556 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_335
timestamp 1586364061
transform 1 0 31924 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_358
timestamp 1586364061
transform 1 0 34040 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_354
timestamp 1586364061
transform 1 0 33672 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_350
timestamp 1586364061
transform 1 0 33304 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33856 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33488 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_362
timestamp 1586364061
transform 1 0 34408 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__296__A
timestamp 1586364061
transform 1 0 34592 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_363
timestamp 1586364061
transform 1 0 34776 0 1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _296_
timestamp 1586364061
transform 1 0 34868 0 1 14688
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36708 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__297__A
timestamp 1586364061
transform 1 0 35880 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__297__B
timestamp 1586364061
transform 1 0 36248 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38088 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_376
timestamp 1586364061
transform 1 0 35696 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_380
timestamp 1586364061
transform 1 0 36064 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_384
timestamp 1586364061
transform 1 0 36432 0 1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_23_396
timestamp 1586364061
transform 1 0 37536 0 1 14688
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 38272 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_407
timestamp 1586364061
transform 1 0 38548 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38732 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_411
timestamp 1586364061
transform 1 0 38916 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39100 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39284 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_418
timestamp 1586364061
transform 1 0 39560 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39744 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_422
timestamp 1586364061
transform 1 0 39928 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__300__B
timestamp 1586364061
transform 1 0 40204 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_364
timestamp 1586364061
transform 1 0 40388 0 1 14688
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41768 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40940 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__300__A
timestamp 1586364061
transform 1 0 41308 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42780 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_431
timestamp 1586364061
transform 1 0 40756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_435
timestamp 1586364061
transform 1 0 41124 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_439
timestamp 1586364061
transform 1 0 41492 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_451
timestamp 1586364061
transform 1 0 42596 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_455
timestamp 1586364061
transform 1 0 42964 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43332 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_461
timestamp 1586364061
transform 1 0 43516 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_473
timestamp 1586364061
transform 1 0 44620 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_365
timestamp 1586364061
transform 1 0 46000 0 1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_23_485
timestamp 1586364061
transform 1 0 45724 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_489
timestamp 1586364061
transform 1 0 46092 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_501
timestamp 1586364061
transform 1 0 47196 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 48852 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_23_513
timestamp 1586364061
transform 1 0 48300 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_366
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10948 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_367
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_6  FILLER_24_99
timestamp 1586364061
transform 1 0 10212 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_116
timestamp 1586364061
transform 1 0 11776 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_133
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_368
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_137
timestamp 1586364061
transform 1 0 13708 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_149
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
timestamp 1586364061
transform 1 0 17848 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_168
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_174
timestamp 1586364061
transform 1 0 17112 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_369
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__375__B
timestamp 1586364061
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_193
timestamp 1586364061
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_197
timestamp 1586364061
transform 1 0 19228 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_204
timestamp 1586364061
transform 1 0 19872 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_212
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22632 0 -1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_15_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22264 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_226
timestamp 1586364061
transform 1 0 21896 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_232
timestamp 1586364061
transform 1 0 22448 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_237
timestamp 1586364061
transform 1 0 22908 0 -1 15776
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_7_.latch
timestamp 1586364061
transform 1 0 24104 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25760 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_249
timestamp 1586364061
transform 1 0 24012 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_261
timestamp 1586364061
transform 1 0 25116 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_265
timestamp 1586364061
transform 1 0 25484 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_274
timestamp 1586364061
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_270
timestamp 1586364061
transform 1 0 25944 0 -1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_370
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_2  FILLER_24_290
timestamp 1586364061
transform 1 0 27784 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_285
timestamp 1586364061
transform 1 0 27324 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27968 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__B
timestamp 1586364061
transform 1 0 27600 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_294
timestamp 1586364061
transform 1 0 28152 0 -1 15776
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
timestamp 1586364061
transform 1 0 28244 0 -1 15776
box -38 -48 1050 592
use scs8hd_nor2_4  _320_
timestamp 1586364061
transform 1 0 30452 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__318__B
timestamp 1586364061
transform 1 0 29624 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30084 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_306
timestamp 1586364061
transform 1 0 29256 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  FILLER_24_312
timestamp 1586364061
transform 1 0 29808 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_317
timestamp 1586364061
transform 1 0 30268 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 32384 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_371
timestamp 1586364061
transform 1 0 32016 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31832 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_328
timestamp 1586364061
transform 1 0 31280 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_3  FILLER_24_337
timestamp 1586364061
transform 1 0 32108 0 -1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34132 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33948 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_351
timestamp 1586364061
transform 1 0 33396 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_8  FILLER_24_368
timestamp 1586364061
transform 1 0 34960 0 -1 15776
box -38 -48 774 592
use scs8hd_nor2_4  _297_
timestamp 1586364061
transform 1 0 35696 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_372
timestamp 1586364061
transform 1 0 37628 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36708 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38088 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37076 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_385
timestamp 1586364061
transform 1 0 36524 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_389
timestamp 1586364061
transform 1 0 36892 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_393
timestamp 1586364061
transform 1 0 37260 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_4  FILLER_24_398
timestamp 1586364061
transform 1 0 37720 0 -1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _300_
timestamp 1586364061
transform 1 0 40480 0 -1 15776
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38272 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40296 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_413
timestamp 1586364061
transform 1 0 39100 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_425
timestamp 1586364061
transform 1 0 40204 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__305__B
timestamp 1586364061
transform 1 0 42228 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41768 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_437
timestamp 1586364061
transform 1 0 41308 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_441
timestamp 1586364061
transform 1 0 41676 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_444
timestamp 1586364061
transform 1 0 41952 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_449
timestamp 1586364061
transform 1 0 42412 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_373
timestamp 1586364061
transform 1 0 43240 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_457
timestamp 1586364061
transform 1 0 43148 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_462
timestamp 1586364061
transform 1 0 43608 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_474
timestamp 1586364061
transform 1 0 44712 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_486
timestamp 1586364061
transform 1 0 45816 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_498
timestamp 1586364061
transform 1 0 46920 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 48852 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_6  FILLER_24_510
timestamp 1586364061
transform 1 0 48024 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_374
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_25_90
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_97
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_101
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_375
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 590 592
use scs8hd_fill_2  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_127
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_140
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_148
timestamp 1586364061
transform 1 0 14720 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_144
timestamp 1586364061
transform 1 0 14352 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_151
timestamp 1586364061
transform 1 0 14996 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15180 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_158
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _374_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_376
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__374__A
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_162
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _180_
timestamp 1586364061
transform 1 0 19872 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 19688 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__375__A
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_193
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_197
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_201
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_25_213
timestamp 1586364061
transform 1 0 20700 0 1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_221
timestamp 1586364061
transform 1 0 21436 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_240
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24012 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_377
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 1 15776
box -38 -48 866 592
use scs8hd_fill_2  FILLER_25_260
timestamp 1586364061
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_264
timestamp 1586364061
transform 1 0 25392 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25208 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25760 0 1 15776
box -38 -48 866 592
use scs8hd_nor2_4  _200_
timestamp 1586364061
transform 1 0 27600 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 27416 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26772 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_277
timestamp 1586364061
transform 1 0 26588 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_281
timestamp 1586364061
transform 1 0 26956 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_285
timestamp 1586364061
transform 1 0 27324 0 1 15776
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 30084 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_378
timestamp 1586364061
transform 1 0 29164 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 29900 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__318__A
timestamp 1586364061
transform 1 0 29532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_297
timestamp 1586364061
transform 1 0 28428 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_301
timestamp 1586364061
transform 1 0 28796 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  FILLER_25_306
timestamp 1586364061
transform 1 0 29256 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_311
timestamp 1586364061
transform 1 0 29716 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31832 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32844 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31648 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_326
timestamp 1586364061
transform 1 0 31096 0 1 15776
box -38 -48 590 592
use scs8hd_fill_2  FILLER_25_343
timestamp 1586364061
transform 1 0 32660 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_347
timestamp 1586364061
transform 1 0 33028 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33212 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33396 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_354
timestamp 1586364061
transform 1 0 33672 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33856 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_358
timestamp 1586364061
transform 1 0 34040 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_362
timestamp 1586364061
transform 1 0 34408 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_367
timestamp 1586364061
transform 1 0 34868 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_379
timestamp 1586364061
transform 1 0 34776 0 1 15776
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35052 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_372
timestamp 1586364061
transform 1 0 35328 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 35512 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 36064 0 1 15776
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38088 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 35880 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37720 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37260 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_376
timestamp 1586364061
transform 1 0 35696 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_391
timestamp 1586364061
transform 1 0 37076 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_395
timestamp 1586364061
transform 1 0 37444 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_400
timestamp 1586364061
transform 1 0 37904 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch
timestamp 1586364061
transform 1 0 40480 0 1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_380
timestamp 1586364061
transform 1 0 40388 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 40204 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__301__A
timestamp 1586364061
transform 1 0 39376 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__301__B
timestamp 1586364061
transform 1 0 39744 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_411
timestamp 1586364061
transform 1 0 38916 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_415
timestamp 1586364061
transform 1 0 39284 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_418
timestamp 1586364061
transform 1 0 39560 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_422
timestamp 1586364061
transform 1 0 39928 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _305_
timestamp 1586364061
transform 1 0 42228 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__305__A
timestamp 1586364061
transform 1 0 42044 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41676 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_439
timestamp 1586364061
transform 1 0 41492 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_443
timestamp 1586364061
transform 1 0 41860 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_456
timestamp 1586364061
transform 1 0 43056 0 1 15776
box -38 -48 314 592
use scs8hd_conb_1  _438_
timestamp 1586364061
transform 1 0 43792 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43332 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44252 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_461
timestamp 1586364061
transform 1 0 43516 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_467
timestamp 1586364061
transform 1 0 44068 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_471
timestamp 1586364061
transform 1 0 44436 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_25_483
timestamp 1586364061
transform 1 0 45540 0 1 15776
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_381
timestamp 1586364061
transform 1 0 46000 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_487
timestamp 1586364061
transform 1 0 45908 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_489
timestamp 1586364061
transform 1 0 46092 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_501
timestamp 1586364061
transform 1 0 47196 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 48852 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_25_513
timestamp 1586364061
transform 1 0 48300 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_382
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_390
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_90
timestamp 1586364061
transform 1 0 9384 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__366__B
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__366__A
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_383
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_94
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
timestamp 1586364061
transform 1 0 9936 0 -1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_26_107
timestamp 1586364061
transform 1 0 10948 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_4  FILLER_27_115
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_109
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_26_115
timestamp 1586364061
transform 1 0 11684 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_119
timestamp 1586364061
transform 1 0 12052 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_123
timestamp 1586364061
transform 1 0 12420 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_391
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_133
timestamp 1586364061
transform 1 0 13340 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_140
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_8  _133_
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_153
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_384
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_157
timestamp 1586364061
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15364 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_8  _134_
timestamp 1586364061
transform 1 0 15916 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_170
timestamp 1586364061
transform 1 0 16744 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_3  FILLER_27_178
timestamp 1586364061
transform 1 0 17480 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_174
timestamp 1586364061
transform 1 0 17112 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_180
timestamp 1586364061
transform 1 0 17664 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__374__B
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_392
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_26_186
timestamp 1586364061
transform 1 0 18216 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_27_199
timestamp 1586364061
transform 1 0 19412 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_195
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _375_
timestamp 1586364061
transform 1 0 18768 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_1  FILLER_27_207
timestamp 1586364061
transform 1 0 20148 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_206
timestamp 1586364061
transform 1 0 20056 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_26_201
timestamp 1586364061
transform 1 0 19596 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__B
timestamp 1586364061
transform 1 0 19872 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch_D
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_13_.latch
timestamp 1586364061
transform 1 0 20424 0 1 16864
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_26_212
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_385
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_221
timestamp 1586364061
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_222
timestamp 1586364061
transform 1 0 21528 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21068 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_15_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21252 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_234
timestamp 1586364061
transform 1 0 22632 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_27_225
timestamp 1586364061
transform 1 0 21804 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_229
timestamp 1586364061
transform 1 0 22172 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_226
timestamp 1586364061
transform 1 0 21896 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22172 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_7_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22264 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22356 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_240
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23276 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_250
timestamp 1586364061
transform 1 0 24104 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_243
timestamp 1586364061
transform 1 0 23460 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_393
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23828 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_27_258
timestamp 1586364061
transform 1 0 24840 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_254
timestamp 1586364061
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_254
timestamp 1586364061
transform 1 0 24472 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24288 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_1  FILLER_27_262
timestamp 1586364061
transform 1 0 25208 0 1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_267
timestamp 1586364061
transform 1 0 25668 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25300 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25484 0 1 16864
box -38 -48 866 592
use scs8hd_fill_1  FILLER_27_280
timestamp 1586364061
transform 1 0 26864 0 1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_274
timestamp 1586364061
transform 1 0 26312 0 1 16864
box -38 -48 590 592
use scs8hd_decap_8  FILLER_26_279
timestamp 1586364061
transform 1 0 26772 0 -1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_386
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_283
timestamp 1586364061
transform 1 0 27140 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_289
timestamp 1586364061
transform 1 0 27692 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26956 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__B
timestamp 1586364061
transform 1 0 27508 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 27324 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
timestamp 1586364061
transform 1 0 27876 0 -1 16864
box -38 -48 1050 592
use scs8hd_nor2_4  _202_
timestamp 1586364061
transform 1 0 27508 0 1 16864
box -38 -48 866 592
use scs8hd_fill_1  FILLER_27_304
timestamp 1586364061
transform 1 0 29072 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_300
timestamp 1586364061
transform 1 0 28704 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_296
timestamp 1586364061
transform 1 0 28336 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_302
timestamp 1586364061
transform 1 0 28888 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28888 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28520 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_394
timestamp 1586364061
transform 1 0 29164 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_313
timestamp 1586364061
transform 1 0 29900 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_309
timestamp 1586364061
transform 1 0 29532 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_308
timestamp 1586364061
transform 1 0 29440 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29256 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__323__A
timestamp 1586364061
transform 1 0 29992 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 16864
box -38 -48 314 592
use scs8hd_nor2_4  _318_
timestamp 1586364061
transform 1 0 29624 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_27_320
timestamp 1586364061
transform 1 0 30544 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_316
timestamp 1586364061
transform 1 0 30176 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_319
timestamp 1586364061
transform 1 0 30452 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__323__B
timestamp 1586364061
transform 1 0 30360 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_328
timestamp 1586364061
transform 1 0 31280 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_26_325
timestamp 1586364061
transform 1 0 31004 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31096 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30912 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31096 0 1 16864
box -38 -48 866 592
use scs8hd_decap_8  FILLER_27_335
timestamp 1586364061
transform 1 0 31924 0 1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_26_337
timestamp 1586364061
transform 1 0 32108 0 -1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_387
timestamp 1586364061
transform 1 0 32016 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32476 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_345
timestamp 1586364061
transform 1 0 32844 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_348
timestamp 1586364061
transform 1 0 33120 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_344
timestamp 1586364061
transform 1 0 32752 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32660 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33028 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_358
timestamp 1586364061
transform 1 0 34040 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_351
timestamp 1586364061
transform 1 0 33396 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33212 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33488 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_367
timestamp 1586364061
transform 1 0 34868 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_362
timestamp 1586364061
transform 1 0 34408 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_361
timestamp 1586364061
transform 1 0 34316 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__298__A
timestamp 1586364061
transform 1 0 34592 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_395
timestamp 1586364061
transform 1 0 34776 0 1 16864
box -38 -48 130 592
use scs8hd_decap_3  FILLER_26_375
timestamp 1586364061
transform 1 0 35604 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_371
timestamp 1586364061
transform 1 0 35236 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35420 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__298__B
timestamp 1586364061
transform 1 0 35052 0 -1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _298_
timestamp 1586364061
transform 1 0 35052 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_382
timestamp 1586364061
transform 1 0 36248 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_378
timestamp 1586364061
transform 1 0 35880 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36064 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36432 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36616 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 35880 0 -1 16864
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_27_395
timestamp 1586364061
transform 1 0 37444 0 1 16864
box -38 -48 406 592
use scs8hd_decap_4  FILLER_26_393
timestamp 1586364061
transform 1 0 37260 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_389
timestamp 1586364061
transform 1 0 36892 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37076 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__303__A
timestamp 1586364061
transform 1 0 37812 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_388
timestamp 1586364061
transform 1 0 37628 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37720 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_401
timestamp 1586364061
transform 1 0 37996 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_401
timestamp 1586364061
transform 1 0 37996 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_409
timestamp 1586364061
transform 1 0 38732 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_405
timestamp 1586364061
transform 1 0 38364 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38916 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__302__B
timestamp 1586364061
transform 1 0 38548 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__303__B
timestamp 1586364061
transform 1 0 38180 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__302__A
timestamp 1586364061
transform 1 0 38272 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _302_
timestamp 1586364061
transform 1 0 38456 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_419
timestamp 1586364061
transform 1 0 39652 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_415
timestamp 1586364061
transform 1 0 39284 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_413
timestamp 1586364061
transform 1 0 39100 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39836 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 39468 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _301_
timestamp 1586364061
transform 1 0 39376 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_423
timestamp 1586364061
transform 1 0 40020 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_425
timestamp 1586364061
transform 1 0 40204 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40480 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_396
timestamp 1586364061
transform 1 0 40388 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40480 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_441
timestamp 1586364061
transform 1 0 41676 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_437
timestamp 1586364061
transform 1 0 41308 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_430
timestamp 1586364061
transform 1 0 40664 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40848 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 41492 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41032 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_445
timestamp 1586364061
transform 1 0 42044 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_451
timestamp 1586364061
transform 1 0 42596 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_6  FILLER_26_443
timestamp 1586364061
transform 1 0 41860 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 41860 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 42412 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 42228 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 42412 0 1 16864
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_26_455
timestamp 1586364061
transform 1 0 42964 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43056 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_464
timestamp 1586364061
transform 1 0 43792 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_460
timestamp 1586364061
transform 1 0 43424 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_468
timestamp 1586364061
transform 1 0 44160 0 -1 16864
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43608 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43976 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_389
timestamp 1586364061
transform 1 0 43240 0 -1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44160 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_6  FILLER_27_481
timestamp 1586364061
transform 1 0 45356 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_477
timestamp 1586364061
transform 1 0 44988 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_480
timestamp 1586364061
transform 1 0 45264 0 -1 16864
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45172 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_397
timestamp 1586364061
transform 1 0 46000 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_492
timestamp 1586364061
transform 1 0 46368 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_504
timestamp 1586364061
transform 1 0 47472 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_487
timestamp 1586364061
transform 1 0 45908 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_489
timestamp 1586364061
transform 1 0 46092 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_501
timestamp 1586364061
transform 1 0 47196 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 48852 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 48852 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_513
timestamp 1586364061
transform 1 0 48300 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_398
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_nor2_4  _366_
timestamp 1586364061
transform 1 0 9752 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_399
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_103
timestamp 1586364061
transform 1 0 10580 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_107
timestamp 1586364061
transform 1 0 10948 0 -1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 17952
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_122
timestamp 1586364061
transform 1 0 12328 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_126
timestamp 1586364061
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_400
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_139
timestamp 1586364061
transform 1 0 13892 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_28_151
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_168
timestamp 1586364061
transform 1 0 16560 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_180
timestamp 1586364061
transform 1 0 17664 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_186
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_401
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 19872 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18400 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_201
timestamp 1586364061
transform 1 0 19596 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_210
timestamp 1586364061
transform 1 0 20424 0 -1 17952
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_LATCH_mem.LATCH_12_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_226
timestamp 1586364061
transform 1 0 21896 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_230
timestamp 1586364061
transform 1 0 22264 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_238
timestamp 1586364061
transform 1 0 23000 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24656 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25668 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_248
timestamp 1586364061
transform 1 0 23920 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_265
timestamp 1586364061
transform 1 0 25484 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26956 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27968 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_402
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27600 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_269
timestamp 1586364061
transform 1 0 25852 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_4  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_280
timestamp 1586364061
transform 1 0 26864 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_284
timestamp 1586364061
transform 1 0 27232 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_290
timestamp 1586364061
transform 1 0 27784 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _323_
timestamp 1586364061
transform 1 0 29992 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_12  FILLER_28_301
timestamp 1586364061
transform 1 0 28796 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_313
timestamp 1586364061
transform 1 0 29900 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_327
timestamp 1586364061
transform 1 0 31188 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_323
timestamp 1586364061
transform 1 0 30820 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31372 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31004 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_335
timestamp 1586364061
transform 1 0 31924 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_331
timestamp 1586364061
transform 1 0 31556 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_403
timestamp 1586364061
transform 1 0 32016 0 -1 17952
box -38 -48 130 592
use scs8hd_conb_1  _436_
timestamp 1586364061
transform 1 0 32108 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_348
timestamp 1586364061
transform 1 0 33120 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_340
timestamp 1586364061
transform 1 0 32384 0 -1 17952
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33396 0 -1 17952
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34960 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33212 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_360
timestamp 1586364061
transform 1 0 34224 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_8  FILLER_28_377
timestamp 1586364061
transform 1 0 35788 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36524 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_392
timestamp 1586364061
transform 1 0 37168 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_388
timestamp 1586364061
transform 1 0 36800 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37352 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36984 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_398
timestamp 1586364061
transform 1 0 37720 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_396
timestamp 1586364061
transform 1 0 37536 0 -1 17952
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_404
timestamp 1586364061
transform 1 0 37628 0 -1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _303_
timestamp 1586364061
transform 1 0 37812 0 -1 17952
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 39376 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40572 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38824 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_408
timestamp 1586364061
transform 1 0 38640 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_412
timestamp 1586364061
transform 1 0 39008 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_427
timestamp 1586364061
transform 1 0 40388 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 41124 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43056 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_431
timestamp 1586364061
transform 1 0 40756 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_8  FILLER_28_446
timestamp 1586364061
transform 1 0 42136 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_454
timestamp 1586364061
transform 1 0 42872 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44896 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_405
timestamp 1586364061
transform 1 0 43240 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_468
timestamp 1586364061
transform 1 0 44160 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_12  FILLER_28_479
timestamp 1586364061
transform 1 0 45172 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_491
timestamp 1586364061
transform 1 0 46276 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_503
timestamp 1586364061
transform 1 0 47380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 48852 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_515
timestamp 1586364061
transform 1 0 48484 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_406
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_nor2_4  _367_
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__367__A
timestamp 1586364061
transform 1 0 9568 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__367__B
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_90
timestamp 1586364061
transform 1 0 9384 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_103
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_107
timestamp 1586364061
transform 1 0 10948 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_407
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_120
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_137
timestamp 1586364061
transform 1 0 13708 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13892 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_141
timestamp 1586364061
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_145
timestamp 1586364061
transform 1 0 14444 0 1 17952
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14536 0 1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_29_153
timestamp 1586364061
transform 1 0 15180 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_149
timestamp 1586364061
transform 1 0 14812 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_163
timestamp 1586364061
transform 1 0 16100 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_187
timestamp 1586364061
transform 1 0 18308 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_408
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_195
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_191
timestamp 1586364061
transform 1 0 18676 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 18492 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_203
timestamp 1586364061
transform 1 0 19780 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_199
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _176_
timestamp 1586364061
transform 1 0 19872 0 1 17952
box -38 -48 866 592
use scs8hd_decap_6  FILLER_29_213
timestamp 1586364061
transform 1 0 20700 0 1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21988 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_219
timestamp 1586364061
transform 1 0 21252 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_222
timestamp 1586364061
transform 1 0 21528 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_236
timestamp 1586364061
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_240
timestamp 1586364061
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_409
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_29_258
timestamp 1586364061
transform 1 0 24840 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_254
timestamp 1586364061
transform 1 0 24472 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 24656 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_262
timestamp 1586364061
transform 1 0 25208 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25392 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25576 0 1 17952
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27416 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 26956 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_275
timestamp 1586364061
transform 1 0 26404 0 1 17952
box -38 -48 590 592
use scs8hd_decap_3  FILLER_29_283
timestamp 1586364061
transform 1 0 27140 0 1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_29_304
timestamp 1586364061
transform 1 0 29072 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_301
timestamp 1586364061
transform 1 0 28796 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_297
timestamp 1586364061
transform 1 0 28428 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__324__A
timestamp 1586364061
transform 1 0 28888 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_410
timestamp 1586364061
transform 1 0 29164 0 1 17952
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_317
timestamp 1586364061
transform 1 0 30268 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_313
timestamp 1586364061
transform 1 0 29900 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_309
timestamp 1586364061
transform 1 0 29532 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30084 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__324__B
timestamp 1586364061
transform 1 0 29716 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 30452 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 30636 0 1 17952
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33120 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32108 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32936 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_332
timestamp 1586364061
transform 1 0 31648 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_336
timestamp 1586364061
transform 1 0 32016 0 1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_29_339
timestamp 1586364061
transform 1 0 32292 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_345
timestamp 1586364061
transform 1 0 32844 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_351
timestamp 1586364061
transform 1 0 33396 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33580 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_355
timestamp 1586364061
transform 1 0 33764 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33948 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_363
timestamp 1586364061
transform 1 0 34500 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_359
timestamp 1586364061
transform 1 0 34132 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34592 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_411
timestamp 1586364061
transform 1 0 34776 0 1 17952
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34868 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_370
timestamp 1586364061
transform 1 0 35144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35328 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_374
timestamp 1586364061
transform 1 0 35512 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_382
timestamp 1586364061
transform 1 0 36248 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_378
timestamp 1586364061
transform 1 0 35880 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35696 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36340 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36524 0 1 17952
box -38 -48 866 592
use scs8hd_fill_2  FILLER_29_394
timestamp 1586364061
transform 1 0 37352 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_398
timestamp 1586364061
transform 1 0 37720 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37536 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37904 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38088 0 1 17952
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40480 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_412
timestamp 1586364061
transform 1 0 40388 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40204 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39836 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39100 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_411
timestamp 1586364061
transform 1 0 38916 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_415
timestamp 1586364061
transform 1 0 39284 0 1 17952
box -38 -48 590 592
use scs8hd_fill_2  FILLER_29_423
timestamp 1586364061
transform 1 0 40020 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42964 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41492 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42780 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41860 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_437
timestamp 1586364061
transform 1 0 41308 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_441
timestamp 1586364061
transform 1 0 41676 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_445
timestamp 1586364061
transform 1 0 42044 0 1 17952
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43976 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_464
timestamp 1586364061
transform 1 0 43792 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_468
timestamp 1586364061
transform 1 0 44160 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_480
timestamp 1586364061
transform 1 0 45264 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_413
timestamp 1586364061
transform 1 0 46000 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_489
timestamp 1586364061
transform 1 0 46092 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_501
timestamp 1586364061
transform 1 0 47196 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 48852 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_513
timestamp 1586364061
transform 1 0 48300 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_414
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10396 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_415
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_104
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_8  _136_
timestamp 1586364061
transform 1 0 11960 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_108
timestamp 1586364061
transform 1 0 11040 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_112
timestamp 1586364061
transform 1 0 11408 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_3  FILLER_30_127
timestamp 1586364061
transform 1 0 12788 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_132
timestamp 1586364061
transform 1 0 13248 0 -1 19040
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_416
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_144
timestamp 1586364061
transform 1 0 14352 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_152
timestamp 1586364061
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_160
timestamp 1586364061
transform 1 0 15824 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_8  _131_
timestamp 1586364061
transform 1 0 16560 0 -1 19040
box -38 -48 866 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 18124 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17940 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_177
timestamp 1586364061
transform 1 0 17388 0 -1 19040
box -38 -48 590 592
use scs8hd_or4_4  _166_
timestamp 1586364061
transform 1 0 19228 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_417
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__406__C
timestamp 1586364061
transform 1 0 19044 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__384__D
timestamp 1586364061
transform 1 0 18676 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__362__D
timestamp 1586364061
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_188
timestamp 1586364061
transform 1 0 18400 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_193
timestamp 1586364061
transform 1 0 18860 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_206
timestamp 1586364061
transform 1 0 20056 0 -1 19040
box -38 -48 590 592
use scs8hd_inv_8  _158_
timestamp 1586364061
transform 1 0 22356 0 -1 19040
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21344 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__362__A
timestamp 1586364061
transform 1 0 21068 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_219
timestamp 1586364061
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_223
timestamp 1586364061
transform 1 0 21620 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_229
timestamp 1586364061
transform 1 0 22172 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_240
timestamp 1586364061
transform 1 0 23184 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_247
timestamp 1586364061
transform 1 0 23828 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_244
timestamp 1586364061
transform 1 0 23552 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l1_in_6_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_8  _157_
timestamp 1586364061
transform 1 0 23920 0 -1 19040
box -38 -48 866 592
use scs8hd_fill_2  FILLER_30_261
timestamp 1586364061
transform 1 0 25116 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_257
timestamp 1586364061
transform 1 0 24748 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24932 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_265
timestamp 1586364061
transform 1 0 25484 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25668 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_8  _156_
timestamp 1586364061
transform 1 0 26956 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_418
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26680 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_269
timestamp 1586364061
transform 1 0 25852 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_280
timestamp 1586364061
transform 1 0 26864 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_290
timestamp 1586364061
transform 1 0 27784 0 -1 19040
box -38 -48 1142 592
use scs8hd_nor2_4  _324_
timestamp 1586364061
transform 1 0 28888 0 -1 19040
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30452 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29900 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30268 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_311
timestamp 1586364061
transform 1 0 29716 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_315
timestamp 1586364061
transform 1 0 30084 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32108 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_419
timestamp 1586364061
transform 1 0 32016 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32844 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_328
timestamp 1586364061
transform 1 0 31280 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_4  FILLER_30_340
timestamp 1586364061
transform 1 0 32384 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_344
timestamp 1586364061
transform 1 0 32752 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_347
timestamp 1586364061
transform 1 0 33028 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35052 0 -1 19040
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33488 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33212 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_351
timestamp 1586364061
transform 1 0 33396 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_361
timestamp 1586364061
transform 1 0 34316 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36616 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38088 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_420
timestamp 1586364061
transform 1 0 37628 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37076 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_378
timestamp 1586364061
transform 1 0 35880 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_389
timestamp 1586364061
transform 1 0 36892 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_393
timestamp 1586364061
transform 1 0 37260 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_4  FILLER_30_398
timestamp 1586364061
transform 1 0 37720 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40388 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40112 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39100 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_411
timestamp 1586364061
transform 1 0 38916 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_415
timestamp 1586364061
transform 1 0 39284 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_30_423
timestamp 1586364061
transform 1 0 40020 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_426
timestamp 1586364061
transform 1 0 40296 0 -1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41400 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42964 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_430
timestamp 1586364061
transform 1 0 40664 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_8  FILLER_30_447
timestamp 1586364061
transform 1 0 42228 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_421
timestamp 1586364061
transform 1 0 43240 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_457
timestamp 1586364061
transform 1 0 43148 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_462
timestamp 1586364061
transform 1 0 43608 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_474
timestamp 1586364061
transform 1 0 44712 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_486
timestamp 1586364061
transform 1 0 45816 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_498
timestamp 1586364061
transform 1 0 46920 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 48852 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_6  FILLER_30_510
timestamp 1586364061
transform 1 0 48024 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_422
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_31_94
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_97
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_101
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_423
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13064 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 590 592
use scs8hd_decap_4  FILLER_31_126
timestamp 1586364061
transform 1 0 12696 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_132
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _435_
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_145
timestamp 1586364061
transform 1 0 14444 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_158
timestamp 1586364061
transform 1 0 15640 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_162
timestamp 1586364061
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use scs8hd_inv_8  _132_
timestamp 1586364061
transform 1 0 16376 0 1 19040
box -38 -48 866 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_187
timestamp 1586364061
transform 1 0 18308 0 1 19040
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_424
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 314 592
use scs8hd_or4_4  _406_
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20792 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__406__A
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__406__B
timestamp 1586364061
transform 1 0 18676 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__384__B
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__384__A
timestamp 1586364061
transform 1 0 20608 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_193
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_206
timestamp 1586364061
transform 1 0 20056 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_210
timestamp 1586364061
transform 1 0 20424 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_217
timestamp 1586364061
transform 1 0 21068 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__362__B
timestamp 1586364061
transform 1 0 21252 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_221
timestamp 1586364061
transform 1 0 21436 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_225
timestamp 1586364061
transform 1 0 21804 0 1 19040
box -38 -48 222 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_1_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 21988 0 1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_31_234
timestamp 1586364061
transform 1 0 22632 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_230
timestamp 1586364061
transform 1 0 22264 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__362__C
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_240
timestamp 1586364061
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25300 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_425
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_254
timestamp 1586364061
transform 1 0 24472 0 1 19040
box -38 -48 406 592
use scs8hd_decap_3  FILLER_31_260
timestamp 1586364061
transform 1 0 25024 0 1 19040
box -38 -48 314 592
use scs8hd_inv_8  _155_
timestamp 1586364061
transform 1 0 27232 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26496 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__290__C
timestamp 1586364061
transform 1 0 28244 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 27048 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_272
timestamp 1586364061
transform 1 0 26128 0 1 19040
box -38 -48 406 592
use scs8hd_decap_4  FILLER_31_278
timestamp 1586364061
transform 1 0 26680 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_293
timestamp 1586364061
transform 1 0 28060 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 29808 0 1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_426
timestamp 1586364061
transform 1 0 29164 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 29624 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28980 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 28612 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_297
timestamp 1586364061
transform 1 0 28428 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_301
timestamp 1586364061
transform 1 0 28796 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_306
timestamp 1586364061
transform 1 0 29256 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_327
timestamp 1586364061
transform 1 0 31188 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_323
timestamp 1586364061
transform 1 0 30820 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31004 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_331
timestamp 1586364061
transform 1 0 31556 0 1 19040
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31372 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_341
timestamp 1586364061
transform 1 0 32476 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_337
timestamp 1586364061
transform 1 0 32108 0 1 19040
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32200 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_345
timestamp 1586364061
transform 1 0 32844 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33028 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32660 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_358
timestamp 1586364061
transform 1 0 34040 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 19040
box -38 -48 866 592
use scs8hd_fill_2  FILLER_31_362
timestamp 1586364061
transform 1 0 34408 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34592 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_427
timestamp 1586364061
transform 1 0 34776 0 1 19040
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34868 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_374
timestamp 1586364061
transform 1 0 35512 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_370
timestamp 1586364061
transform 1 0 35144 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35328 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_382
timestamp 1586364061
transform 1 0 36248 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_378
timestamp 1586364061
transform 1 0 35880 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35696 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36064 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36432 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_395
timestamp 1586364061
transform 1 0 37444 0 1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36616 0 1 19040
box -38 -48 866 592
use scs8hd_fill_2  FILLER_31_402
timestamp 1586364061
transform 1 0 38088 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_399
timestamp 1586364061
transform 1 0 37812 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37904 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_406
timestamp 1586364061
transform 1 0 38456 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__306__B
timestamp 1586364061
transform 1 0 38272 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__306__A
timestamp 1586364061
transform 1 0 38640 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _306_
timestamp 1586364061
transform 1 0 38824 0 1 19040
box -38 -48 866 592
use scs8hd_decap_4  FILLER_31_419
timestamp 1586364061
transform 1 0 39652 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_428
timestamp 1586364061
transform 1 0 40480 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_426
timestamp 1586364061
transform 1 0 40296 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_423
timestamp 1586364061
transform 1 0 40020 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 40112 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_428
timestamp 1586364061
transform 1 0 40388 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_437
timestamp 1586364061
transform 1 0 41308 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_433
timestamp 1586364061
transform 1 0 40940 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41492 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41124 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40664 0 1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 1 19040
box -38 -48 866 592
use scs8hd_fill_2  FILLER_31_454
timestamp 1586364061
transform 1 0 42872 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_450
timestamp 1586364061
transform 1 0 42504 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43056 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42688 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43240 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44896 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43700 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44068 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_461
timestamp 1586364061
transform 1 0 43516 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_465
timestamp 1586364061
transform 1 0 43884 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_469
timestamp 1586364061
transform 1 0 44252 0 1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_475
timestamp 1586364061
transform 1 0 44804 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_478
timestamp 1586364061
transform 1 0 45080 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_429
timestamp 1586364061
transform 1 0 46000 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_486
timestamp 1586364061
transform 1 0 45816 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_489
timestamp 1586364061
transform 1 0 46092 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_501
timestamp 1586364061
transform 1 0 47196 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 48852 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_513
timestamp 1586364061
transform 1 0 48300 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_430
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 9844 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10856 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_431
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_98
timestamp 1586364061
transform 1 0 10120 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_104
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_12  FILLER_32_115
timestamp 1586364061
transform 1 0 11684 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_32_127
timestamp 1586364061
transform 1 0 12788 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_432
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_139
timestamp 1586364061
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_143
timestamp 1586364061
transform 1 0 14260 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_151
timestamp 1586364061
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_163
timestamp 1586364061
transform 1 0 16100 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_167
timestamp 1586364061
transform 1 0 16468 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_175
timestamp 1586364061
transform 1 0 17204 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_171
timestamp 1586364061
transform 1 0 16836 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_179
timestamp 1586364061
transform 1 0 17572 0 -1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17940 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_186
timestamp 1586364061
transform 1 0 18216 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_193
timestamp 1586364061
transform 1 0 18860 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__406__D
timestamp 1586364061
transform 1 0 18676 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__384__C
timestamp 1586364061
transform 1 0 19044 0 -1 20128
box -38 -48 222 592
use scs8hd_or4_4  _384_
timestamp 1586364061
transform 1 0 19228 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_4  FILLER_32_206
timestamp 1586364061
transform 1 0 20056 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_213
timestamp 1586364061
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_210
timestamp 1586364061
transform 1 0 20424 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__330__B
timestamp 1586364061
transform 1 0 20516 0 -1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_433
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_or4_4  _362_
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23184 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_224
timestamp 1586364061
transform 1 0 21712 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_32_236
timestamp 1586364061
transform 1 0 22816 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24564 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l2_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_249
timestamp 1586364061
transform 1 0 24012 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_253
timestamp 1586364061
transform 1 0 24380 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_257
timestamp 1586364061
transform 1 0 24748 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_32_267
timestamp 1586364061
transform 1 0 25668 0 -1 20128
box -38 -48 590 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_0_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 28060 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_434
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__290__B
timestamp 1586364061
transform 1 0 27600 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26220 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_285
timestamp 1586364061
transform 1 0 27324 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_32_290
timestamp 1586364061
transform 1 0 27784 0 -1 20128
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29440 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30452 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__317__D
timestamp 1586364061
transform 1 0 28520 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29900 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_296
timestamp 1586364061
transform 1 0 28336 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_300
timestamp 1586364061
transform 1 0 28704 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_311
timestamp 1586364061
transform 1 0 29716 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_315
timestamp 1586364061
transform 1 0 30084 0 -1 20128
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32568 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_435
timestamp 1586364061
transform 1 0 32016 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_328
timestamp 1586364061
transform 1 0 31280 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_4  FILLER_32_337
timestamp 1586364061
transform 1 0 32108 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_341
timestamp 1586364061
transform 1 0 32476 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_345
timestamp 1586364061
transform 1 0 32844 0 -1 20128
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33580 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33212 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_351
timestamp 1586364061
transform 1 0 33396 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_362
timestamp 1586364061
transform 1 0 34408 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_32_374
timestamp 1586364061
transform 1 0 35512 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36064 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_436
timestamp 1586364061
transform 1 0 37628 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__295__A
timestamp 1586364061
transform 1 0 35696 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37904 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_378
timestamp 1586364061
transform 1 0 35880 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_389
timestamp 1586364061
transform 1 0 36892 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_398
timestamp 1586364061
transform 1 0 37720 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_402
timestamp 1586364061
transform 1 0 38088 0 -1 20128
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 40112 0 -1 20128
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38364 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_414
timestamp 1586364061
transform 1 0 39192 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_422
timestamp 1586364061
transform 1 0 39928 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41860 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41676 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41308 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_435
timestamp 1586364061
transform 1 0 41124 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_439
timestamp 1586364061
transform 1 0 41492 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_446
timestamp 1586364061
transform 1 0 42136 0 -1 20128
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 20128
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44896 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_437
timestamp 1586364061
transform 1 0 43240 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_468
timestamp 1586364061
transform 1 0 44160 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_479
timestamp 1586364061
transform 1 0 45172 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_491
timestamp 1586364061
transform 1 0 46276 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_503
timestamp 1586364061
transform 1 0 47380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 48852 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_32_515
timestamp 1586364061
transform 1 0 48484 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_446
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_438
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 590 592
use scs8hd_decap_8  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_100
timestamp 1586364061
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_96
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_92
timestamp 1586364061
transform 1 0 9568 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_447
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_101
timestamp 1586364061
transform 1 0 10396 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use scs8hd_inv_8  _138_
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 866 592
use scs8hd_inv_8  _137_
timestamp 1586364061
transform 1 0 10488 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_8  FILLER_34_111
timestamp 1586364061
transform 1 0 11316 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_6  FILLER_33_113
timestamp 1586364061
transform 1 0 11500 0 1 20128
box -38 -48 590 592
use scs8hd_decap_4  FILLER_34_124
timestamp 1586364061
transform 1 0 12512 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_119
timestamp 1586364061
transform 1 0 12052 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_127
timestamp 1586364061
transform 1 0 12788 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_119
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_439
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_131
timestamp 1586364061
transform 1 0 13156 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_128
timestamp 1586364061
transform 1 0 12880 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13248 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_8  _135_
timestamp 1586364061
transform 1 0 12972 0 1 20128
box -38 -48 866 592
use scs8hd_decap_12  FILLER_34_139
timestamp 1586364061
transform 1 0 13892 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_34_135
timestamp 1586364061
transform 1 0 13524 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_142
timestamp 1586364061
transform 1 0 14168 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_138
timestamp 1586364061
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13708 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_3.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14536 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_151
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_153
timestamp 1586364061
transform 1 0 15180 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_149
timestamp 1586364061
transform 1 0 14812 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15364 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_448
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_8  FILLER_34_165
timestamp 1586364061
transform 1 0 16284 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_170
timestamp 1586364061
transform 1 0 16744 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_166
timestamp 1586364061
transform 1 0 16376 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_175
timestamp 1586364061
transform 1 0 17204 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_174
timestamp 1586364061
transform 1 0 17112 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17388 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_4  FILLER_34_186
timestamp 1586364061
transform 1 0 18216 0 -1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_440
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_193
timestamp 1586364061
transform 1 0 18860 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_197
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_193
timestamp 1586364061
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19412 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__327__A
timestamp 1586364061
transform 1 0 18676 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_7_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 21216
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_34_206
timestamp 1586364061
transform 1 0 20056 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_4  FILLER_33_205
timestamp 1586364061
transform 1 0 19964 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_201
timestamp 1586364061
transform 1 0 19596 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__330__A
timestamp 1586364061
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _330_
timestamp 1586364061
transform 1 0 20516 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_449
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_224
timestamp 1586364061
transform 1 0 21712 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_224
timestamp 1586364061
transform 1 0 21712 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21528 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_8  FILLER_34_228
timestamp 1586364061
transform 1 0 22080 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_231
timestamp 1586364061
transform 1 0 22356 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22540 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22080 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_236
timestamp 1586364061
transform 1 0 22816 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_239
timestamp 1586364061
transform 1 0 23092 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_235
timestamp 1586364061
transform 1 0 22724 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 22908 0 1 20128
box -38 -48 222 592
use scs8hd_inv_8  _162_
timestamp 1586364061
transform 1 0 22908 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_4  FILLER_34_250
timestamp 1586364061
transform 1 0 24104 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_246
timestamp 1586364061
transform 1 0 23736 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23920 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_441
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l4_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 866 592
use scs8hd_fill_1  FILLER_34_254
timestamp 1586364061
transform 1 0 24472 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_258
timestamp 1586364061
transform 1 0 24840 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_254
timestamp 1586364061
transform 1 0 24472 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.mux_l3_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24564 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_8  FILLER_34_264
timestamp 1586364061
transform 1 0 25392 0 -1 21216
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 25208 0 1 20128
box -38 -48 222 592
use scs8hd_inv_8  _159_
timestamp 1586364061
transform 1 0 25392 0 1 20128
box -38 -48 866 592
use scs8hd_decap_3  FILLER_34_272
timestamp 1586364061
transform 1 0 26128 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_33_277
timestamp 1586364061
transform 1 0 26588 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_273
timestamp 1586364061
transform 1 0 26220 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__290__D
timestamp 1586364061
transform 1 0 26680 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_450
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__290__A
timestamp 1586364061
transform 1 0 27048 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_280
timestamp 1586364061
transform 1 0 26864 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_279
timestamp 1586364061
transform 1 0 26772 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_283
timestamp 1586364061
transform 1 0 27140 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__317__B
timestamp 1586364061
transform 1 0 27416 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__299__A
timestamp 1586364061
transform 1 0 27600 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__317__C
timestamp 1586364061
transform 1 0 27232 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_284
timestamp 1586364061
transform 1 0 27232 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_286
timestamp 1586364061
transform 1 0 27416 0 -1 21216
box -38 -48 222 592
use scs8hd_or4_4  _290_
timestamp 1586364061
transform 1 0 27600 0 1 20128
box -38 -48 866 592
use scs8hd_or4_4  _317_
timestamp 1586364061
transform 1 0 27784 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__317__A
timestamp 1586364061
transform 1 0 28612 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_297
timestamp 1586364061
transform 1 0 28428 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_299
timestamp 1586364061
transform 1 0 28612 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28980 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28796 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_301
timestamp 1586364061
transform 1 0 28796 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_303
timestamp 1586364061
transform 1 0 28980 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_442
timestamp 1586364061
transform 1 0 29164 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__325__B
timestamp 1586364061
transform 1 0 29256 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_306
timestamp 1586364061
transform 1 0 29256 0 1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_34_311
timestamp 1586364061
transform 1 0 29716 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_310
timestamp 1586364061
transform 1 0 29624 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 29716 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29440 0 -1 21216
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 29900 0 1 20128
box -38 -48 1050 592
use scs8hd_nor2_4  _322_
timestamp 1586364061
transform 1 0 30452 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_8  FILLER_34_328
timestamp 1586364061
transform 1 0 31280 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_4  FILLER_33_332
timestamp 1586364061
transform 1 0 31648 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_328
timestamp 1586364061
transform 1 0 31280 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_324
timestamp 1586364061
transform 1 0 30912 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__322__B
timestamp 1586364061
transform 1 0 31464 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__322__A
timestamp 1586364061
transform 1 0 31096 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_345
timestamp 1586364061
transform 1 0 32844 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_341
timestamp 1586364061
transform 1 0 32476 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32016 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 32660 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_451
timestamp 1586364061
transform 1 0 32016 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32200 0 1 20128
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 21216
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_34_348
timestamp 1586364061
transform 1 0 33120 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33028 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_352
timestamp 1586364061
transform 1 0 33488 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_358
timestamp 1586364061
transform 1 0 34040 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33672 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33304 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33856 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_365
timestamp 1586364061
transform 1 0 34684 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_362
timestamp 1586364061
transform 1 0 34408 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34868 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34592 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_443
timestamp 1586364061
transform 1 0 34776 0 1 20128
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34868 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_34_373
timestamp 1586364061
transform 1 0 35420 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_369
timestamp 1586364061
transform 1 0 35052 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_374
timestamp 1586364061
transform 1 0 35512 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_370
timestamp 1586364061
transform 1 0 35144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35236 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35328 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_385
timestamp 1586364061
transform 1 0 36524 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_33_378
timestamp 1586364061
transform 1 0 35880 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 35972 0 1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 36156 0 1 20128
box -38 -48 1050 592
use scs8hd_nor2_4  _295_
timestamp 1586364061
transform 1 0 35696 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36800 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37168 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_392
timestamp 1586364061
transform 1 0 37168 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_390
timestamp 1586364061
transform 1 0 36984 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_452
timestamp 1586364061
transform 1 0 37628 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__295__B
timestamp 1586364061
transform 1 0 37352 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37720 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_396
timestamp 1586364061
transform 1 0 37536 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_394
timestamp 1586364061
transform 1 0 37352 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_34_398
timestamp 1586364061
transform 1 0 37720 0 -1 21216
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37904 0 1 20128
box -38 -48 866 592
use scs8hd_decap_3  FILLER_34_412
timestamp 1586364061
transform 1 0 39008 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_34_407
timestamp 1586364061
transform 1 0 38548 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_413
timestamp 1586364061
transform 1 0 39100 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_409
timestamp 1586364061
transform 1 0 38732 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38824 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39284 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38916 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 39284 0 -1 21216
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 38272 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_424
timestamp 1586364061
transform 1 0 40112 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_33_428
timestamp 1586364061
transform 1 0 40480 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_421
timestamp 1586364061
transform 1 0 39836 0 1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_33_417
timestamp 1586364061
transform 1 0 39468 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39652 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_444
timestamp 1586364061
transform 1 0 40388 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_432
timestamp 1586364061
transform 1 0 40848 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40664 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41032 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41216 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41216 0 1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_34_449
timestamp 1586364061
transform 1 0 42412 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_445
timestamp 1586364061
transform 1 0 42044 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_449
timestamp 1586364061
transform 1 0 42412 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_445
timestamp 1586364061
transform 1 0 42044 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42228 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__307__B
timestamp 1586364061
transform 1 0 42228 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_456
timestamp 1586364061
transform 1 0 43056 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42596 0 1 20128
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42780 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_453
timestamp 1586364061
transform 1 0 43240 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43240 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43608 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_460
timestamp 1586364061
transform 1 0 43424 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_457
timestamp 1586364061
transform 1 0 43148 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43792 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44252 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_467
timestamp 1586364061
transform 1 0 44068 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_468
timestamp 1586364061
transform 1 0 44160 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_12  FILLER_34_472
timestamp 1586364061
transform 1 0 44528 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_471
timestamp 1586364061
transform 1 0 44436 0 1 20128
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44344 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_483
timestamp 1586364061
transform 1 0 45540 0 1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_445
timestamp 1586364061
transform 1 0 46000 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_487
timestamp 1586364061
transform 1 0 45908 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_489
timestamp 1586364061
transform 1 0 46092 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_501
timestamp 1586364061
transform 1 0 47196 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_484
timestamp 1586364061
transform 1 0 45632 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_496
timestamp 1586364061
transform 1 0 46736 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_508
timestamp 1586364061
transform 1 0 47840 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 48852 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 48852 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_33_513
timestamp 1586364061
transform 1 0 48300 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_454
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_35_106
timestamp 1586364061
transform 1 0 10856 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_114
timestamp 1586364061
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__332__B
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__332__A
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12696 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_455
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12880 0 1 21216
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15180 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_139
timestamp 1586364061
transform 1 0 13892 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_143
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_149
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_162
timestamp 1586364061
transform 1 0 16008 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_166
timestamp 1586364061
transform 1 0 16376 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_173
timestamp 1586364061
transform 1 0 17020 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_177
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_181
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_456
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_188
timestamp 1586364061
transform 1 0 18400 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _327_
timestamp 1586364061
transform 1 0 18676 0 1 21216
box -38 -48 866 592
use scs8hd_decap_4  FILLER_35_204
timestamp 1586364061
transform 1 0 19872 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_200
timestamp 1586364061
transform 1 0 19504 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19688 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_211
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20332 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 20700 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 20884 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 22632 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22080 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_226
timestamp 1586364061
transform 1 0 21896 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_230
timestamp 1586364061
transform 1 0 22264 0 1 21216
box -38 -48 406 592
use scs8hd_decap_8  FILLER_35_236
timestamp 1586364061
transform 1 0 22816 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_248
timestamp 1586364061
transform 1 0 23920 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_457
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_260
timestamp 1586364061
transform 1 0 25024 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_256
timestamp 1586364061
transform 1 0 24656 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_252
timestamp 1586364061
transform 1 0 24288 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 24840 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 24472 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 25300 0 1 21216
box -38 -48 222 592
use scs8hd_inv_8  _160_
timestamp 1586364061
transform 1 0 25484 0 1 21216
box -38 -48 866 592
use scs8hd_or4_4  _299_
timestamp 1586364061
transform 1 0 27600 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 26496 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__299__B
timestamp 1586364061
transform 1 0 27416 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__299__C
timestamp 1586364061
transform 1 0 27048 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_274
timestamp 1586364061
transform 1 0 26312 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_278
timestamp 1586364061
transform 1 0 26680 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_284
timestamp 1586364061
transform 1 0 27232 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _325_
timestamp 1586364061
transform 1 0 29256 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_458
timestamp 1586364061
transform 1 0 29164 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__325__A
timestamp 1586364061
transform 1 0 28980 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30728 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_297
timestamp 1586364061
transform 1 0 28428 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_301
timestamp 1586364061
transform 1 0 28796 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_315
timestamp 1586364061
transform 1 0 30084 0 1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_35_321
timestamp 1586364061
transform 1 0 30636 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_331
timestamp 1586364061
transform 1 0 31556 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_327
timestamp 1586364061
transform 1 0 31188 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31372 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30912 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_338
timestamp 1586364061
transform 1 0 32200 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31740 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32384 0 1 21216
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31924 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_342
timestamp 1586364061
transform 1 0 32568 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32752 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32936 0 1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_459
timestamp 1586364061
transform 1 0 34776 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33948 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_355
timestamp 1586364061
transform 1 0 33764 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_359
timestamp 1586364061
transform 1 0 34132 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_363
timestamp 1586364061
transform 1 0 34500 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_384
timestamp 1586364061
transform 1 0 36432 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_380
timestamp 1586364061
transform 1 0 36064 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_376
timestamp 1586364061
transform 1 0 35696 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36248 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36616 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36800 0 1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_35_402
timestamp 1586364061
transform 1 0 38088 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_397
timestamp 1586364061
transform 1 0 37628 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 37904 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_406
timestamp 1586364061
transform 1 0 38456 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38272 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38640 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38824 0 1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_35_419
timestamp 1586364061
transform 1 0 39652 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39836 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_423
timestamp 1586364061
transform 1 0 40020 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40204 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_460
timestamp 1586364061
transform 1 0 40388 0 1 21216
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 21216
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 42136 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 41952 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40940 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__307__A
timestamp 1586364061
transform 1 0 41400 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_431
timestamp 1586364061
transform 1 0 40756 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_435
timestamp 1586364061
transform 1 0 41124 0 1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_35_440
timestamp 1586364061
transform 1 0 41584 0 1 21216
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43884 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43332 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43700 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44896 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_457
timestamp 1586364061
transform 1 0 43148 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_461
timestamp 1586364061
transform 1 0 43516 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_474
timestamp 1586364061
transform 1 0 44712 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_478
timestamp 1586364061
transform 1 0 45080 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_461
timestamp 1586364061
transform 1 0 46000 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_486
timestamp 1586364061
transform 1 0 45816 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_489
timestamp 1586364061
transform 1 0 46092 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_501
timestamp 1586364061
transform 1 0 47196 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 48852 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_513
timestamp 1586364061
transform 1 0 48300 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_462
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_463
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 590 592
use scs8hd_nor2_4  _332_
timestamp 1586364061
transform 1 0 11408 0 -1 22304
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_111
timestamp 1586364061
transform 1 0 11316 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_121
timestamp 1586364061
transform 1 0 12236 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_464
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_140
timestamp 1586364061
transform 1 0 13984 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_146
timestamp 1586364061
transform 1 0 14536 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_149
timestamp 1586364061
transform 1 0 14812 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_8  FILLER_36_163
timestamp 1586364061
transform 1 0 16100 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_171
timestamp 1586364061
transform 1 0 16836 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_182
timestamp 1586364061
transform 1 0 17848 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 -1 22304
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_465
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__327__B
timestamp 1586364061
transform 1 0 19044 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_193
timestamp 1586364061
transform 1 0 18860 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_197
timestamp 1586364061
transform 1 0 19228 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_204
timestamp 1586364061
transform 1 0 19872 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_212
timestamp 1586364061
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_8  _161_
timestamp 1586364061
transform 1 0 22632 0 -1 22304
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 -1 22304
box -38 -48 866 592
use scs8hd_fill_2  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_226
timestamp 1586364061
transform 1 0 21896 0 -1 22304
box -38 -48 774 592
use scs8hd_or2_4  _165_
timestamp 1586364061
transform 1 0 24472 0 -1 22304
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23644 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_243
timestamp 1586364061
transform 1 0 23460 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_247
timestamp 1586364061
transform 1 0 23828 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_253
timestamp 1586364061
transform 1 0 24380 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_261
timestamp 1586364061
transform 1 0 25116 0 -1 22304
box -38 -48 1142 592
use scs8hd_inv_8  _129_
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 28060 0 -1 22304
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_466
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__299__D
timestamp 1586364061
transform 1 0 27600 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_273
timestamp 1586364061
transform 1 0 26220 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_285
timestamp 1586364061
transform 1 0 27324 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_36_290
timestamp 1586364061
transform 1 0 27784 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29716 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30084 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_304
timestamp 1586364061
transform 1 0 29072 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_310
timestamp 1586364061
transform 1 0 29624 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_313
timestamp 1586364061
transform 1 0 29900 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_317
timestamp 1586364061
transform 1 0 30268 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31004 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_36_328
timestamp 1586364061
transform 1 0 31280 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__309__B
timestamp 1586364061
transform 1 0 31556 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_333
timestamp 1586364061
transform 1 0 31740 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_467
timestamp 1586364061
transform 1 0 32016 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_341
timestamp 1586364061
transform 1 0 32476 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_337
timestamp 1586364061
transform 1 0 32108 0 -1 22304
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_0.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32200 0 -1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_36_345
timestamp 1586364061
transform 1 0 32844 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32936 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_348
timestamp 1586364061
transform 1 0 33120 0 -1 22304
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 -1 22304
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35052 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 34500 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34868 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_358
timestamp 1586364061
transform 1 0 34040 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_362
timestamp 1586364061
transform 1 0 34408 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_365
timestamp 1586364061
transform 1 0 34684 0 -1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 37904 0 -1 22304
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36616 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_468
timestamp 1586364061
transform 1 0 37628 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__304__B
timestamp 1586364061
transform 1 0 37076 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_378
timestamp 1586364061
transform 1 0 35880 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_389
timestamp 1586364061
transform 1 0 36892 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_393
timestamp 1586364061
transform 1 0 37260 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_398
timestamp 1586364061
transform 1 0 37720 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 39836 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_8  FILLER_36_411
timestamp 1586364061
transform 1 0 38916 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_419
timestamp 1586364061
transform 1 0 39652 0 -1 22304
box -38 -48 222 592
use scs8hd_nor2_4  _307_
timestamp 1586364061
transform 1 0 41400 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 42412 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_430
timestamp 1586364061
transform 1 0 40664 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_447
timestamp 1586364061
transform 1 0 42228 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_451
timestamp 1586364061
transform 1 0 42596 0 -1 22304
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_469
timestamp 1586364061
transform 1 0 43240 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_457
timestamp 1586364061
transform 1 0 43148 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_468
timestamp 1586364061
transform 1 0 44160 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_480
timestamp 1586364061
transform 1 0 45264 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_492
timestamp 1586364061
transform 1 0 46368 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_504
timestamp 1586364061
transform 1 0 47472 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 48852 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_470
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_471
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__333__A
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__333__B
timestamp 1586364061
transform 1 0 11408 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_114
timestamp 1586364061
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_118
timestamp 1586364061
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_134
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14996 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_144
timestamp 1586364061
transform 1 0 14352 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_148
timestamp 1586364061
transform 1 0 14720 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_160
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_164
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_172
timestamp 1586364061
transform 1 0 16928 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_180
timestamp 1586364061
transform 1 0 17664 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_176
timestamp 1586364061
transform 1 0 17296 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17480 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_472
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_37_188
timestamp 1586364061
transform 1 0 18400 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 1 22304
box -38 -48 866 592
use scs8hd_decap_3  FILLER_37_204
timestamp 1586364061
transform 1 0 19872 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_200
timestamp 1586364061
transform 1 0 19504 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19688 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_213
timestamp 1586364061
transform 1 0 20700 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_209
timestamp 1586364061
transform 1 0 20332 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__356__A
timestamp 1586364061
transform 1 0 22908 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__356__B
timestamp 1586364061
transform 1 0 23276 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_217
timestamp 1586364061
transform 1 0 21068 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_227
timestamp 1586364061
transform 1 0 21988 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_231
timestamp 1586364061
transform 1 0 22356 0 1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_37_239
timestamp 1586364061
transform 1 0 23092 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_248
timestamp 1586364061
transform 1 0 23920 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_243
timestamp 1586364061
transform 1 0 23460 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__216__A
timestamp 1586364061
transform 1 0 24104 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_473
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.lut4_mux_0_.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_252
timestamp 1586364061
transform 1 0 24288 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__216__B
timestamp 1586364061
transform 1 0 24472 0 1 22304
box -38 -48 222 592
use scs8hd_inv_8  _127_
timestamp 1586364061
transform 1 0 24656 0 1 22304
box -38 -48 866 592
use scs8hd_fill_2  FILLER_37_265
timestamp 1586364061
transform 1 0 25484 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 25668 0 1 22304
box -38 -48 222 592
use scs8hd_nor2_4  _311_
timestamp 1586364061
transform 1 0 27324 0 1 22304
box -38 -48 866 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 26220 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__311__A
timestamp 1586364061
transform 1 0 27140 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 26680 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_3_.scs8hd_buf_1_A
timestamp 1586364061
transform 1 0 26036 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_276
timestamp 1586364061
transform 1 0 26496 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_280
timestamp 1586364061
transform 1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_294
timestamp 1586364061
transform 1 0 28152 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_302
timestamp 1586364061
transform 1 0 28888 0 1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_37_298
timestamp 1586364061
transform 1 0 28520 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28980 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 28336 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_474
timestamp 1586364061
transform 1 0 29164 0 1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_37_310
timestamp 1586364061
transform 1 0 29624 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_306
timestamp 1586364061
transform 1 0 29256 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 29440 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29716 0 1 22304
box -38 -48 866 592
use scs8hd_decap_8  FILLER_37_320
timestamp 1586364061
transform 1 0 30544 0 1 22304
box -38 -48 774 592
use scs8hd_nor2_4  _309_
timestamp 1586364061
transform 1 0 31556 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 32568 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__309__A
timestamp 1586364061
transform 1 0 31372 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32936 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_328
timestamp 1586364061
transform 1 0 31280 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_340
timestamp 1586364061
transform 1 0 32384 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_344
timestamp 1586364061
transform 1 0 32752 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_348
timestamp 1586364061
transform 1 0 33120 0 1 22304
box -38 -48 406 592
use scs8hd_decap_4  FILLER_37_358
timestamp 1586364061
transform 1 0 34040 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_352
timestamp 1586364061
transform 1 0 33488 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33580 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33764 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_367
timestamp 1586364061
transform 1 0 34868 0 1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_37_365
timestamp 1586364061
transform 1 0 34684 0 1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_37_362
timestamp 1586364061
transform 1 0 34408 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 34500 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_475
timestamp 1586364061
transform 1 0 34776 0 1 22304
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35144 0 1 22304
box -38 -48 866 592
use scs8hd_nor2_4  _304_
timestamp 1586364061
transform 1 0 36892 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36248 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__304__A
timestamp 1586364061
transform 1 0 36708 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__257__A
timestamp 1586364061
transform 1 0 37904 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_379
timestamp 1586364061
transform 1 0 35972 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_384
timestamp 1586364061
transform 1 0 36432 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_398
timestamp 1586364061
transform 1 0 37720 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_402
timestamp 1586364061
transform 1 0 38088 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_409
timestamp 1586364061
transform 1 0 38732 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__257__B
timestamp 1586364061
transform 1 0 38272 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 38456 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_413
timestamp 1586364061
transform 1 0 39100 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38916 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__255__A
timestamp 1586364061
transform 1 0 39284 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_421
timestamp 1586364061
transform 1 0 39836 0 1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_37_417
timestamp 1586364061
transform 1 0 39468 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__255__B
timestamp 1586364061
transform 1 0 39652 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_476
timestamp 1586364061
transform 1 0 40388 0 1 22304
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_431
timestamp 1586364061
transform 1 0 40756 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 40940 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_439
timestamp 1586364061
transform 1 0 41492 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_435
timestamp 1586364061
transform 1 0 41124 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41308 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_443
timestamp 1586364061
transform 1 0 41860 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 41676 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_447
timestamp 1586364061
transform 1 0 42228 0 1 22304
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42320 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_451
timestamp 1586364061
transform 1 0 42596 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42780 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_455
timestamp 1586364061
transform 1 0 42964 0 1 22304
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43792 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_462
timestamp 1586364061
transform 1 0 43608 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_466
timestamp 1586364061
transform 1 0 43976 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_478
timestamp 1586364061
transform 1 0 45080 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_477
timestamp 1586364061
transform 1 0 46000 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_486
timestamp 1586364061
transform 1 0 45816 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_489
timestamp 1586364061
transform 1 0 46092 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_501
timestamp 1586364061
transform 1 0 47196 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 48852 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_513
timestamp 1586364061
transform 1 0 48300 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_478
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_479
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_nor2_4  _333_
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__346__B
timestamp 1586364061
transform 1 0 12880 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_126
timestamp 1586364061
transform 1 0 12696 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_130
timestamp 1586364061
transform 1 0 13064 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 23392
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_480
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16928 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_38_163
timestamp 1586364061
transform 1 0 16100 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_38_171
timestamp 1586364061
transform 1 0 16836 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_181
timestamp 1586364061
transform 1 0 17756 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18860 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_481
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_189
timestamp 1586364061
transform 1 0 18492 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_nor2_4  _356_
timestamp 1586364061
transform 1 0 22908 0 -1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_12  FILLER_38_224
timestamp 1586364061
transform 1 0 21712 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_236
timestamp 1586364061
transform 1 0 22816 0 -1 23392
box -38 -48 130 592
use scs8hd_nand2_4  _216_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 24472 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23920 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_246
timestamp 1586364061
transform 1 0 23736 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_250
timestamp 1586364061
transform 1 0 24104 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_buf_1  ltile_clb_0.ltile_clb_fle_0.ltile_clb_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_0_.buf4_2_.scs8hd_buf_1
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 27692 0 -1 23392
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_482
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__311__B
timestamp 1586364061
transform 1 0 27324 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26956 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_279
timestamp 1586364061
transform 1 0 26772 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_283
timestamp 1586364061
transform 1 0 27140 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_287
timestamp 1586364061
transform 1 0 27508 0 -1 23392
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 29440 0 -1 23392
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30636 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29256 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_300
timestamp 1586364061
transform 1 0 28704 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_38_319
timestamp 1586364061
transform 1 0 30452 0 -1 23392
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 23392
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_483
timestamp 1586364061
transform 1 0 32016 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_323
timestamp 1586364061
transform 1 0 30820 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_335
timestamp 1586364061
transform 1 0 31924 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_348
timestamp 1586364061
transform 1 0 33120 0 -1 23392
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 34500 0 -1 23392
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_38_360
timestamp 1586364061
transform 1 0 34224 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_38_374
timestamp 1586364061
transform 1 0 35512 0 -1 23392
box -38 -48 222 592
use scs8hd_nor2_4  _257_
timestamp 1586364061
transform 1 0 37720 0 -1 23392
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36248 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_484
timestamp 1586364061
transform 1 0 37628 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__258__B
timestamp 1586364061
transform 1 0 37076 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35696 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_378
timestamp 1586364061
transform 1 0 35880 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_6  FILLER_38_385
timestamp 1586364061
transform 1 0 36524 0 -1 23392
box -38 -48 590 592
use scs8hd_decap_4  FILLER_38_393
timestamp 1586364061
transform 1 0 37260 0 -1 23392
box -38 -48 406 592
use scs8hd_nor2_4  _255_
timestamp 1586364061
transform 1 0 39284 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38732 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39100 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_407
timestamp 1586364061
transform 1 0 38548 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_411
timestamp 1586364061
transform 1 0 38916 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_424
timestamp 1586364061
transform 1 0 40112 0 -1 23392
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_7_.latch
timestamp 1586364061
transform 1 0 40848 0 -1 23392
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42044 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42412 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_443
timestamp 1586364061
transform 1 0 41860 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_447
timestamp 1586364061
transform 1 0 42228 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_451
timestamp 1586364061
transform 1 0 42596 0 -1 23392
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_485
timestamp 1586364061
transform 1 0 43240 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_457
timestamp 1586364061
transform 1 0 43148 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_459
timestamp 1586364061
transform 1 0 43332 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_471
timestamp 1586364061
transform 1 0 44436 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_483
timestamp 1586364061
transform 1 0 45540 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_495
timestamp 1586364061
transform 1 0 46644 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_507
timestamp 1586364061
transform 1 0 47748 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 48852 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_515
timestamp 1586364061
transform 1 0 48484 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_494
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_486
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_495
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__345__A
timestamp 1586364061
transform 1 0 10396 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_39_106
timestamp 1586364061
transform 1 0 10856 0 1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_103
timestamp 1586364061
transform 1 0 10580 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_107
timestamp 1586364061
transform 1 0 10948 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_119
timestamp 1586364061
transform 1 0 12052 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_115
timestamp 1586364061
transform 1 0 11684 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_111
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 11132 0 1 23392
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 11132 0 -1 24480
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_40_125
timestamp 1586364061
transform 1 0 12604 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_40_120
timestamp 1586364061
transform 1 0 12144 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__334__B
timestamp 1586364061
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__334__A
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_487
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_nor2_4  _346_
timestamp 1586364061
transform 1 0 12880 0 -1 24480
box -38 -48 866 592
use scs8hd_nor2_4  _334_
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_39_132
timestamp 1586364061
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__346__A
timestamp 1586364061
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_143
timestamp 1586364061
transform 1 0 14260 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_6  FILLER_40_137
timestamp 1586364061
transform 1 0 13708 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_143
timestamp 1586364061
transform 1 0 14260 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_136
timestamp 1586364061
transform 1 0 13616 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__348__A
timestamp 1586364061
transform 1 0 14352 0 -1 24480
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_152
timestamp 1586364061
transform 1 0 15088 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_6  FILLER_40_146
timestamp 1586364061
transform 1 0 14536 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_496
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14996 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_161
timestamp 1586364061
transform 1 0 15916 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_160
timestamp 1586364061
transform 1 0 15824 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 24480
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15640 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_172
timestamp 1586364061
transform 1 0 16928 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_40_165
timestamp 1586364061
transform 1 0 16284 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_171
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_164
timestamp 1586364061
transform 1 0 16192 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16008 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16652 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_40_180
timestamp 1586364061
transform 1 0 17664 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_179
timestamp 1586364061
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_175
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_488
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 17940 0 -1 24480
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 18216 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_194
timestamp 1586364061
transform 1 0 18952 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_188
timestamp 1586364061
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19136 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_205
timestamp 1586364061
transform 1 0 19964 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_198
timestamp 1586364061
transform 1 0 19320 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_205
timestamp 1586364061
transform 1 0 19964 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_201
timestamp 1586364061
transform 1 0 19596 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20148 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_213
timestamp 1586364061
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_209
timestamp 1586364061
transform 1 0 20332 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_212
timestamp 1586364061
transform 1 0 20608 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_209
timestamp 1586364061
transform 1 0 20332 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__328__A
timestamp 1586364061
transform 1 0 20424 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 20792 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_497
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_40_224
timestamp 1586364061
transform 1 0 21712 0 -1 24480
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch
timestamp 1586364061
transform 1 0 20976 0 1 23392
box -38 -48 1050 592
use scs8hd_nor2_4  _328_
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__328__B
timestamp 1586364061
transform 1 0 22172 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__355__B
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_227
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_231
timestamp 1586364061
transform 1 0 22356 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_229
timestamp 1586364061
transform 1 0 22172 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22540 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_235
timestamp 1586364061
transform 1 0 22724 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_235
timestamp 1586364061
transform 1 0 22724 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_239
timestamp 1586364061
transform 1 0 23092 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23184 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_242
timestamp 1586364061
transform 1 0 23368 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_254
timestamp 1586364061
transform 1 0 24472 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__354__B
timestamp 1586364061
transform 1 0 23644 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__354__A
timestamp 1586364061
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_489
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 23828 0 -1 24480
box -38 -48 1050 592
use scs8hd_nor2_4  _354_
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 866 592
use scs8hd_fill_1  FILLER_40_266
timestamp 1586364061
transform 1 0 25576 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_262
timestamp 1586364061
transform 1 0 25208 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_258
timestamp 1586364061
transform 1 0 24840 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_258
timestamp 1586364061
transform 1 0 24840 0 1 23392
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25668 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 24656 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_269
timestamp 1586364061
transform 1 0 25852 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_277
timestamp 1586364061
transform 1 0 26588 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_274
timestamp 1586364061
transform 1 0 26312 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_270
timestamp 1586364061
transform 1 0 25944 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_498
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_288
timestamp 1586364061
transform 1 0 27600 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_285
timestamp 1586364061
transform 1 0 27324 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_6  FILLER_40_279
timestamp 1586364061
transform 1 0 26772 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_281
timestamp 1586364061
transform 1 0 26956 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__310__B
timestamp 1586364061
transform 1 0 26772 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__310__A
timestamp 1586364061
transform 1 0 27140 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__313__A
timestamp 1586364061
transform 1 0 27416 0 -1 24480
box -38 -48 222 592
use scs8hd_nor2_4  _310_
timestamp 1586364061
transform 1 0 27324 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_292
timestamp 1586364061
transform 1 0 27968 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_294
timestamp 1586364061
transform 1 0 28152 0 1 23392
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28152 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__313__B
timestamp 1586364061
transform 1 0 27784 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_296
timestamp 1586364061
transform 1 0 28336 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_3  FILLER_39_302
timestamp 1586364061
transform 1 0 28888 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__312__A
timestamp 1586364061
transform 1 0 28704 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_490
timestamp 1586364061
transform 1 0 29164 0 1 23392
box -38 -48 130 592
use scs8hd_nor2_4  _312_
timestamp 1586364061
transform 1 0 28704 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_313
timestamp 1586364061
transform 1 0 29900 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_309
timestamp 1586364061
transform 1 0 29532 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_310
timestamp 1586364061
transform 1 0 29624 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_306
timestamp 1586364061
transform 1 0 29256 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29716 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__312__B
timestamp 1586364061
transform 1 0 29440 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29716 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_39_320
timestamp 1586364061
transform 1 0 30544 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30084 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30728 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30268 0 -1 24480
box -38 -48 866 592
use scs8hd_decap_6  FILLER_40_326
timestamp 1586364061
transform 1 0 31096 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_331
timestamp 1586364061
transform 1 0 31556 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_328
timestamp 1586364061
transform 1 0 31280 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_324
timestamp 1586364061
transform 1 0 30912 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31372 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_340
timestamp 1586364061
transform 1 0 32384 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_334
timestamp 1586364061
transform 1 0 31832 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_335
timestamp 1586364061
transform 1 0 31924 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31648 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31740 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32108 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_499
timestamp 1586364061
transform 1 0 32016 0 -1 24480
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32292 0 1 23392
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32108 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_344
timestamp 1586364061
transform 1 0 32752 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_39_348
timestamp 1586364061
transform 1 0 33120 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32568 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_352
timestamp 1586364061
transform 1 0 33488 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_355
timestamp 1586364061
transform 1 0 33764 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_352
timestamp 1586364061
transform 1 0 33488 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__316__B
timestamp 1586364061
transform 1 0 33948 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__316__A
timestamp 1586364061
transform 1 0 33580 0 1 23392
box -38 -48 222 592
use scs8hd_nor2_4  _316_
timestamp 1586364061
transform 1 0 33580 0 -1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_40_366
timestamp 1586364061
transform 1 0 34776 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_362
timestamp 1586364061
transform 1 0 34408 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_367
timestamp 1586364061
transform 1 0 34868 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_39_363
timestamp 1586364061
transform 1 0 34500 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_359
timestamp 1586364061
transform 1 0 34132 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34592 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34960 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_491
timestamp 1586364061
transform 1 0 34776 0 1 23392
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35144 0 -1 24480
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35144 0 1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_40_386
timestamp 1586364061
transform 1 0 36616 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_383
timestamp 1586364061
transform 1 0 36340 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_379
timestamp 1586364061
transform 1 0 35972 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_387
timestamp 1586364061
transform 1 0 36708 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_383
timestamp 1586364061
transform 1 0 36340 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_379
timestamp 1586364061
transform 1 0 35972 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36524 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36156 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36432 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_398
timestamp 1586364061
transform 1 0 37720 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_40_394
timestamp 1586364061
transform 1 0 37352 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__258__A
timestamp 1586364061
transform 1 0 36892 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_500
timestamp 1586364061
transform 1 0 37628 0 -1 24480
box -38 -48 130 592
use scs8hd_nor2_4  _258_
timestamp 1586364061
transform 1 0 37076 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_39_400
timestamp 1586364061
transform 1 0 37904 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 38088 0 1 23392
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 37904 0 -1 24480
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_40_411
timestamp 1586364061
transform 1 0 38916 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_39_404
timestamp 1586364061
transform 1 0 38272 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38456 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38640 0 1 23392
box -38 -48 866 592
use scs8hd_fill_1  FILLER_40_427
timestamp 1586364061
transform 1 0 40388 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_423
timestamp 1586364061
transform 1 0 40020 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_3  FILLER_39_428
timestamp 1586364061
transform 1 0 40480 0 1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_39_417
timestamp 1586364061
transform 1 0 39468 0 1 23392
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40204 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_492
timestamp 1586364061
transform 1 0 40388 0 1 23392
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 40480 0 -1 24480
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_40_439
timestamp 1586364061
transform 1 0 41492 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_438
timestamp 1586364061
transform 1 0 41400 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_434
timestamp 1586364061
transform 1 0 41032 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 41216 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40756 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_40_443
timestamp 1586364061
transform 1 0 41860 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42044 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41676 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41584 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41768 0 1 23392
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42228 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_40_450
timestamp 1586364061
transform 1 0 42504 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_4  FILLER_39_455
timestamp 1586364061
transform 1 0 42964 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_451
timestamp 1586364061
transform 1 0 42596 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42780 0 1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_501
timestamp 1586364061
transform 1 0 43240 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43332 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43700 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_461
timestamp 1586364061
transform 1 0 43516 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_465
timestamp 1586364061
transform 1 0 43884 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_477
timestamp 1586364061
transform 1 0 44988 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_468
timestamp 1586364061
transform 1 0 44160 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_480
timestamp 1586364061
transform 1 0 45264 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_493
timestamp 1586364061
transform 1 0 46000 0 1 23392
box -38 -48 130 592
use scs8hd_decap_3  FILLER_39_485
timestamp 1586364061
transform 1 0 45724 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_489
timestamp 1586364061
transform 1 0 46092 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_501
timestamp 1586364061
transform 1 0 47196 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_492
timestamp 1586364061
transform 1 0 46368 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_504
timestamp 1586364061
transform 1 0 47472 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 48852 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 48852 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_513
timestamp 1586364061
transform 1 0 48300 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_502
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_nor2_4  _345_
timestamp 1586364061
transform 1 0 10396 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__345__B
timestamp 1586364061
transform 1 0 9844 0 1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_41_94
timestamp 1586364061
transform 1 0 9752 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_97
timestamp 1586364061
transform 1 0 10028 0 1 24480
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 12604 0 1 24480
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_503
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_114
timestamp 1586364061
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_140
timestamp 1586364061
transform 1 0 13984 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_136
timestamp 1586364061
transform 1 0 13616 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__348__B
timestamp 1586364061
transform 1 0 13800 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 24480
box -38 -48 222 592
use scs8hd_nor2_4  _348_
timestamp 1586364061
transform 1 0 14352 0 1 24480
box -38 -48 866 592
use scs8hd_fill_2  FILLER_41_153
timestamp 1586364061
transform 1 0 15180 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_157
timestamp 1586364061
transform 1 0 15548 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 24480
box -38 -48 866 592
use scs8hd_nor2_4  _331_
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_504
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__331__A
timestamp 1586364061
transform 1 0 17388 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17020 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_170
timestamp 1586364061
transform 1 0 16744 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_175
timestamp 1586364061
transform 1 0 17204 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_179
timestamp 1586364061
transform 1 0 17572 0 1 24480
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 20148 0 1 24480
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19964 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__331__B
timestamp 1586364061
transform 1 0 19044 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_193
timestamp 1586364061
transform 1 0 18860 0 1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_197
timestamp 1586364061
transform 1 0 19228 0 1 24480
box -38 -48 774 592
use scs8hd_nor2_4  _355_
timestamp 1586364061
transform 1 0 21988 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__355__A
timestamp 1586364061
transform 1 0 21804 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_218
timestamp 1586364061
transform 1 0 21160 0 1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_41_224
timestamp 1586364061
transform 1 0 21712 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_236
timestamp 1586364061
transform 1 0 22816 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_240
timestamp 1586364061
transform 1 0 23184 0 1 24480
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 23920 0 1 24480
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 25668 0 1 24480
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_505
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 25484 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25116 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_259
timestamp 1586364061
transform 1 0 24932 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_263
timestamp 1586364061
transform 1 0 25300 0 1 24480
box -38 -48 222 592
use scs8hd_nor2_4  _313_
timestamp 1586364061
transform 1 0 27416 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26956 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_278
timestamp 1586364061
transform 1 0 26680 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_41_283
timestamp 1586364061
transform 1 0 27140 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_295
timestamp 1586364061
transform 1 0 28244 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_506
timestamp 1586364061
transform 1 0 29164 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 28428 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30268 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_299
timestamp 1586364061
transform 1 0 28612 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_315
timestamp 1586364061
transform 1 0 30084 0 1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_319
timestamp 1586364061
transform 1 0 30452 0 1 24480
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31648 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33028 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31464 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32660 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_327
timestamp 1586364061
transform 1 0 31188 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_341
timestamp 1586364061
transform 1 0 32476 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_345
timestamp 1586364061
transform 1 0 32844 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33212 0 1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_507
timestamp 1586364061
transform 1 0 34776 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33948 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_352
timestamp 1586364061
transform 1 0 33488 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_356
timestamp 1586364061
transform 1 0 33856 0 1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_41_359
timestamp 1586364061
transform 1 0 34132 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_363
timestamp 1586364061
transform 1 0 34500 0 1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_41_387
timestamp 1586364061
transform 1 0 36708 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_380
timestamp 1586364061
transform 1 0 36064 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_376
timestamp 1586364061
transform 1 0 35696 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35880 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36248 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36432 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_394
timestamp 1586364061
transform 1 0 37352 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_391
timestamp 1586364061
transform 1 0 37076 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37168 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 37536 0 1 24480
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 37720 0 1 24480
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_508
timestamp 1586364061
transform 1 0 40388 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38916 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39284 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_409
timestamp 1586364061
transform 1 0 38732 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_413
timestamp 1586364061
transform 1 0 39100 0 1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_417
timestamp 1586364061
transform 1 0 39468 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_425
timestamp 1586364061
transform 1 0 40204 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_428
timestamp 1586364061
transform 1 0 40480 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_439
timestamp 1586364061
transform 1 0 41492 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_435
timestamp 1586364061
transform 1 0 41124 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40664 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41308 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40848 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41676 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41860 0 1 24480
box -38 -48 866 592
use scs8hd_decap_4  FILLER_41_456
timestamp 1586364061
transform 1 0 43056 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_452
timestamp 1586364061
transform 1 0 42688 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42872 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43700 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44160 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44528 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43516 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_460
timestamp 1586364061
transform 1 0 43424 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_466
timestamp 1586364061
transform 1 0 43976 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_470
timestamp 1586364061
transform 1 0 44344 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_474
timestamp 1586364061
transform 1 0 44712 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_509
timestamp 1586364061
transform 1 0 46000 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_486
timestamp 1586364061
transform 1 0 45816 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_489
timestamp 1586364061
transform 1 0 46092 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_501
timestamp 1586364061
transform 1 0 47196 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 48852 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_41_513
timestamp 1586364061
transform 1 0 48300 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_510
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_68
timestamp 1586364061
transform 1 0 7360 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_80
timestamp 1586364061
transform 1 0 8464 0 -1 25568
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10396 0 -1 25568
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_511
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__351__B
timestamp 1586364061
transform 1 0 10028 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_93
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_42_99
timestamp 1586364061
transform 1 0 10212 0 -1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12236 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_112
timestamp 1586364061
transform 1 0 11408 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_42_120
timestamp 1586364061
transform 1 0 12144 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_132
timestamp 1586364061
transform 1 0 13248 0 -1 25568
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 25568
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_512
timestamp 1586364061
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_136
timestamp 1586364061
transform 1 0 13616 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_2  FILLER_42_145
timestamp 1586364061
transform 1 0 14444 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 17940 0 -1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16836 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_165
timestamp 1586364061
transform 1 0 16284 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_169
timestamp 1586364061
transform 1 0 16652 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_173
timestamp 1586364061
transform 1 0 17020 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  FILLER_42_194
timestamp 1586364061
transform 1 0 18952 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__344__C
timestamp 1586364061
transform 1 0 19228 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_203
timestamp 1586364061
transform 1 0 19780 0 -1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__344__D
timestamp 1586364061
transform 1 0 19596 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__329__A
timestamp 1586364061
transform 1 0 20056 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_208
timestamp 1586364061
transform 1 0 20240 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__329__B
timestamp 1586364061
transform 1 0 20424 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_212
timestamp 1586364061
transform 1 0 20608 0 -1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_513
timestamp 1586364061
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23184 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__357__B
timestamp 1586364061
transform 1 0 21620 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22080 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_215
timestamp 1586364061
transform 1 0 20884 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  FILLER_42_225
timestamp 1586364061
transform 1 0 21804 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_238
timestamp 1586364061
transform 1 0 23000 0 -1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24196 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_253
timestamp 1586364061
transform 1 0 24380 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_42_267
timestamp 1586364061
transform 1 0 25668 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_280
timestamp 1586364061
transform 1 0 26864 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_276
timestamp 1586364061
transform 1 0 26496 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_271
timestamp 1586364061
transform 1 0 26036 0 -1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25852 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26680 0 -1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_514
timestamp 1586364061
transform 1 0 26404 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_288
timestamp 1586364061
transform 1 0 27600 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_42_284
timestamp 1586364061
transform 1 0 27232 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__308__D
timestamp 1586364061
transform 1 0 27416 0 -1 25568
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26956 0 -1 25568
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 27968 0 -1 25568
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29716 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29256 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_303
timestamp 1586364061
transform 1 0 28980 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_42_308
timestamp 1586364061
transform 1 0 29440 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_320
timestamp 1586364061
transform 1 0 30544 0 -1 25568
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_515
timestamp 1586364061
transform 1 0 32016 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31004 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31832 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_324
timestamp 1586364061
transform 1 0 30912 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_327
timestamp 1586364061
transform 1 0 31188 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_1  FILLER_42_333
timestamp 1586364061
transform 1 0 31740 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_346
timestamp 1586364061
transform 1 0 32936 0 -1 25568
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33948 0 -1 25568
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34960 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34776 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34408 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_42_354
timestamp 1586364061
transform 1 0 33672 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_42_360
timestamp 1586364061
transform 1 0 34224 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_364
timestamp 1586364061
transform 1 0 34592 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_42_377
timestamp 1586364061
transform 1 0 35788 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_392
timestamp 1586364061
transform 1 0 37168 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_388
timestamp 1586364061
transform 1 0 36800 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36984 0 -1 25568
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36524 0 -1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_42_401
timestamp 1586364061
transform 1 0 37996 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_396
timestamp 1586364061
transform 1 0 37536 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37352 0 -1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_516
timestamp 1586364061
transform 1 0 37628 0 -1 25568
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37720 0 -1 25568
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 -1 25568
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38732 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38180 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_405
timestamp 1586364061
transform 1 0 38364 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_8  FILLER_42_418
timestamp 1586364061
transform 1 0 39560 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_426
timestamp 1586364061
transform 1 0 40296 0 -1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41492 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41308 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_431
timestamp 1586364061
transform 1 0 40756 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_8  FILLER_42_448
timestamp 1586364061
transform 1 0 42320 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_456
timestamp 1586364061
transform 1 0 43056 0 -1 25568
box -38 -48 222 592
use scs8hd_conb_1  _443_
timestamp 1586364061
transform 1 0 45356 0 -1 25568
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43792 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_517
timestamp 1586364061
transform 1 0 43240 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_459
timestamp 1586364061
transform 1 0 43332 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_42_463
timestamp 1586364061
transform 1 0 43700 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_473
timestamp 1586364061
transform 1 0 44620 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_12  FILLER_42_484
timestamp 1586364061
transform 1 0 45632 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_496
timestamp 1586364061
transform 1 0 46736 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_42_508
timestamp 1586364061
transform 1 0 47840 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 48852 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_43_3
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_15
timestamp 1586364061
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_27
timestamp 1586364061
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_39
timestamp 1586364061
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_51
timestamp 1586364061
transform 1 0 5796 0 1 25568
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_518
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_59
timestamp 1586364061
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_43_62
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_74
timestamp 1586364061
transform 1 0 7912 0 1 25568
box -38 -48 1142 592
use scs8hd_nor2_4  _351_
timestamp 1586364061
transform 1 0 10028 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__351__A
timestamp 1586364061
transform 1 0 9844 0 1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_43_86
timestamp 1586364061
transform 1 0 9016 0 1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_43_94
timestamp 1586364061
transform 1 0 9752 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_106
timestamp 1586364061
transform 1 0 10856 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_115
timestamp 1586364061
transform 1 0 11684 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_110
timestamp 1586364061
transform 1 0 11224 0 1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11040 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_127
timestamp 1586364061
transform 1 0 12788 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_123
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_119
timestamp 1586364061
transform 1 0 12052 0 1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_519
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 1 25568
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14720 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14536 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_140
timestamp 1586364061
transform 1 0 13984 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_144
timestamp 1586364061
transform 1 0 14352 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_157
timestamp 1586364061
transform 1 0 15548 0 1 25568
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_520
timestamp 1586364061
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__347__A
timestamp 1586364061
transform 1 0 17480 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__347__B
timestamp 1586364061
transform 1 0 18216 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_162
timestamp 1586364061
transform 1 0 16008 0 1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_43_174
timestamp 1586364061
transform 1 0 17112 0 1 25568
box -38 -48 406 592
use scs8hd_decap_3  FILLER_43_180
timestamp 1586364061
transform 1 0 17664 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_184
timestamp 1586364061
transform 1 0 18032 0 1 25568
box -38 -48 222 592
use scs8hd_nor2_4  _329_
timestamp 1586364061
transform 1 0 20056 0 1 25568
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__344__A
timestamp 1586364061
transform 1 0 19504 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__344__B
timestamp 1586364061
transform 1 0 19872 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_188
timestamp 1586364061
transform 1 0 18400 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_198
timestamp 1586364061
transform 1 0 19320 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_202
timestamp 1586364061
transform 1 0 19688 0 1 25568
box -38 -48 222 592
use scs8hd_nor2_4  _357_
timestamp 1586364061
transform 1 0 21620 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 22632 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__357__A
timestamp 1586364061
transform 1 0 21436 0 1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_43_215
timestamp 1586364061
transform 1 0 20884 0 1 25568
box -38 -48 590 592
use scs8hd_fill_2  FILLER_43_232
timestamp 1586364061
transform 1 0 22448 0 1 25568
box -38 -48 222 592
use scs8hd_decap_8  FILLER_43_236
timestamp 1586364061
transform 1 0 22816 0 1 25568
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25024 0 1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_521
timestamp 1586364061
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24472 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_245
timestamp 1586364061
transform 1 0 23644 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_249
timestamp 1586364061
transform 1 0 24012 0 1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_43_253
timestamp 1586364061
transform 1 0 24380 0 1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_43_256
timestamp 1586364061
transform 1 0 24656 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_273
timestamp 1586364061
transform 1 0 26220 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_269
timestamp 1586364061
transform 1 0 25852 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26036 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__308__C
timestamp 1586364061
transform 1 0 26404 0 1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26588 0 1 25568
box -38 -48 866 592
use scs8hd_fill_2  FILLER_43_286
timestamp 1586364061
transform 1 0 27416 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__308__A
timestamp 1586364061
transform 1 0 27600 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_290
timestamp 1586364061
transform 1 0 27784 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__308__B
timestamp 1586364061
transform 1 0 27968 0 1 25568
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28152 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_301
timestamp 1586364061
transform 1 0 28796 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_297
timestamp 1586364061
transform 1 0 28428 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28612 0 1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_522
timestamp 1586364061
transform 1 0 29164 0 1 25568
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_43_317
timestamp 1586364061
transform 1 0 30268 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_313
timestamp 1586364061
transform 1 0 29900 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_309
timestamp 1586364061
transform 1 0 29532 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30084 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29716 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 30544 0 1 25568
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 30728 0 1 25568
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32476 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32292 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31924 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_333
timestamp 1586364061
transform 1 0 31740 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_337
timestamp 1586364061
transform 1 0 32108 0 1 25568
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 34868 0 1 25568
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_523
timestamp 1586364061
transform 1 0 34776 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33948 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 34592 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33488 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_350
timestamp 1586364061
transform 1 0 33304 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_354
timestamp 1586364061
transform 1 0 33672 0 1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_43_359
timestamp 1586364061
transform 1 0 34132 0 1 25568
box -38 -48 406 592
use scs8hd_fill_1  FILLER_43_363
timestamp 1586364061
transform 1 0 34500 0 1 25568
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36616 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 37996 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36432 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36064 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37628 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_378
timestamp 1586364061
transform 1 0 35880 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_382
timestamp 1586364061
transform 1 0 36248 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_395
timestamp 1586364061
transform 1 0 37444 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_399
timestamp 1586364061
transform 1 0 37812 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_407
timestamp 1586364061
transform 1 0 38548 0 1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_43_403
timestamp 1586364061
transform 1 0 38180 0 1 25568
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38640 0 1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38824 0 1 25568
box -38 -48 866 592
use scs8hd_fill_2  FILLER_43_419
timestamp 1586364061
transform 1 0 39652 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__261__A
timestamp 1586364061
transform 1 0 39836 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_428
timestamp 1586364061
transform 1 0 40480 0 1 25568
box -38 -48 314 592
use scs8hd_fill_2  FILLER_43_423
timestamp 1586364061
transform 1 0 40020 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__261__B
timestamp 1586364061
transform 1 0 40204 0 1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_524
timestamp 1586364061
transform 1 0 40388 0 1 25568
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42872 0 1 25568
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41308 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41124 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42320 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40756 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_433
timestamp 1586364061
transform 1 0 40940 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_446
timestamp 1586364061
transform 1 0 42136 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_450
timestamp 1586364061
transform 1 0 42504 0 1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_43_461
timestamp 1586364061
transform 1 0 43516 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_457
timestamp 1586364061
transform 1 0 43148 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43700 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43332 0 1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43884 0 1 25568
box -38 -48 866 592
use scs8hd_fill_2  FILLER_43_474
timestamp 1586364061
transform 1 0 44712 0 1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_43_482
timestamp 1586364061
transform 1 0 45448 0 1 25568
box -38 -48 590 592
use scs8hd_fill_2  FILLER_43_478
timestamp 1586364061
transform 1 0 45080 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45264 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44896 0 1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_525
timestamp 1586364061
transform 1 0 46000 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_489
timestamp 1586364061
transform 1 0 46092 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_501
timestamp 1586364061
transform 1 0 47196 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 48852 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_43_513
timestamp 1586364061
transform 1 0 48300 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_15
timestamp 1586364061
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_526
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_4  FILLER_44_27
timestamp 1586364061
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_12  FILLER_44_32
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_44
timestamp 1586364061
transform 1 0 5152 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_56
timestamp 1586364061
transform 1 0 6256 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_68
timestamp 1586364061
transform 1 0 7360 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_80
timestamp 1586364061
transform 1 0 8464 0 -1 26656
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10488 0 -1 26656
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_527
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__350__A
timestamp 1586364061
transform 1 0 10028 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_93
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_3  FILLER_44_99
timestamp 1586364061
transform 1 0 10212 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_8  FILLER_44_105
timestamp 1586364061
transform 1 0 10764 0 -1 26656
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13064 0 -1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 26656
box -38 -48 866 592
use scs8hd_decap_8  FILLER_44_122
timestamp 1586364061
transform 1 0 12328 0 -1 26656
box -38 -48 774 592
use scs8hd_decap_8  FILLER_44_133
timestamp 1586364061
transform 1 0 13340 0 -1 26656
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14076 0 -1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_528
timestamp 1586364061
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15456 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_44_144
timestamp 1586364061
transform 1 0 14352 0 -1 26656
box -38 -48 590 592
use scs8hd_fill_1  FILLER_44_152
timestamp 1586364061
transform 1 0 15088 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_44_154
timestamp 1586364061
transform 1 0 15272 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_158
timestamp 1586364061
transform 1 0 15640 0 -1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _347_
timestamp 1586364061
transform 1 0 17480 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_169
timestamp 1586364061
transform 1 0 16652 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_3  FILLER_44_175
timestamp 1586364061
transform 1 0 17204 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_3  FILLER_44_187
timestamp 1586364061
transform 1 0 18308 0 -1 26656
box -38 -48 314 592
use scs8hd_or4_4  _344_
timestamp 1586364061
transform 1 0 19228 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_529
timestamp 1586364061
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__326__D
timestamp 1586364061
transform 1 0 20240 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18584 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18952 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_192
timestamp 1586364061
transform 1 0 18768 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_44_196
timestamp 1586364061
transform 1 0 19136 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_44_206
timestamp 1586364061
transform 1 0 20056 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_210
timestamp 1586364061
transform 1 0 20424 0 -1 26656
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 22080 0 -1 26656
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__360__B
timestamp 1586364061
transform 1 0 21068 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21804 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_215
timestamp 1586364061
transform 1 0 20884 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_44_219
timestamp 1586364061
transform 1 0 21252 0 -1 26656
box -38 -48 590 592
use scs8hd_fill_1  FILLER_44_227
timestamp 1586364061
transform 1 0 21988 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_8  FILLER_44_239
timestamp 1586364061
transform 1 0 23092 0 -1 26656
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23828 0 -1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_44_250
timestamp 1586364061
transform 1 0 24104 0 -1 26656
box -38 -48 590 592
use scs8hd_decap_8  FILLER_44_267
timestamp 1586364061
transform 1 0 25668 0 -1 26656
box -38 -48 774 592
use scs8hd_or4_4  _308_
timestamp 1586364061
transform 1 0 27232 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_530
timestamp 1586364061
transform 1 0 26404 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__254__C
timestamp 1586364061
transform 1 0 27048 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26680 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28244 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_276
timestamp 1586364061
transform 1 0 26496 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_280
timestamp 1586364061
transform 1 0 26864 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_293
timestamp 1586364061
transform 1 0 28060 0 -1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29164 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30728 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_44_297
timestamp 1586364061
transform 1 0 28428 0 -1 26656
box -38 -48 774 592
use scs8hd_decap_8  FILLER_44_314
timestamp 1586364061
transform 1 0 29992 0 -1 26656
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31004 0 -1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32108 0 -1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_531
timestamp 1586364061
transform 1 0 32016 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_1  FILLER_44_324
timestamp 1586364061
transform 1 0 30912 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_8  FILLER_44_328
timestamp 1586364061
transform 1 0 31280 0 -1 26656
box -38 -48 774 592
use scs8hd_decap_3  FILLER_44_346
timestamp 1586364061
transform 1 0 32936 0 -1 26656
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33948 0 -1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34960 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__314__B
timestamp 1586364061
transform 1 0 33212 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_1_in_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 34776 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_44_351
timestamp 1586364061
transform 1 0 33396 0 -1 26656
box -38 -48 590 592
use scs8hd_decap_6  FILLER_44_360
timestamp 1586364061
transform 1 0 34224 0 -1 26656
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_6_.latch
timestamp 1586364061
transform 1 0 37996 0 -1 26656
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36524 0 -1 26656
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_532
timestamp 1586364061
transform 1 0 37628 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__256__B
timestamp 1586364061
transform 1 0 36984 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37444 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_44_377
timestamp 1586364061
transform 1 0 35788 0 -1 26656
box -38 -48 774 592
use scs8hd_fill_2  FILLER_44_388
timestamp 1586364061
transform 1 0 36800 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_44_392
timestamp 1586364061
transform 1 0 37168 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_3  FILLER_44_398
timestamp 1586364061
transform 1 0 37720 0 -1 26656
box -38 -48 314 592
use scs8hd_nor2_4  _261_
timestamp 1586364061
transform 1 0 39744 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39192 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_412
timestamp 1586364061
transform 1 0 39008 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_416
timestamp 1586364061
transform 1 0 39376 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_6  FILLER_44_429
timestamp 1586364061
transform 1 0 40572 0 -1 26656
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 41124 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43056 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_437
timestamp 1586364061
transform 1 0 41308 0 -1 26656
box -38 -48 406 592
use scs8hd_decap_6  FILLER_44_450
timestamp 1586364061
transform 1 0 42504 0 -1 26656
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44344 0 -1 26656
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 26656
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_533
timestamp 1586364061
transform 1 0 43240 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43884 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_44_462
timestamp 1586364061
transform 1 0 43608 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_3  FILLER_44_467
timestamp 1586364061
transform 1 0 44068 0 -1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_44_473
timestamp 1586364061
transform 1 0 44620 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_485
timestamp 1586364061
transform 1 0 45724 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_497
timestamp 1586364061
transform 1 0 46828 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_44_509
timestamp 1586364061
transform 1 0 47932 0 -1 26656
box -38 -48 590 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 48852 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_1  FILLER_44_515
timestamp 1586364061
transform 1 0 48484 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_decap_12  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_15
timestamp 1586364061
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_27
timestamp 1586364061
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_39
timestamp 1586364061
transform 1 0 4692 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_45_51
timestamp 1586364061
transform 1 0 5796 0 1 26656
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_534
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_45_59
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_62
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_74
timestamp 1586364061
transform 1 0 7912 0 1 26656
box -38 -48 1142 592
use scs8hd_nor2_4  _350_
timestamp 1586364061
transform 1 0 10028 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9844 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__350__B
timestamp 1586364061
transform 1 0 9476 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_86
timestamp 1586364061
transform 1 0 9016 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_90
timestamp 1586364061
transform 1 0 9384 0 1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_45_93
timestamp 1586364061
transform 1 0 9660 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_106
timestamp 1586364061
transform 1 0 10856 0 1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_535
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11040 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11408 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_110
timestamp 1586364061
transform 1 0 11224 0 1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_45_114
timestamp 1586364061
transform 1 0 11592 0 1 26656
box -38 -48 590 592
use scs8hd_fill_2  FILLER_45_132
timestamp 1586364061
transform 1 0 13248 0 1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14904 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_136
timestamp 1586364061
transform 1 0 13616 0 1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_45_140
timestamp 1586364061
transform 1 0 13984 0 1 26656
box -38 -48 774 592
use scs8hd_fill_2  FILLER_45_159
timestamp 1586364061
transform 1 0 15732 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_170
timestamp 1586364061
transform 1 0 16744 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_163
timestamp 1586364061
transform 1 0 16100 0 1 26656
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16468 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  FILLER_45_178
timestamp 1586364061
transform 1 0 17480 0 1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_45_174
timestamp 1586364061
transform 1 0 17112 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17296 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16928 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__349__A
timestamp 1586364061
transform 1 0 17756 0 1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_536
timestamp 1586364061
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use scs8hd_nor2_4  _349_
timestamp 1586364061
transform 1 0 18032 0 1 26656
box -38 -48 866 592
use scs8hd_or4_4  _326_
timestamp 1586364061
transform 1 0 19872 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__326__A
timestamp 1586364061
transform 1 0 19688 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__326__C
timestamp 1586364061
transform 1 0 19320 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_193
timestamp 1586364061
transform 1 0 18860 0 1 26656
box -38 -48 406 592
use scs8hd_fill_1  FILLER_45_197
timestamp 1586364061
transform 1 0 19228 0 1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_45_200
timestamp 1586364061
transform 1 0 19504 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_213
timestamp 1586364061
transform 1 0 20700 0 1 26656
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21804 0 1 26656
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__360__A
timestamp 1586364061
transform 1 0 21068 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_219
timestamp 1586364061
transform 1 0 21252 0 1 26656
box -38 -48 406 592
use scs8hd_fill_2  FILLER_45_236
timestamp 1586364061
transform 1 0 22816 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_240
timestamp 1586364061
transform 1 0 23184 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_251
timestamp 1586364061
transform 1 0 24196 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_45_245
timestamp 1586364061
transform 1 0 23644 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_537
timestamp 1586364061
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23920 0 1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_45_255
timestamp 1586364061
transform 1 0 24564 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24748 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24380 0 1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24932 0 1 26656
box -38 -48 866 592
use scs8hd_fill_2  FILLER_45_268
timestamp 1586364061
transform 1 0 25760 0 1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 1 26656
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28060 0 1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__254__A
timestamp 1586364061
transform 1 0 27508 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__254__B
timestamp 1586364061
transform 1 0 27876 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__254__D
timestamp 1586364061
transform 1 0 26312 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25944 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_272
timestamp 1586364061
transform 1 0 26128 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_285
timestamp 1586364061
transform 1 0 27324 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_289
timestamp 1586364061
transform 1 0 27692 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_303
timestamp 1586364061
transform 1 0 28980 0 1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_45_300
timestamp 1586364061
transform 1 0 28704 0 1 26656
box -38 -48 130 592
use scs8hd_decap_4  FILLER_45_296
timestamp 1586364061
transform 1 0 28336 0 1 26656
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__339__A
timestamp 1586364061
transform 1 0 28796 0 1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_538
timestamp 1586364061
transform 1 0 29164 0 1 26656
box -38 -48 130 592
use scs8hd_decap_3  FILLER_45_310
timestamp 1586364061
transform 1 0 29624 0 1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_45_306
timestamp 1586364061
transform 1 0 29256 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__339__B
timestamp 1586364061
transform 1 0 29440 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__315__A
timestamp 1586364061
transform 1 0 29900 0 1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _315_
timestamp 1586364061
transform 1 0 30084 0 1 26656
box -38 -48 866 592
use scs8hd_fill_2  FILLER_45_324
timestamp 1586364061
transform 1 0 30912 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31096 0 1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_45_328
timestamp 1586364061
transform 1 0 31280 0 1 26656
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__336__B
timestamp 1586364061
transform 1 0 31648 0 1 26656
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31832 0 1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_45_341
timestamp 1586364061
transform 1 0 32476 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_337
timestamp 1586364061
transform 1 0 32108 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32292 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_345
timestamp 1586364061
transform 1 0 32844 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__336__A
timestamp 1586364061
transform 1 0 32660 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__314__A
timestamp 1586364061
transform 1 0 33028 0 1 26656
box -38 -48 222 592
use scs8hd_nor2_4  _314_
timestamp 1586364061
transform 1 0 33212 0 1 26656
box -38 -48 866 592
use scs8hd_conb_1  _437_
timestamp 1586364061
transform 1 0 34868 0 1 26656
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_539
timestamp 1586364061
transform 1 0 34776 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34592 0 1 26656
box -38 -48 222 592
use scs8hd_decap_6  FILLER_45_358
timestamp 1586364061
transform 1 0 34040 0 1 26656
box -38 -48 590 592
use scs8hd_decap_6  FILLER_45_370
timestamp 1586364061
transform 1 0 35144 0 1 26656
box -38 -48 590 592
use scs8hd_nor2_4  _256_
timestamp 1586364061
transform 1 0 36616 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 37720 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__259__A
timestamp 1586364061
transform 1 0 36064 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__256__A
timestamp 1586364061
transform 1 0 36432 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__259__B
timestamp 1586364061
transform 1 0 35696 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_378
timestamp 1586364061
transform 1 0 35880 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_382
timestamp 1586364061
transform 1 0 36248 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_45_395
timestamp 1586364061
transform 1 0 37444 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  FILLER_45_400
timestamp 1586364061
transform 1 0 37904 0 1 26656
box -38 -48 314 592
use scs8hd_decap_4  FILLER_45_412
timestamp 1586364061
transform 1 0 39008 0 1 26656
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38180 0 1 26656
box -38 -48 866 592
use scs8hd_fill_2  FILLER_45_419
timestamp 1586364061
transform 1 0 39652 0 1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_45_416
timestamp 1586364061
transform 1 0 39376 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39836 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39468 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_423
timestamp 1586364061
transform 1 0 40020 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__260__A
timestamp 1586364061
transform 1 0 40204 0 1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_540
timestamp 1586364061
transform 1 0 40388 0 1 26656
box -38 -48 130 592
use scs8hd_nor2_4  _260_
timestamp 1586364061
transform 1 0 40480 0 1 26656
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42044 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 41492 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41860 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_437
timestamp 1586364061
transform 1 0 41308 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_441
timestamp 1586364061
transform 1 0 41676 0 1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_45_454
timestamp 1586364061
transform 1 0 42872 0 1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_45_463
timestamp 1586364061
transform 1 0 43700 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_459
timestamp 1586364061
transform 1 0 43332 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43148 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43516 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43884 0 1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44068 0 1 26656
box -38 -48 866 592
use scs8hd_fill_2  FILLER_45_483
timestamp 1586364061
transform 1 0 45540 0 1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_45_480
timestamp 1586364061
transform 1 0 45264 0 1 26656
box -38 -48 130 592
use scs8hd_decap_4  FILLER_45_476
timestamp 1586364061
transform 1 0 44896 0 1 26656
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45356 0 1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_541
timestamp 1586364061
transform 1 0 46000 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45724 0 1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_45_487
timestamp 1586364061
transform 1 0 45908 0 1 26656
box -38 -48 130 592
use scs8hd_decap_12  FILLER_45_489
timestamp 1586364061
transform 1 0 46092 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_45_501
timestamp 1586364061
transform 1 0 47196 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 48852 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  FILLER_45_513
timestamp 1586364061
transform 1 0 48300 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_15
timestamp 1586364061
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_15
timestamp 1586364061
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_542
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_27
timestamp 1586364061
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use scs8hd_decap_12  FILLER_46_32
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_44
timestamp 1586364061
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_27
timestamp 1586364061
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_39
timestamp 1586364061
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_47_51
timestamp 1586364061
transform 1 0 5796 0 1 27744
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_550
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_56
timestamp 1586364061
transform 1 0 6256 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_68
timestamp 1586364061
transform 1 0 7360 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_46_80
timestamp 1586364061
transform 1 0 8464 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_59
timestamp 1586364061
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_62
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_74
timestamp 1586364061
transform 1 0 7912 0 1 27744
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_47_90
timestamp 1586364061
transform 1 0 9384 0 1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_47_86
timestamp 1586364061
transform 1 0 9016 0 1 27744
box -38 -48 406 592
use scs8hd_decap_8  FILLER_46_84
timestamp 1586364061
transform 1 0 8832 0 -1 27744
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_543
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9476 0 1 27744
box -38 -48 314 592
use scs8hd_conb_1  _433_
timestamp 1586364061
transform 1 0 8556 0 -1 27744
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9844 0 -1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9936 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_93
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_98
timestamp 1586364061
transform 1 0 10120 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_94
timestamp 1586364061
transform 1 0 9752 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_98
timestamp 1586364061
transform 1 0 10120 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__352__A
timestamp 1586364061
transform 1 0 10304 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__352__B
timestamp 1586364061
transform 1 0 10672 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_102
timestamp 1586364061
transform 1 0 10488 0 -1 27744
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10488 0 1 27744
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10856 0 -1 27744
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_47_117
timestamp 1586364061
transform 1 0 11868 0 1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_47_113
timestamp 1586364061
transform 1 0 11500 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_46_117
timestamp 1586364061
transform 1 0 11868 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_127
timestamp 1586364061
transform 1 0 12788 0 1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_47_123
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_120
timestamp 1586364061
transform 1 0 12144 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_125
timestamp 1586364061
transform 1 0 12604 0 -1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_46_121
timestamp 1586364061
transform 1 0 12236 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11960 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_551
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_46_132
timestamp 1586364061
transform 1 0 13248 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_129
timestamp 1586364061
transform 1 0 12972 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12880 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 -1 27744
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 1 27744
box -38 -48 866 592
use scs8hd_decap_4  FILLER_47_144
timestamp 1586364061
transform 1 0 14352 0 1 27744
box -38 -48 406 592
use scs8hd_decap_3  FILLER_47_139
timestamp 1586364061
transform 1 0 13892 0 1 27744
box -38 -48 314 592
use scs8hd_decap_8  FILLER_46_143
timestamp 1586364061
transform 1 0 14260 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_148
timestamp 1586364061
transform 1 0 14720 0 1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_544
timestamp 1586364061
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14996 0 1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_160
timestamp 1586364061
transform 1 0 15824 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_168
timestamp 1586364061
transform 1 0 16560 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_164
timestamp 1586364061
transform 1 0 16192 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_171
timestamp 1586364061
transform 1 0 16836 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_163
timestamp 1586364061
transform 1 0 16100 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 27744
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_47_184
timestamp 1586364061
transform 1 0 18032 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_179
timestamp 1586364061
transform 1 0 17572 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_175
timestamp 1586364061
transform 1 0 17204 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_182
timestamp 1586364061
transform 1 0 17848 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__349__B
timestamp 1586364061
transform 1 0 18032 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_552
timestamp 1586364061
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_46_186
timestamp 1586364061
transform 1 0 18216 0 -1 27744
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18124 0 1 27744
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_47_196
timestamp 1586364061
transform 1 0 19136 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 27744
box -38 -48 866 592
use scs8hd_decap_3  FILLER_47_205
timestamp 1586364061
transform 1 0 19964 0 1 27744
box -38 -48 314 592
use scs8hd_decap_3  FILLER_47_200
timestamp 1586364061
transform 1 0 19504 0 1 27744
box -38 -48 314 592
use scs8hd_decap_4  FILLER_46_206
timestamp 1586364061
transform 1 0 20056 0 -1 27744
box -38 -48 406 592
use scs8hd_fill_1  FILLER_46_203
timestamp 1586364061
transform 1 0 19780 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_199
timestamp 1586364061
transform 1 0 19412 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__326__B
timestamp 1586364061
transform 1 0 19872 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19320 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_212
timestamp 1586364061
transform 1 0 20608 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__361__B
timestamp 1586364061
transform 1 0 20424 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__361__A
timestamp 1586364061
transform 1 0 20240 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_545
timestamp 1586364061
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use scs8hd_nor2_4  _361_
timestamp 1586364061
transform 1 0 20424 0 1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_223
timestamp 1586364061
transform 1 0 21620 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_219
timestamp 1586364061
transform 1 0 21252 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_215
timestamp 1586364061
transform 1 0 20884 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21436 0 1 27744
box -38 -48 222 592
use scs8hd_nor2_4  _360_
timestamp 1586364061
transform 1 0 21068 0 -1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_233
timestamp 1586364061
transform 1 0 22540 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_47_227
timestamp 1586364061
transform 1 0 21988 0 1 27744
box -38 -48 314 592
use scs8hd_decap_8  FILLER_46_226
timestamp 1586364061
transform 1 0 21896 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21804 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 27744
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22264 0 1 27744
box -38 -48 314 592
use scs8hd_decap_3  FILLER_47_241
timestamp 1586364061
transform 1 0 23276 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_237
timestamp 1586364061
transform 1 0 22908 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23092 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_249
timestamp 1586364061
transform 1 0 24012 0 1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_47_245
timestamp 1586364061
transform 1 0 23644 0 1 27744
box -38 -48 406 592
use scs8hd_decap_8  FILLER_46_247
timestamp 1586364061
transform 1 0 23828 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_46_243
timestamp 1586364061
transform 1 0 23460 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24104 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_553
timestamp 1586364061
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_259
timestamp 1586364061
transform 1 0 24932 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_255
timestamp 1586364061
transform 1 0 24564 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_259
timestamp 1586364061
transform 1 0 24932 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_255
timestamp 1586364061
transform 1 0 24564 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25116 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25116 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24748 0 1 27744
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 -1 27744
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24288 0 1 27744
box -38 -48 314 592
use scs8hd_decap_8  FILLER_46_267
timestamp 1586364061
transform 1 0 25668 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_46_263
timestamp 1586364061
transform 1 0 25300 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25484 0 -1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25300 0 1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_278
timestamp 1586364061
transform 1 0 26680 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_47_272
timestamp 1586364061
transform 1 0 26128 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_46_276
timestamp 1586364061
transform 1 0 26496 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26680 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26496 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_546
timestamp 1586364061
transform 1 0 26404 0 -1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_287
timestamp 1586364061
transform 1 0 27508 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_283
timestamp 1586364061
transform 1 0 27140 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_280
timestamp 1586364061
transform 1 0 26864 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27324 0 1 27744
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26864 0 1 27744
box -38 -48 314 592
use scs8hd_or4_4  _254_
timestamp 1586364061
transform 1 0 27232 0 -1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_294
timestamp 1586364061
transform 1 0 28152 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_293
timestamp 1586364061
transform 1 0 28060 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__337__B
timestamp 1586364061
transform 1 0 28244 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__337__A
timestamp 1586364061
transform 1 0 27692 0 1 27744
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27876 0 1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_47_302
timestamp 1586364061
transform 1 0 28888 0 1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_47_298
timestamp 1586364061
transform 1 0 28520 0 1 27744
box -38 -48 406 592
use scs8hd_decap_4  FILLER_46_297
timestamp 1586364061
transform 1 0 28428 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28336 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_554
timestamp 1586364061
transform 1 0 29164 0 1 27744
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 29256 0 1 27744
box -38 -48 1050 592
use scs8hd_nor2_4  _339_
timestamp 1586364061
transform 1 0 28796 0 -1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_317
timestamp 1586364061
transform 1 0 30268 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_317
timestamp 1586364061
transform 1 0 30268 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_1  FILLER_46_314
timestamp 1586364061
transform 1 0 29992 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_310
timestamp 1586364061
transform 1 0 29624 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__315__B
timestamp 1586364061
transform 1 0 30084 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_321
timestamp 1586364061
transform 1 0 30636 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 30452 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_333
timestamp 1586364061
transform 1 0 31740 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_329
timestamp 1586364061
transform 1 0 31372 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_325
timestamp 1586364061
transform 1 0 31004 0 1 27744
box -38 -48 130 592
use scs8hd_decap_8  FILLER_46_328
timestamp 1586364061
transform 1 0 31280 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30820 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31556 0 1 27744
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31096 0 1 27744
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31004 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_346
timestamp 1586364061
transform 1 0 32936 0 -1 27744
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 31924 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_547
timestamp 1586364061
transform 1 0 32016 0 -1 27744
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch
timestamp 1586364061
transform 1 0 32108 0 1 27744
box -38 -48 1050 592
use scs8hd_nor2_4  _336_
timestamp 1586364061
transform 1 0 32108 0 -1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_348
timestamp 1586364061
transform 1 0 33120 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_47_356
timestamp 1586364061
transform 1 0 33856 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_352
timestamp 1586364061
transform 1 0 33488 0 1 27744
box -38 -48 222 592
use scs8hd_decap_6  FILLER_46_358
timestamp 1586364061
transform 1 0 34040 0 -1 27744
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33672 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 33304 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_362
timestamp 1586364061
transform 1 0 34408 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_367
timestamp 1586364061
transform 1 0 34868 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_555
timestamp 1586364061
transform 1 0 34776 0 1 27744
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_1_in_1.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34592 0 -1 27744
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 27744
box -38 -48 866 592
use scs8hd_decap_8  FILLER_46_371
timestamp 1586364061
transform 1 0 35236 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35052 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_6  FILLER_47_380
timestamp 1586364061
transform 1 0 36064 0 1 27744
box -38 -48 590 592
use scs8hd_fill_2  FILLER_47_376
timestamp 1586364061
transform 1 0 35696 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_379
timestamp 1586364061
transform 1 0 35972 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35880 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36616 0 1 27744
box -38 -48 222 592
use scs8hd_nor2_4  _259_
timestamp 1586364061
transform 1 0 36064 0 -1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_396
timestamp 1586364061
transform 1 0 37536 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_47_388
timestamp 1586364061
transform 1 0 36800 0 1 27744
box -38 -48 314 592
use scs8hd_decap_6  FILLER_46_389
timestamp 1586364061
transform 1 0 36892 0 -1 27744
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37444 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37076 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37720 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_548
timestamp 1586364061
transform 1 0 37628 0 -1 27744
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37260 0 1 27744
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 37720 0 -1 27744
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_47_400
timestamp 1586364061
transform 1 0 37904 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38088 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_409
timestamp 1586364061
transform 1 0 38732 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38916 0 -1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38272 0 1 27744
box -38 -48 866 592
use scs8hd_decap_4  FILLER_47_421
timestamp 1586364061
transform 1 0 39836 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_417
timestamp 1586364061
transform 1 0 39468 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_413
timestamp 1586364061
transform 1 0 39100 0 1 27744
box -38 -48 222 592
use scs8hd_decap_4  FILLER_46_413
timestamp 1586364061
transform 1 0 39100 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39652 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39284 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 39468 0 -1 27744
box -38 -48 866 592
use scs8hd_fill_2  FILLER_47_428
timestamp 1586364061
transform 1 0 40480 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_426
timestamp 1586364061
transform 1 0 40296 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__260__B
timestamp 1586364061
transform 1 0 40480 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__262__B
timestamp 1586364061
transform 1 0 40204 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_556
timestamp 1586364061
transform 1 0 40388 0 1 27744
box -38 -48 130 592
use scs8hd_decap_3  FILLER_47_432
timestamp 1586364061
transform 1 0 40848 0 1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_46_434
timestamp 1586364061
transform 1 0 41032 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_430
timestamp 1586364061
transform 1 0 40664 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__262__A
timestamp 1586364061
transform 1 0 40664 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 41124 0 1 27744
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 41308 0 1 27744
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 41124 0 -1 27744
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_47_452
timestamp 1586364061
transform 1 0 42688 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_448
timestamp 1586364061
transform 1 0 42320 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_450
timestamp 1586364061
transform 1 0 42504 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_46_446
timestamp 1586364061
transform 1 0 42136 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42320 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42504 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42964 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_461
timestamp 1586364061
transform 1 0 43516 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_457
timestamp 1586364061
transform 1 0 43148 0 1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_46_459
timestamp 1586364061
transform 1 0 43332 0 -1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43608 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43332 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_549
timestamp 1586364061
transform 1 0 43240 0 -1 27744
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43792 0 -1 27744
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43608 0 1 27744
box -38 -48 866 592
use scs8hd_decap_12  FILLER_47_475
timestamp 1586364061
transform 1 0 44804 0 1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_471
timestamp 1586364061
transform 1 0 44436 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_473
timestamp 1586364061
transform 1 0 44620 0 -1 27744
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44620 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 45356 0 -1 27744
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_557
timestamp 1586364061
transform 1 0 46000 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_490
timestamp 1586364061
transform 1 0 46184 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_502
timestamp 1586364061
transform 1 0 47288 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_47_487
timestamp 1586364061
transform 1 0 45908 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_47_489
timestamp 1586364061
transform 1 0 46092 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_501
timestamp 1586364061
transform 1 0 47196 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 48852 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 48852 0 1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_46_514
timestamp 1586364061
transform 1 0 48392 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_47_513
timestamp 1586364061
transform 1 0 48300 0 1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_3
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_15
timestamp 1586364061
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_558
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_4  FILLER_48_27
timestamp 1586364061
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_12  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_44
timestamp 1586364061
transform 1 0 5152 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_56
timestamp 1586364061
transform 1 0 6256 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_68
timestamp 1586364061
transform 1 0 7360 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_80
timestamp 1586364061
transform 1 0 8464 0 -1 28832
box -38 -48 1142 592
use scs8hd_nor2_4  _352_
timestamp 1586364061
transform 1 0 10304 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_559
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9844 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_93
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_97
timestamp 1586364061
transform 1 0 10028 0 -1 28832
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11960 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11316 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_109
timestamp 1586364061
transform 1 0 11132 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_113
timestamp 1586364061
transform 1 0 11500 0 -1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_48_117
timestamp 1586364061
transform 1 0 11868 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_48_127
timestamp 1586364061
transform 1 0 12788 0 -1 28832
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 28832
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_560
timestamp 1586364061
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_139
timestamp 1586364061
transform 1 0 13892 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_6  FILLER_48_145
timestamp 1586364061
transform 1 0 14444 0 -1 28832
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__220__B
timestamp 1586364061
transform 1 0 16376 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18124 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_163
timestamp 1586364061
transform 1 0 16100 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_6  FILLER_48_168
timestamp 1586364061
transform 1 0 16560 0 -1 28832
box -38 -48 590 592
use scs8hd_fill_2  FILLER_48_183
timestamp 1586364061
transform 1 0 17940 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_187
timestamp 1586364061
transform 1 0 18308 0 -1 28832
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 28832
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18676 0 -1 28832
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_561
timestamp 1586364061
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__353__D
timestamp 1586364061
transform 1 0 20240 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_48_194
timestamp 1586364061
transform 1 0 18952 0 -1 28832
box -38 -48 774 592
use scs8hd_fill_1  FILLER_48_202
timestamp 1586364061
transform 1 0 19688 0 -1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_48_206
timestamp 1586364061
transform 1 0 20056 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_210
timestamp 1586364061
transform 1 0 20424 0 -1 28832
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21160 0 -1 28832
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22908 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22356 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_215
timestamp 1586364061
transform 1 0 20884 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_48_229
timestamp 1586364061
transform 1 0 22172 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_233
timestamp 1586364061
transform 1 0 22540 0 -1 28832
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24656 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_48_246
timestamp 1586364061
transform 1 0 23736 0 -1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_48_254
timestamp 1586364061
transform 1 0 24472 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_48_267
timestamp 1586364061
transform 1 0 25668 0 -1 28832
box -38 -48 774 592
use scs8hd_nor2_4  _337_
timestamp 1586364061
transform 1 0 28152 0 -1 28832
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_562
timestamp 1586364061
transform 1 0 26404 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_48_285
timestamp 1586364061
transform 1 0 27324 0 -1 28832
box -38 -48 774 592
use scs8hd_fill_1  FILLER_48_293
timestamp 1586364061
transform 1 0 28060 0 -1 28832
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 29716 0 -1 28832
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29256 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_303
timestamp 1586364061
transform 1 0 28980 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_48_308
timestamp 1586364061
transform 1 0 29440 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_48_322
timestamp 1586364061
transform 1 0 30728 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_330
timestamp 1586364061
transform 1 0 31464 0 -1 28832
box -38 -48 406 592
use scs8hd_fill_2  FILLER_48_326
timestamp 1586364061
transform 1 0 31096 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31280 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30912 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_341
timestamp 1586364061
transform 1 0 32476 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_48_337
timestamp 1586364061
transform 1 0 32108 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31832 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32292 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32752 0 -1 28832
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_563
timestamp 1586364061
transform 1 0 32016 0 -1 28832
box -38 -48 130 592
use scs8hd_fill_1  FILLER_48_346
timestamp 1586364061
transform 1 0 32936 0 -1 28832
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 33028 0 -1 28832
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34776 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34224 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_358
timestamp 1586364061
transform 1 0 34040 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_48_362
timestamp 1586364061
transform 1 0 34408 0 -1 28832
box -38 -48 406 592
use scs8hd_decap_8  FILLER_48_375
timestamp 1586364061
transform 1 0 35604 0 -1 28832
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37904 0 -1 28832
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36616 0 -1 28832
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_564
timestamp 1586364061
transform 1 0 37628 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__267__B
timestamp 1586364061
transform 1 0 37076 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37444 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_383
timestamp 1586364061
transform 1 0 36340 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_48_389
timestamp 1586364061
transform 1 0 36892 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_393
timestamp 1586364061
transform 1 0 37260 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_398
timestamp 1586364061
transform 1 0 37720 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_407
timestamp 1586364061
transform 1 0 38548 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_403
timestamp 1586364061
transform 1 0 38180 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38732 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38364 0 -1 28832
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 38916 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_6  FILLER_48_419
timestamp 1586364061
transform 1 0 39652 0 -1 28832
box -38 -48 590 592
use scs8hd_decap_3  FILLER_48_414
timestamp 1586364061
transform 1 0 39192 0 -1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 39468 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_48_425
timestamp 1586364061
transform 1 0 40204 0 -1 28832
box -38 -48 130 592
use scs8hd_nor2_4  _262_
timestamp 1586364061
transform 1 0 40296 0 -1 28832
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41860 0 -1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__271__B
timestamp 1586364061
transform 1 0 42320 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 41308 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 41676 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_435
timestamp 1586364061
transform 1 0 41124 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_439
timestamp 1586364061
transform 1 0 41492 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_446
timestamp 1586364061
transform 1 0 42136 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_48_450
timestamp 1586364061
transform 1 0 42504 0 -1 28832
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44344 0 -1 28832
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 43332 0 -1 28832
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_565
timestamp 1586364061
transform 1 0 43240 0 -1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43792 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 44160 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_462
timestamp 1586364061
transform 1 0 43608 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_466
timestamp 1586364061
transform 1 0 43976 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_48_473
timestamp 1586364061
transform 1 0 44620 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_485
timestamp 1586364061
transform 1 0 45724 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_497
timestamp 1586364061
transform 1 0 46828 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_48_509
timestamp 1586364061
transform 1 0 47932 0 -1 28832
box -38 -48 590 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 48852 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_1  FILLER_48_515
timestamp 1586364061
transform 1 0 48484 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_15
timestamp 1586364061
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_27
timestamp 1586364061
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_39
timestamp 1586364061
transform 1 0 4692 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_49_51
timestamp 1586364061
transform 1 0 5796 0 1 28832
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_566
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_49_59
timestamp 1586364061
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_62
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_74
timestamp 1586364061
transform 1 0 7912 0 1 28832
box -38 -48 1142 592
use scs8hd_nor2_4  _224_
timestamp 1586364061
transform 1 0 10212 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__224__A
timestamp 1586364061
transform 1 0 10028 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__224__B
timestamp 1586364061
transform 1 0 9660 0 1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_49_86
timestamp 1586364061
transform 1 0 9016 0 1 28832
box -38 -48 590 592
use scs8hd_fill_1  FILLER_49_92
timestamp 1586364061
transform 1 0 9568 0 1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_49_95
timestamp 1586364061
transform 1 0 9844 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_116
timestamp 1586364061
transform 1 0 11776 0 1 28832
box -38 -48 406 592
use scs8hd_fill_2  FILLER_49_112
timestamp 1586364061
transform 1 0 11408 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_108
timestamp 1586364061
transform 1 0 11040 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11592 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11224 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__219__A
timestamp 1586364061
transform 1 0 12144 0 1 28832
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_567
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_nor2_4  _219_
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 866 592
use scs8hd_fill_2  FILLER_49_132
timestamp 1586364061
transform 1 0 13248 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_49_140
timestamp 1586364061
transform 1 0 13984 0 1 28832
box -38 -48 590 592
use scs8hd_fill_2  FILLER_49_136
timestamp 1586364061
transform 1 0 13616 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_151
timestamp 1586364061
transform 1 0 14996 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15180 0 1 28832
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14720 0 1 28832
box -38 -48 314 592
use scs8hd_decap_4  FILLER_49_159
timestamp 1586364061
transform 1 0 15732 0 1 28832
box -38 -48 406 592
use scs8hd_fill_2  FILLER_49_155
timestamp 1586364061
transform 1 0 15364 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_49_163
timestamp 1586364061
transform 1 0 16100 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__220__A
timestamp 1586364061
transform 1 0 16192 0 1 28832
box -38 -48 222 592
use scs8hd_nor2_4  _220_
timestamp 1586364061
transform 1 0 16376 0 1 28832
box -38 -48 866 592
use scs8hd_fill_2  FILLER_49_179
timestamp 1586364061
transform 1 0 17572 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_175
timestamp 1586364061
transform 1 0 17204 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_187
timestamp 1586364061
transform 1 0 18308 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 28832
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_568
timestamp 1586364061
transform 1 0 17940 0 1 28832
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_49_195
timestamp 1586364061
transform 1 0 19044 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_191
timestamp 1586364061
transform 1 0 18676 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18860 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_1.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_203
timestamp 1586364061
transform 1 0 19780 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_199
timestamp 1586364061
transform 1 0 19412 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__353__C
timestamp 1586364061
transform 1 0 19596 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__353__A
timestamp 1586364061
transform 1 0 19964 0 1 28832
box -38 -48 222 592
use scs8hd_or4_4  _353_
timestamp 1586364061
transform 1 0 20148 0 1 28832
box -38 -48 866 592
use scs8hd_nor2_4  _358_
timestamp 1586364061
transform 1 0 21712 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21160 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 22724 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__358__A
timestamp 1586364061
transform 1 0 21528 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_216
timestamp 1586364061
transform 1 0 20976 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_220
timestamp 1586364061
transform 1 0 21344 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_233
timestamp 1586364061
transform 1 0 22540 0 1 28832
box -38 -48 222 592
use scs8hd_decap_6  FILLER_49_237
timestamp 1586364061
transform 1 0 22908 0 1 28832
box -38 -48 590 592
use scs8hd_fill_2  FILLER_49_250
timestamp 1586364061
transform 1 0 24104 0 1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_49_245
timestamp 1586364061
transform 1 0 23644 0 1 28832
box -38 -48 314 592
use scs8hd_fill_1  FILLER_49_243
timestamp 1586364061
transform 1 0 23460 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 1 28832
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_569
timestamp 1586364061
transform 1 0 23552 0 1 28832
box -38 -48 130 592
use scs8hd_decap_6  FILLER_49_257
timestamp 1586364061
transform 1 0 24748 0 1 28832
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24288 0 1 28832
box -38 -48 222 592
use scs8hd_conb_1  _432_
timestamp 1586364061
transform 1 0 24472 0 1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25300 0 1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25484 0 1 28832
box -38 -48 866 592
use scs8hd_inv_8  _130_
timestamp 1586364061
transform 1 0 27048 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 26864 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26496 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__338__A
timestamp 1586364061
transform 1 0 28152 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_274
timestamp 1586364061
transform 1 0 26312 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_278
timestamp 1586364061
transform 1 0 26680 0 1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_49_291
timestamp 1586364061
transform 1 0 27876 0 1 28832
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch
timestamp 1586364061
transform 1 0 29256 0 1 28832
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_570
timestamp 1586364061
transform 1 0 29164 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__338__B
timestamp 1586364061
transform 1 0 28520 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30452 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_296
timestamp 1586364061
transform 1 0 28336 0 1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_49_300
timestamp 1586364061
transform 1 0 28704 0 1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_49_317
timestamp 1586364061
transform 1 0 30268 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_321
timestamp 1586364061
transform 1 0 30636 0 1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31004 0 1 28832
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32752 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__342__A
timestamp 1586364061
transform 1 0 32108 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__342__B
timestamp 1586364061
transform 1 0 32476 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30820 0 1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_49_334
timestamp 1586364061
transform 1 0 31832 0 1 28832
box -38 -48 314 592
use scs8hd_fill_2  FILLER_49_339
timestamp 1586364061
transform 1 0 32292 0 1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_49_343
timestamp 1586364061
transform 1 0 32660 0 1 28832
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_571
timestamp 1586364061
transform 1 0 34776 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33948 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_353
timestamp 1586364061
transform 1 0 33580 0 1 28832
box -38 -48 406 592
use scs8hd_decap_4  FILLER_49_359
timestamp 1586364061
transform 1 0 34132 0 1 28832
box -38 -48 406 592
use scs8hd_fill_1  FILLER_49_363
timestamp 1586364061
transform 1 0 34500 0 1 28832
box -38 -48 130 592
use scs8hd_nor2_4  _267_
timestamp 1586364061
transform 1 0 36616 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 37720 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36432 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35880 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_376
timestamp 1586364061
transform 1 0 35696 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_380
timestamp 1586364061
transform 1 0 36064 0 1 28832
box -38 -48 406 592
use scs8hd_decap_3  FILLER_49_395
timestamp 1586364061
transform 1 0 37444 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_49_400
timestamp 1586364061
transform 1 0 37904 0 1 28832
box -38 -48 314 592
use scs8hd_decap_4  FILLER_49_412
timestamp 1586364061
transform 1 0 39008 0 1 28832
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38180 0 1 28832
box -38 -48 866 592
use scs8hd_fill_2  FILLER_49_419
timestamp 1586364061
transform 1 0 39652 0 1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_49_416
timestamp 1586364061
transform 1 0 39376 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__264__B
timestamp 1586364061
transform 1 0 39836 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 39468 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_423
timestamp 1586364061
transform 1 0 40020 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__264__A
timestamp 1586364061
transform 1 0 40204 0 1 28832
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_572
timestamp 1586364061
transform 1 0 40388 0 1 28832
box -38 -48 130 592
use scs8hd_nor2_4  _264_
timestamp 1586364061
transform 1 0 40480 0 1 28832
box -38 -48 866 592
use scs8hd_nor2_4  _271_
timestamp 1586364061
transform 1 0 42044 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 41492 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__271__A
timestamp 1586364061
transform 1 0 41860 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_437
timestamp 1586364061
transform 1 0 41308 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_441
timestamp 1586364061
transform 1 0 41676 0 1 28832
box -38 -48 222 592
use scs8hd_decap_4  FILLER_49_454
timestamp 1586364061
transform 1 0 42872 0 1 28832
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43700 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 43332 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 45080 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44712 0 1 28832
box -38 -48 222 592
use scs8hd_fill_1  FILLER_49_458
timestamp 1586364061
transform 1 0 43240 0 1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_49_461
timestamp 1586364061
transform 1 0 43516 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_472
timestamp 1586364061
transform 1 0 44528 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_476
timestamp 1586364061
transform 1 0 44896 0 1 28832
box -38 -48 222 592
use scs8hd_decap_8  FILLER_49_480
timestamp 1586364061
transform 1 0 45264 0 1 28832
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_573
timestamp 1586364061
transform 1 0 46000 0 1 28832
box -38 -48 130 592
use scs8hd_decap_12  FILLER_49_489
timestamp 1586364061
transform 1 0 46092 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_501
timestamp 1586364061
transform 1 0 47196 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 48852 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_49_513
timestamp 1586364061
transform 1 0 48300 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_3
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_15
timestamp 1586364061
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_574
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_50_27
timestamp 1586364061
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_12  FILLER_50_32
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_44
timestamp 1586364061
transform 1 0 5152 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_56
timestamp 1586364061
transform 1 0 6256 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_68
timestamp 1586364061
transform 1 0 7360 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_80
timestamp 1586364061
transform 1 0 8464 0 -1 29920
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10856 0 -1 29920
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9844 0 -1 29920
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_575
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__218__A
timestamp 1586364061
transform 1 0 10304 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_93
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_98
timestamp 1586364061
transform 1 0 10120 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_102
timestamp 1586364061
transform 1 0 10488 0 -1 29920
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_6_.latch
timestamp 1586364061
transform 1 0 12972 0 -1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__219__B
timestamp 1586364061
transform 1 0 12420 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_50_117
timestamp 1586364061
transform 1 0 11868 0 -1 29920
box -38 -48 590 592
use scs8hd_decap_4  FILLER_50_125
timestamp 1586364061
transform 1 0 12604 0 -1 29920
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_576
timestamp 1586364061
transform 1 0 15180 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_50_140
timestamp 1586364061
transform 1 0 13984 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_3  FILLER_50_148
timestamp 1586364061
transform 1 0 14720 0 -1 29920
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16928 0 -1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18124 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_50_163
timestamp 1586364061
transform 1 0 16100 0 -1 29920
box -38 -48 774 592
use scs8hd_fill_1  FILLER_50_171
timestamp 1586364061
transform 1 0 16836 0 -1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_50_183
timestamp 1586364061
transform 1 0 17940 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_187
timestamp 1586364061
transform 1 0 18308 0 -1 29920
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_577
timestamp 1586364061
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__353__B
timestamp 1586364061
transform 1 0 20148 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18492 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_50_200
timestamp 1586364061
transform 1 0 19504 0 -1 29920
box -38 -48 590 592
use scs8hd_fill_1  FILLER_50_206
timestamp 1586364061
transform 1 0 20056 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_50_209
timestamp 1586364061
transform 1 0 20332 0 -1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_50_213
timestamp 1586364061
transform 1 0 20700 0 -1 29920
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 22172 0 -1 29920
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 -1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__359__B
timestamp 1586364061
transform 1 0 21620 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__358__B
timestamp 1586364061
transform 1 0 21988 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_50_215
timestamp 1586364061
transform 1 0 20884 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_50_221
timestamp 1586364061
transform 1 0 21436 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_225
timestamp 1586364061
transform 1 0 21804 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_50_240
timestamp 1586364061
transform 1 0 23184 0 -1 29920
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23920 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25484 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24932 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_257
timestamp 1586364061
transform 1 0 24748 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_261
timestamp 1586364061
transform 1 0 25116 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_6  FILLER_50_267
timestamp 1586364061
transform 1 0 25668 0 -1 29920
box -38 -48 590 592
use scs8hd_nor2_4  _338_
timestamp 1586364061
transform 1 0 28152 0 -1 29920
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 29920
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_578
timestamp 1586364061
transform 1 0 26404 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__335__C
timestamp 1586364061
transform 1 0 27048 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__335__D
timestamp 1586364061
transform 1 0 27416 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_50_279
timestamp 1586364061
transform 1 0 26772 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_50_284
timestamp 1586364061
transform 1 0 27232 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_50_288
timestamp 1586364061
transform 1 0 27600 0 -1 29920
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30176 0 -1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29256 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29992 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_3  FILLER_50_303
timestamp 1586364061
transform 1 0 28980 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_6  FILLER_50_308
timestamp 1586364061
transform 1 0 29440 0 -1 29920
box -38 -48 590 592
use scs8hd_nor2_4  _342_
timestamp 1586364061
transform 1 0 32108 0 -1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_579
timestamp 1586364061
transform 1 0 32016 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31188 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_325
timestamp 1586364061
transform 1 0 31004 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_50_329
timestamp 1586364061
transform 1 0 31372 0 -1 29920
box -38 -48 590 592
use scs8hd_fill_1  FILLER_50_335
timestamp 1586364061
transform 1 0 31924 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_3  FILLER_50_346
timestamp 1586364061
transform 1 0 32936 0 -1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_50_355
timestamp 1586364061
transform 1 0 33764 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_351
timestamp 1586364061
transform 1 0 33396 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33580 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33212 0 -1 29920
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33948 0 -1 29920
box -38 -48 866 592
use scs8hd_fill_2  FILLER_50_366
timestamp 1586364061
transform 1 0 34776 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34960 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_370
timestamp 1586364061
transform 1 0 35144 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35328 0 -1 29920
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35512 0 -1 29920
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 37720 0 -1 29920
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36524 0 -1 29920
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_580
timestamp 1586364061
transform 1 0 37628 0 -1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__267__A
timestamp 1586364061
transform 1 0 36984 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37352 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_50_377
timestamp 1586364061
transform 1 0 35788 0 -1 29920
box -38 -48 774 592
use scs8hd_fill_2  FILLER_50_388
timestamp 1586364061
transform 1 0 36800 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_50_392
timestamp 1586364061
transform 1 0 37168 0 -1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_50_396
timestamp 1586364061
transform 1 0 37536 0 -1 29920
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_6_.latch
timestamp 1586364061
transform 1 0 39468 0 -1 29920
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_50_409
timestamp 1586364061
transform 1 0 38732 0 -1 29920
box -38 -48 774 592
use scs8hd_fill_2  FILLER_50_428
timestamp 1586364061
transform 1 0 40480 0 -1 29920
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_7_.latch
timestamp 1586364061
transform 1 0 41216 0 -1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43056 0 -1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40664 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_50_432
timestamp 1586364061
transform 1 0 40848 0 -1 29920
box -38 -48 406 592
use scs8hd_decap_8  FILLER_50_447
timestamp 1586364061
transform 1 0 42228 0 -1 29920
box -38 -48 774 592
use scs8hd_fill_1  FILLER_50_455
timestamp 1586364061
transform 1 0 42964 0 -1 29920
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 43332 0 -1 29920
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 45080 0 -1 29920
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_581
timestamp 1586364061
transform 1 0 43240 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_8  FILLER_50_470
timestamp 1586364061
transform 1 0 44344 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_12  FILLER_50_481
timestamp 1586364061
transform 1 0 45356 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_493
timestamp 1586364061
transform 1 0 46460 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_50_505
timestamp 1586364061
transform 1 0 47564 0 -1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 48852 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_50_513
timestamp 1586364061
transform 1 0 48300 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_51_3
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_15
timestamp 1586364061
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_27
timestamp 1586364061
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_39
timestamp 1586364061
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_51
timestamp 1586364061
transform 1 0 5796 0 1 29920
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_582
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_59
timestamp 1586364061
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_51_62
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_74
timestamp 1586364061
transform 1 0 7912 0 1 29920
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch
timestamp 1586364061
transform 1 0 10580 0 1 29920
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9568 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__218__B
timestamp 1586364061
transform 1 0 9384 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_86
timestamp 1586364061
transform 1 0 9016 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_95
timestamp 1586364061
transform 1 0 9844 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_99
timestamp 1586364061
transform 1 0 10212 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_114
timestamp 1586364061
transform 1 0 11592 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_118
timestamp 1586364061
transform 1 0 11960 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 29920
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_583
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_51_128
timestamp 1586364061
transform 1 0 12880 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13064 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_132
timestamp 1586364061
transform 1 0 13248 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 29920
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15180 0 1 29920
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_145
timestamp 1586364061
transform 1 0 14444 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_149
timestamp 1586364061
transform 1 0 14812 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_162
timestamp 1586364061
transform 1 0 16008 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_166
timestamp 1586364061
transform 1 0 16376 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 1 29920
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_51_173
timestamp 1586364061
transform 1 0 17020 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17204 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_177
timestamp 1586364061
transform 1 0 17388 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17572 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_184
timestamp 1586364061
transform 1 0 18032 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_181
timestamp 1586364061
transform 1 0 17756 0 1 29920
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_584
timestamp 1586364061
transform 1 0 17940 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__221__A
timestamp 1586364061
transform 1 0 18216 0 1 29920
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18768 0 1 29920
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20792 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 18584 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__359__A
timestamp 1586364061
transform 1 0 20608 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__221__B
timestamp 1586364061
transform 1 0 19964 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_188
timestamp 1586364061
transform 1 0 18400 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_203
timestamp 1586364061
transform 1 0 19780 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_207
timestamp 1586364061
transform 1 0 20148 0 1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_51_211
timestamp 1586364061
transform 1 0 20516 0 1 29920
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 21804 0 1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21252 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_217
timestamp 1586364061
transform 1 0 21068 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_221
timestamp 1586364061
transform 1 0 21436 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_236
timestamp 1586364061
transform 1 0 22816 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_240
timestamp 1586364061
transform 1 0 23184 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_248
timestamp 1586364061
transform 1 0 23920 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 29920
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_585
timestamp 1586364061
transform 1 0 23552 0 1 29920
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_51_252
timestamp 1586364061
transform 1 0 24288 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24472 0 1 29920
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24656 0 1 29920
box -38 -48 866 592
use scs8hd_fill_2  FILLER_51_265
timestamp 1586364061
transform 1 0 25484 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25668 0 1 29920
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26220 0 1 29920
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28152 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__335__A
timestamp 1586364061
transform 1 0 27232 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__335__B
timestamp 1586364061
transform 1 0 27600 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26036 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_269
timestamp 1586364061
transform 1 0 25852 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_282
timestamp 1586364061
transform 1 0 27048 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_286
timestamp 1586364061
transform 1 0 27416 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_290
timestamp 1586364061
transform 1 0 27784 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_301
timestamp 1586364061
transform 1 0 28796 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_297
timestamp 1586364061
transform 1 0 28428 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28980 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28612 0 1 29920
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_586
timestamp 1586364061
transform 1 0 29164 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_313
timestamp 1586364061
transform 1 0 29900 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_306
timestamp 1586364061
transform 1 0 29256 0 1 29920
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29624 0 1 29920
box -38 -48 314 592
use scs8hd_fill_1  FILLER_51_321
timestamp 1586364061
transform 1 0 30636 0 1 29920
box -38 -48 130 592
use scs8hd_fill_2  FILLER_51_317
timestamp 1586364061
transform 1 0 30268 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30452 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30084 0 1 29920
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30728 0 1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32936 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32568 0 1 29920
box -38 -48 222 592
use scs8hd_decap_8  FILLER_51_331
timestamp 1586364061
transform 1 0 31556 0 1 29920
box -38 -48 774 592
use scs8hd_decap_3  FILLER_51_339
timestamp 1586364061
transform 1 0 32292 0 1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_51_344
timestamp 1586364061
transform 1 0 32752 0 1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_51_348
timestamp 1586364061
transform 1 0 33120 0 1 29920
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 29920
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 29920
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_587
timestamp 1586364061
transform 1 0 34776 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34500 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_358
timestamp 1586364061
transform 1 0 34040 0 1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_51_362
timestamp 1586364061
transform 1 0 34408 0 1 29920
box -38 -48 130 592
use scs8hd_fill_1  FILLER_51_365
timestamp 1586364061
transform 1 0 34684 0 1 29920
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 37352 0 1 29920
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 37168 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36064 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_376
timestamp 1586364061
transform 1 0 35696 0 1 29920
box -38 -48 406 592
use scs8hd_decap_8  FILLER_51_382
timestamp 1586364061
transform 1 0 36248 0 1 29920
box -38 -48 774 592
use scs8hd_fill_2  FILLER_51_390
timestamp 1586364061
transform 1 0 36984 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_405
timestamp 1586364061
transform 1 0 38364 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38548 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_409
timestamp 1586364061
transform 1 0 38732 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38916 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_416
timestamp 1586364061
transform 1 0 39376 0 1 29920
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39100 0 1 29920
box -38 -48 314 592
use scs8hd_decap_4  FILLER_51_420
timestamp 1586364061
transform 1 0 39744 0 1 29920
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39560 0 1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_51_424
timestamp 1586364061
transform 1 0 40112 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_428
timestamp 1586364061
transform 1 0 40480 0 1 29920
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_588
timestamp 1586364061
transform 1 0 40388 0 1 29920
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42688 0 1 29920
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41124 0 1 29920
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42228 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40940 0 1 29920
box -38 -48 222 592
use scs8hd_fill_1  FILLER_51_432
timestamp 1586364061
transform 1 0 40848 0 1 29920
box -38 -48 130 592
use scs8hd_decap_3  FILLER_51_444
timestamp 1586364061
transform 1 0 41952 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_51_449
timestamp 1586364061
transform 1 0 42412 0 1 29920
box -38 -48 314 592
use scs8hd_fill_2  FILLER_51_455
timestamp 1586364061
transform 1 0 42964 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_459
timestamp 1586364061
transform 1 0 43332 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43516 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43148 0 1 29920
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43700 0 1 29920
box -38 -48 866 592
use scs8hd_fill_2  FILLER_51_472
timestamp 1586364061
transform 1 0 44528 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44712 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_480
timestamp 1586364061
transform 1 0 45264 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_476
timestamp 1586364061
transform 1 0 44896 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 45448 0 1 29920
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 45080 0 1 29920
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 46092 0 1 29920
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_589
timestamp 1586364061
transform 1 0 46000 0 1 29920
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 46552 0 1 29920
box -38 -48 222 592
use scs8hd_decap_4  FILLER_51_484
timestamp 1586364061
transform 1 0 45632 0 1 29920
box -38 -48 406 592
use scs8hd_fill_2  FILLER_51_492
timestamp 1586364061
transform 1 0 46368 0 1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_51_496
timestamp 1586364061
transform 1 0 46736 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_508
timestamp 1586364061
transform 1 0 47840 0 1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 48852 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_15
timestamp 1586364061
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_15
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_590
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_27
timestamp 1586364061
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_52_32
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_44
timestamp 1586364061
transform 1 0 5152 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_27
timestamp 1586364061
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_39
timestamp 1586364061
transform 1 0 4692 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_51
timestamp 1586364061
transform 1 0 5796 0 1 31008
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_598
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_56
timestamp 1586364061
transform 1 0 6256 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_68
timestamp 1586364061
transform 1 0 7360 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_80
timestamp 1586364061
transform 1 0 8464 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_59
timestamp 1586364061
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_53_62
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_74
timestamp 1586364061
transform 1 0 7912 0 1 31008
box -38 -48 1142 592
use scs8hd_nor2_4  _218_
timestamp 1586364061
transform 1 0 10212 0 -1 31008
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_591
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__223__A
timestamp 1586364061
transform 1 0 10396 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__223__B
timestamp 1586364061
transform 1 0 10764 0 1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_52_93
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 590 592
use scs8hd_decap_12  FILLER_53_86
timestamp 1586364061
transform 1 0 9016 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_53_98
timestamp 1586364061
transform 1 0 10120 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_103
timestamp 1586364061
transform 1 0 10580 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_53_107
timestamp 1586364061
transform 1 0 10948 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_114
timestamp 1586364061
transform 1 0 11592 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_108
timestamp 1586364061
transform 1 0 11040 0 -1 31008
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11776 0 -1 31008
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_118
timestamp 1586364061
transform 1 0 11960 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_125
timestamp 1586364061
transform 1 0 12604 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_599
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_132
timestamp 1586364061
transform 1 0 13248 0 1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_52_129
timestamp 1586364061
transform 1 0 12972 0 -1 31008
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_53_144
timestamp 1586364061
transform 1 0 14352 0 1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_53_140
timestamp 1586364061
transform 1 0 13984 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_136
timestamp 1586364061
transform 1 0 13616 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_138
timestamp 1586364061
transform 1 0 13800 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_52_135
timestamp 1586364061
transform 1 0 13524 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 31008
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_152
timestamp 1586364061
transform 1 0 15088 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_148
timestamp 1586364061
transform 1 0 14720 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_145
timestamp 1586364061
transform 1 0 14444 0 -1 31008
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14904 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_592
timestamp 1586364061
transform 1 0 15180 0 -1 31008
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14444 0 1 31008
box -38 -48 314 592
use scs8hd_decap_4  FILLER_53_160
timestamp 1586364061
transform 1 0 15824 0 1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_156
timestamp 1586364061
transform 1 0 15456 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 31008
box -38 -48 866 592
use scs8hd_decap_4  FILLER_52_168
timestamp 1586364061
transform 1 0 16560 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_3  FILLER_52_163
timestamp 1586364061
transform 1 0 16100 0 -1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__222__B
timestamp 1586364061
transform 1 0 16376 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__222__A
timestamp 1586364061
transform 1 0 16192 0 1 31008
box -38 -48 222 592
use scs8hd_nor2_4  _222_
timestamp 1586364061
transform 1 0 16376 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_179
timestamp 1586364061
transform 1 0 17572 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_175
timestamp 1586364061
transform 1 0 17204 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_175
timestamp 1586364061
transform 1 0 17204 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_52_172
timestamp 1586364061
transform 1 0 16928 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17388 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_1  FILLER_53_184
timestamp 1586364061
transform 1 0 18032 0 1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_52_186
timestamp 1586364061
transform 1 0 18216 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 17756 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_600
timestamp 1586364061
transform 1 0 17940 0 1 31008
box -38 -48 130 592
use scs8hd_or2_4  _163_
timestamp 1586364061
transform 1 0 18124 0 1 31008
box -38 -48 682 592
use scs8hd_fill_2  FILLER_53_196
timestamp 1586364061
transform 1 0 19136 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_192
timestamp 1586364061
transform 1 0 18768 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_190
timestamp 1586364061
transform 1 0 18584 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__217__C
timestamp 1586364061
transform 1 0 18768 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__217__A
timestamp 1586364061
transform 1 0 18952 0 1 31008
box -38 -48 222 592
use scs8hd_nor2_4  _221_
timestamp 1586364061
transform 1 0 18952 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_52_207
timestamp 1586364061
transform 1 0 20148 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_203
timestamp 1586364061
transform 1 0 19780 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__B
timestamp 1586364061
transform 1 0 19964 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 19320 0 1 31008
box -38 -48 222 592
use scs8hd_or4_4  _226_
timestamp 1586364061
transform 1 0 19504 0 1 31008
box -38 -48 866 592
use scs8hd_fill_1  FILLER_53_213
timestamp 1586364061
transform 1 0 20700 0 1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_53_209
timestamp 1586364061
transform 1 0 20332 0 1 31008
box -38 -48 406 592
use scs8hd_decap_3  FILLER_52_211
timestamp 1586364061
transform 1 0 20516 0 -1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__226__C
timestamp 1586364061
transform 1 0 20332 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20792 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_593
timestamp 1586364061
transform 1 0 20792 0 -1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_216
timestamp 1586364061
transform 1 0 20976 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_52_215
timestamp 1586364061
transform 1 0 20884 0 -1 31008
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 21160 0 1 31008
box -38 -48 222 592
use scs8hd_nor2_4  _359_
timestamp 1586364061
transform 1 0 21160 0 -1 31008
box -38 -48 866 592
use scs8hd_or2_4  _164_
timestamp 1586364061
transform 1 0 21344 0 1 31008
box -38 -48 682 592
use scs8hd_fill_2  FILLER_53_231
timestamp 1586364061
transform 1 0 22356 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_227
timestamp 1586364061
transform 1 0 21988 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_231
timestamp 1586364061
transform 1 0 22356 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_52_227
timestamp 1586364061
transform 1 0 21988 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22172 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__253__A
timestamp 1586364061
transform 1 0 22540 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 22172 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_53_239
timestamp 1586364061
transform 1 0 23092 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_235
timestamp 1586364061
transform 1 0 22724 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__253__B
timestamp 1586364061
transform 1 0 22908 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22724 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_52_251
timestamp 1586364061
transform 1 0 24196 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_52_248
timestamp 1586364061
transform 1 0 23920 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_244
timestamp 1586364061
transform 1 0 23552 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24012 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__215__A
timestamp 1586364061
transform 1 0 23368 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_601
timestamp 1586364061
transform 1 0 23552 0 1 31008
box -38 -48 130 592
use scs8hd_or2_4  _215_
timestamp 1586364061
transform 1 0 23644 0 1 31008
box -38 -48 682 592
use scs8hd_fill_2  FILLER_53_260
timestamp 1586364061
transform 1 0 25024 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_256
timestamp 1586364061
transform 1 0 24656 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_252
timestamp 1586364061
transform 1 0 24288 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_52_255
timestamp 1586364061
transform 1 0 24564 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__236__B
timestamp 1586364061
transform 1 0 24380 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 24840 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__215__B
timestamp 1586364061
transform 1 0 24472 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24656 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_52_265
timestamp 1586364061
transform 1 0 25484 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25668 0 -1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25208 0 1 31008
box -38 -48 866 592
use scs8hd_decap_4  FILLER_53_278
timestamp 1586364061
transform 1 0 26680 0 1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_53_275
timestamp 1586364061
transform 1 0 26404 0 1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_53_271
timestamp 1586364061
transform 1 0 26036 0 1 31008
box -38 -48 406 592
use scs8hd_decap_6  FILLER_52_276
timestamp 1586364061
transform 1 0 26496 0 -1 31008
box -38 -48 590 592
use scs8hd_decap_6  FILLER_52_269
timestamp 1586364061
transform 1 0 25852 0 -1 31008
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26496 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_594
timestamp 1586364061
transform 1 0 26404 0 -1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_284
timestamp 1586364061
transform 1 0 27232 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__281__B
timestamp 1586364061
transform 1 0 27048 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__281__A
timestamp 1586364061
transform 1 0 27416 0 1 31008
box -38 -48 222 592
use scs8hd_nor2_4  _340_
timestamp 1586364061
transform 1 0 27600 0 1 31008
box -38 -48 866 592
use scs8hd_or4_4  _335_
timestamp 1586364061
transform 1 0 27048 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_52_295
timestamp 1586364061
transform 1 0 28244 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_291
timestamp 1586364061
transform 1 0 27876 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__281__D
timestamp 1586364061
transform 1 0 28060 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__340__A
timestamp 1586364061
transform 1 0 28612 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__281__C
timestamp 1586364061
transform 1 0 28428 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_299
timestamp 1586364061
transform 1 0 28612 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_53_297
timestamp 1586364061
transform 1 0 28428 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_301
timestamp 1586364061
transform 1 0 28796 0 1 31008
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28980 0 -1 31008
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_602
timestamp 1586364061
transform 1 0 29164 0 1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_306
timestamp 1586364061
transform 1 0 29256 0 -1 31008
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 29256 0 1 31008
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_53_317
timestamp 1586364061
transform 1 0 30268 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_52_313
timestamp 1586364061
transform 1 0 29900 0 -1 31008
box -38 -48 130 592
use scs8hd_fill_1  FILLER_52_310
timestamp 1586364061
transform 1 0 29624 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29716 0 -1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29992 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_321
timestamp 1586364061
transform 1 0 30636 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30452 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_333
timestamp 1586364061
transform 1 0 31740 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_53_328
timestamp 1586364061
transform 1 0 31280 0 1 31008
box -38 -48 314 592
use scs8hd_decap_8  FILLER_52_327
timestamp 1586364061
transform 1 0 31188 0 -1 31008
box -38 -48 774 592
use scs8hd_fill_2  FILLER_52_323
timestamp 1586364061
transform 1 0 30820 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31004 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30820 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 31556 0 1 31008
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31004 0 1 31008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_52_345
timestamp 1586364061
transform 1 0 32844 0 -1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_52_341
timestamp 1586364061
transform 1 0 32476 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_337
timestamp 1586364061
transform 1 0 32108 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_52_335
timestamp 1586364061
transform 1 0 31924 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32660 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32292 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 31924 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_595
timestamp 1586364061
transform 1 0 32016 0 -1 31008
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 32108 0 1 31008
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_53_348
timestamp 1586364061
transform 1 0 33120 0 1 31008
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32936 0 -1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_358
timestamp 1586364061
transform 1 0 34040 0 1 31008
box -38 -48 222 592
use scs8hd_decap_6  FILLER_52_355
timestamp 1586364061
transform 1 0 33764 0 -1 31008
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33856 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_362
timestamp 1586364061
transform 1 0 34408 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34316 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_603
timestamp 1586364061
transform 1 0 34776 0 1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34500 0 -1 31008
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_52_372
timestamp 1586364061
transform 1 0 35328 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35512 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_53_385
timestamp 1586364061
transform 1 0 36524 0 1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_53_381
timestamp 1586364061
transform 1 0 36156 0 1 31008
box -38 -48 406 592
use scs8hd_decap_3  FILLER_53_376
timestamp 1586364061
transform 1 0 35696 0 1 31008
box -38 -48 314 592
use scs8hd_decap_4  FILLER_52_383
timestamp 1586364061
transform 1 0 36340 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_52_376
timestamp 1586364061
transform 1 0 35696 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35880 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35972 0 1 31008
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36064 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_6  FILLER_52_390
timestamp 1586364061
transform 1 0 36984 0 -1 31008
box -38 -48 590 592
use scs8hd_fill_1  FILLER_52_387
timestamp 1586364061
transform 1 0 36708 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__266__B
timestamp 1586364061
transform 1 0 36800 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__266__A
timestamp 1586364061
transform 1 0 36616 0 1 31008
box -38 -48 222 592
use scs8hd_nor2_4  _266_
timestamp 1586364061
transform 1 0 36800 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_402
timestamp 1586364061
transform 1 0 38088 0 1 31008
box -38 -48 222 592
use scs8hd_decap_3  FILLER_53_397
timestamp 1586364061
transform 1 0 37628 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_52_402
timestamp 1586364061
transform 1 0 38088 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_398
timestamp 1586364061
transform 1 0 37720 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_52_396
timestamp 1586364061
transform 1 0 37536 0 -1 31008
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37904 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37904 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_596
timestamp 1586364061
transform 1 0 37628 0 -1 31008
box -38 -48 130 592
use scs8hd_fill_2  FILLER_53_406
timestamp 1586364061
transform 1 0 38456 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_52_413
timestamp 1586364061
transform 1 0 39100 0 -1 31008
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__265__B
timestamp 1586364061
transform 1 0 38272 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__265__A
timestamp 1586364061
transform 1 0 38640 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38272 0 -1 31008
box -38 -48 866 592
use scs8hd_nor2_4  _265_
timestamp 1586364061
transform 1 0 38824 0 1 31008
box -38 -48 866 592
use scs8hd_fill_2  FILLER_53_423
timestamp 1586364061
transform 1 0 40020 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_419
timestamp 1586364061
transform 1 0 39652 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39836 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_604
timestamp 1586364061
transform 1 0 40388 0 1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40204 0 -1 31008
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_435
timestamp 1586364061
transform 1 0 41124 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_431
timestamp 1586364061
transform 1 0 40756 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_438
timestamp 1586364061
transform 1 0 41400 0 -1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_52_434
timestamp 1586364061
transform 1 0 41032 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41216 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40940 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41308 0 1 31008
box -38 -48 222 592
use scs8hd_fill_1  FILLER_53_446
timestamp 1586364061
transform 1 0 42136 0 1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_53_442
timestamp 1586364061
transform 1 0 41768 0 1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_52_446
timestamp 1586364061
transform 1 0 42136 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_4  FILLER_52_442
timestamp 1586364061
transform 1 0 41768 0 -1 31008
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41584 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42228 0 1 31008
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41492 0 1 31008
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42228 0 -1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_453
timestamp 1586364061
transform 1 0 42780 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_449
timestamp 1586364061
transform 1 0 42412 0 1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_52_450
timestamp 1586364061
transform 1 0 42504 0 -1 31008
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42596 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42964 0 1 31008
box -38 -48 222 592
use scs8hd_fill_2  FILLER_53_457
timestamp 1586364061
transform 1 0 43148 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43332 0 1 31008
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_597
timestamp 1586364061
transform 1 0 43240 0 -1 31008
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43332 0 -1 31008
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43516 0 1 31008
box -38 -48 866 592
use scs8hd_decap_3  FILLER_53_474
timestamp 1586364061
transform 1 0 44712 0 1 31008
box -38 -48 314 592
use scs8hd_fill_2  FILLER_53_470
timestamp 1586364061
transform 1 0 44344 0 1 31008
box -38 -48 222 592
use scs8hd_decap_4  FILLER_52_472
timestamp 1586364061
transform 1 0 44528 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_2  FILLER_52_468
timestamp 1586364061
transform 1 0 44160 0 -1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44528 0 1 31008
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44344 0 -1 31008
box -38 -48 222 592
use scs8hd_decap_8  FILLER_53_479
timestamp 1586364061
transform 1 0 45172 0 1 31008
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 44988 0 1 31008
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 44896 0 -1 31008
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_605
timestamp 1586364061
transform 1 0 46000 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_485
timestamp 1586364061
transform 1 0 45724 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_497
timestamp 1586364061
transform 1 0 46828 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_52_509
timestamp 1586364061
transform 1 0 47932 0 -1 31008
box -38 -48 590 592
use scs8hd_fill_1  FILLER_53_487
timestamp 1586364061
transform 1 0 45908 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_53_489
timestamp 1586364061
transform 1 0 46092 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_501
timestamp 1586364061
transform 1 0 47196 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 48852 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 48852 0 1 31008
box -38 -48 314 592
use scs8hd_fill_1  FILLER_52_515
timestamp 1586364061
transform 1 0 48484 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_3  FILLER_53_513
timestamp 1586364061
transform 1 0 48300 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_606
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_4  FILLER_54_27
timestamp 1586364061
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_54_32
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_44
timestamp 1586364061
transform 1 0 5152 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_56
timestamp 1586364061
transform 1 0 6256 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_68
timestamp 1586364061
transform 1 0 7360 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_80
timestamp 1586364061
transform 1 0 8464 0 -1 32096
box -38 -48 1142 592
use scs8hd_nor2_4  _223_
timestamp 1586364061
transform 1 0 10396 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_607
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_8  FILLER_54_93
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 774 592
use scs8hd_decap_4  FILLER_54_114
timestamp 1586364061
transform 1 0 11592 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_54_110
timestamp 1586364061
transform 1 0 11224 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11408 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_126
timestamp 1586364061
transform 1 0 12696 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_122
timestamp 1586364061
transform 1 0 12328 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_54_118
timestamp 1586364061
transform 1 0 11960 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12512 0 -1 32096
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12052 0 -1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 32096
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 -1 32096
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_608
timestamp 1586364061
transform 1 0 15180 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_54_139
timestamp 1586364061
transform 1 0 13892 0 -1 32096
box -38 -48 774 592
use scs8hd_decap_4  FILLER_54_149
timestamp 1586364061
transform 1 0 14812 0 -1 32096
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 18124 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_54_163
timestamp 1586364061
transform 1 0 16100 0 -1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_54_168
timestamp 1586364061
transform 1 0 16560 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_54_172
timestamp 1586364061
transform 1 0 16928 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  FILLER_54_182
timestamp 1586364061
transform 1 0 17848 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_4  FILLER_54_187
timestamp 1586364061
transform 1 0 18308 0 -1 32096
box -38 -48 406 592
use scs8hd_or4_4  _217_
timestamp 1586364061
transform 1 0 19228 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_609
timestamp 1586364061
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__217__B
timestamp 1586364061
transform 1 0 19044 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__D
timestamp 1586364061
transform 1 0 20240 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__217__D
timestamp 1586364061
transform 1 0 18676 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_193
timestamp 1586364061
transform 1 0 18860 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_206
timestamp 1586364061
transform 1 0 20056 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_210
timestamp 1586364061
transform 1 0 20424 0 -1 32096
box -38 -48 406 592
use scs8hd_nand2_4  _253_
timestamp 1586364061
transform 1 0 22080 0 -1 32096
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21068 0 -1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__244__D
timestamp 1586364061
transform 1 0 21528 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 23276 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_215
timestamp 1586364061
transform 1 0 20884 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_220
timestamp 1586364061
transform 1 0 21344 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_224
timestamp 1586364061
transform 1 0 21712 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_4  FILLER_54_237
timestamp 1586364061
transform 1 0 22908 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_54_251
timestamp 1586364061
transform 1 0 24196 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_247
timestamp 1586364061
transform 1 0 23828 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_243
timestamp 1586364061
transform 1 0 23460 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__C
timestamp 1586364061
transform 1 0 24012 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__B
timestamp 1586364061
transform 1 0 23644 0 -1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _236_
timestamp 1586364061
transform 1 0 24380 0 -1 32096
box -38 -48 866 592
use scs8hd_fill_2  FILLER_54_266
timestamp 1586364061
transform 1 0 25576 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_262
timestamp 1586364061
transform 1 0 25208 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25760 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25392 0 -1 32096
box -38 -48 222 592
use scs8hd_or4_4  _281_
timestamp 1586364061
transform 1 0 27692 0 -1 32096
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_0.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 32096
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_610
timestamp 1586364061
transform 1 0 26404 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__340__B
timestamp 1586364061
transform 1 0 27508 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26956 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_54_270
timestamp 1586364061
transform 1 0 25944 0 -1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_54_279
timestamp 1586364061
transform 1 0 26772 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_283
timestamp 1586364061
transform 1 0 27140 0 -1 32096
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29716 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__272__D
timestamp 1586364061
transform 1 0 28704 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__282__B
timestamp 1586364061
transform 1 0 30728 0 -1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_0_in_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29256 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_298
timestamp 1586364061
transform 1 0 28520 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_302
timestamp 1586364061
transform 1 0 28888 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_3  FILLER_54_308
timestamp 1586364061
transform 1 0 29440 0 -1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_54_320
timestamp 1586364061
transform 1 0 30544 0 -1 32096
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_0_in_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 32096
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_611
timestamp 1586364061
transform 1 0 32016 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__341__B
timestamp 1586364061
transform 1 0 31372 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_324
timestamp 1586364061
transform 1 0 30912 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_54_328
timestamp 1586364061
transform 1 0 31280 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_4  FILLER_54_331
timestamp 1586364061
transform 1 0 31556 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_54_335
timestamp 1586364061
transform 1 0 31924 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_348
timestamp 1586364061
transform 1 0 33120 0 -1 32096
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34408 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35420 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_360
timestamp 1586364061
transform 1 0 34224 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_371
timestamp 1586364061
transform 1 0 35236 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_375
timestamp 1586364061
transform 1 0 35604 0 -1 32096
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35972 0 -1 32096
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37904 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_612
timestamp 1586364061
transform 1 0 37628 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_8  FILLER_54_388
timestamp 1586364061
transform 1 0 36800 0 -1 32096
box -38 -48 774 592
use scs8hd_fill_1  FILLER_54_396
timestamp 1586364061
transform 1 0 37536 0 -1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_54_398
timestamp 1586364061
transform 1 0 37720 0 -1 32096
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39652 0 -1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38916 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_409
timestamp 1586364061
transform 1 0 38732 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_6  FILLER_54_413
timestamp 1586364061
transform 1 0 39100 0 -1 32096
box -38 -48 590 592
use scs8hd_decap_8  FILLER_54_422
timestamp 1586364061
transform 1 0 39928 0 -1 32096
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42228 0 -1 32096
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40664 0 -1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41676 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_54_439
timestamp 1586364061
transform 1 0 41492 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_443
timestamp 1586364061
transform 1 0 41860 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_8  FILLER_54_450
timestamp 1586364061
transform 1 0 42504 0 -1 32096
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 44988 0 -1 32096
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43424 0 -1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_613
timestamp 1586364061
transform 1 0 43240 0 -1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 44436 0 -1 32096
box -38 -48 222 592
use scs8hd_fill_1  FILLER_54_459
timestamp 1586364061
transform 1 0 43332 0 -1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_54_469
timestamp 1586364061
transform 1 0 44252 0 -1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_54_473
timestamp 1586364061
transform 1 0 44620 0 -1 32096
box -38 -48 406 592
use scs8hd_decap_12  FILLER_54_480
timestamp 1586364061
transform 1 0 45264 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_492
timestamp 1586364061
transform 1 0 46368 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_504
timestamp 1586364061
transform 1 0 47472 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 48852 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_15
timestamp 1586364061
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_27
timestamp 1586364061
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_39
timestamp 1586364061
transform 1 0 4692 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_55_51
timestamp 1586364061
transform 1 0 5796 0 1 32096
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_614
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_59
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_62
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_74
timestamp 1586364061
transform 1 0 7912 0 1 32096
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10580 0 1 32096
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10028 0 1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_55_86
timestamp 1586364061
transform 1 0 9016 0 1 32096
box -38 -48 774 592
use scs8hd_decap_3  FILLER_55_94
timestamp 1586364061
transform 1 0 9752 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_99
timestamp 1586364061
transform 1 0 10212 0 1 32096
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_615
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_114
timestamp 1586364061
transform 1 0 11592 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_118
timestamp 1586364061
transform 1 0 11960 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_132
timestamp 1586364061
transform 1 0 13248 0 1 32096
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14628 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15640 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_136
timestamp 1586364061
transform 1 0 13616 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_140
timestamp 1586364061
transform 1 0 13984 0 1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_55_144
timestamp 1586364061
transform 1 0 14352 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_156
timestamp 1586364061
transform 1 0 15456 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_160
timestamp 1586364061
transform 1 0 15824 0 1 32096
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 32096
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_616
timestamp 1586364061
transform 1 0 17940 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_175
timestamp 1586364061
transform 1 0 17204 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_179
timestamp 1586364061
transform 1 0 17572 0 1 32096
box -38 -48 222 592
use scs8hd_inv_8  _128_
timestamp 1586364061
transform 1 0 19596 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 19412 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__244__C
timestamp 1586364061
transform 1 0 20700 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__245__A
timestamp 1586364061
transform 1 0 19044 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_193
timestamp 1586364061
transform 1 0 18860 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_197
timestamp 1586364061
transform 1 0 19228 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_210
timestamp 1586364061
transform 1 0 20424 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_215
timestamp 1586364061
transform 1 0 20884 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__244__A
timestamp 1586364061
transform 1 0 21068 0 1 32096
box -38 -48 222 592
use scs8hd_or4_4  _244_
timestamp 1586364061
transform 1 0 21252 0 1 32096
box -38 -48 866 592
use scs8hd_fill_2  FILLER_55_232
timestamp 1586364061
transform 1 0 22448 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_228
timestamp 1586364061
transform 1 0 22080 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__B
timestamp 1586364061
transform 1 0 22632 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 22264 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_240
timestamp 1586364061
transform 1 0 23184 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_236
timestamp 1586364061
transform 1 0 22816 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 32096
box -38 -48 222 592
use scs8hd_or4_4  _235_
timestamp 1586364061
transform 1 0 23644 0 1 32096
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 25208 0 1 32096
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_617
timestamp 1586364061
transform 1 0 23552 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 23368 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 25024 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__D
timestamp 1586364061
transform 1 0 24656 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_254
timestamp 1586364061
transform 1 0 24472 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_258
timestamp 1586364061
transform 1 0 24840 0 1 32096
box -38 -48 222 592
use scs8hd_or4_4  _263_
timestamp 1586364061
transform 1 0 27600 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__263__A
timestamp 1586364061
transform 1 0 27416 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__263__D
timestamp 1586364061
transform 1 0 27048 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__263__C
timestamp 1586364061
transform 1 0 26680 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_273
timestamp 1586364061
transform 1 0 26220 0 1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_55_277
timestamp 1586364061
transform 1 0 26588 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_280
timestamp 1586364061
transform 1 0 26864 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_284
timestamp 1586364061
transform 1 0 27232 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_301
timestamp 1586364061
transform 1 0 28796 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_297
timestamp 1586364061
transform 1 0 28428 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__272__B
timestamp 1586364061
transform 1 0 28980 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__272__A
timestamp 1586364061
transform 1 0 28612 0 1 32096
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_618
timestamp 1586364061
transform 1 0 29164 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_310
timestamp 1586364061
transform 1 0 29624 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_306
timestamp 1586364061
transform 1 0 29256 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__272__C
timestamp 1586364061
transform 1 0 29440 0 1 32096
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29808 0 1 32096
box -38 -48 866 592
use scs8hd_fill_2  FILLER_55_321
timestamp 1586364061
transform 1 0 30636 0 1 32096
box -38 -48 222 592
use scs8hd_nor2_4  _341_
timestamp 1586364061
transform 1 0 31372 0 1 32096
box -38 -48 866 592
use scs8hd_conb_1  _434_
timestamp 1586364061
transform 1 0 32936 0 1 32096
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__282__A
timestamp 1586364061
transform 1 0 30820 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__341__A
timestamp 1586364061
transform 1 0 31188 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__343__A
timestamp 1586364061
transform 1 0 32384 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__343__B
timestamp 1586364061
transform 1 0 32752 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_325
timestamp 1586364061
transform 1 0 31004 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_338
timestamp 1586364061
transform 1 0 32200 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_342
timestamp 1586364061
transform 1 0 32568 0 1 32096
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 32096
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_619
timestamp 1586364061
transform 1 0 34776 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34132 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 32096
box -38 -48 222 592
use scs8hd_decap_8  FILLER_55_349
timestamp 1586364061
transform 1 0 33212 0 1 32096
box -38 -48 774 592
use scs8hd_fill_2  FILLER_55_357
timestamp 1586364061
transform 1 0 33948 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_361
timestamp 1586364061
transform 1 0 34316 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_382
timestamp 1586364061
transform 1 0 36248 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_376
timestamp 1586364061
transform 1 0 35696 0 1 32096
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__268__A
timestamp 1586364061
transform 1 0 36064 0 1 32096
box -38 -48 222 592
use scs8hd_decap_6  FILLER_55_386
timestamp 1586364061
transform 1 0 36616 0 1 32096
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__268__B
timestamp 1586364061
transform 1 0 36432 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37168 0 1 32096
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37352 0 1 32096
box -38 -48 314 592
use scs8hd_fill_2  FILLER_55_401
timestamp 1586364061
transform 1 0 37996 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_397
timestamp 1586364061
transform 1 0 37628 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 37812 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38180 0 1 32096
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38364 0 1 32096
box -38 -48 866 592
use scs8hd_fill_2  FILLER_55_422
timestamp 1586364061
transform 1 0 39928 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_418
timestamp 1586364061
transform 1 0 39560 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_414
timestamp 1586364061
transform 1 0 39192 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 39376 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 39744 0 1 32096
box -38 -48 222 592
use scs8hd_decap_3  FILLER_55_428
timestamp 1586364061
transform 1 0 40480 0 1 32096
box -38 -48 314 592
use scs8hd_fill_1  FILLER_55_426
timestamp 1586364061
transform 1 0 40296 0 1 32096
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40112 0 1 32096
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_620
timestamp 1586364061
transform 1 0 40388 0 1 32096
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42688 0 1 32096
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40940 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40756 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41952 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 42504 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_442
timestamp 1586364061
transform 1 0 41768 0 1 32096
box -38 -48 222 592
use scs8hd_decap_4  FILLER_55_446
timestamp 1586364061
transform 1 0 42136 0 1 32096
box -38 -48 406 592
use scs8hd_fill_2  FILLER_55_455
timestamp 1586364061
transform 1 0 42964 0 1 32096
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43700 0 1 32096
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43148 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 43516 0 1 32096
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 44712 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_459
timestamp 1586364061
transform 1 0 43332 0 1 32096
box -38 -48 222 592
use scs8hd_fill_2  FILLER_55_472
timestamp 1586364061
transform 1 0 44528 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_476
timestamp 1586364061
transform 1 0 44896 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_621
timestamp 1586364061
transform 1 0 46000 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_489
timestamp 1586364061
transform 1 0 46092 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_501
timestamp 1586364061
transform 1 0 47196 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 48852 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_55_513
timestamp 1586364061
transform 1 0 48300 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_15
timestamp 1586364061
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_622
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_56_27
timestamp 1586364061
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_12  FILLER_56_32
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_44
timestamp 1586364061
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_56
timestamp 1586364061
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_68
timestamp 1586364061
transform 1 0 7360 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_80
timestamp 1586364061
transform 1 0 8464 0 -1 33184
box -38 -48 1142 592
use scs8hd_conb_1  _447_
timestamp 1586364061
transform 1 0 10120 0 -1 33184
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_623
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__225__B
timestamp 1586364061
transform 1 0 10580 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_56_93
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_56_97
timestamp 1586364061
transform 1 0 10028 0 -1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_56_101
timestamp 1586364061
transform 1 0 10396 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_56_105
timestamp 1586364061
transform 1 0 10764 0 -1 33184
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11132 0 -1 33184
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_56_120
timestamp 1586364061
transform 1 0 12144 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_8  FILLER_56_125
timestamp 1586364061
transform 1 0 12604 0 -1 33184
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 33184
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_624
timestamp 1586364061
transform 1 0 15180 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_56_142
timestamp 1586364061
transform 1 0 14168 0 -1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_56_146
timestamp 1586364061
transform 1 0 14536 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_56_149
timestamp 1586364061
transform 1 0 14812 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_12  FILLER_56_157
timestamp 1586364061
transform 1 0 15548 0 -1 33184
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 16744 0 -1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__248__A
timestamp 1586364061
transform 1 0 18308 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17940 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_56_169
timestamp 1586364061
transform 1 0 16652 0 -1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_56_181
timestamp 1586364061
transform 1 0 17756 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_185
timestamp 1586364061
transform 1 0 18124 0 -1 33184
box -38 -48 222 592
use scs8hd_nor2_4  _245_
timestamp 1586364061
transform 1 0 18952 0 -1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_625
timestamp 1586364061
transform 1 0 20792 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__245__B
timestamp 1586364061
transform 1 0 18768 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_56_189
timestamp 1586364061
transform 1 0 18492 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_8  FILLER_56_203
timestamp 1586364061
transform 1 0 19780 0 -1 33184
box -38 -48 774 592
use scs8hd_decap_3  FILLER_56_211
timestamp 1586364061
transform 1 0 20516 0 -1 33184
box -38 -48 314 592
use scs8hd_nor2_4  _239_
timestamp 1586364061
transform 1 0 21896 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__244__B
timestamp 1586364061
transform 1 0 21252 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_56_215
timestamp 1586364061
transform 1 0 20884 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_4  FILLER_56_221
timestamp 1586364061
transform 1 0 21436 0 -1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_56_225
timestamp 1586364061
transform 1 0 21804 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_8  FILLER_56_235
timestamp 1586364061
transform 1 0 22724 0 -1 33184
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 23460 0 -1 33184
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 -1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__241__B
timestamp 1586364061
transform 1 0 24840 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25668 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_56_254
timestamp 1586364061
transform 1 0 24472 0 -1 33184
box -38 -48 406 592
use scs8hd_fill_2  FILLER_56_260
timestamp 1586364061
transform 1 0 25024 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_265
timestamp 1586364061
transform 1 0 25484 0 -1 33184
box -38 -48 222 592
use scs8hd_or4_4  _272_
timestamp 1586364061
transform 1 0 28060 0 -1 33184
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_626
timestamp 1586364061
transform 1 0 26404 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__263__B
timestamp 1586364061
transform 1 0 27600 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26036 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_269
timestamp 1586364061
transform 1 0 25852 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_273
timestamp 1586364061
transform 1 0 26220 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_56_285
timestamp 1586364061
transform 1 0 27324 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_56_290
timestamp 1586364061
transform 1 0 27784 0 -1 33184
box -38 -48 314 592
use scs8hd_nor2_4  _282_
timestamp 1586364061
transform 1 0 30176 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__285__B
timestamp 1586364061
transform 1 0 29256 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29808 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_56_302
timestamp 1586364061
transform 1 0 28888 0 -1 33184
box -38 -48 406 592
use scs8hd_decap_4  FILLER_56_308
timestamp 1586364061
transform 1 0 29440 0 -1 33184
box -38 -48 406 592
use scs8hd_fill_2  FILLER_56_314
timestamp 1586364061
transform 1 0 29992 0 -1 33184
box -38 -48 222 592
use scs8hd_nor2_4  _343_
timestamp 1586364061
transform 1 0 32108 0 -1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_627
timestamp 1586364061
transform 1 0 32016 0 -1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 31188 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31556 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33120 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_325
timestamp 1586364061
transform 1 0 31004 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_329
timestamp 1586364061
transform 1 0 31372 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_56_333
timestamp 1586364061
transform 1 0 31740 0 -1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_56_346
timestamp 1586364061
transform 1 0 32936 0 -1 33184
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34132 0 -1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34868 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_56_350
timestamp 1586364061
transform 1 0 33304 0 -1 33184
box -38 -48 774 592
use scs8hd_fill_1  FILLER_56_358
timestamp 1586364061
transform 1 0 34040 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_4  FILLER_56_362
timestamp 1586364061
transform 1 0 34408 0 -1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_56_366
timestamp 1586364061
transform 1 0 34776 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_8  FILLER_56_369
timestamp 1586364061
transform 1 0 35052 0 -1 33184
box -38 -48 774 592
use scs8hd_nor2_4  _268_
timestamp 1586364061
transform 1 0 36064 0 -1 33184
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 37720 0 -1 33184
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_628
timestamp 1586364061
transform 1 0 37628 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_3  FILLER_56_377
timestamp 1586364061
transform 1 0 35788 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_8  FILLER_56_389
timestamp 1586364061
transform 1 0 36892 0 -1 33184
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 39744 0 -1 33184
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__270__B
timestamp 1586364061
transform 1 0 39008 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_56_409
timestamp 1586364061
transform 1 0 38732 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_6  FILLER_56_414
timestamp 1586364061
transform 1 0 39192 0 -1 33184
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41492 0 -1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40940 0 -1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41308 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_431
timestamp 1586364061
transform 1 0 40756 0 -1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_56_435
timestamp 1586364061
transform 1 0 41124 0 -1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_56_448
timestamp 1586364061
transform 1 0 42320 0 -1 33184
box -38 -48 774 592
use scs8hd_fill_2  FILLER_56_456
timestamp 1586364061
transform 1 0 43056 0 -1 33184
box -38 -48 222 592
use scs8hd_conb_1  _442_
timestamp 1586364061
transform 1 0 45080 0 -1 33184
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 43332 0 -1 33184
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_629
timestamp 1586364061
transform 1 0 43240 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_8  FILLER_56_470
timestamp 1586364061
transform 1 0 44344 0 -1 33184
box -38 -48 774 592
use scs8hd_decap_12  FILLER_56_481
timestamp 1586364061
transform 1 0 45356 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_493
timestamp 1586364061
transform 1 0 46460 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_56_505
timestamp 1586364061
transform 1 0 47564 0 -1 33184
box -38 -48 774 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 48852 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_56_513
timestamp 1586364061
transform 1 0 48300 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_15
timestamp 1586364061
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_27
timestamp 1586364061
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_39
timestamp 1586364061
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_57_51
timestamp 1586364061
transform 1 0 5796 0 1 33184
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_630
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_57_59
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_57_62
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_74
timestamp 1586364061
transform 1 0 7912 0 1 33184
box -38 -48 1142 592
use scs8hd_nor2_4  _225_
timestamp 1586364061
transform 1 0 10580 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__225__A
timestamp 1586364061
transform 1 0 10396 0 1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_57_86
timestamp 1586364061
transform 1 0 9016 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_57_98
timestamp 1586364061
transform 1 0 10120 0 1 33184
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_631
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11868 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_112
timestamp 1586364061
transform 1 0 11408 0 1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_57_116
timestamp 1586364061
transform 1 0 11776 0 1 33184
box -38 -48 130 592
use scs8hd_decap_3  FILLER_57_119
timestamp 1586364061
transform 1 0 12052 0 1 33184
box -38 -48 314 592
use scs8hd_decap_4  FILLER_57_132
timestamp 1586364061
transform 1 0 13248 0 1 33184
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14628 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 13616 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__230__B
timestamp 1586364061
transform 1 0 13984 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_138
timestamp 1586364061
transform 1 0 13800 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_57_142
timestamp 1586364061
transform 1 0 14168 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_156
timestamp 1586364061
transform 1 0 15456 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_160
timestamp 1586364061
transform 1 0 15824 0 1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_57_164
timestamp 1586364061
transform 1 0 16192 0 1 33184
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16008 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_179
timestamp 1586364061
transform 1 0 17572 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_175
timestamp 1586364061
transform 1 0 17204 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 33184
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_57_184
timestamp 1586364061
transform 1 0 18032 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 33184
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_632
timestamp 1586364061
transform 1 0 17940 0 1 33184
box -38 -48 130 592
use scs8hd_nor2_4  _248_
timestamp 1586364061
transform 1 0 18308 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 19320 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__250__A
timestamp 1586364061
transform 1 0 20700 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__250__B
timestamp 1586364061
transform 1 0 20332 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19688 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_196
timestamp 1586364061
transform 1 0 19136 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_200
timestamp 1586364061
transform 1 0 19504 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_204
timestamp 1586364061
transform 1 0 19872 0 1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_57_208
timestamp 1586364061
transform 1 0 20240 0 1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_57_211
timestamp 1586364061
transform 1 0 20516 0 1 33184
box -38 -48 222 592
use scs8hd_nor2_4  _250_
timestamp 1586364061
transform 1 0 20884 0 1 33184
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22908 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 21896 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22264 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_224
timestamp 1586364061
transform 1 0 21712 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_228
timestamp 1586364061
transform 1 0 22080 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_235
timestamp 1586364061
transform 1 0 22724 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_239
timestamp 1586364061
transform 1 0 23092 0 1 33184
box -38 -48 406 592
use scs8hd_fill_2  FILLER_57_250
timestamp 1586364061
transform 1 0 24104 0 1 33184
box -38 -48 222 592
use scs8hd_decap_3  FILLER_57_245
timestamp 1586364061
transform 1 0 23644 0 1 33184
box -38 -48 314 592
use scs8hd_fill_1  FILLER_57_243
timestamp 1586364061
transform 1 0 23460 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23920 0 1 33184
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_633
timestamp 1586364061
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24288 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24472 0 1 33184
box -38 -48 866 592
use scs8hd_fill_2  FILLER_57_267
timestamp 1586364061
transform 1 0 25668 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_263
timestamp 1586364061
transform 1 0 25300 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 25484 0 1 33184
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 26036 0 1 33184
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27784 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28244 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 25852 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27232 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27600 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_282
timestamp 1586364061
transform 1 0 27048 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_286
timestamp 1586364061
transform 1 0 27416 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_293
timestamp 1586364061
transform 1 0 28060 0 1 33184
box -38 -48 222 592
use scs8hd_nor2_4  _285_
timestamp 1586364061
transform 1 0 29256 0 1 33184
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_634
timestamp 1586364061
transform 1 0 29164 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 30268 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__285__A
timestamp 1586364061
transform 1 0 28980 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28612 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_297
timestamp 1586364061
transform 1 0 28428 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_301
timestamp 1586364061
transform 1 0 28796 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_315
timestamp 1586364061
transform 1 0 30084 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_319
timestamp 1586364061
transform 1 0 30452 0 1 33184
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 31096 0 1 33184
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32844 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 30912 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 32292 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32660 0 1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_57_323
timestamp 1586364061
transform 1 0 30820 0 1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_57_337
timestamp 1586364061
transform 1 0 32108 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_341
timestamp 1586364061
transform 1 0 32476 0 1 33184
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_635
timestamp 1586364061
transform 1 0 34776 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 35512 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33856 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_354
timestamp 1586364061
transform 1 0 33672 0 1 33184
box -38 -48 222 592
use scs8hd_decap_8  FILLER_57_358
timestamp 1586364061
transform 1 0 34040 0 1 33184
box -38 -48 774 592
use scs8hd_decap_6  FILLER_57_367
timestamp 1586364061
transform 1 0 34868 0 1 33184
box -38 -48 590 592
use scs8hd_fill_1  FILLER_57_373
timestamp 1586364061
transform 1 0 35420 0 1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_57_384
timestamp 1586364061
transform 1 0 36432 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_380
timestamp 1586364061
transform 1 0 36064 0 1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_57_376
timestamp 1586364061
transform 1 0 35696 0 1 33184
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36248 0 1 33184
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35788 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_395
timestamp 1586364061
transform 1 0 37444 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_391
timestamp 1586364061
transform 1 0 37076 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36616 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37260 0 1 33184
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36800 0 1 33184
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37628 0 1 33184
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37812 0 1 33184
box -38 -48 866 592
use scs8hd_fill_2  FILLER_57_408
timestamp 1586364061
transform 1 0 38640 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38824 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_412
timestamp 1586364061
transform 1 0 39008 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__270__A
timestamp 1586364061
transform 1 0 39192 0 1 33184
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39376 0 1 33184
box -38 -48 314 592
use scs8hd_fill_2  FILLER_57_419
timestamp 1586364061
transform 1 0 39652 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39836 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_423
timestamp 1586364061
transform 1 0 40020 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40204 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_428
timestamp 1586364061
transform 1 0 40480 0 1 33184
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_636
timestamp 1586364061
transform 1 0 40388 0 1 33184
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42228 0 1 33184
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40664 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__269__A
timestamp 1586364061
transform 1 0 41676 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__269__B
timestamp 1586364061
transform 1 0 42044 0 1 33184
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42688 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_439
timestamp 1586364061
transform 1 0 41492 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_443
timestamp 1586364061
transform 1 0 41860 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_450
timestamp 1586364061
transform 1 0 42504 0 1 33184
box -38 -48 222 592
use scs8hd_decap_4  FILLER_57_454
timestamp 1586364061
transform 1 0 42872 0 1 33184
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 43516 0 1 33184
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 43332 0 1 33184
box -38 -48 222 592
use scs8hd_fill_1  FILLER_57_458
timestamp 1586364061
transform 1 0 43240 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_470
timestamp 1586364061
transform 1 0 44344 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_57_482
timestamp 1586364061
transform 1 0 45448 0 1 33184
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_637
timestamp 1586364061
transform 1 0 46000 0 1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_57_489
timestamp 1586364061
transform 1 0 46092 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_501
timestamp 1586364061
transform 1 0 47196 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 48852 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_57_513
timestamp 1586364061
transform 1 0 48300 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_638
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_44
timestamp 1586364061
transform 1 0 5152 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_56
timestamp 1586364061
transform 1 0 6256 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_68
timestamp 1586364061
transform 1 0 7360 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_80
timestamp 1586364061
transform 1 0 8464 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_639
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__227__B
timestamp 1586364061
transform 1 0 10580 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10948 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_58_93
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 774 592
use scs8hd_fill_2  FILLER_58_101
timestamp 1586364061
transform 1 0 10396 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_105
timestamp 1586364061
transform 1 0 10764 0 -1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11868 0 -1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_58_109
timestamp 1586364061
transform 1 0 11132 0 -1 34272
box -38 -48 774 592
use scs8hd_decap_3  FILLER_58_120
timestamp 1586364061
transform 1 0 12144 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_8  FILLER_58_125
timestamp 1586364061
transform 1 0 12604 0 -1 34272
box -38 -48 774 592
use scs8hd_decap_3  FILLER_58_133
timestamp 1586364061
transform 1 0 13340 0 -1 34272
box -38 -48 314 592
use scs8hd_nor2_4  _230_
timestamp 1586364061
transform 1 0 13616 0 -1 34272
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 34272
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_640
timestamp 1586364061
transform 1 0 15180 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_145
timestamp 1586364061
transform 1 0 14444 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_149
timestamp 1586364061
transform 1 0 14812 0 -1 34272
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17848 0 -1 34272
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__248__B
timestamp 1586364061
transform 1 0 18308 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_163
timestamp 1586364061
transform 1 0 16100 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_167
timestamp 1586364061
transform 1 0 16468 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_58_174
timestamp 1586364061
transform 1 0 17112 0 -1 34272
box -38 -48 774 592
use scs8hd_fill_2  FILLER_58_185
timestamp 1586364061
transform 1 0 18124 0 -1 34272
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18860 0 -1 34272
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_641
timestamp 1586364061
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20056 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_189
timestamp 1586364061
transform 1 0 18492 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_58_204
timestamp 1586364061
transform 1 0 19872 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_58_208
timestamp 1586364061
transform 1 0 20240 0 -1 34272
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 21436 0 -1 34272
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22632 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21068 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_215
timestamp 1586364061
transform 1 0 20884 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_219
timestamp 1586364061
transform 1 0 21252 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_232
timestamp 1586364061
transform 1 0 22448 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_58_236
timestamp 1586364061
transform 1 0 22816 0 -1 34272
box -38 -48 774 592
use scs8hd_nor2_4  _241_
timestamp 1586364061
transform 1 0 24840 0 -1 34272
box -38 -48 866 592
use scs8hd_conb_1  _445_
timestamp 1586364061
transform 1 0 23828 0 -1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24288 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_58_244
timestamp 1586364061
transform 1 0 23552 0 -1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_58_250
timestamp 1586364061
transform 1 0 24104 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_254
timestamp 1586364061
transform 1 0 24472 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_8  FILLER_58_267
timestamp 1586364061
transform 1 0 25668 0 -1 34272
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27140 0 -1 34272
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_642
timestamp 1586364061
transform 1 0 26404 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26956 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_276
timestamp 1586364061
transform 1 0 26496 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_58_280
timestamp 1586364061
transform 1 0 26864 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_292
timestamp 1586364061
transform 1 0 27968 0 -1 34272
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 29440 0 -1 34272
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__287__B
timestamp 1586364061
transform 1 0 30636 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_304
timestamp 1586364061
transform 1 0 29072 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_58_319
timestamp 1586364061
transform 1 0 30452 0 -1 34272
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 34272
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_643
timestamp 1586364061
transform 1 0 32016 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31004 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_323
timestamp 1586364061
transform 1 0 30820 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_58_327
timestamp 1586364061
transform 1 0 31188 0 -1 34272
box -38 -48 774 592
use scs8hd_fill_1  FILLER_58_335
timestamp 1586364061
transform 1 0 31924 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_58_348
timestamp 1586364061
transform 1 0 33120 0 -1 34272
box -38 -48 774 592
use scs8hd_conb_1  _440_
timestamp 1586364061
transform 1 0 33856 0 -1 34272
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 35512 0 -1 34272
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__276__B
timestamp 1586364061
transform 1 0 34960 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__275__B
timestamp 1586364061
transform 1 0 34500 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_359
timestamp 1586364061
transform 1 0 34132 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_3  FILLER_58_365
timestamp 1586364061
transform 1 0 34684 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_4  FILLER_58_370
timestamp 1586364061
transform 1 0 35144 0 -1 34272
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37996 0 -1 34272
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_644
timestamp 1586364061
transform 1 0 37628 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__273__B
timestamp 1586364061
transform 1 0 36708 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37076 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_385
timestamp 1586364061
transform 1 0 36524 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_389
timestamp 1586364061
transform 1 0 36892 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_393
timestamp 1586364061
transform 1 0 37260 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_3  FILLER_58_398
timestamp 1586364061
transform 1 0 37720 0 -1 34272
box -38 -48 314 592
use scs8hd_nor2_4  _270_
timestamp 1586364061
transform 1 0 39008 0 -1 34272
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40572 0 -1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__278__B
timestamp 1586364061
transform 1 0 38824 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 40388 0 -1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38456 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_404
timestamp 1586364061
transform 1 0 38272 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_408
timestamp 1586364061
transform 1 0 38640 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_58_421
timestamp 1586364061
transform 1 0 39836 0 -1 34272
box -38 -48 590 592
use scs8hd_nor2_4  _269_
timestamp 1586364061
transform 1 0 41676 0 -1 34272
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41308 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_58_432
timestamp 1586364061
transform 1 0 40848 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_58_436
timestamp 1586364061
transform 1 0 41216 0 -1 34272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_58_439
timestamp 1586364061
transform 1 0 41492 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_58_450
timestamp 1586364061
transform 1 0 42504 0 -1 34272
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_645
timestamp 1586364061
transform 1 0 43240 0 -1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 43516 0 -1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_58_459
timestamp 1586364061
transform 1 0 43332 0 -1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_58_463
timestamp 1586364061
transform 1 0 43700 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_475
timestamp 1586364061
transform 1 0 44804 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_487
timestamp 1586364061
transform 1 0 45908 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_499
timestamp 1586364061
transform 1 0 47012 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 48852 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_4  FILLER_58_511
timestamp 1586364061
transform 1 0 48116 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_58_515
timestamp 1586364061
transform 1 0 48484 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_59_3
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_15
timestamp 1586364061
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_15
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_654
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_27
timestamp 1586364061
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_39
timestamp 1586364061
transform 1 0 4692 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_59_51
timestamp 1586364061
transform 1 0 5796 0 1 34272
box -38 -48 774 592
use scs8hd_decap_4  FILLER_60_27
timestamp 1586364061
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_12  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_44
timestamp 1586364061
transform 1 0 5152 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_646
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_59
timestamp 1586364061
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_62
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_74
timestamp 1586364061
transform 1 0 7912 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_56
timestamp 1586364061
transform 1 0 6256 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_68
timestamp 1586364061
transform 1 0 7360 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_80
timestamp 1586364061
transform 1 0 8464 0 -1 35360
box -38 -48 1142 592
use scs8hd_nor2_4  _227_
timestamp 1586364061
transform 1 0 10580 0 1 34272
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10856 0 -1 35360
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_655
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 10396 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__B
timestamp 1586364061
transform 1 0 10396 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_86
timestamp 1586364061
transform 1 0 9016 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_59_98
timestamp 1586364061
transform 1 0 10120 0 1 34272
box -38 -48 314 592
use scs8hd_decap_8  FILLER_60_93
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_3  FILLER_60_103
timestamp 1586364061
transform 1 0 10580 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_60_117
timestamp 1586364061
transform 1 0 11868 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_116
timestamp 1586364061
transform 1 0 11776 0 1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_112
timestamp 1586364061
transform 1 0 11408 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11592 0 1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 1 34272
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_647
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12144 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_59_123
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_60_121
timestamp 1586364061
transform 1 0 12236 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_127
timestamp 1586364061
transform 1 0 12788 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_131
timestamp 1586364061
transform 1 0 13156 0 1 34272
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch
timestamp 1586364061
transform 1 0 12604 0 -1 35360
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 13340 0 1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13524 0 1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_138
timestamp 1586364061
transform 1 0 13800 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14260 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_142
timestamp 1586364061
transform 1 0 14168 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_60_142
timestamp 1586364061
transform 1 0 14168 0 -1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_60_145
timestamp 1586364061
transform 1 0 14444 0 -1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14536 0 1 34272
box -38 -48 866 592
use scs8hd_decap_6  FILLER_60_136
timestamp 1586364061
transform 1 0 13616 0 -1 35360
box -38 -48 590 592
use scs8hd_decap_3  FILLER_60_154
timestamp 1586364061
transform 1 0 15272 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_4  FILLER_60_149
timestamp 1586364061
transform 1 0 14812 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_155
timestamp 1586364061
transform 1 0 15364 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15548 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_656
timestamp 1586364061
transform 1 0 15180 0 -1 35360
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15548 0 -1 35360
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_59_159
timestamp 1586364061
transform 1 0 15732 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15916 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_60_168
timestamp 1586364061
transform 1 0 16560 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 -1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 1 34272
box -38 -48 866 592
use scs8hd_decap_4  FILLER_60_172
timestamp 1586364061
transform 1 0 16928 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_178
timestamp 1586364061
transform 1 0 17480 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_172
timestamp 1586364061
transform 1 0 16928 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__229__B
timestamp 1586364061
transform 1 0 17664 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 17296 0 1 34272
box -38 -48 222 592
use scs8hd_nor2_4  _229_
timestamp 1586364061
transform 1 0 17296 0 -1 35360
box -38 -48 866 592
use scs8hd_decap_8  FILLER_60_185
timestamp 1586364061
transform 1 0 18124 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_59_187
timestamp 1586364061
transform 1 0 18308 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_59_182
timestamp 1586364061
transform 1 0 17848 0 1 34272
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_648
timestamp 1586364061
transform 1 0 17940 0 1 34272
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_60_193
timestamp 1586364061
transform 1 0 18860 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_197
timestamp 1586364061
transform 1 0 19228 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_191
timestamp 1586364061
transform 1 0 18676 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_3.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 19412 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 35360
box -38 -48 866 592
use scs8hd_decap_8  FILLER_60_206
timestamp 1586364061
transform 1 0 20056 0 -1 35360
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_7_.latch
timestamp 1586364061
transform 1 0 19596 0 1 34272
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_59_212
timestamp 1586364061
transform 1 0 20608 0 1 34272
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_657
timestamp 1586364061
transform 1 0 20792 0 -1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_60_224
timestamp 1586364061
transform 1 0 21712 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_222
timestamp 1586364061
transform 1 0 21528 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_59_217
timestamp 1586364061
transform 1 0 21068 0 1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 35360
box -38 -48 866 592
use scs8hd_decap_4  FILLER_60_228
timestamp 1586364061
transform 1 0 22080 0 -1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22448 0 -1 35360
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21896 0 1 34272
box -38 -48 866 592
use scs8hd_decap_4  FILLER_60_241
timestamp 1586364061
transform 1 0 23276 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_3  FILLER_59_239
timestamp 1586364061
transform 1 0 23092 0 1 34272
box -38 -48 314 592
use scs8hd_fill_2  FILLER_59_235
timestamp 1586364061
transform 1 0 22724 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22908 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_60_248
timestamp 1586364061
transform 1 0 23920 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_60_245
timestamp 1586364061
transform 1 0 23644 0 -1 35360
box -38 -48 130 592
use scs8hd_fill_1  FILLER_59_245
timestamp 1586364061
transform 1 0 23644 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__238__B
timestamp 1586364061
transform 1 0 23736 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 23368 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_649
timestamp 1586364061
transform 1 0 23552 0 1 34272
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 24288 0 -1 35360
box -38 -48 1050 592
use scs8hd_nor2_4  _238_
timestamp 1586364061
transform 1 0 23736 0 1 34272
box -38 -48 866 592
use scs8hd_fill_2  FILLER_60_263
timestamp 1586364061
transform 1 0 25300 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_259
timestamp 1586364061
transform 1 0 24932 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_255
timestamp 1586364061
transform 1 0 24564 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25484 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25116 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 24748 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25300 0 1 34272
box -38 -48 866 592
use scs8hd_decap_4  FILLER_60_267
timestamp 1586364061
transform 1 0 25668 0 -1 35360
box -38 -48 406 592
use scs8hd_decap_6  FILLER_60_276
timestamp 1586364061
transform 1 0 26496 0 -1 35360
box -38 -48 590 592
use scs8hd_fill_2  FILLER_60_273
timestamp 1586364061
transform 1 0 26220 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_1  FILLER_59_276
timestamp 1586364061
transform 1 0 26496 0 1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_59_272
timestamp 1586364061
transform 1 0 26128 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26036 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26588 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_658
timestamp 1586364061
transform 1 0 26404 0 -1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_279
timestamp 1586364061
transform 1 0 26772 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26956 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27140 0 1 34272
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27048 0 -1 35360
box -38 -48 866 592
use scs8hd_decap_6  FILLER_60_295
timestamp 1586364061
transform 1 0 28244 0 -1 35360
box -38 -48 590 592
use scs8hd_fill_2  FILLER_60_291
timestamp 1586364061
transform 1 0 27876 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_292
timestamp 1586364061
transform 1 0 27968 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28060 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28152 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_60_301
timestamp 1586364061
transform 1 0 28796 0 -1 35360
box -38 -48 130 592
use scs8hd_fill_1  FILLER_59_304
timestamp 1586364061
transform 1 0 29072 0 1 34272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_300
timestamp 1586364061
transform 1 0 28704 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_296
timestamp 1586364061
transform 1 0 28336 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__284__B
timestamp 1586364061
transform 1 0 28520 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__284__A
timestamp 1586364061
transform 1 0 28888 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_650
timestamp 1586364061
transform 1 0 29164 0 1 34272
box -38 -48 130 592
use scs8hd_nor2_4  _284_
timestamp 1586364061
transform 1 0 28888 0 -1 35360
box -38 -48 866 592
use scs8hd_decap_8  FILLER_60_311
timestamp 1586364061
transform 1 0 29716 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_4  FILLER_59_313
timestamp 1586364061
transform 1 0 29900 0 1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_309
timestamp 1586364061
transform 1 0 29532 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29716 0 1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 34272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_59_317
timestamp 1586364061
transform 1 0 30268 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__287__A
timestamp 1586364061
transform 1 0 30360 0 1 34272
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30544 0 1 34272
box -38 -48 866 592
use scs8hd_nor2_4  _287_
timestamp 1586364061
transform 1 0 30452 0 -1 35360
box -38 -48 866 592
use scs8hd_decap_8  FILLER_60_328
timestamp 1586364061
transform 1 0 31280 0 -1 35360
box -38 -48 774 592
use scs8hd_fill_2  FILLER_59_329
timestamp 1586364061
transform 1 0 31372 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31556 0 1 34272
box -38 -48 222 592
use scs8hd_decap_3  FILLER_60_341
timestamp 1586364061
transform 1 0 32476 0 -1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_60_337
timestamp 1586364061
transform 1 0 32108 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_333
timestamp 1586364061
transform 1 0 31740 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32292 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32108 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_659
timestamp 1586364061
transform 1 0 32016 0 -1 35360
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32292 0 1 34272
box -38 -48 866 592
use scs8hd_fill_2  FILLER_59_348
timestamp 1586364061
transform 1 0 33120 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32752 0 -1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32936 0 -1 35360
box -38 -48 866 592
use scs8hd_decap_8  FILLER_60_355
timestamp 1586364061
transform 1 0 33764 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_4  FILLER_59_356
timestamp 1586364061
transform 1 0 33856 0 1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_352
timestamp 1586364061
transform 1 0 33488 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33672 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33304 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_59_367
timestamp 1586364061
transform 1 0 34868 0 1 34272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_362
timestamp 1586364061
transform 1 0 34408 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__275__A
timestamp 1586364061
transform 1 0 34224 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__276__A
timestamp 1586364061
transform 1 0 34592 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_651
timestamp 1586364061
transform 1 0 34776 0 1 34272
box -38 -48 130 592
use scs8hd_nor2_4  _276_
timestamp 1586364061
transform 1 0 34960 0 1 34272
box -38 -48 866 592
use scs8hd_nor2_4  _275_
timestamp 1586364061
transform 1 0 34500 0 -1 35360
box -38 -48 866 592
use scs8hd_decap_4  FILLER_60_372
timestamp 1586364061
transform 1 0 35328 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_60_379
timestamp 1586364061
transform 1 0 35972 0 -1 35360
box -38 -48 130 592
use scs8hd_fill_1  FILLER_60_376
timestamp 1586364061
transform 1 0 35696 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_3  FILLER_59_382
timestamp 1586364061
transform 1 0 36248 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  FILLER_59_377
timestamp 1586364061
transform 1 0 35788 0 1 34272
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__273__A
timestamp 1586364061
transform 1 0 36064 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 35788 0 -1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36524 0 1 34272
box -38 -48 866 592
use scs8hd_nor2_4  _273_
timestamp 1586364061
transform 1 0 36064 0 -1 35360
box -38 -48 866 592
use scs8hd_fill_2  FILLER_60_393
timestamp 1586364061
transform 1 0 37260 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_60_389
timestamp 1586364061
transform 1 0 36892 0 -1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_394
timestamp 1586364061
transform 1 0 37352 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37444 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37076 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch_D
timestamp 1586364061
transform 1 0 37720 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_660
timestamp 1586364061
transform 1 0 37628 0 -1 35360
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch
timestamp 1586364061
transform 1 0 37720 0 -1 35360
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_59_400
timestamp 1586364061
transform 1 0 37904 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_7_.latch_SLEEPB
timestamp 1586364061
transform 1 0 38088 0 1 34272
box -38 -48 222 592
use scs8hd_decap_8  FILLER_60_409
timestamp 1586364061
transform 1 0 38732 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_4  FILLER_59_404
timestamp 1586364061
transform 1 0 38272 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__278__A
timestamp 1586364061
transform 1 0 38640 0 1 34272
box -38 -48 222 592
use scs8hd_nor2_4  _278_
timestamp 1586364061
transform 1 0 38824 0 1 34272
box -38 -48 866 592
use scs8hd_fill_1  FILLER_60_417
timestamp 1586364061
transform 1 0 39468 0 -1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_423
timestamp 1586364061
transform 1 0 40020 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_419
timestamp 1586364061
transform 1 0 39652 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40204 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 39836 0 1 34272
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 39560 0 -1 35360
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_60_429
timestamp 1586364061
transform 1 0 40572 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_428
timestamp 1586364061
transform 1 0 40480 0 1 34272
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_652
timestamp 1586364061
transform 1 0 40388 0 1 34272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_60_433
timestamp 1586364061
transform 1 0 40940 0 -1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_439
timestamp 1586364061
transform 1 0 41492 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_433
timestamp 1586364061
transform 1 0 40940 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41124 0 -1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41308 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40756 0 -1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41308 0 -1 35360
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41676 0 1 34272
box -38 -48 314 592
use scs8hd_conb_1  _441_
timestamp 1586364061
transform 1 0 40664 0 1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_60_446
timestamp 1586364061
transform 1 0 42136 0 -1 35360
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_59_455
timestamp 1586364061
transform 1 0 42964 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_448
timestamp 1586364061
transform 1 0 42320 0 1 34272
box -38 -48 406 592
use scs8hd_fill_2  FILLER_59_444
timestamp 1586364061
transform 1 0 41952 0 1 34272
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42136 0 1 34272
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 42688 0 1 34272
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_661
timestamp 1586364061
transform 1 0 43240 0 -1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 43148 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_459
timestamp 1586364061
transform 1 0 43332 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_471
timestamp 1586364061
transform 1 0 44436 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_59_483
timestamp 1586364061
transform 1 0 45540 0 1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_60_459
timestamp 1586364061
transform 1 0 43332 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_471
timestamp 1586364061
transform 1 0 44436 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_483
timestamp 1586364061
transform 1 0 45540 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_653
timestamp 1586364061
transform 1 0 46000 0 1 34272
box -38 -48 130 592
use scs8hd_fill_1  FILLER_59_487
timestamp 1586364061
transform 1 0 45908 0 1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_59_489
timestamp 1586364061
transform 1 0 46092 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_501
timestamp 1586364061
transform 1 0 47196 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_495
timestamp 1586364061
transform 1 0 46644 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_60_507
timestamp 1586364061
transform 1 0 47748 0 -1 35360
box -38 -48 774 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 48852 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 48852 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_59_513
timestamp 1586364061
transform 1 0 48300 0 1 34272
box -38 -48 314 592
use scs8hd_fill_1  FILLER_60_515
timestamp 1586364061
transform 1 0 48484 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_3
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_15
timestamp 1586364061
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_27
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_39
timestamp 1586364061
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_51
timestamp 1586364061
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_662
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_59
timestamp 1586364061
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_62
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_74
timestamp 1586364061
transform 1 0 7912 0 1 35360
box -38 -48 1142 592
use scs8hd_nor2_4  _228_
timestamp 1586364061
transform 1 0 10764 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 10396 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 10028 0 1 35360
box -38 -48 222 592
use scs8hd_decap_8  FILLER_61_86
timestamp 1586364061
transform 1 0 9016 0 1 35360
box -38 -48 774 592
use scs8hd_decap_3  FILLER_61_94
timestamp 1586364061
transform 1 0 9752 0 1 35360
box -38 -48 314 592
use scs8hd_fill_2  FILLER_61_99
timestamp 1586364061
transform 1 0 10212 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_103
timestamp 1586364061
transform 1 0 10580 0 1 35360
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch
timestamp 1586364061
transform 1 0 12512 0 1 35360
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_663
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__B
timestamp 1586364061
transform 1 0 11776 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_114
timestamp 1586364061
transform 1 0 11592 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_118
timestamp 1586364061
transform 1 0 11960 0 1 35360
box -38 -48 222 592
use scs8hd_fill_1  FILLER_61_123
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13708 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_135
timestamp 1586364061
transform 1 0 13524 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_139
timestamp 1586364061
transform 1 0 13892 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_152
timestamp 1586364061
transform 1 0 15088 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_156
timestamp 1586364061
transform 1 0 15456 0 1 35360
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 35360
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_664
timestamp 1586364061
transform 1 0 17940 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 16192 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18308 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_162
timestamp 1586364061
transform 1 0 16008 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_175
timestamp 1586364061
transform 1 0 17204 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_179
timestamp 1586364061
transform 1 0 17572 0 1 35360
box -38 -48 406 592
use scs8hd_decap_3  FILLER_61_184
timestamp 1586364061
transform 1 0 18032 0 1 35360
box -38 -48 314 592
use scs8hd_conb_1  _444_
timestamp 1586364061
transform 1 0 18492 0 1 35360
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19504 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 18952 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_192
timestamp 1586364061
transform 1 0 18768 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_196
timestamp 1586364061
transform 1 0 19136 0 1 35360
box -38 -48 222 592
use scs8hd_decap_6  FILLER_61_209
timestamp 1586364061
transform 1 0 20332 0 1 35360
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21804 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__237__B
timestamp 1586364061
transform 1 0 23000 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21620 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21252 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20884 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_217
timestamp 1586364061
transform 1 0 21068 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_221
timestamp 1586364061
transform 1 0 21436 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_234
timestamp 1586364061
transform 1 0 22632 0 1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_61_240
timestamp 1586364061
transform 1 0 23184 0 1 35360
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 24288 0 1 35360
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_665
timestamp 1586364061
transform 1 0 23552 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 24104 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25484 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 23368 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_245
timestamp 1586364061
transform 1 0 23644 0 1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_61_249
timestamp 1586364061
transform 1 0 24012 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_263
timestamp 1586364061
transform 1 0 25300 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_267
timestamp 1586364061
transform 1 0 25668 0 1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 1 35360
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26036 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27048 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__283__B
timestamp 1586364061
transform 1 0 27416 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25852 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_280
timestamp 1586364061
transform 1 0 26864 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_284
timestamp 1586364061
transform 1 0 27232 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_301
timestamp 1586364061
transform 1 0 28796 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_297
timestamp 1586364061
transform 1 0 28428 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28980 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__283__A
timestamp 1586364061
transform 1 0 28612 0 1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_666
timestamp 1586364061
transform 1 0 29164 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_313
timestamp 1586364061
transform 1 0 29900 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_309
timestamp 1586364061
transform 1 0 29532 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29716 0 1 35360
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_61_317
timestamp 1586364061
transform 1 0 30268 0 1 35360
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 30084 0 1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30544 0 1 35360
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32844 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32660 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32292 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31924 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31556 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_329
timestamp 1586364061
transform 1 0 31372 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_333
timestamp 1586364061
transform 1 0 31740 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_337
timestamp 1586364061
transform 1 0 32108 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_341
timestamp 1586364061
transform 1 0 32476 0 1 35360
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch
timestamp 1586364061
transform 1 0 35512 0 1 35360
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_667
timestamp 1586364061
transform 1 0 34776 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34316 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 35328 0 1 35360
box -38 -48 222 592
use scs8hd_decap_6  FILLER_61_354
timestamp 1586364061
transform 1 0 33672 0 1 35360
box -38 -48 590 592
use scs8hd_fill_1  FILLER_61_360
timestamp 1586364061
transform 1 0 34224 0 1 35360
box -38 -48 130 592
use scs8hd_decap_3  FILLER_61_363
timestamp 1586364061
transform 1 0 34500 0 1 35360
box -38 -48 314 592
use scs8hd_decap_4  FILLER_61_367
timestamp 1586364061
transform 1 0 34868 0 1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_61_371
timestamp 1586364061
transform 1 0 35236 0 1 35360
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38088 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37720 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36708 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37352 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_385
timestamp 1586364061
transform 1 0 36524 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_389
timestamp 1586364061
transform 1 0 36892 0 1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_61_393
timestamp 1586364061
transform 1 0 37260 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_396
timestamp 1586364061
transform 1 0 37536 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_400
timestamp 1586364061
transform 1 0 37904 0 1 35360
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_668
timestamp 1586364061
transform 1 0 40388 0 1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39652 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39100 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_411
timestamp 1586364061
transform 1 0 38916 0 1 35360
box -38 -48 222 592
use scs8hd_decap_4  FILLER_61_415
timestamp 1586364061
transform 1 0 39284 0 1 35360
box -38 -48 406 592
use scs8hd_decap_4  FILLER_61_421
timestamp 1586364061
transform 1 0 39836 0 1 35360
box -38 -48 406 592
use scs8hd_fill_2  FILLER_61_428
timestamp 1586364061
transform 1 0 40480 0 1 35360
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40664 0 1 35360
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42228 0 1 35360
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42044 0 1 35360
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41676 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_439
timestamp 1586364061
transform 1 0 41492 0 1 35360
box -38 -48 222 592
use scs8hd_fill_2  FILLER_61_443
timestamp 1586364061
transform 1 0 41860 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_456
timestamp 1586364061
transform 1 0 43056 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_468
timestamp 1586364061
transform 1 0 44160 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_480
timestamp 1586364061
transform 1 0 45264 0 1 35360
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_669
timestamp 1586364061
transform 1 0 46000 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_489
timestamp 1586364061
transform 1 0 46092 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_501
timestamp 1586364061
transform 1 0 47196 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 48852 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_61_513
timestamp 1586364061
transform 1 0 48300 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_670
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_12  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_56
timestamp 1586364061
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_68
timestamp 1586364061
transform 1 0 7360 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_80
timestamp 1586364061
transform 1 0 8464 0 -1 36448
box -38 -48 1142 592
use scs8hd_nor2_4  _232_
timestamp 1586364061
transform 1 0 10396 0 -1 36448
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_671
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_8  FILLER_62_93
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 -1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12052 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_8  FILLER_62_110
timestamp 1586364061
transform 1 0 11224 0 -1 36448
box -38 -48 774 592
use scs8hd_fill_1  FILLER_62_118
timestamp 1586364061
transform 1 0 11960 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_3  FILLER_62_121
timestamp 1586364061
transform 1 0 12236 0 -1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_62_133
timestamp 1586364061
transform 1 0 13340 0 -1 36448
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 36448
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 36448
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_672
timestamp 1586364061
transform 1 0 15180 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13524 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13892 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_137
timestamp 1586364061
transform 1 0 13708 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_62_141
timestamp 1586364061
transform 1 0 14076 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_8  FILLER_62_145
timestamp 1586364061
transform 1 0 14444 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_8  FILLER_62_157
timestamp 1586364061
transform 1 0 15548 0 -1 36448
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16376 0 -1 36448
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__247__B
timestamp 1586364061
transform 1 0 18124 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_62_165
timestamp 1586364061
transform 1 0 16284 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_8  FILLER_62_177
timestamp 1586364061
transform 1 0 17388 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_3  FILLER_62_187
timestamp 1586364061
transform 1 0 18308 0 -1 36448
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 18584 0 -1 36448
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_673
timestamp 1586364061
transform 1 0 20792 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19780 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_201
timestamp 1586364061
transform 1 0 19596 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_205
timestamp 1586364061
transform 1 0 19964 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_62_209
timestamp 1586364061
transform 1 0 20332 0 -1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_62_212
timestamp 1586364061
transform 1 0 20608 0 -1 36448
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21804 0 -1 36448
box -38 -48 866 592
use scs8hd_decap_8  FILLER_62_215
timestamp 1586364061
transform 1 0 20884 0 -1 36448
box -38 -48 774 592
use scs8hd_fill_2  FILLER_62_223
timestamp 1586364061
transform 1 0 21620 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_62_234
timestamp 1586364061
transform 1 0 22632 0 -1 36448
box -38 -48 1142 592
use scs8hd_nor2_4  _237_
timestamp 1586364061
transform 1 0 23736 0 -1 36448
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 36448
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24748 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_255
timestamp 1586364061
transform 1 0 24564 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_259
timestamp 1586364061
transform 1 0 24932 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_62_263
timestamp 1586364061
transform 1 0 25300 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_6  FILLER_62_267
timestamp 1586364061
transform 1 0 25668 0 -1 36448
box -38 -48 590 592
use scs8hd_fill_2  FILLER_62_276
timestamp 1586364061
transform 1 0 26496 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 36448
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_674
timestamp 1586364061
transform 1 0 26404 0 -1 36448
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26680 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_62_285
timestamp 1586364061
transform 1 0 27324 0 -1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_62_281
timestamp 1586364061
transform 1 0 26956 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27600 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27140 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_290
timestamp 1586364061
transform 1 0 27784 0 -1 36448
box -38 -48 222 592
use scs8hd_nor2_4  _283_
timestamp 1586364061
transform 1 0 27968 0 -1 36448
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 29532 0 -1 36448
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30728 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28980 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_301
timestamp 1586364061
transform 1 0 28796 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_305
timestamp 1586364061
transform 1 0 29164 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_2  FILLER_62_320
timestamp 1586364061
transform 1 0 30544 0 -1 36448
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32752 0 -1 36448
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_675
timestamp 1586364061
transform 1 0 32016 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32292 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31280 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_324
timestamp 1586364061
transform 1 0 30912 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_6  FILLER_62_330
timestamp 1586364061
transform 1 0 31464 0 -1 36448
box -38 -48 590 592
use scs8hd_fill_2  FILLER_62_337
timestamp 1586364061
transform 1 0 32108 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_3  FILLER_62_341
timestamp 1586364061
transform 1 0 32476 0 -1 36448
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_0_in_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34316 0 -1 36448
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__274__B
timestamp 1586364061
transform 1 0 34868 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35512 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_8  FILLER_62_353
timestamp 1586364061
transform 1 0 33580 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_3  FILLER_62_364
timestamp 1586364061
transform 1 0 34592 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_4  FILLER_62_369
timestamp 1586364061
transform 1 0 35052 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_62_373
timestamp 1586364061
transform 1 0 35420 0 -1 36448
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 35788 0 -1 36448
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 37720 0 -1 36448
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_676
timestamp 1586364061
transform 1 0 37628 0 -1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36984 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_62_376
timestamp 1586364061
transform 1 0 35696 0 -1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_62_388
timestamp 1586364061
transform 1 0 36800 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_392
timestamp 1586364061
transform 1 0 37168 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_62_396
timestamp 1586364061
transform 1 0 37536 0 -1 36448
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39652 0 -1 36448
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 40112 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_62_407
timestamp 1586364061
transform 1 0 38548 0 -1 36448
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_62_422
timestamp 1586364061
transform 1 0 39928 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_426
timestamp 1586364061
transform 1 0 40296 0 -1 36448
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40664 0 -1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42228 0 -1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41676 0 -1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_62_439
timestamp 1586364061
transform 1 0 41492 0 -1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_62_443
timestamp 1586364061
transform 1 0 41860 0 -1 36448
box -38 -48 406 592
use scs8hd_decap_8  FILLER_62_449
timestamp 1586364061
transform 1 0 42412 0 -1 36448
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_677
timestamp 1586364061
transform 1 0 43240 0 -1 36448
box -38 -48 130 592
use scs8hd_fill_1  FILLER_62_457
timestamp 1586364061
transform 1 0 43148 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_459
timestamp 1586364061
transform 1 0 43332 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_471
timestamp 1586364061
transform 1 0 44436 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_483
timestamp 1586364061
transform 1 0 45540 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_495
timestamp 1586364061
transform 1 0 46644 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_62_507
timestamp 1586364061
transform 1 0 47748 0 -1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 48852 0 -1 36448
box -38 -48 314 592
use scs8hd_fill_1  FILLER_62_515
timestamp 1586364061
transform 1 0 48484 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_51
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_678
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_59
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_74
timestamp 1586364061
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_86
timestamp 1586364061
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_98
timestamp 1586364061
transform 1 0 10120 0 1 36448
box -38 -48 774 592
use scs8hd_fill_2  FILLER_63_106
timestamp 1586364061
transform 1 0 10856 0 1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_63_110
timestamp 1586364061
transform 1 0 11224 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11040 0 1 36448
box -38 -48 222 592
use scs8hd_conb_1  _446_
timestamp 1586364061
transform 1 0 11316 0 1 36448
box -38 -48 314 592
use scs8hd_decap_4  FILLER_63_114
timestamp 1586364061
transform 1 0 11592 0 1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_63_121
timestamp 1586364061
transform 1 0 12236 0 1 36448
box -38 -48 130 592
use scs8hd_fill_1  FILLER_63_118
timestamp 1586364061
transform 1 0 11960 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_679
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_63_131
timestamp 1586364061
transform 1 0 13156 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_127
timestamp 1586364061
transform 1 0 12788 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_14_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13340 0 1 36448
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15088 0 1 36448
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14904 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_144
timestamp 1586364061
transform 1 0 14352 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_148
timestamp 1586364061
transform 1 0 14720 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_161
timestamp 1586364061
transform 1 0 15916 0 1 36448
box -38 -48 222 592
use scs8hd_decap_3  FILLER_63_165
timestamp 1586364061
transform 1 0 16284 0 1 36448
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16100 0 1 36448
box -38 -48 222 592
use scs8hd_decap_6  FILLER_63_174
timestamp 1586364061
transform 1 0 17112 0 1 36448
box -38 -48 590 592
use scs8hd_fill_2  FILLER_63_170
timestamp 1586364061
transform 1 0 16744 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__246__B
timestamp 1586364061
transform 1 0 16928 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__246__A
timestamp 1586364061
transform 1 0 16560 0 1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_63_180
timestamp 1586364061
transform 1 0 17664 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__247__A
timestamp 1586364061
transform 1 0 17756 0 1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_63_184
timestamp 1586364061
transform 1 0 18032 0 1 36448
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_680
timestamp 1586364061
transform 1 0 17940 0 1 36448
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18676 0 1 36448
box -38 -48 1050 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20424 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 18492 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19872 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20240 0 1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_63_188
timestamp 1586364061
transform 1 0 18400 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_202
timestamp 1586364061
transform 1 0 19688 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_206
timestamp 1586364061
transform 1 0 20056 0 1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_63_219
timestamp 1586364061
transform 1 0 21252 0 1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_63_223
timestamp 1586364061
transform 1 0 21620 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_63_226
timestamp 1586364061
transform 1 0 21896 0 1 36448
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21988 0 1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_63_234
timestamp 1586364061
transform 1 0 22632 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_230
timestamp 1586364061
transform 1 0 22264 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_63_238
timestamp 1586364061
transform 1 0 23000 0 1 36448
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22816 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__242__B
timestamp 1586364061
transform 1 0 23368 0 1 36448
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_681
timestamp 1586364061
transform 1 0 23552 0 1 36448
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_63_248
timestamp 1586364061
transform 1 0 23920 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_63_256
timestamp 1586364061
transform 1 0 24656 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_252
timestamp 1586364061
transform 1 0 24288 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 24472 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_260
timestamp 1586364061
transform 1 0 25024 0 1 36448
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24748 0 1 36448
box -38 -48 314 592
use scs8hd_decap_4  FILLER_63_264
timestamp 1586364061
transform 1 0 25392 0 1 36448
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25208 0 1 36448
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25760 0 1 36448
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26772 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26220 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26588 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27784 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_271
timestamp 1586364061
transform 1 0 26036 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_275
timestamp 1586364061
transform 1 0 26404 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_288
timestamp 1586364061
transform 1 0 27600 0 1 36448
box -38 -48 222 592
use scs8hd_decap_4  FILLER_63_292
timestamp 1586364061
transform 1 0 27968 0 1 36448
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch
timestamp 1586364061
transform 1 0 29532 0 1 36448
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_682
timestamp 1586364061
transform 1 0 29164 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__288__A
timestamp 1586364061
transform 1 0 30728 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28980 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28428 0 1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_63_296
timestamp 1586364061
transform 1 0 28336 0 1 36448
box -38 -48 130 592
use scs8hd_decap_4  FILLER_63_299
timestamp 1586364061
transform 1 0 28612 0 1 36448
box -38 -48 406 592
use scs8hd_decap_3  FILLER_63_306
timestamp 1586364061
transform 1 0 29256 0 1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_63_320
timestamp 1586364061
transform 1 0 30544 0 1 36448
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32844 0 1 36448
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31280 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 32292 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__288__B
timestamp 1586364061
transform 1 0 31096 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32660 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_324
timestamp 1586364061
transform 1 0 30912 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_337
timestamp 1586364061
transform 1 0 32108 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_341
timestamp 1586364061
transform 1 0 32476 0 1 36448
box -38 -48 222 592
use scs8hd_nor2_4  _274_
timestamp 1586364061
transform 1 0 34868 0 1 36448
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_683
timestamp 1586364061
transform 1 0 34776 0 1 36448
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__274__A
timestamp 1586364061
transform 1 0 34592 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33856 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34224 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_354
timestamp 1586364061
transform 1 0 33672 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_358
timestamp 1586364061
transform 1 0 34040 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_362
timestamp 1586364061
transform 1 0 34408 0 1 36448
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36524 0 1 36448
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__277__A
timestamp 1586364061
transform 1 0 35880 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__279__B
timestamp 1586364061
transform 1 0 37996 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__277__B
timestamp 1586364061
transform 1 0 36248 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_376
timestamp 1586364061
transform 1 0 35696 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_380
timestamp 1586364061
transform 1 0 36064 0 1 36448
box -38 -48 222 592
use scs8hd_fill_1  FILLER_63_384
timestamp 1586364061
transform 1 0 36432 0 1 36448
box -38 -48 130 592
use scs8hd_decap_6  FILLER_63_394
timestamp 1586364061
transform 1 0 37352 0 1 36448
box -38 -48 590 592
use scs8hd_fill_1  FILLER_63_400
timestamp 1586364061
transform 1 0 37904 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_406
timestamp 1586364061
transform 1 0 38456 0 1 36448
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 38180 0 1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_63_410
timestamp 1586364061
transform 1 0 38824 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38640 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__279__A
timestamp 1586364061
transform 1 0 39008 0 1 36448
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39192 0 1 36448
box -38 -48 314 592
use scs8hd_fill_2  FILLER_63_417
timestamp 1586364061
transform 1 0 39468 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_421
timestamp 1586364061
transform 1 0 39836 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39652 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_425
timestamp 1586364061
transform 1 0 40204 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 40020 0 1 36448
box -38 -48 222 592
use scs8hd_decap_3  FILLER_63_428
timestamp 1586364061
transform 1 0 40480 0 1 36448
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_684
timestamp 1586364061
transform 1 0 40388 0 1 36448
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40756 0 1 36448
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41768 0 1 36448
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41216 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 42228 0 1 36448
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 41584 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_434
timestamp 1586364061
transform 1 0 41032 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_438
timestamp 1586364061
transform 1 0 41400 0 1 36448
box -38 -48 222 592
use scs8hd_fill_2  FILLER_63_445
timestamp 1586364061
transform 1 0 42044 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_449
timestamp 1586364061
transform 1 0 42412 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_461
timestamp 1586364061
transform 1 0 43516 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_473
timestamp 1586364061
transform 1 0 44620 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_685
timestamp 1586364061
transform 1 0 46000 0 1 36448
box -38 -48 130 592
use scs8hd_decap_3  FILLER_63_485
timestamp 1586364061
transform 1 0 45724 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_489
timestamp 1586364061
transform 1 0 46092 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_501
timestamp 1586364061
transform 1 0 47196 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 48852 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_63_513
timestamp 1586364061
transform 1 0 48300 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_686
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_68
timestamp 1586364061
transform 1 0 7360 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_80
timestamp 1586364061
transform 1 0 8464 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_687
timestamp 1586364061
transform 1 0 9568 0 -1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__233__B
timestamp 1586364061
transform 1 0 10764 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_64_93
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_64_107
timestamp 1586364061
transform 1 0 10948 0 -1 37536
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 -1 37536
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11500 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_111
timestamp 1586364061
transform 1 0 11316 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_64_115
timestamp 1586364061
transform 1 0 11684 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_8  FILLER_64_128
timestamp 1586364061
transform 1 0 12880 0 -1 37536
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13616 0 -1 37536
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 37536
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_688
timestamp 1586364061
transform 1 0 15180 0 -1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_64_139
timestamp 1586364061
transform 1 0 13892 0 -1 37536
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_64_151
timestamp 1586364061
transform 1 0 14996 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_157
timestamp 1586364061
transform 1 0 15548 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_161
timestamp 1586364061
transform 1 0 15916 0 -1 37536
box -38 -48 222 592
use scs8hd_nor2_4  _246_
timestamp 1586364061
transform 1 0 16560 0 -1 37536
box -38 -48 866 592
use scs8hd_nor2_4  _247_
timestamp 1586364061
transform 1 0 18124 0 -1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17572 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16100 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_3  FILLER_64_165
timestamp 1586364061
transform 1 0 16284 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_2  FILLER_64_177
timestamp 1586364061
transform 1 0 17388 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_64_181
timestamp 1586364061
transform 1 0 17756 0 -1 37536
box -38 -48 406 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 37536
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_689
timestamp 1586364061
transform 1 0 20792 0 -1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__251__B
timestamp 1586364061
transform 1 0 19136 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19504 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_194
timestamp 1586364061
transform 1 0 18952 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_198
timestamp 1586364061
transform 1 0 19320 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_1  FILLER_64_202
timestamp 1586364061
transform 1 0 19688 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_206
timestamp 1586364061
transform 1 0 20056 0 -1 37536
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21712 0 -1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23276 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_8  FILLER_64_215
timestamp 1586364061
transform 1 0 20884 0 -1 37536
box -38 -48 774 592
use scs8hd_fill_1  FILLER_64_223
timestamp 1586364061
transform 1 0 21620 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_8  FILLER_64_233
timestamp 1586364061
transform 1 0 22540 0 -1 37536
box -38 -48 774 592
use scs8hd_nor2_4  _242_
timestamp 1586364061
transform 1 0 24012 0 -1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 25024 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__243__B
timestamp 1586364061
transform 1 0 25392 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_6  FILLER_64_243
timestamp 1586364061
transform 1 0 23460 0 -1 37536
box -38 -48 590 592
use scs8hd_fill_2  FILLER_64_258
timestamp 1586364061
transform 1 0 24840 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_262
timestamp 1586364061
transform 1 0 25208 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_8  FILLER_64_266
timestamp 1586364061
transform 1 0 25576 0 -1 37536
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26864 0 -1 37536
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_690
timestamp 1586364061
transform 1 0 26404 0 -1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26680 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_1  FILLER_64_274
timestamp 1586364061
transform 1 0 26312 0 -1 37536
box -38 -48 130 592
use scs8hd_fill_2  FILLER_64_276
timestamp 1586364061
transform 1 0 26496 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_8  FILLER_64_289
timestamp 1586364061
transform 1 0 27692 0 -1 37536
box -38 -48 774 592
use scs8hd_nor2_4  _288_
timestamp 1586364061
transform 1 0 30360 0 -1 37536
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28428 0 -1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_6_.latch_D
timestamp 1586364061
transform 1 0 29532 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__289__B
timestamp 1586364061
transform 1 0 29992 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_3  FILLER_64_306
timestamp 1586364061
transform 1 0 29256 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_3  FILLER_64_311
timestamp 1586364061
transform 1 0 29716 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_2  FILLER_64_316
timestamp 1586364061
transform 1 0 30176 0 -1 37536
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 37536
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_691
timestamp 1586364061
transform 1 0 32016 0 -1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31832 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31372 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_327
timestamp 1586364061
transform 1 0 31188 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_3  FILLER_64_331
timestamp 1586364061
transform 1 0 31556 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_2  FILLER_64_348
timestamp 1586364061
transform 1 0 33120 0 -1 37536
box -38 -48 222 592
use scs8hd_nor2_4  _277_
timestamp 1586364061
transform 1 0 35420 0 -1 37536
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33856 0 -1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 35236 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33304 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33672 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_352
timestamp 1586364061
transform 1 0 33488 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_6  FILLER_64_365
timestamp 1586364061
transform 1 0 34684 0 -1 37536
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_692
timestamp 1586364061
transform 1 0 37628 0 -1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36432 0 -1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36800 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_382
timestamp 1586364061
transform 1 0 36248 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_386
timestamp 1586364061
transform 1 0 36616 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_6  FILLER_64_390
timestamp 1586364061
transform 1 0 36984 0 -1 37536
box -38 -48 590 592
use scs8hd_fill_1  FILLER_64_396
timestamp 1586364061
transform 1 0 37536 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_398
timestamp 1586364061
transform 1 0 37720 0 -1 37536
box -38 -48 590 592
use scs8hd_nor2_4  _279_
timestamp 1586364061
transform 1 0 38364 0 -1 37536
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 39928 0 -1 37536
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_64_404
timestamp 1586364061
transform 1 0 38272 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_8  FILLER_64_414
timestamp 1586364061
transform 1 0 39192 0 -1 37536
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 41676 0 -1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41124 0 -1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_64_433
timestamp 1586364061
transform 1 0 40940 0 -1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_64_437
timestamp 1586364061
transform 1 0 41308 0 -1 37536
box -38 -48 406 592
use scs8hd_decap_8  FILLER_64_450
timestamp 1586364061
transform 1 0 42504 0 -1 37536
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_693
timestamp 1586364061
transform 1 0 43240 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_459
timestamp 1586364061
transform 1 0 43332 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_471
timestamp 1586364061
transform 1 0 44436 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_483
timestamp 1586364061
transform 1 0 45540 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_495
timestamp 1586364061
transform 1 0 46644 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_64_507
timestamp 1586364061
transform 1 0 47748 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 48852 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_64_515
timestamp 1586364061
transform 1 0 48484 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_3  PHY_130
timestamp 1586364061
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_65_3
timestamp 1586364061
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_15
timestamp 1586364061
transform 1 0 2484 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_27
timestamp 1586364061
transform 1 0 3588 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_39
timestamp 1586364061
transform 1 0 4692 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_65_51
timestamp 1586364061
transform 1 0 5796 0 1 37536
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_694
timestamp 1586364061
transform 1 0 6716 0 1 37536
box -38 -48 130 592
use scs8hd_fill_2  FILLER_65_59
timestamp 1586364061
transform 1 0 6532 0 1 37536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_65_62
timestamp 1586364061
transform 1 0 6808 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_74
timestamp 1586364061
transform 1 0 7912 0 1 37536
box -38 -48 1142 592
use scs8hd_nor2_4  _233_
timestamp 1586364061
transform 1 0 10764 0 1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 10580 0 1 37536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_65_86
timestamp 1586364061
transform 1 0 9016 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_65_98
timestamp 1586364061
transform 1 0 10120 0 1 37536
box -38 -48 406 592
use scs8hd_fill_1  FILLER_65_102
timestamp 1586364061
transform 1 0 10488 0 1 37536
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 37536
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_695
timestamp 1586364061
transform 1 0 12328 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_114
timestamp 1586364061
transform 1 0 11592 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_118
timestamp 1586364061
transform 1 0 11960 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_132
timestamp 1586364061
transform 1 0 13248 0 1 37536
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 1 37536
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15180 0 1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_136
timestamp 1586364061
transform 1 0 13616 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_140
timestamp 1586364061
transform 1 0 13984 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_145
timestamp 1586364061
transform 1 0 14444 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_149
timestamp 1586364061
transform 1 0 14812 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_162
timestamp 1586364061
transform 1 0 16008 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_166
timestamp 1586364061
transform 1 0 16376 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 1 37536
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16744 0 1 37536
box -38 -48 314 592
use scs8hd_fill_2  FILLER_65_173
timestamp 1586364061
transform 1 0 17020 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17204 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_177
timestamp 1586364061
transform 1 0 17388 0 1 37536
box -38 -48 406 592
use scs8hd_decap_4  FILLER_65_184
timestamp 1586364061
transform 1 0 18032 0 1 37536
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__249__B
timestamp 1586364061
transform 1 0 17756 0 1 37536
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_696
timestamp 1586364061
transform 1 0 17940 0 1 37536
box -38 -48 130 592
use scs8hd_nor2_4  _251_
timestamp 1586364061
transform 1 0 19044 0 1 37536
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20608 0 1 37536
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20424 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__249__A
timestamp 1586364061
transform 1 0 18400 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__251__A
timestamp 1586364061
transform 1 0 18860 0 1 37536
box -38 -48 222 592
use scs8hd_decap_3  FILLER_65_190
timestamp 1586364061
transform 1 0 18584 0 1 37536
box -38 -48 314 592
use scs8hd_decap_6  FILLER_65_204
timestamp 1586364061
transform 1 0 19872 0 1 37536
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22356 0 1 37536
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22816 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23276 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21804 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_223
timestamp 1586364061
transform 1 0 21620 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_227
timestamp 1586364061
transform 1 0 21988 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_234
timestamp 1586364061
transform 1 0 22632 0 1 37536
box -38 -48 222 592
use scs8hd_decap_3  FILLER_65_238
timestamp 1586364061
transform 1 0 23000 0 1 37536
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 24840 0 1 37536
box -38 -48 1050 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 37536
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_697
timestamp 1586364061
transform 1 0 23552 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 24656 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 37536
box -38 -48 222 592
use scs8hd_fill_1  FILLER_65_243
timestamp 1586364061
transform 1 0 23460 0 1 37536
box -38 -48 130 592
use scs8hd_fill_2  FILLER_65_248
timestamp 1586364061
transform 1 0 23920 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_252
timestamp 1586364061
transform 1 0 24288 0 1 37536
box -38 -48 406 592
use scs8hd_decap_3  FILLER_65_273
timestamp 1586364061
transform 1 0 26220 0 1 37536
box -38 -48 314 592
use scs8hd_fill_2  FILLER_65_269
timestamp 1586364061
transform 1 0 25852 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26036 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26496 0 1 37536
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26680 0 1 37536
box -38 -48 866 592
use scs8hd_fill_2  FILLER_65_287
timestamp 1586364061
transform 1 0 27508 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_295
timestamp 1586364061
transform 1 0 28244 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_291
timestamp 1586364061
transform 1 0 27876 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28060 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27692 0 1 37536
box -38 -48 222 592
use scs8hd_nor2_4  _289_
timestamp 1586364061
transform 1 0 29992 0 1 37536
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_698
timestamp 1586364061
transform 1 0 29164 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28428 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__289__A
timestamp 1586364061
transform 1 0 29808 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29440 0 1 37536
box -38 -48 222 592
use scs8hd_decap_6  FILLER_65_299
timestamp 1586364061
transform 1 0 28612 0 1 37536
box -38 -48 590 592
use scs8hd_fill_2  FILLER_65_306
timestamp 1586364061
transform 1 0 29256 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_310
timestamp 1586364061
transform 1 0 29624 0 1 37536
box -38 -48 222 592
use scs8hd_decap_3  FILLER_65_327
timestamp 1586364061
transform 1 0 31188 0 1 37536
box -38 -48 314 592
use scs8hd_fill_2  FILLER_65_323
timestamp 1586364061
transform 1 0 30820 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31004 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31464 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_339
timestamp 1586364061
transform 1 0 32292 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_335
timestamp 1586364061
transform 1 0 31924 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32476 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32108 0 1 37536
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31648 0 1 37536
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32660 0 1 37536
box -38 -48 866 592
use scs8hd_decap_4  FILLER_65_352
timestamp 1586364061
transform 1 0 33488 0 1 37536
box -38 -48 406 592
use scs8hd_decap_6  FILLER_65_359
timestamp 1586364061
transform 1 0 34132 0 1 37536
box -38 -48 590 592
use scs8hd_fill_1  FILLER_65_356
timestamp 1586364061
transform 1 0 33856 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33948 0 1 37536
box -38 -48 222 592
use scs8hd_decap_3  FILLER_65_367
timestamp 1586364061
transform 1 0 34868 0 1 37536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_65_365
timestamp 1586364061
transform 1 0 34684 0 1 37536
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_699
timestamp 1586364061
transform 1 0 34776 0 1 37536
box -38 -48 130 592
use scs8hd_fill_2  FILLER_65_373
timestamp 1586364061
transform 1 0 35420 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 35604 0 1 37536
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35144 0 1 37536
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36156 0 1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 37720 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35972 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 37352 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_377
timestamp 1586364061
transform 1 0 35788 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_390
timestamp 1586364061
transform 1 0 36984 0 1 37536
box -38 -48 406 592
use scs8hd_fill_2  FILLER_65_396
timestamp 1586364061
transform 1 0 37536 0 1 37536
box -38 -48 222 592
use scs8hd_decap_4  FILLER_65_400
timestamp 1586364061
transform 1 0 37904 0 1 37536
box -38 -48 406 592
use scs8hd_fill_1  FILLER_65_404
timestamp 1586364061
transform 1 0 38272 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38364 0 1 37536
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38548 0 1 37536
box -38 -48 866 592
use scs8hd_decap_4  FILLER_65_420
timestamp 1586364061
transform 1 0 39744 0 1 37536
box -38 -48 406 592
use scs8hd_fill_2  FILLER_65_416
timestamp 1586364061
transform 1 0 39376 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 39560 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_428
timestamp 1586364061
transform 1 0 40480 0 1 37536
box -38 -48 222 592
use scs8hd_fill_1  FILLER_65_424
timestamp 1586364061
transform 1 0 40112 0 1 37536
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40204 0 1 37536
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_700
timestamp 1586364061
transform 1 0 40388 0 1 37536
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 42412 0 1 37536
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40848 0 1 37536
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 40664 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 42228 0 1 37536
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 41860 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_441
timestamp 1586364061
transform 1 0 41676 0 1 37536
box -38 -48 222 592
use scs8hd_fill_2  FILLER_65_445
timestamp 1586364061
transform 1 0 42044 0 1 37536
box -38 -48 222 592
use scs8hd_decap_12  FILLER_65_458
timestamp 1586364061
transform 1 0 43240 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_470
timestamp 1586364061
transform 1 0 44344 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_65_482
timestamp 1586364061
transform 1 0 45448 0 1 37536
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_701
timestamp 1586364061
transform 1 0 46000 0 1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_65_489
timestamp 1586364061
transform 1 0 46092 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_65_501
timestamp 1586364061
transform 1 0 47196 0 1 37536
box -38 -48 1142 592
use scs8hd_decap_3  PHY_131
timestamp 1586364061
transform -1 0 48852 0 1 37536
box -38 -48 314 592
use scs8hd_decap_3  FILLER_65_513
timestamp 1586364061
transform 1 0 48300 0 1 37536
box -38 -48 314 592
use scs8hd_decap_3  PHY_132
timestamp 1586364061
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_3  PHY_134
timestamp 1586364061
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use scs8hd_decap_12  FILLER_66_3
timestamp 1586364061
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_15
timestamp 1586364061
transform 1 0 2484 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_3
timestamp 1586364061
transform 1 0 1380 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_15
timestamp 1586364061
transform 1 0 2484 0 1 38624
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_702
timestamp 1586364061
transform 1 0 3956 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_4  FILLER_66_27
timestamp 1586364061
transform 1 0 3588 0 -1 38624
box -38 -48 406 592
use scs8hd_decap_12  FILLER_66_32
timestamp 1586364061
transform 1 0 4048 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_44
timestamp 1586364061
transform 1 0 5152 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_27
timestamp 1586364061
transform 1 0 3588 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_39
timestamp 1586364061
transform 1 0 4692 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_67_51
timestamp 1586364061
transform 1 0 5796 0 1 38624
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_710
timestamp 1586364061
transform 1 0 6716 0 1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_56
timestamp 1586364061
transform 1 0 6256 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_68
timestamp 1586364061
transform 1 0 7360 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_80
timestamp 1586364061
transform 1 0 8464 0 -1 38624
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_67_59
timestamp 1586364061
transform 1 0 6532 0 1 38624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_67_62
timestamp 1586364061
transform 1 0 6808 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_74
timestamp 1586364061
transform 1 0 7912 0 1 38624
box -38 -48 1142 592
use scs8hd_nor2_4  _234_
timestamp 1586364061
transform 1 0 10764 0 1 38624
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_703
timestamp 1586364061
transform 1 0 9568 0 -1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 10580 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__234__B
timestamp 1586364061
transform 1 0 10764 0 -1 38624
box -38 -48 222 592
use scs8hd_decap_12  FILLER_66_93
timestamp 1586364061
transform 1 0 9660 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_66_107
timestamp 1586364061
transform 1 0 10948 0 -1 38624
box -38 -48 406 592
use scs8hd_decap_12  FILLER_67_86
timestamp 1586364061
transform 1 0 9016 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_67_98
timestamp 1586364061
transform 1 0 10120 0 1 38624
box -38 -48 406 592
use scs8hd_fill_1  FILLER_67_102
timestamp 1586364061
transform 1 0 10488 0 1 38624
box -38 -48 130 592
use scs8hd_fill_2  FILLER_67_118
timestamp 1586364061
transform 1 0 11960 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_114
timestamp 1586364061
transform 1 0 11592 0 1 38624
box -38 -48 222 592
use scs8hd_fill_1  FILLER_66_111
timestamp 1586364061
transform 1 0 11316 0 -1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 38624
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 38624
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_66_127
timestamp 1586364061
transform 1 0 12788 0 -1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_66_123
timestamp 1586364061
transform 1 0 12420 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_711
timestamp 1586364061
transform 1 0 12328 0 1 38624
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 38624
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12420 0 1 38624
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_67_134
timestamp 1586364061
transform 1 0 13432 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_142
timestamp 1586364061
transform 1 0 14168 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_138
timestamp 1586364061
transform 1 0 13800 0 1 38624
box -38 -48 222 592
use scs8hd_decap_6  FILLER_66_140
timestamp 1586364061
transform 1 0 13984 0 -1 38624
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 38624
box -38 -48 222 592
use scs8hd_fill_1  FILLER_66_152
timestamp 1586364061
transform 1 0 15088 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_4  FILLER_66_148
timestamp 1586364061
transform 1 0 14720 0 -1 38624
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_704
timestamp 1586364061
transform 1 0 15180 0 -1 38624
box -38 -48 130 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14536 0 1 38624
box -38 -48 866 592
use scs8hd_decap_3  FILLER_67_159
timestamp 1586364061
transform 1 0 15732 0 1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_155
timestamp 1586364061
transform 1 0 15364 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 38624
box -38 -48 866 592
use scs8hd_fill_1  FILLER_66_170
timestamp 1586364061
transform 1 0 16744 0 -1 38624
box -38 -48 130 592
use scs8hd_fill_1  FILLER_66_167
timestamp 1586364061
transform 1 0 16468 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_4  FILLER_66_163
timestamp 1586364061
transform 1 0 16100 0 -1 38624
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 38624
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 16192 0 1 38624
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_67_184
timestamp 1586364061
transform 1 0 18032 0 1 38624
box -38 -48 406 592
use scs8hd_fill_2  FILLER_67_179
timestamp 1586364061
transform 1 0 17572 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_175
timestamp 1586364061
transform 1 0 17204 0 1 38624
box -38 -48 222 592
use scs8hd_decap_8  FILLER_66_180
timestamp 1586364061
transform 1 0 17664 0 -1 38624
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_712
timestamp 1586364061
transform 1 0 17940 0 1 38624
box -38 -48 130 592
use scs8hd_fill_2  FILLER_67_191
timestamp 1586364061
transform 1 0 18676 0 1 38624
box -38 -48 222 592
use scs8hd_fill_1  FILLER_67_188
timestamp 1586364061
transform 1 0 18400 0 1 38624
box -38 -48 130 592
use scs8hd_fill_2  FILLER_66_197
timestamp 1586364061
transform 1 0 19228 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__252__B
timestamp 1586364061
transform 1 0 19412 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 18492 0 1 38624
box -38 -48 222 592
use scs8hd_nor2_4  _252_
timestamp 1586364061
transform 1 0 18860 0 1 38624
box -38 -48 866 592
use scs8hd_nor2_4  _249_
timestamp 1586364061
transform 1 0 18400 0 -1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_67_206
timestamp 1586364061
transform 1 0 20056 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_202
timestamp 1586364061
transform 1 0 19688 0 1 38624
box -38 -48 222 592
use scs8hd_fill_1  FILLER_66_209
timestamp 1586364061
transform 1 0 20332 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_8  FILLER_66_201
timestamp 1586364061
transform 1 0 19596 0 -1 38624
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20424 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__252__A
timestamp 1586364061
transform 1 0 19872 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20240 0 1 38624
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 20424 0 1 38624
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_66_212
timestamp 1586364061
transform 1 0 20608 0 -1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_705
timestamp 1586364061
transform 1 0 20792 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_3  FILLER_67_221
timestamp 1586364061
transform 1 0 21436 0 1 38624
box -38 -48 314 592
use scs8hd_fill_1  FILLER_66_223
timestamp 1586364061
transform 1 0 21620 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_8  FILLER_66_215
timestamp 1586364061
transform 1 0 20884 0 -1 38624
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21712 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21712 0 -1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_67_232
timestamp 1586364061
transform 1 0 22448 0 1 38624
box -38 -48 222 592
use scs8hd_decap_3  FILLER_67_226
timestamp 1586364061
transform 1 0 21896 0 1 38624
box -38 -48 314 592
use scs8hd_decap_8  FILLER_66_233
timestamp 1586364061
transform 1 0 22540 0 -1 38624
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22632 0 1 38624
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22172 0 1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_240
timestamp 1586364061
transform 1 0 23184 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_236
timestamp 1586364061
transform 1 0 22816 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23276 0 -1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_66_250
timestamp 1586364061
transform 1 0 24104 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24288 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 23368 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_713
timestamp 1586364061
transform 1 0 23552 0 1 38624
box -38 -48 130 592
use scs8hd_nor2_4  _240_
timestamp 1586364061
transform 1 0 23644 0 1 38624
box -38 -48 866 592
use scs8hd_fill_2  FILLER_67_258
timestamp 1586364061
transform 1 0 24840 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_254
timestamp 1586364061
transform 1 0 24472 0 1 38624
box -38 -48 222 592
use scs8hd_decap_4  FILLER_66_254
timestamp 1586364061
transform 1 0 24472 0 -1 38624
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 25024 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 24656 0 1 38624
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 25208 0 1 38624
box -38 -48 1050 592
use scs8hd_nor2_4  _243_
timestamp 1586364061
transform 1 0 24840 0 -1 38624
box -38 -48 866 592
use scs8hd_decap_8  FILLER_66_267
timestamp 1586364061
transform 1 0 25668 0 -1 38624
box -38 -48 774 592
use scs8hd_fill_2  FILLER_67_277
timestamp 1586364061
transform 1 0 26588 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_273
timestamp 1586364061
transform 1 0 26220 0 1 38624
box -38 -48 222 592
use scs8hd_decap_4  FILLER_66_276
timestamp 1586364061
transform 1 0 26496 0 -1 38624
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26404 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_706
timestamp 1586364061
transform 1 0 26404 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_6  FILLER_67_288
timestamp 1586364061
transform 1 0 27600 0 1 38624
box -38 -48 590 592
use scs8hd_fill_2  FILLER_67_284
timestamp 1586364061
transform 1 0 27232 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26772 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27416 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26864 0 -1 38624
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26956 0 1 38624
box -38 -48 314 592
use scs8hd_fill_1  FILLER_67_294
timestamp 1586364061
transform 1 0 28152 0 1 38624
box -38 -48 130 592
use scs8hd_decap_8  FILLER_66_289
timestamp 1586364061
transform 1 0 27692 0 -1 38624
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28244 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_301
timestamp 1586364061
transform 1 0 28796 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_297
timestamp 1586364061
transform 1 0 28428 0 1 38624
box -38 -48 222 592
use scs8hd_decap_6  FILLER_66_300
timestamp 1586364061
transform 1 0 28704 0 -1 38624
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__286__B
timestamp 1586364061
transform 1 0 28612 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_714
timestamp 1586364061
transform 1 0 29164 0 1 38624
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28428 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_6  FILLER_66_308
timestamp 1586364061
transform 1 0 29440 0 -1 38624
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__286__A
timestamp 1586364061
transform 1 0 29256 0 -1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29992 0 -1 38624
box -38 -48 866 592
use scs8hd_nor2_4  _286_
timestamp 1586364061
transform 1 0 29256 0 1 38624
box -38 -48 866 592
use scs8hd_decap_6  FILLER_67_315
timestamp 1586364061
transform 1 0 30084 0 1 38624
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 30636 0 1 38624
box -38 -48 222 592
use scs8hd_decap_8  FILLER_66_327
timestamp 1586364061
transform 1 0 31188 0 -1 38624
box -38 -48 774 592
use scs8hd_fill_2  FILLER_66_323
timestamp 1586364061
transform 1 0 30820 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31004 0 -1 38624
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 30820 0 1 38624
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_707
timestamp 1586364061
transform 1 0 32016 0 -1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32292 0 1 38624
box -38 -48 222 592
use scs8hd_fill_1  FILLER_66_335
timestamp 1586364061
transform 1 0 31924 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_3  FILLER_66_337
timestamp 1586364061
transform 1 0 32108 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_4  FILLER_67_334
timestamp 1586364061
transform 1 0 31832 0 1 38624
box -38 -48 406 592
use scs8hd_fill_1  FILLER_67_338
timestamp 1586364061
transform 1 0 32200 0 1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32660 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_341
timestamp 1586364061
transform 1 0 32476 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32384 0 -1 38624
box -38 -48 866 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32844 0 1 38624
box -38 -48 866 592
use scs8hd_decap_3  FILLER_67_358
timestamp 1586364061
transform 1 0 34040 0 1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_354
timestamp 1586364061
transform 1 0 33672 0 1 38624
box -38 -48 222 592
use scs8hd_decap_8  FILLER_66_360
timestamp 1586364061
transform 1 0 34224 0 -1 38624
box -38 -48 774 592
use scs8hd_decap_4  FILLER_66_353
timestamp 1586364061
transform 1 0 33580 0 -1 38624
box -38 -48 406 592
use scs8hd_fill_2  FILLER_66_349
timestamp 1586364061
transform 1 0 33212 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33396 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33856 0 1 38624
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33948 0 -1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_372
timestamp 1586364061
transform 1 0 35328 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_367
timestamp 1586364061
transform 1 0 34868 0 1 38624
box -38 -48 222 592
use scs8hd_decap_3  FILLER_67_363
timestamp 1586364061
transform 1 0 34500 0 1 38624
box -38 -48 314 592
use scs8hd_decap_3  FILLER_66_368
timestamp 1586364061
transform 1 0 34960 0 -1 38624
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34316 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_715
timestamp 1586364061
transform 1 0 34776 0 1 38624
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35052 0 1 38624
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 35236 0 -1 38624
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35512 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_376
timestamp 1586364061
transform 1 0 35696 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_66_386
timestamp 1586364061
transform 1 0 36616 0 -1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_66_382
timestamp 1586364061
transform 1 0 36248 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36432 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36064 0 1 38624
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37076 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36800 0 -1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_389
timestamp 1586364061
transform 1 0 36892 0 1 38624
box -38 -48 222 592
use scs8hd_decap_4  FILLER_67_393
timestamp 1586364061
transform 1 0 37260 0 1 38624
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_708
timestamp 1586364061
transform 1 0 37628 0 -1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 37628 0 1 38624
box -38 -48 222 592
use scs8hd_fill_1  FILLER_66_396
timestamp 1586364061
transform 1 0 37536 0 -1 38624
box -38 -48 130 592
use scs8hd_fill_2  FILLER_67_399
timestamp 1586364061
transform 1 0 37812 0 1 38624
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 37720 0 -1 38624
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_66_390
timestamp 1586364061
transform 1 0 36984 0 -1 38624
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 37996 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_403
timestamp 1586364061
transform 1 0 38180 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_66_409
timestamp 1586364061
transform 1 0 38732 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 38916 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38364 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38548 0 1 38624
box -38 -48 866 592
use scs8hd_decap_6  FILLER_67_420
timestamp 1586364061
transform 1 0 39744 0 1 38624
box -38 -48 590 592
use scs8hd_fill_2  FILLER_67_416
timestamp 1586364061
transform 1 0 39376 0 1 38624
box -38 -48 222 592
use scs8hd_decap_8  FILLER_66_420
timestamp 1586364061
transform 1 0 39744 0 -1 38624
box -38 -48 774 592
use scs8hd_decap_4  FILLER_66_413
timestamp 1586364061
transform 1 0 39100 0 -1 38624
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39560 0 1 38624
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 39468 0 -1 38624
box -38 -48 314 592
use scs8hd_fill_1  FILLER_67_426
timestamp 1586364061
transform 1 0 40296 0 1 38624
box -38 -48 130 592
use scs8hd_decap_3  FILLER_66_428
timestamp 1586364061
transform 1 0 40480 0 -1 38624
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_716
timestamp 1586364061
transform 1 0 40388 0 1 38624
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40480 0 1 38624
box -38 -48 314 592
use scs8hd_fill_2  FILLER_67_442
timestamp 1586364061
transform 1 0 41768 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_435
timestamp 1586364061
transform 1 0 41124 0 1 38624
box -38 -48 222 592
use scs8hd_fill_2  FILLER_67_431
timestamp 1586364061
transform 1 0 40756 0 1 38624
box -38 -48 222 592
use scs8hd_decap_8  FILLER_66_440
timestamp 1586364061
transform 1 0 41584 0 -1 38624
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41308 0 1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 40940 0 1 38624
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 40756 0 -1 38624
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 41492 0 1 38624
box -38 -48 314 592
use scs8hd_decap_12  FILLER_67_446
timestamp 1586364061
transform 1 0 42136 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_66_451
timestamp 1586364061
transform 1 0 42596 0 -1 38624
box -38 -48 590 592
use scs8hd_fill_1  FILLER_66_448
timestamp 1586364061
transform 1 0 42320 0 -1 38624
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 42412 0 -1 38624
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 41952 0 1 38624
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_709
timestamp 1586364061
transform 1 0 43240 0 -1 38624
box -38 -48 130 592
use scs8hd_fill_1  FILLER_66_457
timestamp 1586364061
transform 1 0 43148 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_459
timestamp 1586364061
transform 1 0 43332 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_471
timestamp 1586364061
transform 1 0 44436 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_66_483
timestamp 1586364061
transform 1 0 45540 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_458
timestamp 1586364061
transform 1 0 43240 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_470
timestamp 1586364061
transform 1 0 44344 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_67_482
timestamp 1586364061
transform 1 0 45448 0 1 38624
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_717
timestamp 1586364061
transform 1 0 46000 0 1 38624
box -38 -48 130 592
use scs8hd_decap_12  FILLER_66_495
timestamp 1586364061
transform 1 0 46644 0 -1 38624
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_66_507
timestamp 1586364061
transform 1 0 47748 0 -1 38624
box -38 -48 774 592
use scs8hd_decap_12  FILLER_67_489
timestamp 1586364061
transform 1 0 46092 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_67_501
timestamp 1586364061
transform 1 0 47196 0 1 38624
box -38 -48 1142 592
use scs8hd_decap_3  PHY_133
timestamp 1586364061
transform -1 0 48852 0 -1 38624
box -38 -48 314 592
use scs8hd_decap_3  PHY_135
timestamp 1586364061
transform -1 0 48852 0 1 38624
box -38 -48 314 592
use scs8hd_fill_1  FILLER_66_515
timestamp 1586364061
transform 1 0 48484 0 -1 38624
box -38 -48 130 592
use scs8hd_decap_3  FILLER_67_513
timestamp 1586364061
transform 1 0 48300 0 1 38624
box -38 -48 314 592
use scs8hd_decap_3  PHY_136
timestamp 1586364061
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_12  FILLER_68_3
timestamp 1586364061
transform 1 0 1380 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_15
timestamp 1586364061
transform 1 0 2484 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_718
timestamp 1586364061
transform 1 0 3956 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_4  FILLER_68_27
timestamp 1586364061
transform 1 0 3588 0 -1 39712
box -38 -48 406 592
use scs8hd_decap_12  FILLER_68_32
timestamp 1586364061
transform 1 0 4048 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_44
timestamp 1586364061
transform 1 0 5152 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_56
timestamp 1586364061
transform 1 0 6256 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_68
timestamp 1586364061
transform 1 0 7360 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_80
timestamp 1586364061
transform 1 0 8464 0 -1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_719
timestamp 1586364061
transform 1 0 9568 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_93
timestamp 1586364061
transform 1 0 9660 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_105
timestamp 1586364061
transform 1 0 10764 0 -1 39712
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 39712
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13248 0 -1 39712
box -38 -48 866 592
use scs8hd_decap_4  FILLER_68_117
timestamp 1586364061
transform 1 0 11868 0 -1 39712
box -38 -48 406 592
use scs8hd_decap_8  FILLER_68_124
timestamp 1586364061
transform 1 0 12512 0 -1 39712
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 -1 39712
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_720
timestamp 1586364061
transform 1 0 15180 0 -1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14536 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_68_141
timestamp 1586364061
transform 1 0 14076 0 -1 39712
box -38 -48 406 592
use scs8hd_fill_1  FILLER_68_145
timestamp 1586364061
transform 1 0 14444 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_4  FILLER_68_148
timestamp 1586364061
transform 1 0 14720 0 -1 39712
box -38 -48 406 592
use scs8hd_fill_1  FILLER_68_152
timestamp 1586364061
transform 1 0 15088 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_3  FILLER_68_154
timestamp 1586364061
transform 1 0 15272 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_4  FILLER_68_160
timestamp 1586364061
transform 1 0 15824 0 -1 39712
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16560 0 -1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 -1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_68_166
timestamp 1586364061
transform 1 0 16376 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_68_177
timestamp 1586364061
transform 1 0 17388 0 -1 39712
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18492 0 -1 39712
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_721
timestamp 1586364061
transform 1 0 20792 0 -1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19688 0 -1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 -1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_68_200
timestamp 1586364061
transform 1 0 19504 0 -1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_68_204
timestamp 1586364061
transform 1 0 19872 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_6  FILLER_68_208
timestamp 1586364061
transform 1 0 20240 0 -1 39712
box -38 -48 590 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21712 0 -1 39712
box -38 -48 866 592
use scs8hd_decap_8  FILLER_68_215
timestamp 1586364061
transform 1 0 20884 0 -1 39712
box -38 -48 774 592
use scs8hd_fill_1  FILLER_68_223
timestamp 1586364061
transform 1 0 21620 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_233
timestamp 1586364061
transform 1 0 22540 0 -1 39712
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_3_in_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 23920 0 -1 39712
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__240__B
timestamp 1586364061
transform 1 0 23644 0 -1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_3_in_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25208 0 -1 39712
box -38 -48 222 592
use scs8hd_fill_1  FILLER_68_247
timestamp 1586364061
transform 1 0 23828 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_3  FILLER_68_259
timestamp 1586364061
transform 1 0 24932 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_8  FILLER_68_264
timestamp 1586364061
transform 1 0 25392 0 -1 39712
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26864 0 -1 39712
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_722
timestamp 1586364061
transform 1 0 26404 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_3  FILLER_68_272
timestamp 1586364061
transform 1 0 26128 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_4  FILLER_68_276
timestamp 1586364061
transform 1 0 26496 0 -1 39712
box -38 -48 406 592
use scs8hd_decap_12  FILLER_68_289
timestamp 1586364061
transform 1 0 27692 0 -1 39712
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  ltile_clb_0.mem_fle_2_in_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 29164 0 -1 39712
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30360 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_68_301
timestamp 1586364061
transform 1 0 28796 0 -1 39712
box -38 -48 406 592
use scs8hd_fill_2  FILLER_68_316
timestamp 1586364061
transform 1 0 30176 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_3  FILLER_68_320
timestamp 1586364061
transform 1 0 30544 0 -1 39712
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31004 0 -1 39712
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32752 0 -1 39712
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_723
timestamp 1586364061
transform 1 0 32016 0 -1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mem_fle_2_in_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30820 0 -1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 32384 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_8  FILLER_68_328
timestamp 1586364061
transform 1 0 31280 0 -1 39712
box -38 -48 774 592
use scs8hd_decap_3  FILLER_68_337
timestamp 1586364061
transform 1 0 32108 0 -1 39712
box -38 -48 314 592
use scs8hd_fill_2  FILLER_68_342
timestamp 1586364061
transform 1 0 32568 0 -1 39712
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34316 0 -1 39712
box -38 -48 314 592
use scs8hd_decap_8  FILLER_68_353
timestamp 1586364061
transform 1 0 33580 0 -1 39712
box -38 -48 774 592
use scs8hd_decap_12  FILLER_68_364
timestamp 1586364061
transform 1 0 34592 0 -1 39712
box -38 -48 1142 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36064 0 -1 39712
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_724
timestamp 1586364061
transform 1 0 37628 0 -1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35880 0 -1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_68_376
timestamp 1586364061
transform 1 0 35696 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_8  FILLER_68_389
timestamp 1586364061
transform 1 0 36892 0 -1 39712
box -38 -48 774 592
use scs8hd_decap_8  FILLER_68_398
timestamp 1586364061
transform 1 0 37720 0 -1 39712
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 40572 0 -1 39712
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38640 0 -1 39712
box -38 -48 866 592
use scs8hd_fill_2  FILLER_68_406
timestamp 1586364061
transform 1 0 38456 0 -1 39712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_68_417
timestamp 1586364061
transform 1 0 39468 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_432
timestamp 1586364061
transform 1 0 40848 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_444
timestamp 1586364061
transform 1 0 41952 0 -1 39712
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_68_456
timestamp 1586364061
transform 1 0 43056 0 -1 39712
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_725
timestamp 1586364061
transform 1 0 43240 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_68_459
timestamp 1586364061
transform 1 0 43332 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_471
timestamp 1586364061
transform 1 0 44436 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_483
timestamp 1586364061
transform 1 0 45540 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_68_495
timestamp 1586364061
transform 1 0 46644 0 -1 39712
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_68_507
timestamp 1586364061
transform 1 0 47748 0 -1 39712
box -38 -48 774 592
use scs8hd_decap_3  PHY_137
timestamp 1586364061
transform -1 0 48852 0 -1 39712
box -38 -48 314 592
use scs8hd_fill_1  FILLER_68_515
timestamp 1586364061
transform 1 0 48484 0 -1 39712
box -38 -48 130 592
use scs8hd_decap_3  PHY_138
timestamp 1586364061
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use scs8hd_decap_12  FILLER_69_3
timestamp 1586364061
transform 1 0 1380 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_15
timestamp 1586364061
transform 1 0 2484 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_27
timestamp 1586364061
transform 1 0 3588 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_39
timestamp 1586364061
transform 1 0 4692 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_69_51
timestamp 1586364061
transform 1 0 5796 0 1 39712
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_726
timestamp 1586364061
transform 1 0 6716 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_59
timestamp 1586364061
transform 1 0 6532 0 1 39712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_69_62
timestamp 1586364061
transform 1 0 6808 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_74
timestamp 1586364061
transform 1 0 7912 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_86
timestamp 1586364061
transform 1 0 9016 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_98
timestamp 1586364061
transform 1 0 10120 0 1 39712
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12880 0 1 39712
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_727
timestamp 1586364061
transform 1 0 12328 0 1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13340 0 1 39712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_69_110
timestamp 1586364061
transform 1 0 11224 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_69_123
timestamp 1586364061
transform 1 0 12420 0 1 39712
box -38 -48 406 592
use scs8hd_fill_1  FILLER_69_127
timestamp 1586364061
transform 1 0 12788 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_131
timestamp 1586364061
transform 1 0 13156 0 1 39712
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14536 0 1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 39712
box -38 -48 222 592
use scs8hd_decap_6  FILLER_69_135
timestamp 1586364061
transform 1 0 13524 0 1 39712
box -38 -48 590 592
use scs8hd_fill_1  FILLER_69_141
timestamp 1586364061
transform 1 0 14076 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_144
timestamp 1586364061
transform 1 0 14352 0 1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_69_155
timestamp 1586364061
transform 1 0 15364 0 1 39712
box -38 -48 406 592
use scs8hd_fill_1  FILLER_69_159
timestamp 1586364061
transform 1 0 15732 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_162
timestamp 1586364061
transform 1 0 16008 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 39712
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 39712
box -38 -48 866 592
use scs8hd_fill_2  FILLER_69_179
timestamp 1586364061
transform 1 0 17572 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_175
timestamp 1586364061
transform 1 0 17204 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_184
timestamp 1586364061
transform 1 0 18032 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 39712
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_728
timestamp 1586364061
transform 1 0 17940 0 1 39712
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 1 39712
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18676 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20700 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_189
timestamp 1586364061
transform 1 0 18492 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_193
timestamp 1586364061
transform 1 0 18860 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_206
timestamp 1586364061
transform 1 0 20056 0 1 39712
box -38 -48 222 592
use scs8hd_decap_3  FILLER_69_210
timestamp 1586364061
transform 1 0 20424 0 1 39712
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21620 0 1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23184 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21068 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22632 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_215
timestamp 1586364061
transform 1 0 20884 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_219
timestamp 1586364061
transform 1 0 21252 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_232
timestamp 1586364061
transform 1 0 22448 0 1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_69_236
timestamp 1586364061
transform 1 0 22816 0 1 39712
box -38 -48 406 592
use scs8hd_fill_2  FILLER_69_251
timestamp 1586364061
transform 1 0 24196 0 1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_69_245
timestamp 1586364061
transform 1 0 23644 0 1 39712
box -38 -48 406 592
use scs8hd_fill_2  FILLER_69_242
timestamp 1586364061
transform 1 0 23368 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24012 0 1 39712
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_729
timestamp 1586364061
transform 1 0 23552 0 1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24380 0 1 39712
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24564 0 1 39712
box -38 -48 866 592
use scs8hd_fill_2  FILLER_69_268
timestamp 1586364061
transform 1 0 25760 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_264
timestamp 1586364061
transform 1 0 25392 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25576 0 1 39712
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26864 0 1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26680 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26312 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25944 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27876 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_272
timestamp 1586364061
transform 1 0 26128 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_276
timestamp 1586364061
transform 1 0 26496 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_289
timestamp 1586364061
transform 1 0 27692 0 1 39712
box -38 -48 222 592
use scs8hd_decap_8  FILLER_69_293
timestamp 1586364061
transform 1 0 28060 0 1 39712
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29992 0 1 39712
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_730
timestamp 1586364061
transform 1 0 29164 0 1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28980 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29808 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29440 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_301
timestamp 1586364061
transform 1 0 28796 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_306
timestamp 1586364061
transform 1 0 29256 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_310
timestamp 1586364061
transform 1 0 29624 0 1 39712
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32476 0 1 39712
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 32292 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31924 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31004 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31556 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_323
timestamp 1586364061
transform 1 0 30820 0 1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_69_327
timestamp 1586364061
transform 1 0 31188 0 1 39712
box -38 -48 406 592
use scs8hd_fill_2  FILLER_69_333
timestamp 1586364061
transform 1 0 31740 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_337
timestamp 1586364061
transform 1 0 32108 0 1 39712
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_731
timestamp 1586364061
transform 1 0 34776 0 1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35052 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33948 0 1 39712
box -38 -48 222 592
use scs8hd_decap_6  FILLER_69_350
timestamp 1586364061
transform 1 0 33304 0 1 39712
box -38 -48 590 592
use scs8hd_fill_1  FILLER_69_356
timestamp 1586364061
transform 1 0 33856 0 1 39712
box -38 -48 130 592
use scs8hd_decap_6  FILLER_69_359
timestamp 1586364061
transform 1 0 34132 0 1 39712
box -38 -48 590 592
use scs8hd_fill_1  FILLER_69_365
timestamp 1586364061
transform 1 0 34684 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_367
timestamp 1586364061
transform 1 0 34868 0 1 39712
box -38 -48 222 592
use scs8hd_decap_6  FILLER_69_371
timestamp 1586364061
transform 1 0 35236 0 1 39712
box -38 -48 590 592
use scs8hd_nor2_4  _280_
timestamp 1586364061
transform 1 0 36984 0 1 39712
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35788 0 1 39712
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36248 0 1 39712
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__280__A
timestamp 1586364061
transform 1 0 36800 0 1 39712
box -38 -48 222 592
use scs8hd_fill_2  FILLER_69_380
timestamp 1586364061
transform 1 0 36064 0 1 39712
box -38 -48 222 592
use scs8hd_decap_4  FILLER_69_384
timestamp 1586364061
transform 1 0 36432 0 1 39712
box -38 -48 406 592
use scs8hd_decap_4  FILLER_69_399
timestamp 1586364061
transform 1 0 37812 0 1 39712
box -38 -48 406 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 38640 0 1 39712
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_732
timestamp 1586364061
transform 1 0 40388 0 1 39712
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 38272 0 1 39712
box -38 -48 222 592
use scs8hd_fill_1  FILLER_69_403
timestamp 1586364061
transform 1 0 38180 0 1 39712
box -38 -48 130 592
use scs8hd_fill_2  FILLER_69_406
timestamp 1586364061
transform 1 0 38456 0 1 39712
box -38 -48 222 592
use scs8hd_decap_8  FILLER_69_417
timestamp 1586364061
transform 1 0 39468 0 1 39712
box -38 -48 774 592
use scs8hd_fill_2  FILLER_69_425
timestamp 1586364061
transform 1 0 40204 0 1 39712
box -38 -48 222 592
use scs8hd_decap_12  FILLER_69_428
timestamp 1586364061
transform 1 0 40480 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_440
timestamp 1586364061
transform 1 0 41584 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_452
timestamp 1586364061
transform 1 0 42688 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_464
timestamp 1586364061
transform 1 0 43792 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_476
timestamp 1586364061
transform 1 0 44896 0 1 39712
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_733
timestamp 1586364061
transform 1 0 46000 0 1 39712
box -38 -48 130 592
use scs8hd_decap_12  FILLER_69_489
timestamp 1586364061
transform 1 0 46092 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_69_501
timestamp 1586364061
transform 1 0 47196 0 1 39712
box -38 -48 1142 592
use scs8hd_decap_3  PHY_139
timestamp 1586364061
transform -1 0 48852 0 1 39712
box -38 -48 314 592
use scs8hd_decap_3  FILLER_69_513
timestamp 1586364061
transform 1 0 48300 0 1 39712
box -38 -48 314 592
use scs8hd_decap_3  PHY_140
timestamp 1586364061
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_70_3
timestamp 1586364061
transform 1 0 1380 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_15
timestamp 1586364061
transform 1 0 2484 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_734
timestamp 1586364061
transform 1 0 3956 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_4  FILLER_70_27
timestamp 1586364061
transform 1 0 3588 0 -1 40800
box -38 -48 406 592
use scs8hd_decap_12  FILLER_70_32
timestamp 1586364061
transform 1 0 4048 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_44
timestamp 1586364061
transform 1 0 5152 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_56
timestamp 1586364061
transform 1 0 6256 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_68
timestamp 1586364061
transform 1 0 7360 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_80
timestamp 1586364061
transform 1 0 8464 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_735
timestamp 1586364061
transform 1 0 9568 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_70_93
timestamp 1586364061
transform 1 0 9660 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_105
timestamp 1586364061
transform 1 0 10764 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_117
timestamp 1586364061
transform 1 0 11868 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_129
timestamp 1586364061
transform 1 0 12972 0 -1 40800
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 40800
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_736
timestamp 1586364061
transform 1 0 15180 0 -1 40800
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_1  FILLER_70_141
timestamp 1586364061
transform 1 0 14076 0 -1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_70_145
timestamp 1586364061
transform 1 0 14444 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_4  FILLER_70_149
timestamp 1586364061
transform 1 0 14812 0 -1 40800
box -38 -48 406 592
use scs8hd_decap_8  FILLER_70_154
timestamp 1586364061
transform 1 0 15272 0 -1 40800
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 -1 40800
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16468 0 -1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_3  FILLER_70_162
timestamp 1586364061
transform 1 0 16008 0 -1 40800
box -38 -48 314 592
use scs8hd_decap_8  FILLER_70_176
timestamp 1586364061
transform 1 0 17296 0 -1 40800
box -38 -48 774 592
use scs8hd_decap_8  FILLER_70_187
timestamp 1586364061
transform 1 0 18308 0 -1 40800
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 40800
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_737
timestamp 1586364061
transform 1 0 20792 0 -1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_70_195
timestamp 1586364061
transform 1 0 19044 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_8  FILLER_70_206
timestamp 1586364061
transform 1 0 20056 0 -1 40800
box -38 -48 774 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23184 0 -1 40800
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21620 0 -1 40800
box -38 -48 866 592
use scs8hd_decap_8  FILLER_70_215
timestamp 1586364061
transform 1 0 20884 0 -1 40800
box -38 -48 774 592
use scs8hd_decap_8  FILLER_70_232
timestamp 1586364061
transform 1 0 22448 0 -1 40800
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 -1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24564 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_70_243
timestamp 1586364061
transform 1 0 23460 0 -1 40800
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_70_257
timestamp 1586364061
transform 1 0 24748 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_8  FILLER_70_267
timestamp 1586364061
transform 1 0 25668 0 -1 40800
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26864 0 -1 40800
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_738
timestamp 1586364061
transform 1 0 26404 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_4  FILLER_70_276
timestamp 1586364061
transform 1 0 26496 0 -1 40800
box -38 -48 406 592
use scs8hd_decap_12  FILLER_70_289
timestamp 1586364061
transform 1 0 27692 0 -1 40800
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 28980 0 -1 40800
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29992 0 -1 40800
box -38 -48 866 592
use scs8hd_fill_2  FILLER_70_301
timestamp 1586364061
transform 1 0 28796 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_8  FILLER_70_306
timestamp 1586364061
transform 1 0 29256 0 -1 40800
box -38 -48 774 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32384 0 -1 40800
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_739
timestamp 1586364061
transform 1 0 32016 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_70_323
timestamp 1586364061
transform 1 0 30820 0 -1 40800
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_70_335
timestamp 1586364061
transform 1 0 31924 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_3  FILLER_70_337
timestamp 1586364061
transform 1 0 32108 0 -1 40800
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_10_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34960 0 -1 40800
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_13_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33948 0 -1 40800
box -38 -48 314 592
use scs8hd_decap_8  FILLER_70_349
timestamp 1586364061
transform 1 0 33212 0 -1 40800
box -38 -48 774 592
use scs8hd_decap_8  FILLER_70_360
timestamp 1586364061
transform 1 0 34224 0 -1 40800
box -38 -48 774 592
use scs8hd_decap_12  FILLER_70_371
timestamp 1586364061
transform 1 0 35236 0 -1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_740
timestamp 1586364061
transform 1 0 37628 0 -1 40800
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__280__B
timestamp 1586364061
transform 1 0 36984 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_6  FILLER_70_383
timestamp 1586364061
transform 1 0 36340 0 -1 40800
box -38 -48 590 592
use scs8hd_fill_1  FILLER_70_389
timestamp 1586364061
transform 1 0 36892 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_4  FILLER_70_392
timestamp 1586364061
transform 1 0 37168 0 -1 40800
box -38 -48 406 592
use scs8hd_fill_1  FILLER_70_396
timestamp 1586364061
transform 1 0 37536 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_6  FILLER_70_398
timestamp 1586364061
transform 1 0 37720 0 -1 40800
box -38 -48 590 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 38272 0 -1 40800
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 38732 0 -1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 39100 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_70_407
timestamp 1586364061
transform 1 0 38548 0 -1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_70_411
timestamp 1586364061
transform 1 0 38916 0 -1 40800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_70_415
timestamp 1586364061
transform 1 0 39284 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_427
timestamp 1586364061
transform 1 0 40388 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_439
timestamp 1586364061
transform 1 0 41492 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_70_451
timestamp 1586364061
transform 1 0 42596 0 -1 40800
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_741
timestamp 1586364061
transform 1 0 43240 0 -1 40800
box -38 -48 130 592
use scs8hd_fill_1  FILLER_70_457
timestamp 1586364061
transform 1 0 43148 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_70_459
timestamp 1586364061
transform 1 0 43332 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_471
timestamp 1586364061
transform 1 0 44436 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_483
timestamp 1586364061
transform 1 0 45540 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_70_495
timestamp 1586364061
transform 1 0 46644 0 -1 40800
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_70_507
timestamp 1586364061
transform 1 0 47748 0 -1 40800
box -38 -48 774 592
use scs8hd_decap_3  PHY_141
timestamp 1586364061
transform -1 0 48852 0 -1 40800
box -38 -48 314 592
use scs8hd_fill_1  FILLER_70_515
timestamp 1586364061
transform 1 0 48484 0 -1 40800
box -38 -48 130 592
use scs8hd_decap_3  PHY_142
timestamp 1586364061
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use scs8hd_decap_12  FILLER_71_3
timestamp 1586364061
transform 1 0 1380 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_15
timestamp 1586364061
transform 1 0 2484 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_27
timestamp 1586364061
transform 1 0 3588 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_39
timestamp 1586364061
transform 1 0 4692 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_71_51
timestamp 1586364061
transform 1 0 5796 0 1 40800
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_742
timestamp 1586364061
transform 1 0 6716 0 1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_71_59
timestamp 1586364061
transform 1 0 6532 0 1 40800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_71_62
timestamp 1586364061
transform 1 0 6808 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_74
timestamp 1586364061
transform 1 0 7912 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_86
timestamp 1586364061
transform 1 0 9016 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_98
timestamp 1586364061
transform 1 0 10120 0 1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_743
timestamp 1586364061
transform 1 0 12328 0 1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_71_110
timestamp 1586364061
transform 1 0 11224 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_123
timestamp 1586364061
transform 1 0 12420 0 1 40800
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14352 0 1 40800
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 1 40800
box -38 -48 222 592
use scs8hd_decap_8  FILLER_71_135
timestamp 1586364061
transform 1 0 13524 0 1 40800
box -38 -48 774 592
use scs8hd_fill_1  FILLER_71_143
timestamp 1586364061
transform 1 0 14260 0 1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_71_147
timestamp 1586364061
transform 1 0 14628 0 1 40800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_71_151
timestamp 1586364061
transform 1 0 14996 0 1 40800
box -38 -48 1142 592
use scs8hd_nor2_4  _231_
timestamp 1586364061
transform 1 0 16376 0 1 40800
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 1 40800
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_744
timestamp 1586364061
transform 1 0 17940 0 1 40800
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 16192 0 1 40800
box -38 -48 222 592
use scs8hd_fill_1  FILLER_71_163
timestamp 1586364061
transform 1 0 16100 0 1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_71_175
timestamp 1586364061
transform 1 0 17204 0 1 40800
box -38 -48 222 592
use scs8hd_decap_4  FILLER_71_179
timestamp 1586364061
transform 1 0 17572 0 1 40800
box -38 -48 406 592
use scs8hd_fill_2  FILLER_71_184
timestamp 1586364061
transform 1 0 18032 0 1 40800
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18676 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19044 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_189
timestamp 1586364061
transform 1 0 18492 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_193
timestamp 1586364061
transform 1 0 18860 0 1 40800
box -38 -48 222 592
use scs8hd_decap_6  FILLER_71_206
timestamp 1586364061
transform 1 0 20056 0 1 40800
box -38 -48 590 592
use scs8hd_fill_2  FILLER_71_214
timestamp 1586364061
transform 1 0 20792 0 1 40800
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 1 40800
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22540 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_218
timestamp 1586364061
transform 1 0 21160 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_231
timestamp 1586364061
transform 1 0 22356 0 1 40800
box -38 -48 222 592
use scs8hd_decap_6  FILLER_71_235
timestamp 1586364061
transform 1 0 22724 0 1 40800
box -38 -48 590 592
use scs8hd_fill_1  FILLER_71_241
timestamp 1586364061
transform 1 0 23276 0 1 40800
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 40800
box -38 -48 314 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24840 0 1 40800
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_745
timestamp 1586364061
transform 1 0 23552 0 1 40800
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24196 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 40800
box -38 -48 222 592
use scs8hd_decap_3  FILLER_71_248
timestamp 1586364061
transform 1 0 23920 0 1 40800
box -38 -48 314 592
use scs8hd_decap_3  FILLER_71_253
timestamp 1586364061
transform 1 0 24380 0 1 40800
box -38 -48 314 592
use scs8hd_fill_2  FILLER_71_267
timestamp 1586364061
transform 1 0 25668 0 1 40800
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26588 0 1 40800
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25852 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27048 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27416 0 1 40800
box -38 -48 222 592
use scs8hd_decap_6  FILLER_71_271
timestamp 1586364061
transform 1 0 26036 0 1 40800
box -38 -48 590 592
use scs8hd_fill_2  FILLER_71_280
timestamp 1586364061
transform 1 0 26864 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_284
timestamp 1586364061
transform 1 0 27232 0 1 40800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_71_288
timestamp 1586364061
transform 1 0 27600 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_71_300
timestamp 1586364061
transform 1 0 28704 0 1 40800
box -38 -48 406 592
use scs8hd_decap_4  FILLER_71_306
timestamp 1586364061
transform 1 0 29256 0 1 40800
box -38 -48 406 592
use scs8hd_fill_1  FILLER_71_304
timestamp 1586364061
transform 1 0 29072 0 1 40800
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_746
timestamp 1586364061
transform 1 0 29164 0 1 40800
box -38 -48 130 592
use scs8hd_fill_2  FILLER_71_313
timestamp 1586364061
transform 1 0 29900 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30084 0 1 40800
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29624 0 1 40800
box -38 -48 314 592
use scs8hd_decap_6  FILLER_71_321
timestamp 1586364061
transform 1 0 30636 0 1 40800
box -38 -48 590 592
use scs8hd_fill_2  FILLER_71_317
timestamp 1586364061
transform 1 0 30268 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30452 0 1 40800
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31188 0 1 40800
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32200 0 1 40800
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31648 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32660 0 1 40800
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_8_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33028 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_330
timestamp 1586364061
transform 1 0 31464 0 1 40800
box -38 -48 222 592
use scs8hd_decap_4  FILLER_71_334
timestamp 1586364061
transform 1 0 31832 0 1 40800
box -38 -48 406 592
use scs8hd_fill_2  FILLER_71_341
timestamp 1586364061
transform 1 0 32476 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_345
timestamp 1586364061
transform 1 0 32844 0 1 40800
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33212 0 1 40800
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_747
timestamp 1586364061
transform 1 0 34776 0 1 40800
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_2_in_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33672 0 1 40800
box -38 -48 222 592
use scs8hd_fill_2  FILLER_71_352
timestamp 1586364061
transform 1 0 33488 0 1 40800
box -38 -48 222 592
use scs8hd_decap_8  FILLER_71_356
timestamp 1586364061
transform 1 0 33856 0 1 40800
box -38 -48 774 592
use scs8hd_fill_2  FILLER_71_364
timestamp 1586364061
transform 1 0 34592 0 1 40800
box -38 -48 222 592
use scs8hd_decap_12  FILLER_71_367
timestamp 1586364061
transform 1 0 34868 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_379
timestamp 1586364061
transform 1 0 35972 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_391
timestamp 1586364061
transform 1 0 37076 0 1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_748
timestamp 1586364061
transform 1 0 40388 0 1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_71_403
timestamp 1586364061
transform 1 0 38180 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_415
timestamp 1586364061
transform 1 0 39284 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_428
timestamp 1586364061
transform 1 0 40480 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_440
timestamp 1586364061
transform 1 0 41584 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_452
timestamp 1586364061
transform 1 0 42688 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_464
timestamp 1586364061
transform 1 0 43792 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_476
timestamp 1586364061
transform 1 0 44896 0 1 40800
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_749
timestamp 1586364061
transform 1 0 46000 0 1 40800
box -38 -48 130 592
use scs8hd_decap_12  FILLER_71_489
timestamp 1586364061
transform 1 0 46092 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_71_501
timestamp 1586364061
transform 1 0 47196 0 1 40800
box -38 -48 1142 592
use scs8hd_decap_3  PHY_143
timestamp 1586364061
transform -1 0 48852 0 1 40800
box -38 -48 314 592
use scs8hd_decap_3  FILLER_71_513
timestamp 1586364061
transform 1 0 48300 0 1 40800
box -38 -48 314 592
use scs8hd_decap_3  PHY_144
timestamp 1586364061
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use scs8hd_decap_3  PHY_146
timestamp 1586364061
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use scs8hd_decap_12  FILLER_72_3
timestamp 1586364061
transform 1 0 1380 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_15
timestamp 1586364061
transform 1 0 2484 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_3
timestamp 1586364061
transform 1 0 1380 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_15
timestamp 1586364061
transform 1 0 2484 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_750
timestamp 1586364061
transform 1 0 3956 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_4  FILLER_72_27
timestamp 1586364061
transform 1 0 3588 0 -1 41888
box -38 -48 406 592
use scs8hd_decap_12  FILLER_72_32
timestamp 1586364061
transform 1 0 4048 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_44
timestamp 1586364061
transform 1 0 5152 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_27
timestamp 1586364061
transform 1 0 3588 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_39
timestamp 1586364061
transform 1 0 4692 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_73_51
timestamp 1586364061
transform 1 0 5796 0 1 41888
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_758
timestamp 1586364061
transform 1 0 6716 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_56
timestamp 1586364061
transform 1 0 6256 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_68
timestamp 1586364061
transform 1 0 7360 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_80
timestamp 1586364061
transform 1 0 8464 0 -1 41888
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_73_59
timestamp 1586364061
transform 1 0 6532 0 1 41888
box -38 -48 222 592
use scs8hd_decap_12  FILLER_73_62
timestamp 1586364061
transform 1 0 6808 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_74
timestamp 1586364061
transform 1 0 7912 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_751
timestamp 1586364061
transform 1 0 9568 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_93
timestamp 1586364061
transform 1 0 9660 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_105
timestamp 1586364061
transform 1 0 10764 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_86
timestamp 1586364061
transform 1 0 9016 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_98
timestamp 1586364061
transform 1 0 10120 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_759
timestamp 1586364061
transform 1 0 12328 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_117
timestamp 1586364061
transform 1 0 11868 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_129
timestamp 1586364061
transform 1 0 12972 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_110
timestamp 1586364061
transform 1 0 11224 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_123
timestamp 1586364061
transform 1 0 12420 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_752
timestamp 1586364061
transform 1 0 15180 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_141
timestamp 1586364061
transform 1 0 14076 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_154
timestamp 1586364061
transform 1 0 15272 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_135
timestamp 1586364061
transform 1 0 13524 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_147
timestamp 1586364061
transform 1 0 14628 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_159
timestamp 1586364061
transform 1 0 15732 0 1 41888
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_2.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 -1 41888
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_760
timestamp 1586364061
transform 1 0 17940 0 1 41888
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__231__B
timestamp 1586364061
transform 1 0 16376 0 -1 41888
box -38 -48 222 592
use scs8hd_decap_12  FILLER_72_171
timestamp 1586364061
transform 1 0 16836 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_72_183
timestamp 1586364061
transform 1 0 17940 0 -1 41888
box -38 -48 774 592
use scs8hd_decap_12  FILLER_73_171
timestamp 1586364061
transform 1 0 16836 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_184
timestamp 1586364061
transform 1 0 18032 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_196
timestamp 1586364061
transform 1 0 19136 0 1 41888
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_72_200
timestamp 1586364061
transform 1 0 19504 0 -1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_72_196
timestamp 1586364061
transform 1 0 19136 0 -1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_72_191
timestamp 1586364061
transform 1 0 18676 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 -1 41888
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18860 0 -1 41888
box -38 -48 314 592
use scs8hd_decap_12  FILLER_73_208
timestamp 1586364061
transform 1 0 20240 0 1 41888
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_72_212
timestamp 1586364061
transform 1 0 20608 0 -1 41888
box -38 -48 222 592
use scs8hd_decap_8  FILLER_72_204
timestamp 1586364061
transform 1 0 19872 0 -1 41888
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 -1 41888
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_753
timestamp 1586364061
transform 1 0 20792 0 -1 41888
box -38 -48 130 592
use scs8hd_fill_2  FILLER_73_227
timestamp 1586364061
transform 1 0 21988 0 1 41888
box -38 -48 222 592
use scs8hd_fill_2  FILLER_73_223
timestamp 1586364061
transform 1 0 21620 0 1 41888
box -38 -48 222 592
use scs8hd_fill_1  FILLER_72_221
timestamp 1586364061
transform 1 0 21436 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_6  FILLER_72_215
timestamp 1586364061
transform 1 0 20884 0 -1 41888
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21804 0 1 41888
box -38 -48 222 592
use scs8hd_ebufn_2  ltile_clb_0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 -1 41888
box -38 -48 866 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21344 0 1 41888
box -38 -48 314 592
use scs8hd_decap_12  FILLER_73_231
timestamp 1586364061
transform 1 0 22356 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_231
timestamp 1586364061
transform 1 0 22356 0 -1 41888
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22172 0 1 41888
box -38 -48 222 592
use scs8hd_decap_8  FILLER_73_245
timestamp 1586364061
transform 1 0 23644 0 1 41888
box -38 -48 774 592
use scs8hd_fill_1  FILLER_73_243
timestamp 1586364061
transform 1 0 23460 0 1 41888
box -38 -48 130 592
use scs8hd_decap_4  FILLER_72_254
timestamp 1586364061
transform 1 0 24472 0 -1 41888
box -38 -48 406 592
use scs8hd_decap_8  FILLER_72_243
timestamp 1586364061
transform 1 0 23460 0 -1 41888
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_761
timestamp 1586364061
transform 1 0 23552 0 1 41888
box -38 -48 130 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24380 0 1 41888
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24196 0 -1 41888
box -38 -48 314 592
use scs8hd_decap_12  FILLER_73_260
timestamp 1586364061
transform 1 0 25024 0 1 41888
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_73_256
timestamp 1586364061
transform 1 0 24656 0 1 41888
box -38 -48 222 592
use scs8hd_decap_8  FILLER_72_265
timestamp 1586364061
transform 1 0 25484 0 -1 41888
box -38 -48 774 592
use scs8hd_fill_2  FILLER_72_260
timestamp 1586364061
transform 1 0 25024 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24840 0 -1 41888
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_ltile_clb_0.mux_fle_3_in_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24840 0 1 41888
box -38 -48 222 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25208 0 -1 41888
box -38 -48 314 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_1.INVTX1_8_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26588 0 -1 41888
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_754
timestamp 1586364061
transform 1 0 26404 0 -1 41888
box -38 -48 130 592
use scs8hd_fill_2  FILLER_72_273
timestamp 1586364061
transform 1 0 26220 0 -1 41888
box -38 -48 222 592
use scs8hd_fill_1  FILLER_72_276
timestamp 1586364061
transform 1 0 26496 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_280
timestamp 1586364061
transform 1 0 26864 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_292
timestamp 1586364061
transform 1 0 27968 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_272
timestamp 1586364061
transform 1 0 26128 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_284
timestamp 1586364061
transform 1 0 27232 0 1 41888
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_11_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29624 0 -1 41888
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_762
timestamp 1586364061
transform 1 0 29164 0 1 41888
box -38 -48 130 592
use scs8hd_decap_6  FILLER_72_304
timestamp 1586364061
transform 1 0 29072 0 -1 41888
box -38 -48 590 592
use scs8hd_decap_12  FILLER_72_313
timestamp 1586364061
transform 1 0 29900 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_73_296
timestamp 1586364061
transform 1 0 28336 0 1 41888
box -38 -48 774 592
use scs8hd_fill_1  FILLER_73_304
timestamp 1586364061
transform 1 0 29072 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_73_306
timestamp 1586364061
transform 1 0 29256 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_318
timestamp 1586364061
transform 1 0 30360 0 1 41888
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_2_in_0.INVTX1_12_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32476 0 -1 41888
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_755
timestamp 1586364061
transform 1 0 32016 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_8  FILLER_72_325
timestamp 1586364061
transform 1 0 31004 0 -1 41888
box -38 -48 774 592
use scs8hd_decap_3  FILLER_72_333
timestamp 1586364061
transform 1 0 31740 0 -1 41888
box -38 -48 314 592
use scs8hd_decap_4  FILLER_72_337
timestamp 1586364061
transform 1 0 32108 0 -1 41888
box -38 -48 406 592
use scs8hd_decap_12  FILLER_72_344
timestamp 1586364061
transform 1 0 32752 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_330
timestamp 1586364061
transform 1 0 31464 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_342
timestamp 1586364061
transform 1 0 32568 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_763
timestamp 1586364061
transform 1 0 34776 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_356
timestamp 1586364061
transform 1 0 33856 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_368
timestamp 1586364061
transform 1 0 34960 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_354
timestamp 1586364061
transform 1 0 33672 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_367
timestamp 1586364061
transform 1 0 34868 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_756
timestamp 1586364061
transform 1 0 37628 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_380
timestamp 1586364061
transform 1 0 36064 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_72_392
timestamp 1586364061
transform 1 0 37168 0 -1 41888
box -38 -48 406 592
use scs8hd_fill_1  FILLER_72_396
timestamp 1586364061
transform 1 0 37536 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_398
timestamp 1586364061
transform 1 0 37720 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_379
timestamp 1586364061
transform 1 0 35972 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_391
timestamp 1586364061
transform 1 0 37076 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_764
timestamp 1586364061
transform 1 0 40388 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_410
timestamp 1586364061
transform 1 0 38824 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_422
timestamp 1586364061
transform 1 0 39928 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_403
timestamp 1586364061
transform 1 0 38180 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_415
timestamp 1586364061
transform 1 0 39284 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_428
timestamp 1586364061
transform 1 0 40480 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_434
timestamp 1586364061
transform 1 0 41032 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_446
timestamp 1586364061
transform 1 0 42136 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_440
timestamp 1586364061
transform 1 0 41584 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_452
timestamp 1586364061
transform 1 0 42688 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_757
timestamp 1586364061
transform 1 0 43240 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_459
timestamp 1586364061
transform 1 0 43332 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_471
timestamp 1586364061
transform 1 0 44436 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_72_483
timestamp 1586364061
transform 1 0 45540 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_464
timestamp 1586364061
transform 1 0 43792 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_476
timestamp 1586364061
transform 1 0 44896 0 1 41888
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_765
timestamp 1586364061
transform 1 0 46000 0 1 41888
box -38 -48 130 592
use scs8hd_decap_12  FILLER_72_495
timestamp 1586364061
transform 1 0 46644 0 -1 41888
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_72_507
timestamp 1586364061
transform 1 0 47748 0 -1 41888
box -38 -48 774 592
use scs8hd_decap_12  FILLER_73_489
timestamp 1586364061
transform 1 0 46092 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_73_501
timestamp 1586364061
transform 1 0 47196 0 1 41888
box -38 -48 1142 592
use scs8hd_decap_3  PHY_145
timestamp 1586364061
transform -1 0 48852 0 -1 41888
box -38 -48 314 592
use scs8hd_decap_3  PHY_147
timestamp 1586364061
transform -1 0 48852 0 1 41888
box -38 -48 314 592
use scs8hd_fill_1  FILLER_72_515
timestamp 1586364061
transform 1 0 48484 0 -1 41888
box -38 -48 130 592
use scs8hd_decap_3  FILLER_73_513
timestamp 1586364061
transform 1 0 48300 0 1 41888
box -38 -48 314 592
use scs8hd_decap_3  PHY_148
timestamp 1586364061
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_74_3
timestamp 1586364061
transform 1 0 1380 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_15
timestamp 1586364061
transform 1 0 2484 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_766
timestamp 1586364061
transform 1 0 3956 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_4  FILLER_74_27
timestamp 1586364061
transform 1 0 3588 0 -1 42976
box -38 -48 406 592
use scs8hd_decap_12  FILLER_74_32
timestamp 1586364061
transform 1 0 4048 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_44
timestamp 1586364061
transform 1 0 5152 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_56
timestamp 1586364061
transform 1 0 6256 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_68
timestamp 1586364061
transform 1 0 7360 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_80
timestamp 1586364061
transform 1 0 8464 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_767
timestamp 1586364061
transform 1 0 9568 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_93
timestamp 1586364061
transform 1 0 9660 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_105
timestamp 1586364061
transform 1 0 10764 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_117
timestamp 1586364061
transform 1 0 11868 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_129
timestamp 1586364061
transform 1 0 12972 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_768
timestamp 1586364061
transform 1 0 15180 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_141
timestamp 1586364061
transform 1 0 14076 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_154
timestamp 1586364061
transform 1 0 15272 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_166
timestamp 1586364061
transform 1 0 16376 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_178
timestamp 1586364061
transform 1 0 17480 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_769
timestamp 1586364061
transform 1 0 20792 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_190
timestamp 1586364061
transform 1 0 18584 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_202
timestamp 1586364061
transform 1 0 19688 0 -1 42976
box -38 -48 1142 592
use scs8hd_inv_1  ltile_clb_0.mux_fle_3_in_0.INVTX1_9_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21252 0 -1 42976
box -38 -48 314 592
use scs8hd_decap_4  FILLER_74_215
timestamp 1586364061
transform 1 0 20884 0 -1 42976
box -38 -48 406 592
use scs8hd_decap_12  FILLER_74_222
timestamp 1586364061
transform 1 0 21528 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_234
timestamp 1586364061
transform 1 0 22632 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_246
timestamp 1586364061
transform 1 0 23736 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_258
timestamp 1586364061
transform 1 0 24840 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_770
timestamp 1586364061
transform 1 0 26404 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_4  FILLER_74_270
timestamp 1586364061
transform 1 0 25944 0 -1 42976
box -38 -48 406 592
use scs8hd_fill_1  FILLER_74_274
timestamp 1586364061
transform 1 0 26312 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_276
timestamp 1586364061
transform 1 0 26496 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_288
timestamp 1586364061
transform 1 0 27600 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_300
timestamp 1586364061
transform 1 0 28704 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_312
timestamp 1586364061
transform 1 0 29808 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_771
timestamp 1586364061
transform 1 0 32016 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_324
timestamp 1586364061
transform 1 0 30912 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_337
timestamp 1586364061
transform 1 0 32108 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_349
timestamp 1586364061
transform 1 0 33212 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_361
timestamp 1586364061
transform 1 0 34316 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_373
timestamp 1586364061
transform 1 0 35420 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_772
timestamp 1586364061
transform 1 0 37628 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_385
timestamp 1586364061
transform 1 0 36524 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_398
timestamp 1586364061
transform 1 0 37720 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_410
timestamp 1586364061
transform 1 0 38824 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_422
timestamp 1586364061
transform 1 0 39928 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_434
timestamp 1586364061
transform 1 0 41032 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_446
timestamp 1586364061
transform 1 0 42136 0 -1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_773
timestamp 1586364061
transform 1 0 43240 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_74_459
timestamp 1586364061
transform 1 0 43332 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_471
timestamp 1586364061
transform 1 0 44436 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_483
timestamp 1586364061
transform 1 0 45540 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_74_495
timestamp 1586364061
transform 1 0 46644 0 -1 42976
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_74_507
timestamp 1586364061
transform 1 0 47748 0 -1 42976
box -38 -48 774 592
use scs8hd_decap_3  PHY_149
timestamp 1586364061
transform -1 0 48852 0 -1 42976
box -38 -48 314 592
use scs8hd_fill_1  FILLER_74_515
timestamp 1586364061
transform 1 0 48484 0 -1 42976
box -38 -48 130 592
use scs8hd_decap_3  PHY_150
timestamp 1586364061
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use scs8hd_decap_12  FILLER_75_3
timestamp 1586364061
transform 1 0 1380 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_15
timestamp 1586364061
transform 1 0 2484 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_27
timestamp 1586364061
transform 1 0 3588 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_39
timestamp 1586364061
transform 1 0 4692 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_75_51
timestamp 1586364061
transform 1 0 5796 0 1 42976
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_774
timestamp 1586364061
transform 1 0 6716 0 1 42976
box -38 -48 130 592
use scs8hd_fill_2  FILLER_75_59
timestamp 1586364061
transform 1 0 6532 0 1 42976
box -38 -48 222 592
use scs8hd_decap_12  FILLER_75_62
timestamp 1586364061
transform 1 0 6808 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_74
timestamp 1586364061
transform 1 0 7912 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_86
timestamp 1586364061
transform 1 0 9016 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_98
timestamp 1586364061
transform 1 0 10120 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_775
timestamp 1586364061
transform 1 0 12328 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_110
timestamp 1586364061
transform 1 0 11224 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_123
timestamp 1586364061
transform 1 0 12420 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_135
timestamp 1586364061
transform 1 0 13524 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_147
timestamp 1586364061
transform 1 0 14628 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_159
timestamp 1586364061
transform 1 0 15732 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_776
timestamp 1586364061
transform 1 0 17940 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_171
timestamp 1586364061
transform 1 0 16836 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_184
timestamp 1586364061
transform 1 0 18032 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_196
timestamp 1586364061
transform 1 0 19136 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_208
timestamp 1586364061
transform 1 0 20240 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_220
timestamp 1586364061
transform 1 0 21344 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_232
timestamp 1586364061
transform 1 0 22448 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_777
timestamp 1586364061
transform 1 0 23552 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_245
timestamp 1586364061
transform 1 0 23644 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_257
timestamp 1586364061
transform 1 0 24748 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_269
timestamp 1586364061
transform 1 0 25852 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_281
timestamp 1586364061
transform 1 0 26956 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_293
timestamp 1586364061
transform 1 0 28060 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_778
timestamp 1586364061
transform 1 0 29164 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_306
timestamp 1586364061
transform 1 0 29256 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_318
timestamp 1586364061
transform 1 0 30360 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_330
timestamp 1586364061
transform 1 0 31464 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_342
timestamp 1586364061
transform 1 0 32568 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_779
timestamp 1586364061
transform 1 0 34776 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_354
timestamp 1586364061
transform 1 0 33672 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_367
timestamp 1586364061
transform 1 0 34868 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_379
timestamp 1586364061
transform 1 0 35972 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_391
timestamp 1586364061
transform 1 0 37076 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_780
timestamp 1586364061
transform 1 0 40388 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_403
timestamp 1586364061
transform 1 0 38180 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_415
timestamp 1586364061
transform 1 0 39284 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_428
timestamp 1586364061
transform 1 0 40480 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_440
timestamp 1586364061
transform 1 0 41584 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_452
timestamp 1586364061
transform 1 0 42688 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_464
timestamp 1586364061
transform 1 0 43792 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_476
timestamp 1586364061
transform 1 0 44896 0 1 42976
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_781
timestamp 1586364061
transform 1 0 46000 0 1 42976
box -38 -48 130 592
use scs8hd_decap_12  FILLER_75_489
timestamp 1586364061
transform 1 0 46092 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_75_501
timestamp 1586364061
transform 1 0 47196 0 1 42976
box -38 -48 1142 592
use scs8hd_decap_3  PHY_151
timestamp 1586364061
transform -1 0 48852 0 1 42976
box -38 -48 314 592
use scs8hd_decap_3  FILLER_75_513
timestamp 1586364061
transform 1 0 48300 0 1 42976
box -38 -48 314 592
use scs8hd_decap_3  PHY_152
timestamp 1586364061
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_76_3
timestamp 1586364061
transform 1 0 1380 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_15
timestamp 1586364061
transform 1 0 2484 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_782
timestamp 1586364061
transform 1 0 3956 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_4  FILLER_76_27
timestamp 1586364061
transform 1 0 3588 0 -1 44064
box -38 -48 406 592
use scs8hd_decap_12  FILLER_76_32
timestamp 1586364061
transform 1 0 4048 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_44
timestamp 1586364061
transform 1 0 5152 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_56
timestamp 1586364061
transform 1 0 6256 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_68
timestamp 1586364061
transform 1 0 7360 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_80
timestamp 1586364061
transform 1 0 8464 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_783
timestamp 1586364061
transform 1 0 9568 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_93
timestamp 1586364061
transform 1 0 9660 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_105
timestamp 1586364061
transform 1 0 10764 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_117
timestamp 1586364061
transform 1 0 11868 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_129
timestamp 1586364061
transform 1 0 12972 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_784
timestamp 1586364061
transform 1 0 15180 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_141
timestamp 1586364061
transform 1 0 14076 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_154
timestamp 1586364061
transform 1 0 15272 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_166
timestamp 1586364061
transform 1 0 16376 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_178
timestamp 1586364061
transform 1 0 17480 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_785
timestamp 1586364061
transform 1 0 20792 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_190
timestamp 1586364061
transform 1 0 18584 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_202
timestamp 1586364061
transform 1 0 19688 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_215
timestamp 1586364061
transform 1 0 20884 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_227
timestamp 1586364061
transform 1 0 21988 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_239
timestamp 1586364061
transform 1 0 23092 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_251
timestamp 1586364061
transform 1 0 24196 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_263
timestamp 1586364061
transform 1 0 25300 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_786
timestamp 1586364061
transform 1 0 26404 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_276
timestamp 1586364061
transform 1 0 26496 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_288
timestamp 1586364061
transform 1 0 27600 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_300
timestamp 1586364061
transform 1 0 28704 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_312
timestamp 1586364061
transform 1 0 29808 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_787
timestamp 1586364061
transform 1 0 32016 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_324
timestamp 1586364061
transform 1 0 30912 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_337
timestamp 1586364061
transform 1 0 32108 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_349
timestamp 1586364061
transform 1 0 33212 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_361
timestamp 1586364061
transform 1 0 34316 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_373
timestamp 1586364061
transform 1 0 35420 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_788
timestamp 1586364061
transform 1 0 37628 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_385
timestamp 1586364061
transform 1 0 36524 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_398
timestamp 1586364061
transform 1 0 37720 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_410
timestamp 1586364061
transform 1 0 38824 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_422
timestamp 1586364061
transform 1 0 39928 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_434
timestamp 1586364061
transform 1 0 41032 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_446
timestamp 1586364061
transform 1 0 42136 0 -1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_789
timestamp 1586364061
transform 1 0 43240 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_76_459
timestamp 1586364061
transform 1 0 43332 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_471
timestamp 1586364061
transform 1 0 44436 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_483
timestamp 1586364061
transform 1 0 45540 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_76_495
timestamp 1586364061
transform 1 0 46644 0 -1 44064
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_76_507
timestamp 1586364061
transform 1 0 47748 0 -1 44064
box -38 -48 774 592
use scs8hd_decap_3  PHY_153
timestamp 1586364061
transform -1 0 48852 0 -1 44064
box -38 -48 314 592
use scs8hd_fill_1  FILLER_76_515
timestamp 1586364061
transform 1 0 48484 0 -1 44064
box -38 -48 130 592
use scs8hd_decap_3  PHY_154
timestamp 1586364061
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use scs8hd_decap_12  FILLER_77_3
timestamp 1586364061
transform 1 0 1380 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_15
timestamp 1586364061
transform 1 0 2484 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_27
timestamp 1586364061
transform 1 0 3588 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_39
timestamp 1586364061
transform 1 0 4692 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_77_51
timestamp 1586364061
transform 1 0 5796 0 1 44064
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_790
timestamp 1586364061
transform 1 0 6716 0 1 44064
box -38 -48 130 592
use scs8hd_fill_2  FILLER_77_59
timestamp 1586364061
transform 1 0 6532 0 1 44064
box -38 -48 222 592
use scs8hd_decap_12  FILLER_77_62
timestamp 1586364061
transform 1 0 6808 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_74
timestamp 1586364061
transform 1 0 7912 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_86
timestamp 1586364061
transform 1 0 9016 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_98
timestamp 1586364061
transform 1 0 10120 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_791
timestamp 1586364061
transform 1 0 12328 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_110
timestamp 1586364061
transform 1 0 11224 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_123
timestamp 1586364061
transform 1 0 12420 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_135
timestamp 1586364061
transform 1 0 13524 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_147
timestamp 1586364061
transform 1 0 14628 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_159
timestamp 1586364061
transform 1 0 15732 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_792
timestamp 1586364061
transform 1 0 17940 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_171
timestamp 1586364061
transform 1 0 16836 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_184
timestamp 1586364061
transform 1 0 18032 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_196
timestamp 1586364061
transform 1 0 19136 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_208
timestamp 1586364061
transform 1 0 20240 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_220
timestamp 1586364061
transform 1 0 21344 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_232
timestamp 1586364061
transform 1 0 22448 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_793
timestamp 1586364061
transform 1 0 23552 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_245
timestamp 1586364061
transform 1 0 23644 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_257
timestamp 1586364061
transform 1 0 24748 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_269
timestamp 1586364061
transform 1 0 25852 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_281
timestamp 1586364061
transform 1 0 26956 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_293
timestamp 1586364061
transform 1 0 28060 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_794
timestamp 1586364061
transform 1 0 29164 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_306
timestamp 1586364061
transform 1 0 29256 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_318
timestamp 1586364061
transform 1 0 30360 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_330
timestamp 1586364061
transform 1 0 31464 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_342
timestamp 1586364061
transform 1 0 32568 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_795
timestamp 1586364061
transform 1 0 34776 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_354
timestamp 1586364061
transform 1 0 33672 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_367
timestamp 1586364061
transform 1 0 34868 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_379
timestamp 1586364061
transform 1 0 35972 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_391
timestamp 1586364061
transform 1 0 37076 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_796
timestamp 1586364061
transform 1 0 40388 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_403
timestamp 1586364061
transform 1 0 38180 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_415
timestamp 1586364061
transform 1 0 39284 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_428
timestamp 1586364061
transform 1 0 40480 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_440
timestamp 1586364061
transform 1 0 41584 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_452
timestamp 1586364061
transform 1 0 42688 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_464
timestamp 1586364061
transform 1 0 43792 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_476
timestamp 1586364061
transform 1 0 44896 0 1 44064
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_797
timestamp 1586364061
transform 1 0 46000 0 1 44064
box -38 -48 130 592
use scs8hd_decap_12  FILLER_77_489
timestamp 1586364061
transform 1 0 46092 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_77_501
timestamp 1586364061
transform 1 0 47196 0 1 44064
box -38 -48 1142 592
use scs8hd_decap_3  PHY_155
timestamp 1586364061
transform -1 0 48852 0 1 44064
box -38 -48 314 592
use scs8hd_decap_3  FILLER_77_513
timestamp 1586364061
transform 1 0 48300 0 1 44064
box -38 -48 314 592
use scs8hd_decap_3  PHY_156
timestamp 1586364061
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use scs8hd_decap_12  FILLER_78_3
timestamp 1586364061
transform 1 0 1380 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_15
timestamp 1586364061
transform 1 0 2484 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_798
timestamp 1586364061
transform 1 0 3956 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_4  FILLER_78_27
timestamp 1586364061
transform 1 0 3588 0 -1 45152
box -38 -48 406 592
use scs8hd_decap_12  FILLER_78_32
timestamp 1586364061
transform 1 0 4048 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_44
timestamp 1586364061
transform 1 0 5152 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_56
timestamp 1586364061
transform 1 0 6256 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_68
timestamp 1586364061
transform 1 0 7360 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_80
timestamp 1586364061
transform 1 0 8464 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_799
timestamp 1586364061
transform 1 0 9568 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_93
timestamp 1586364061
transform 1 0 9660 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_105
timestamp 1586364061
transform 1 0 10764 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_117
timestamp 1586364061
transform 1 0 11868 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_129
timestamp 1586364061
transform 1 0 12972 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_800
timestamp 1586364061
transform 1 0 15180 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_141
timestamp 1586364061
transform 1 0 14076 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_154
timestamp 1586364061
transform 1 0 15272 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_166
timestamp 1586364061
transform 1 0 16376 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_178
timestamp 1586364061
transform 1 0 17480 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_801
timestamp 1586364061
transform 1 0 20792 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_190
timestamp 1586364061
transform 1 0 18584 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_202
timestamp 1586364061
transform 1 0 19688 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_215
timestamp 1586364061
transform 1 0 20884 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_227
timestamp 1586364061
transform 1 0 21988 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_239
timestamp 1586364061
transform 1 0 23092 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_251
timestamp 1586364061
transform 1 0 24196 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_263
timestamp 1586364061
transform 1 0 25300 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_802
timestamp 1586364061
transform 1 0 26404 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_276
timestamp 1586364061
transform 1 0 26496 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_288
timestamp 1586364061
transform 1 0 27600 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_300
timestamp 1586364061
transform 1 0 28704 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_312
timestamp 1586364061
transform 1 0 29808 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_803
timestamp 1586364061
transform 1 0 32016 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_324
timestamp 1586364061
transform 1 0 30912 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_337
timestamp 1586364061
transform 1 0 32108 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_349
timestamp 1586364061
transform 1 0 33212 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_361
timestamp 1586364061
transform 1 0 34316 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_373
timestamp 1586364061
transform 1 0 35420 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_804
timestamp 1586364061
transform 1 0 37628 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_385
timestamp 1586364061
transform 1 0 36524 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_398
timestamp 1586364061
transform 1 0 37720 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_410
timestamp 1586364061
transform 1 0 38824 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_422
timestamp 1586364061
transform 1 0 39928 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_434
timestamp 1586364061
transform 1 0 41032 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_446
timestamp 1586364061
transform 1 0 42136 0 -1 45152
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_805
timestamp 1586364061
transform 1 0 43240 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_78_459
timestamp 1586364061
transform 1 0 43332 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_471
timestamp 1586364061
transform 1 0 44436 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_483
timestamp 1586364061
transform 1 0 45540 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_78_495
timestamp 1586364061
transform 1 0 46644 0 -1 45152
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_78_507
timestamp 1586364061
transform 1 0 47748 0 -1 45152
box -38 -48 774 592
use scs8hd_decap_3  PHY_157
timestamp 1586364061
transform -1 0 48852 0 -1 45152
box -38 -48 314 592
use scs8hd_fill_1  FILLER_78_515
timestamp 1586364061
transform 1 0 48484 0 -1 45152
box -38 -48 130 592
use scs8hd_decap_3  PHY_158
timestamp 1586364061
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use scs8hd_decap_3  PHY_160
timestamp 1586364061
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use scs8hd_decap_12  FILLER_79_3
timestamp 1586364061
transform 1 0 1380 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_15
timestamp 1586364061
transform 1 0 2484 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_3
timestamp 1586364061
transform 1 0 1380 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_15
timestamp 1586364061
transform 1 0 2484 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_814
timestamp 1586364061
transform 1 0 3956 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_27
timestamp 1586364061
transform 1 0 3588 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_39
timestamp 1586364061
transform 1 0 4692 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_79_51
timestamp 1586364061
transform 1 0 5796 0 1 45152
box -38 -48 774 592
use scs8hd_decap_4  FILLER_80_27
timestamp 1586364061
transform 1 0 3588 0 -1 46240
box -38 -48 406 592
use scs8hd_decap_12  FILLER_80_32
timestamp 1586364061
transform 1 0 4048 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_44
timestamp 1586364061
transform 1 0 5152 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_806
timestamp 1586364061
transform 1 0 6716 0 1 45152
box -38 -48 130 592
use scs8hd_fill_2  FILLER_79_59
timestamp 1586364061
transform 1 0 6532 0 1 45152
box -38 -48 222 592
use scs8hd_decap_12  FILLER_79_62
timestamp 1586364061
transform 1 0 6808 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_74
timestamp 1586364061
transform 1 0 7912 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_56
timestamp 1586364061
transform 1 0 6256 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_68
timestamp 1586364061
transform 1 0 7360 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_80
timestamp 1586364061
transform 1 0 8464 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_815
timestamp 1586364061
transform 1 0 9568 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_86
timestamp 1586364061
transform 1 0 9016 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_98
timestamp 1586364061
transform 1 0 10120 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_93
timestamp 1586364061
transform 1 0 9660 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_105
timestamp 1586364061
transform 1 0 10764 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_807
timestamp 1586364061
transform 1 0 12328 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_110
timestamp 1586364061
transform 1 0 11224 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_123
timestamp 1586364061
transform 1 0 12420 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_117
timestamp 1586364061
transform 1 0 11868 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_129
timestamp 1586364061
transform 1 0 12972 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_816
timestamp 1586364061
transform 1 0 15180 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_135
timestamp 1586364061
transform 1 0 13524 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_147
timestamp 1586364061
transform 1 0 14628 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_159
timestamp 1586364061
transform 1 0 15732 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_141
timestamp 1586364061
transform 1 0 14076 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_154
timestamp 1586364061
transform 1 0 15272 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_808
timestamp 1586364061
transform 1 0 17940 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_171
timestamp 1586364061
transform 1 0 16836 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_184
timestamp 1586364061
transform 1 0 18032 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_166
timestamp 1586364061
transform 1 0 16376 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_178
timestamp 1586364061
transform 1 0 17480 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_817
timestamp 1586364061
transform 1 0 20792 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_196
timestamp 1586364061
transform 1 0 19136 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_208
timestamp 1586364061
transform 1 0 20240 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_190
timestamp 1586364061
transform 1 0 18584 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_202
timestamp 1586364061
transform 1 0 19688 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_220
timestamp 1586364061
transform 1 0 21344 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_232
timestamp 1586364061
transform 1 0 22448 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_215
timestamp 1586364061
transform 1 0 20884 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_227
timestamp 1586364061
transform 1 0 21988 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_239
timestamp 1586364061
transform 1 0 23092 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_809
timestamp 1586364061
transform 1 0 23552 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_245
timestamp 1586364061
transform 1 0 23644 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_257
timestamp 1586364061
transform 1 0 24748 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_251
timestamp 1586364061
transform 1 0 24196 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_263
timestamp 1586364061
transform 1 0 25300 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_818
timestamp 1586364061
transform 1 0 26404 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_269
timestamp 1586364061
transform 1 0 25852 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_281
timestamp 1586364061
transform 1 0 26956 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_293
timestamp 1586364061
transform 1 0 28060 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_276
timestamp 1586364061
transform 1 0 26496 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_288
timestamp 1586364061
transform 1 0 27600 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_810
timestamp 1586364061
transform 1 0 29164 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_306
timestamp 1586364061
transform 1 0 29256 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_318
timestamp 1586364061
transform 1 0 30360 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_300
timestamp 1586364061
transform 1 0 28704 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_312
timestamp 1586364061
transform 1 0 29808 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_819
timestamp 1586364061
transform 1 0 32016 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_330
timestamp 1586364061
transform 1 0 31464 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_342
timestamp 1586364061
transform 1 0 32568 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_324
timestamp 1586364061
transform 1 0 30912 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_337
timestamp 1586364061
transform 1 0 32108 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_811
timestamp 1586364061
transform 1 0 34776 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_354
timestamp 1586364061
transform 1 0 33672 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_367
timestamp 1586364061
transform 1 0 34868 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_349
timestamp 1586364061
transform 1 0 33212 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_361
timestamp 1586364061
transform 1 0 34316 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_373
timestamp 1586364061
transform 1 0 35420 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_820
timestamp 1586364061
transform 1 0 37628 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_379
timestamp 1586364061
transform 1 0 35972 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_391
timestamp 1586364061
transform 1 0 37076 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_385
timestamp 1586364061
transform 1 0 36524 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_398
timestamp 1586364061
transform 1 0 37720 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_812
timestamp 1586364061
transform 1 0 40388 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_403
timestamp 1586364061
transform 1 0 38180 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_415
timestamp 1586364061
transform 1 0 39284 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_428
timestamp 1586364061
transform 1 0 40480 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_410
timestamp 1586364061
transform 1 0 38824 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_422
timestamp 1586364061
transform 1 0 39928 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_440
timestamp 1586364061
transform 1 0 41584 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_452
timestamp 1586364061
transform 1 0 42688 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_434
timestamp 1586364061
transform 1 0 41032 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_446
timestamp 1586364061
transform 1 0 42136 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_821
timestamp 1586364061
transform 1 0 43240 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_464
timestamp 1586364061
transform 1 0 43792 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_476
timestamp 1586364061
transform 1 0 44896 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_459
timestamp 1586364061
transform 1 0 43332 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_471
timestamp 1586364061
transform 1 0 44436 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_483
timestamp 1586364061
transform 1 0 45540 0 -1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_813
timestamp 1586364061
transform 1 0 46000 0 1 45152
box -38 -48 130 592
use scs8hd_decap_12  FILLER_79_489
timestamp 1586364061
transform 1 0 46092 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_79_501
timestamp 1586364061
transform 1 0 47196 0 1 45152
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_80_495
timestamp 1586364061
transform 1 0 46644 0 -1 46240
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_80_507
timestamp 1586364061
transform 1 0 47748 0 -1 46240
box -38 -48 774 592
use scs8hd_decap_3  PHY_159
timestamp 1586364061
transform -1 0 48852 0 1 45152
box -38 -48 314 592
use scs8hd_decap_3  PHY_161
timestamp 1586364061
transform -1 0 48852 0 -1 46240
box -38 -48 314 592
use scs8hd_decap_3  FILLER_79_513
timestamp 1586364061
transform 1 0 48300 0 1 45152
box -38 -48 314 592
use scs8hd_fill_1  FILLER_80_515
timestamp 1586364061
transform 1 0 48484 0 -1 46240
box -38 -48 130 592
use scs8hd_decap_3  PHY_162
timestamp 1586364061
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use scs8hd_decap_12  FILLER_81_3
timestamp 1586364061
transform 1 0 1380 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_15
timestamp 1586364061
transform 1 0 2484 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_27
timestamp 1586364061
transform 1 0 3588 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_39
timestamp 1586364061
transform 1 0 4692 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_81_51
timestamp 1586364061
transform 1 0 5796 0 1 46240
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_822
timestamp 1586364061
transform 1 0 6716 0 1 46240
box -38 -48 130 592
use scs8hd_fill_2  FILLER_81_59
timestamp 1586364061
transform 1 0 6532 0 1 46240
box -38 -48 222 592
use scs8hd_decap_12  FILLER_81_62
timestamp 1586364061
transform 1 0 6808 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_74
timestamp 1586364061
transform 1 0 7912 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_86
timestamp 1586364061
transform 1 0 9016 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_98
timestamp 1586364061
transform 1 0 10120 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_823
timestamp 1586364061
transform 1 0 12328 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_110
timestamp 1586364061
transform 1 0 11224 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_123
timestamp 1586364061
transform 1 0 12420 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_135
timestamp 1586364061
transform 1 0 13524 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_147
timestamp 1586364061
transform 1 0 14628 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_159
timestamp 1586364061
transform 1 0 15732 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_824
timestamp 1586364061
transform 1 0 17940 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_171
timestamp 1586364061
transform 1 0 16836 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_184
timestamp 1586364061
transform 1 0 18032 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_196
timestamp 1586364061
transform 1 0 19136 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_208
timestamp 1586364061
transform 1 0 20240 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_220
timestamp 1586364061
transform 1 0 21344 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_232
timestamp 1586364061
transform 1 0 22448 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_825
timestamp 1586364061
transform 1 0 23552 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_245
timestamp 1586364061
transform 1 0 23644 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_257
timestamp 1586364061
transform 1 0 24748 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_269
timestamp 1586364061
transform 1 0 25852 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_281
timestamp 1586364061
transform 1 0 26956 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_293
timestamp 1586364061
transform 1 0 28060 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_826
timestamp 1586364061
transform 1 0 29164 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_306
timestamp 1586364061
transform 1 0 29256 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_318
timestamp 1586364061
transform 1 0 30360 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_330
timestamp 1586364061
transform 1 0 31464 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_342
timestamp 1586364061
transform 1 0 32568 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_827
timestamp 1586364061
transform 1 0 34776 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_354
timestamp 1586364061
transform 1 0 33672 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_367
timestamp 1586364061
transform 1 0 34868 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_379
timestamp 1586364061
transform 1 0 35972 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_391
timestamp 1586364061
transform 1 0 37076 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_828
timestamp 1586364061
transform 1 0 40388 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_403
timestamp 1586364061
transform 1 0 38180 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_415
timestamp 1586364061
transform 1 0 39284 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_428
timestamp 1586364061
transform 1 0 40480 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_440
timestamp 1586364061
transform 1 0 41584 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_452
timestamp 1586364061
transform 1 0 42688 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_464
timestamp 1586364061
transform 1 0 43792 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_476
timestamp 1586364061
transform 1 0 44896 0 1 46240
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_829
timestamp 1586364061
transform 1 0 46000 0 1 46240
box -38 -48 130 592
use scs8hd_decap_12  FILLER_81_489
timestamp 1586364061
transform 1 0 46092 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_81_501
timestamp 1586364061
transform 1 0 47196 0 1 46240
box -38 -48 1142 592
use scs8hd_decap_3  PHY_163
timestamp 1586364061
transform -1 0 48852 0 1 46240
box -38 -48 314 592
use scs8hd_decap_3  FILLER_81_513
timestamp 1586364061
transform 1 0 48300 0 1 46240
box -38 -48 314 592
use scs8hd_decap_3  PHY_164
timestamp 1586364061
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use scs8hd_decap_12  FILLER_82_3
timestamp 1586364061
transform 1 0 1380 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_15
timestamp 1586364061
transform 1 0 2484 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_830
timestamp 1586364061
transform 1 0 3956 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_4  FILLER_82_27
timestamp 1586364061
transform 1 0 3588 0 -1 47328
box -38 -48 406 592
use scs8hd_decap_12  FILLER_82_32
timestamp 1586364061
transform 1 0 4048 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_44
timestamp 1586364061
transform 1 0 5152 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_831
timestamp 1586364061
transform 1 0 6808 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_56
timestamp 1586364061
transform 1 0 6256 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_63
timestamp 1586364061
transform 1 0 6900 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_75
timestamp 1586364061
transform 1 0 8004 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_832
timestamp 1586364061
transform 1 0 9660 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_87
timestamp 1586364061
transform 1 0 9108 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_94
timestamp 1586364061
transform 1 0 9752 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_106
timestamp 1586364061
transform 1 0 10856 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_833
timestamp 1586364061
transform 1 0 12512 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_118
timestamp 1586364061
transform 1 0 11960 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_125
timestamp 1586364061
transform 1 0 12604 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_834
timestamp 1586364061
transform 1 0 15364 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_137
timestamp 1586364061
transform 1 0 13708 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_149
timestamp 1586364061
transform 1 0 14812 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_156
timestamp 1586364061
transform 1 0 15456 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_835
timestamp 1586364061
transform 1 0 18216 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_168
timestamp 1586364061
transform 1 0 16560 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_180
timestamp 1586364061
transform 1 0 17664 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_187
timestamp 1586364061
transform 1 0 18308 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_199
timestamp 1586364061
transform 1 0 19412 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_211
timestamp 1586364061
transform 1 0 20516 0 -1 47328
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_836
timestamp 1586364061
transform 1 0 21068 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_218
timestamp 1586364061
transform 1 0 21160 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_230
timestamp 1586364061
transform 1 0 22264 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_837
timestamp 1586364061
transform 1 0 23920 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_242
timestamp 1586364061
transform 1 0 23368 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_249
timestamp 1586364061
transform 1 0 24012 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_261
timestamp 1586364061
transform 1 0 25116 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_838
timestamp 1586364061
transform 1 0 26772 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_273
timestamp 1586364061
transform 1 0 26220 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_280
timestamp 1586364061
transform 1 0 26864 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_292
timestamp 1586364061
transform 1 0 27968 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_839
timestamp 1586364061
transform 1 0 29624 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_304
timestamp 1586364061
transform 1 0 29072 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_311
timestamp 1586364061
transform 1 0 29716 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_840
timestamp 1586364061
transform 1 0 32476 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_323
timestamp 1586364061
transform 1 0 30820 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_335
timestamp 1586364061
transform 1 0 31924 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_342
timestamp 1586364061
transform 1 0 32568 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_841
timestamp 1586364061
transform 1 0 35328 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_354
timestamp 1586364061
transform 1 0 33672 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_366
timestamp 1586364061
transform 1 0 34776 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_373
timestamp 1586364061
transform 1 0 35420 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_385
timestamp 1586364061
transform 1 0 36524 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_397
timestamp 1586364061
transform 1 0 37628 0 -1 47328
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_842
timestamp 1586364061
transform 1 0 38180 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_404
timestamp 1586364061
transform 1 0 38272 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_416
timestamp 1586364061
transform 1 0 39376 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_428
timestamp 1586364061
transform 1 0 40480 0 -1 47328
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_843
timestamp 1586364061
transform 1 0 41032 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_12  FILLER_82_435
timestamp 1586364061
transform 1 0 41124 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_447
timestamp 1586364061
transform 1 0 42228 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_844
timestamp 1586364061
transform 1 0 43884 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_459
timestamp 1586364061
transform 1 0 43332 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_466
timestamp 1586364061
transform 1 0 43976 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_82_478
timestamp 1586364061
transform 1 0 45080 0 -1 47328
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_845
timestamp 1586364061
transform 1 0 46736 0 -1 47328
box -38 -48 130 592
use scs8hd_decap_6  FILLER_82_490
timestamp 1586364061
transform 1 0 46184 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_12  FILLER_82_497
timestamp 1586364061
transform 1 0 46828 0 -1 47328
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_82_509
timestamp 1586364061
transform 1 0 47932 0 -1 47328
box -38 -48 590 592
use scs8hd_decap_3  PHY_165
timestamp 1586364061
transform -1 0 48852 0 -1 47328
box -38 -48 314 592
use scs8hd_fill_1  FILLER_82_515
timestamp 1586364061
transform 1 0 48484 0 -1 47328
box -38 -48 130 592
<< labels >>
rlabel metal2 s 12438 0 12494 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 16026 0 16082 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 19522 0 19578 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 23110 0 23166 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 26698 0 26754 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 2778 49520 2834 50000 6 address[5]
port 5 nsew default input
rlabel metal2 s 8298 49520 8354 50000 6 address[6]
port 6 nsew default input
rlabel metal3 s 0 8304 480 8424 6 address[7]
port 7 nsew default input
rlabel metal2 s 13818 49520 13874 50000 6 address[8]
port 8 nsew default input
rlabel metal2 s 19430 49520 19486 50000 6 address[9]
port 9 nsew default input
rlabel metal3 s 49520 31288 50000 31408 6 bottom_width_0_height_0__pin_10_
port 10 nsew default tristate
rlabel metal2 s 37370 0 37426 480 6 bottom_width_0_height_0__pin_14_
port 11 nsew default input
rlabel metal2 s 30286 0 30342 480 6 bottom_width_0_height_0__pin_2_
port 12 nsew default input
rlabel metal2 s 33874 0 33930 480 6 bottom_width_0_height_0__pin_6_
port 13 nsew default input
rlabel metal2 s 8850 0 8906 480 6 clk
port 14 nsew default input
rlabel metal3 s 49520 18776 50000 18896 6 data_in
port 15 nsew default input
rlabel metal3 s 49520 6264 50000 6384 6 enable
port 16 nsew default input
rlabel metal3 s 49520 43800 50000 43920 6 left_width_0_height_0__pin_11_
port 17 nsew default tristate
rlabel metal2 s 24950 49520 25006 50000 6 left_width_0_height_0__pin_3_
port 18 nsew default input
rlabel metal2 s 30470 49520 30526 50000 6 left_width_0_height_0__pin_7_
port 19 nsew default input
rlabel metal2 s 5262 0 5318 480 6 reset
port 20 nsew default input
rlabel metal3 s 0 24896 480 25016 6 right_width_0_height_0__pin_13_
port 21 nsew default tristate
rlabel metal2 s 40958 0 41014 480 6 right_width_0_height_0__pin_1_
port 22 nsew default input
rlabel metal2 s 36082 49520 36138 50000 6 right_width_0_height_0__pin_5_
port 23 nsew default input
rlabel metal2 s 41602 49520 41658 50000 6 right_width_0_height_0__pin_9_
port 24 nsew default input
rlabel metal2 s 1766 0 1822 480 6 set
port 25 nsew default input
rlabel metal2 s 44546 0 44602 480 6 top_width_0_height_0__pin_0_
port 26 nsew default input
rlabel metal2 s 48134 0 48190 480 6 top_width_0_height_0__pin_12_
port 27 nsew default tristate
rlabel metal2 s 47122 49520 47178 50000 6 top_width_0_height_0__pin_4_
port 28 nsew default input
rlabel metal3 s 0 41624 480 41744 6 top_width_0_height_0__pin_8_
port 29 nsew default input
rlabel metal4 s 4208 2128 4528 47376 6 vpwr
port 30 nsew default input
rlabel metal4 s 19568 2128 19888 47376 6 vgnd
port 31 nsew default input
<< end >>
