magic
tech EFS8A
magscale 1 2
timestamp 1604427683
<< viali >>
rect 15201 18921 15235 18955
rect 15130 18785 15164 18819
rect 13407 18377 13441 18411
rect 13867 18377 13901 18411
rect 15155 18377 15189 18411
rect 13223 18173 13257 18207
rect 22883 10965 22917 10999
rect 24263 10761 24297 10795
rect 10187 10693 10221 10727
rect 10003 10557 10037 10591
rect 22883 10557 22917 10591
rect 23150 10557 23184 10591
rect 10555 10421 10589 10455
rect 22975 10217 23009 10251
rect 20491 2601 20525 2635
rect 22055 2601 22089 2635
rect 20307 2465 20341 2499
rect 20951 2465 20985 2499
rect 21411 2465 21445 2499
rect 21595 2329 21629 2363
<< metal1 >>
rect 23788 21904 23794 21956
rect 23846 21944 23852 21956
rect 25076 21944 25082 21956
rect 23846 21916 25082 21944
rect 23846 21904 23852 21916
rect 25076 21904 25082 21916
rect 25134 21904 25140 21956
rect 38 21786 27822 21808
rect 38 21734 4916 21786
rect 4968 21734 4980 21786
rect 5032 21734 5044 21786
rect 5096 21734 5108 21786
rect 5160 21734 14916 21786
rect 14968 21734 14980 21786
rect 15032 21734 15044 21786
rect 15096 21734 15108 21786
rect 15160 21734 24916 21786
rect 24968 21734 24980 21786
rect 25032 21734 25044 21786
rect 25096 21734 25108 21786
rect 25160 21734 27822 21786
rect 38 21712 27822 21734
rect 38 21242 27822 21264
rect 38 21190 9916 21242
rect 9968 21190 9980 21242
rect 10032 21190 10044 21242
rect 10096 21190 10108 21242
rect 10160 21190 19916 21242
rect 19968 21190 19980 21242
rect 20032 21190 20044 21242
rect 20096 21190 20108 21242
rect 20160 21190 27822 21242
rect 38 21168 27822 21190
rect 38 20698 27822 20720
rect 38 20646 4916 20698
rect 4968 20646 4980 20698
rect 5032 20646 5044 20698
rect 5096 20646 5108 20698
rect 5160 20646 14916 20698
rect 14968 20646 14980 20698
rect 15032 20646 15044 20698
rect 15096 20646 15108 20698
rect 15160 20646 24916 20698
rect 24968 20646 24980 20698
rect 25032 20646 25044 20698
rect 25096 20646 25108 20698
rect 25160 20646 27822 20698
rect 38 20624 27822 20646
rect 38 20154 27822 20176
rect 38 20102 9916 20154
rect 9968 20102 9980 20154
rect 10032 20102 10044 20154
rect 10096 20102 10108 20154
rect 10160 20102 19916 20154
rect 19968 20102 19980 20154
rect 20032 20102 20044 20154
rect 20096 20102 20108 20154
rect 20160 20102 27822 20154
rect 38 20080 27822 20102
rect 38 19610 27822 19632
rect 38 19558 4916 19610
rect 4968 19558 4980 19610
rect 5032 19558 5044 19610
rect 5096 19558 5108 19610
rect 5160 19558 14916 19610
rect 14968 19558 14980 19610
rect 15032 19558 15044 19610
rect 15096 19558 15108 19610
rect 15160 19558 24916 19610
rect 24968 19558 24980 19610
rect 25032 19558 25044 19610
rect 25096 19558 25108 19610
rect 25160 19558 27822 19610
rect 38 19536 27822 19558
rect 38 19066 27822 19088
rect 38 19014 9916 19066
rect 9968 19014 9980 19066
rect 10032 19014 10044 19066
rect 10096 19014 10108 19066
rect 10160 19014 19916 19066
rect 19968 19014 19980 19066
rect 20032 19014 20044 19066
rect 20096 19014 20108 19066
rect 20160 19014 27822 19066
rect 38 18992 27822 19014
rect 15189 18955 15247 18961
rect 15189 18921 15201 18955
rect 15235 18952 15247 18955
rect 15324 18952 15330 18964
rect 15235 18924 15330 18952
rect 15235 18921 15247 18924
rect 15189 18915 15247 18921
rect 15324 18912 15330 18924
rect 15382 18912 15388 18964
rect 15140 18825 15146 18828
rect 15118 18819 15146 18825
rect 15118 18785 15130 18819
rect 15118 18779 15146 18785
rect 15140 18776 15146 18779
rect 15198 18776 15204 18828
rect 38 18522 27822 18544
rect 38 18470 4916 18522
rect 4968 18470 4980 18522
rect 5032 18470 5044 18522
rect 5096 18470 5108 18522
rect 5160 18470 14916 18522
rect 14968 18470 14980 18522
rect 15032 18470 15044 18522
rect 15096 18470 15108 18522
rect 15160 18470 24916 18522
rect 24968 18470 24980 18522
rect 25032 18470 25044 18522
rect 25096 18470 25108 18522
rect 25160 18470 27822 18522
rect 38 18448 27822 18470
rect 13392 18408 13398 18420
rect 13353 18380 13398 18408
rect 13392 18368 13398 18380
rect 13450 18368 13456 18420
rect 13855 18411 13913 18417
rect 13855 18377 13867 18411
rect 13901 18408 13913 18411
rect 15143 18411 15201 18417
rect 15143 18408 15155 18411
rect 13901 18380 15155 18408
rect 13901 18377 13913 18380
rect 13855 18371 13913 18377
rect 15143 18377 15155 18380
rect 15189 18408 15201 18411
rect 15232 18408 15238 18420
rect 15189 18380 15238 18408
rect 15189 18377 15201 18380
rect 15143 18371 15201 18377
rect 13211 18207 13269 18213
rect 13211 18173 13223 18207
rect 13257 18204 13269 18207
rect 13870 18204 13898 18371
rect 15232 18368 15238 18380
rect 15290 18368 15296 18420
rect 13257 18176 13898 18204
rect 13257 18173 13269 18176
rect 13211 18167 13269 18173
rect 38 17978 27822 18000
rect 38 17926 9916 17978
rect 9968 17926 9980 17978
rect 10032 17926 10044 17978
rect 10096 17926 10108 17978
rect 10160 17926 19916 17978
rect 19968 17926 19980 17978
rect 20032 17926 20044 17978
rect 20096 17926 20108 17978
rect 20160 17926 27822 17978
rect 38 17904 27822 17926
rect 38 17434 27822 17456
rect 38 17382 4916 17434
rect 4968 17382 4980 17434
rect 5032 17382 5044 17434
rect 5096 17382 5108 17434
rect 5160 17382 14916 17434
rect 14968 17382 14980 17434
rect 15032 17382 15044 17434
rect 15096 17382 15108 17434
rect 15160 17382 24916 17434
rect 24968 17382 24980 17434
rect 25032 17382 25044 17434
rect 25096 17382 25108 17434
rect 25160 17382 27822 17434
rect 38 17360 27822 17382
rect 38 16890 27822 16912
rect 38 16838 9916 16890
rect 9968 16838 9980 16890
rect 10032 16838 10044 16890
rect 10096 16838 10108 16890
rect 10160 16838 19916 16890
rect 19968 16838 19980 16890
rect 20032 16838 20044 16890
rect 20096 16838 20108 16890
rect 20160 16838 27822 16890
rect 38 16816 27822 16838
rect 38 16346 27822 16368
rect 38 16294 4916 16346
rect 4968 16294 4980 16346
rect 5032 16294 5044 16346
rect 5096 16294 5108 16346
rect 5160 16294 14916 16346
rect 14968 16294 14980 16346
rect 15032 16294 15044 16346
rect 15096 16294 15108 16346
rect 15160 16294 24916 16346
rect 24968 16294 24980 16346
rect 25032 16294 25044 16346
rect 25096 16294 25108 16346
rect 25160 16294 27822 16346
rect 38 16272 27822 16294
rect 38 15802 27822 15824
rect 38 15750 9916 15802
rect 9968 15750 9980 15802
rect 10032 15750 10044 15802
rect 10096 15750 10108 15802
rect 10160 15750 19916 15802
rect 19968 15750 19980 15802
rect 20032 15750 20044 15802
rect 20096 15750 20108 15802
rect 20160 15750 27822 15802
rect 38 15728 27822 15750
rect 38 15258 27822 15280
rect 38 15206 4916 15258
rect 4968 15206 4980 15258
rect 5032 15206 5044 15258
rect 5096 15206 5108 15258
rect 5160 15206 14916 15258
rect 14968 15206 14980 15258
rect 15032 15206 15044 15258
rect 15096 15206 15108 15258
rect 15160 15206 24916 15258
rect 24968 15206 24980 15258
rect 25032 15206 25044 15258
rect 25096 15206 25108 15258
rect 25160 15206 27822 15258
rect 38 15184 27822 15206
rect 38 14714 27822 14736
rect 38 14662 9916 14714
rect 9968 14662 9980 14714
rect 10032 14662 10044 14714
rect 10096 14662 10108 14714
rect 10160 14662 19916 14714
rect 19968 14662 19980 14714
rect 20032 14662 20044 14714
rect 20096 14662 20108 14714
rect 20160 14662 27822 14714
rect 38 14640 27822 14662
rect 38 14170 27822 14192
rect 38 14118 4916 14170
rect 4968 14118 4980 14170
rect 5032 14118 5044 14170
rect 5096 14118 5108 14170
rect 5160 14118 14916 14170
rect 14968 14118 14980 14170
rect 15032 14118 15044 14170
rect 15096 14118 15108 14170
rect 15160 14118 24916 14170
rect 24968 14118 24980 14170
rect 25032 14118 25044 14170
rect 25096 14118 25108 14170
rect 25160 14118 27822 14170
rect 38 14096 27822 14118
rect 38 13626 27822 13648
rect 38 13574 9916 13626
rect 9968 13574 9980 13626
rect 10032 13574 10044 13626
rect 10096 13574 10108 13626
rect 10160 13574 19916 13626
rect 19968 13574 19980 13626
rect 20032 13574 20044 13626
rect 20096 13574 20108 13626
rect 20160 13574 27822 13626
rect 38 13552 27822 13574
rect 38 13082 27822 13104
rect 38 13030 4916 13082
rect 4968 13030 4980 13082
rect 5032 13030 5044 13082
rect 5096 13030 5108 13082
rect 5160 13030 14916 13082
rect 14968 13030 14980 13082
rect 15032 13030 15044 13082
rect 15096 13030 15108 13082
rect 15160 13030 24916 13082
rect 24968 13030 24980 13082
rect 25032 13030 25044 13082
rect 25096 13030 25108 13082
rect 25160 13030 27822 13082
rect 38 13008 27822 13030
rect 38 12538 27822 12560
rect 38 12486 9916 12538
rect 9968 12486 9980 12538
rect 10032 12486 10044 12538
rect 10096 12486 10108 12538
rect 10160 12486 19916 12538
rect 19968 12486 19980 12538
rect 20032 12486 20044 12538
rect 20096 12486 20108 12538
rect 20160 12486 27822 12538
rect 38 12464 27822 12486
rect 38 11994 27822 12016
rect 38 11942 4916 11994
rect 4968 11942 4980 11994
rect 5032 11942 5044 11994
rect 5096 11942 5108 11994
rect 5160 11942 14916 11994
rect 14968 11942 14980 11994
rect 15032 11942 15044 11994
rect 15096 11942 15108 11994
rect 15160 11942 24916 11994
rect 24968 11942 24980 11994
rect 25032 11942 25044 11994
rect 25096 11942 25108 11994
rect 25160 11942 27822 11994
rect 38 11920 27822 11942
rect 38 11450 27822 11472
rect 38 11398 9916 11450
rect 9968 11398 9980 11450
rect 10032 11398 10044 11450
rect 10096 11398 10108 11450
rect 10160 11398 19916 11450
rect 19968 11398 19980 11450
rect 20032 11398 20044 11450
rect 20096 11398 20108 11450
rect 20160 11398 27822 11450
rect 38 11376 27822 11398
rect 22868 10996 22874 11008
rect 22829 10968 22874 10996
rect 22868 10956 22874 10968
rect 22926 10956 22932 11008
rect 38 10906 27822 10928
rect 38 10854 4916 10906
rect 4968 10854 4980 10906
rect 5032 10854 5044 10906
rect 5096 10854 5108 10906
rect 5160 10854 14916 10906
rect 14968 10854 14980 10906
rect 15032 10854 15044 10906
rect 15096 10854 15108 10906
rect 15160 10854 24916 10906
rect 24968 10854 24980 10906
rect 25032 10854 25044 10906
rect 25096 10854 25108 10906
rect 25160 10854 27822 10906
rect 38 10832 27822 10854
rect 24251 10795 24309 10801
rect 24251 10761 24263 10795
rect 24297 10792 24309 10795
rect 24432 10792 24438 10804
rect 24297 10764 24438 10792
rect 24297 10761 24309 10764
rect 24251 10755 24309 10761
rect 24432 10752 24438 10764
rect 24490 10752 24496 10804
rect 10172 10724 10178 10736
rect 10133 10696 10178 10724
rect 10172 10684 10178 10696
rect 10230 10684 10236 10736
rect 9991 10591 10049 10597
rect 9991 10557 10003 10591
rect 10037 10588 10049 10591
rect 22868 10588 22874 10600
rect 10037 10560 10586 10588
rect 22829 10560 22874 10588
rect 10037 10557 10049 10560
rect 9991 10551 10049 10557
rect 10558 10464 10586 10560
rect 22868 10548 22874 10560
rect 22926 10548 22932 10600
rect 22960 10548 22966 10600
rect 23018 10588 23024 10600
rect 23138 10591 23196 10597
rect 23138 10588 23150 10591
rect 23018 10560 23150 10588
rect 23018 10548 23024 10560
rect 23138 10557 23150 10560
rect 23184 10588 23196 10591
rect 23880 10588 23886 10600
rect 23184 10560 23886 10588
rect 23184 10557 23196 10560
rect 23138 10551 23196 10557
rect 23880 10548 23886 10560
rect 23938 10548 23944 10600
rect 10540 10452 10546 10464
rect 10501 10424 10546 10452
rect 10540 10412 10546 10424
rect 10598 10412 10604 10464
rect 38 10362 27822 10384
rect 38 10310 9916 10362
rect 9968 10310 9980 10362
rect 10032 10310 10044 10362
rect 10096 10310 10108 10362
rect 10160 10310 19916 10362
rect 19968 10310 19980 10362
rect 20032 10310 20044 10362
rect 20096 10310 20108 10362
rect 20160 10310 27822 10362
rect 38 10288 27822 10310
rect 22960 10248 22966 10260
rect 22921 10220 22966 10248
rect 22960 10208 22966 10220
rect 23018 10208 23024 10260
rect 38 9818 27822 9840
rect 38 9766 4916 9818
rect 4968 9766 4980 9818
rect 5032 9766 5044 9818
rect 5096 9766 5108 9818
rect 5160 9766 14916 9818
rect 14968 9766 14980 9818
rect 15032 9766 15044 9818
rect 15096 9766 15108 9818
rect 15160 9766 24916 9818
rect 24968 9766 24980 9818
rect 25032 9766 25044 9818
rect 25096 9766 25108 9818
rect 25160 9766 27822 9818
rect 38 9744 27822 9766
rect 38 9274 27822 9296
rect 38 9222 9916 9274
rect 9968 9222 9980 9274
rect 10032 9222 10044 9274
rect 10096 9222 10108 9274
rect 10160 9222 19916 9274
rect 19968 9222 19980 9274
rect 20032 9222 20044 9274
rect 20096 9222 20108 9274
rect 20160 9222 27822 9274
rect 38 9200 27822 9222
rect 38 8730 27822 8752
rect 38 8678 4916 8730
rect 4968 8678 4980 8730
rect 5032 8678 5044 8730
rect 5096 8678 5108 8730
rect 5160 8678 14916 8730
rect 14968 8678 14980 8730
rect 15032 8678 15044 8730
rect 15096 8678 15108 8730
rect 15160 8678 24916 8730
rect 24968 8678 24980 8730
rect 25032 8678 25044 8730
rect 25096 8678 25108 8730
rect 25160 8678 27822 8730
rect 38 8656 27822 8678
rect 38 8186 27822 8208
rect 38 8134 9916 8186
rect 9968 8134 9980 8186
rect 10032 8134 10044 8186
rect 10096 8134 10108 8186
rect 10160 8134 19916 8186
rect 19968 8134 19980 8186
rect 20032 8134 20044 8186
rect 20096 8134 20108 8186
rect 20160 8134 27822 8186
rect 38 8112 27822 8134
rect 38 7642 27822 7664
rect 38 7590 4916 7642
rect 4968 7590 4980 7642
rect 5032 7590 5044 7642
rect 5096 7590 5108 7642
rect 5160 7590 14916 7642
rect 14968 7590 14980 7642
rect 15032 7590 15044 7642
rect 15096 7590 15108 7642
rect 15160 7590 24916 7642
rect 24968 7590 24980 7642
rect 25032 7590 25044 7642
rect 25096 7590 25108 7642
rect 25160 7590 27822 7642
rect 38 7568 27822 7590
rect 38 7098 27822 7120
rect 38 7046 9916 7098
rect 9968 7046 9980 7098
rect 10032 7046 10044 7098
rect 10096 7046 10108 7098
rect 10160 7046 19916 7098
rect 19968 7046 19980 7098
rect 20032 7046 20044 7098
rect 20096 7046 20108 7098
rect 20160 7046 27822 7098
rect 38 7024 27822 7046
rect 38 6554 27822 6576
rect 38 6502 4916 6554
rect 4968 6502 4980 6554
rect 5032 6502 5044 6554
rect 5096 6502 5108 6554
rect 5160 6502 14916 6554
rect 14968 6502 14980 6554
rect 15032 6502 15044 6554
rect 15096 6502 15108 6554
rect 15160 6502 24916 6554
rect 24968 6502 24980 6554
rect 25032 6502 25044 6554
rect 25096 6502 25108 6554
rect 25160 6502 27822 6554
rect 38 6480 27822 6502
rect 38 6010 27822 6032
rect 38 5958 9916 6010
rect 9968 5958 9980 6010
rect 10032 5958 10044 6010
rect 10096 5958 10108 6010
rect 10160 5958 19916 6010
rect 19968 5958 19980 6010
rect 20032 5958 20044 6010
rect 20096 5958 20108 6010
rect 20160 5958 27822 6010
rect 38 5936 27822 5958
rect 38 5466 27822 5488
rect 38 5414 4916 5466
rect 4968 5414 4980 5466
rect 5032 5414 5044 5466
rect 5096 5414 5108 5466
rect 5160 5414 14916 5466
rect 14968 5414 14980 5466
rect 15032 5414 15044 5466
rect 15096 5414 15108 5466
rect 15160 5414 24916 5466
rect 24968 5414 24980 5466
rect 25032 5414 25044 5466
rect 25096 5414 25108 5466
rect 25160 5414 27822 5466
rect 38 5392 27822 5414
rect 38 4922 27822 4944
rect 38 4870 9916 4922
rect 9968 4870 9980 4922
rect 10032 4870 10044 4922
rect 10096 4870 10108 4922
rect 10160 4870 19916 4922
rect 19968 4870 19980 4922
rect 20032 4870 20044 4922
rect 20096 4870 20108 4922
rect 20160 4870 27822 4922
rect 38 4848 27822 4870
rect 38 4378 27822 4400
rect 38 4326 4916 4378
rect 4968 4326 4980 4378
rect 5032 4326 5044 4378
rect 5096 4326 5108 4378
rect 5160 4326 14916 4378
rect 14968 4326 14980 4378
rect 15032 4326 15044 4378
rect 15096 4326 15108 4378
rect 15160 4326 24916 4378
rect 24968 4326 24980 4378
rect 25032 4326 25044 4378
rect 25096 4326 25108 4378
rect 25160 4326 27822 4378
rect 38 4304 27822 4326
rect 38 3834 27822 3856
rect 38 3782 9916 3834
rect 9968 3782 9980 3834
rect 10032 3782 10044 3834
rect 10096 3782 10108 3834
rect 10160 3782 19916 3834
rect 19968 3782 19980 3834
rect 20032 3782 20044 3834
rect 20096 3782 20108 3834
rect 20160 3782 27822 3834
rect 38 3760 27822 3782
rect 38 3290 27822 3312
rect 38 3238 4916 3290
rect 4968 3238 4980 3290
rect 5032 3238 5044 3290
rect 5096 3238 5108 3290
rect 5160 3238 14916 3290
rect 14968 3238 14980 3290
rect 15032 3238 15044 3290
rect 15096 3238 15108 3290
rect 15160 3238 24916 3290
rect 24968 3238 24980 3290
rect 25032 3238 25044 3290
rect 25096 3238 25108 3290
rect 25160 3238 27822 3290
rect 38 3216 27822 3238
rect 38 2746 27822 2768
rect 38 2694 9916 2746
rect 9968 2694 9980 2746
rect 10032 2694 10044 2746
rect 10096 2694 10108 2746
rect 10160 2694 19916 2746
rect 19968 2694 19980 2746
rect 20032 2694 20044 2746
rect 20096 2694 20108 2746
rect 20160 2694 27822 2746
rect 38 2672 27822 2694
rect 20476 2632 20482 2644
rect 20437 2604 20482 2632
rect 20476 2592 20482 2604
rect 20534 2592 20540 2644
rect 22040 2632 22046 2644
rect 22001 2604 22046 2632
rect 22040 2592 22046 2604
rect 22098 2592 22104 2644
rect 20295 2499 20353 2505
rect 20295 2465 20307 2499
rect 20341 2496 20353 2499
rect 20939 2499 20997 2505
rect 20939 2496 20951 2499
rect 20341 2468 20951 2496
rect 20341 2465 20353 2468
rect 20295 2459 20353 2465
rect 20939 2465 20951 2468
rect 20985 2496 20997 2499
rect 21399 2499 21457 2505
rect 21399 2496 21411 2499
rect 20985 2468 21411 2496
rect 20985 2465 20997 2468
rect 20939 2459 20997 2465
rect 21399 2465 21411 2468
rect 21445 2496 21457 2499
rect 22058 2496 22086 2592
rect 21445 2468 22086 2496
rect 21445 2465 21457 2468
rect 21399 2459 21457 2465
rect 21583 2363 21641 2369
rect 21583 2329 21595 2363
rect 21629 2360 21641 2363
rect 23880 2360 23886 2372
rect 21629 2332 23886 2360
rect 21629 2329 21641 2332
rect 21583 2323 21641 2329
rect 23880 2320 23886 2332
rect 23938 2320 23944 2372
rect 38 2202 27822 2224
rect 38 2150 4916 2202
rect 4968 2150 4980 2202
rect 5032 2150 5044 2202
rect 5096 2150 5108 2202
rect 5160 2150 14916 2202
rect 14968 2150 14980 2202
rect 15032 2150 15044 2202
rect 15096 2150 15108 2202
rect 15160 2150 24916 2202
rect 24968 2150 24980 2202
rect 25032 2150 25044 2202
rect 25096 2150 25108 2202
rect 25160 2150 27822 2202
rect 38 2128 27822 2150
<< via1 >>
rect 23794 21904 23846 21956
rect 25082 21904 25134 21956
rect 4916 21734 4968 21786
rect 4980 21734 5032 21786
rect 5044 21734 5096 21786
rect 5108 21734 5160 21786
rect 14916 21734 14968 21786
rect 14980 21734 15032 21786
rect 15044 21734 15096 21786
rect 15108 21734 15160 21786
rect 24916 21734 24968 21786
rect 24980 21734 25032 21786
rect 25044 21734 25096 21786
rect 25108 21734 25160 21786
rect 9916 21190 9968 21242
rect 9980 21190 10032 21242
rect 10044 21190 10096 21242
rect 10108 21190 10160 21242
rect 19916 21190 19968 21242
rect 19980 21190 20032 21242
rect 20044 21190 20096 21242
rect 20108 21190 20160 21242
rect 4916 20646 4968 20698
rect 4980 20646 5032 20698
rect 5044 20646 5096 20698
rect 5108 20646 5160 20698
rect 14916 20646 14968 20698
rect 14980 20646 15032 20698
rect 15044 20646 15096 20698
rect 15108 20646 15160 20698
rect 24916 20646 24968 20698
rect 24980 20646 25032 20698
rect 25044 20646 25096 20698
rect 25108 20646 25160 20698
rect 9916 20102 9968 20154
rect 9980 20102 10032 20154
rect 10044 20102 10096 20154
rect 10108 20102 10160 20154
rect 19916 20102 19968 20154
rect 19980 20102 20032 20154
rect 20044 20102 20096 20154
rect 20108 20102 20160 20154
rect 4916 19558 4968 19610
rect 4980 19558 5032 19610
rect 5044 19558 5096 19610
rect 5108 19558 5160 19610
rect 14916 19558 14968 19610
rect 14980 19558 15032 19610
rect 15044 19558 15096 19610
rect 15108 19558 15160 19610
rect 24916 19558 24968 19610
rect 24980 19558 25032 19610
rect 25044 19558 25096 19610
rect 25108 19558 25160 19610
rect 9916 19014 9968 19066
rect 9980 19014 10032 19066
rect 10044 19014 10096 19066
rect 10108 19014 10160 19066
rect 19916 19014 19968 19066
rect 19980 19014 20032 19066
rect 20044 19014 20096 19066
rect 20108 19014 20160 19066
rect 15330 18912 15382 18964
rect 15146 18819 15198 18828
rect 15146 18785 15164 18819
rect 15164 18785 15198 18819
rect 15146 18776 15198 18785
rect 4916 18470 4968 18522
rect 4980 18470 5032 18522
rect 5044 18470 5096 18522
rect 5108 18470 5160 18522
rect 14916 18470 14968 18522
rect 14980 18470 15032 18522
rect 15044 18470 15096 18522
rect 15108 18470 15160 18522
rect 24916 18470 24968 18522
rect 24980 18470 25032 18522
rect 25044 18470 25096 18522
rect 25108 18470 25160 18522
rect 13398 18411 13450 18420
rect 13398 18377 13407 18411
rect 13407 18377 13441 18411
rect 13441 18377 13450 18411
rect 13398 18368 13450 18377
rect 15238 18368 15290 18420
rect 9916 17926 9968 17978
rect 9980 17926 10032 17978
rect 10044 17926 10096 17978
rect 10108 17926 10160 17978
rect 19916 17926 19968 17978
rect 19980 17926 20032 17978
rect 20044 17926 20096 17978
rect 20108 17926 20160 17978
rect 4916 17382 4968 17434
rect 4980 17382 5032 17434
rect 5044 17382 5096 17434
rect 5108 17382 5160 17434
rect 14916 17382 14968 17434
rect 14980 17382 15032 17434
rect 15044 17382 15096 17434
rect 15108 17382 15160 17434
rect 24916 17382 24968 17434
rect 24980 17382 25032 17434
rect 25044 17382 25096 17434
rect 25108 17382 25160 17434
rect 9916 16838 9968 16890
rect 9980 16838 10032 16890
rect 10044 16838 10096 16890
rect 10108 16838 10160 16890
rect 19916 16838 19968 16890
rect 19980 16838 20032 16890
rect 20044 16838 20096 16890
rect 20108 16838 20160 16890
rect 4916 16294 4968 16346
rect 4980 16294 5032 16346
rect 5044 16294 5096 16346
rect 5108 16294 5160 16346
rect 14916 16294 14968 16346
rect 14980 16294 15032 16346
rect 15044 16294 15096 16346
rect 15108 16294 15160 16346
rect 24916 16294 24968 16346
rect 24980 16294 25032 16346
rect 25044 16294 25096 16346
rect 25108 16294 25160 16346
rect 9916 15750 9968 15802
rect 9980 15750 10032 15802
rect 10044 15750 10096 15802
rect 10108 15750 10160 15802
rect 19916 15750 19968 15802
rect 19980 15750 20032 15802
rect 20044 15750 20096 15802
rect 20108 15750 20160 15802
rect 4916 15206 4968 15258
rect 4980 15206 5032 15258
rect 5044 15206 5096 15258
rect 5108 15206 5160 15258
rect 14916 15206 14968 15258
rect 14980 15206 15032 15258
rect 15044 15206 15096 15258
rect 15108 15206 15160 15258
rect 24916 15206 24968 15258
rect 24980 15206 25032 15258
rect 25044 15206 25096 15258
rect 25108 15206 25160 15258
rect 9916 14662 9968 14714
rect 9980 14662 10032 14714
rect 10044 14662 10096 14714
rect 10108 14662 10160 14714
rect 19916 14662 19968 14714
rect 19980 14662 20032 14714
rect 20044 14662 20096 14714
rect 20108 14662 20160 14714
rect 4916 14118 4968 14170
rect 4980 14118 5032 14170
rect 5044 14118 5096 14170
rect 5108 14118 5160 14170
rect 14916 14118 14968 14170
rect 14980 14118 15032 14170
rect 15044 14118 15096 14170
rect 15108 14118 15160 14170
rect 24916 14118 24968 14170
rect 24980 14118 25032 14170
rect 25044 14118 25096 14170
rect 25108 14118 25160 14170
rect 9916 13574 9968 13626
rect 9980 13574 10032 13626
rect 10044 13574 10096 13626
rect 10108 13574 10160 13626
rect 19916 13574 19968 13626
rect 19980 13574 20032 13626
rect 20044 13574 20096 13626
rect 20108 13574 20160 13626
rect 4916 13030 4968 13082
rect 4980 13030 5032 13082
rect 5044 13030 5096 13082
rect 5108 13030 5160 13082
rect 14916 13030 14968 13082
rect 14980 13030 15032 13082
rect 15044 13030 15096 13082
rect 15108 13030 15160 13082
rect 24916 13030 24968 13082
rect 24980 13030 25032 13082
rect 25044 13030 25096 13082
rect 25108 13030 25160 13082
rect 9916 12486 9968 12538
rect 9980 12486 10032 12538
rect 10044 12486 10096 12538
rect 10108 12486 10160 12538
rect 19916 12486 19968 12538
rect 19980 12486 20032 12538
rect 20044 12486 20096 12538
rect 20108 12486 20160 12538
rect 4916 11942 4968 11994
rect 4980 11942 5032 11994
rect 5044 11942 5096 11994
rect 5108 11942 5160 11994
rect 14916 11942 14968 11994
rect 14980 11942 15032 11994
rect 15044 11942 15096 11994
rect 15108 11942 15160 11994
rect 24916 11942 24968 11994
rect 24980 11942 25032 11994
rect 25044 11942 25096 11994
rect 25108 11942 25160 11994
rect 9916 11398 9968 11450
rect 9980 11398 10032 11450
rect 10044 11398 10096 11450
rect 10108 11398 10160 11450
rect 19916 11398 19968 11450
rect 19980 11398 20032 11450
rect 20044 11398 20096 11450
rect 20108 11398 20160 11450
rect 22874 10999 22926 11008
rect 22874 10965 22883 10999
rect 22883 10965 22917 10999
rect 22917 10965 22926 10999
rect 22874 10956 22926 10965
rect 4916 10854 4968 10906
rect 4980 10854 5032 10906
rect 5044 10854 5096 10906
rect 5108 10854 5160 10906
rect 14916 10854 14968 10906
rect 14980 10854 15032 10906
rect 15044 10854 15096 10906
rect 15108 10854 15160 10906
rect 24916 10854 24968 10906
rect 24980 10854 25032 10906
rect 25044 10854 25096 10906
rect 25108 10854 25160 10906
rect 24438 10752 24490 10804
rect 10178 10727 10230 10736
rect 10178 10693 10187 10727
rect 10187 10693 10221 10727
rect 10221 10693 10230 10727
rect 10178 10684 10230 10693
rect 22874 10591 22926 10600
rect 22874 10557 22883 10591
rect 22883 10557 22917 10591
rect 22917 10557 22926 10591
rect 22874 10548 22926 10557
rect 22966 10548 23018 10600
rect 23886 10548 23938 10600
rect 10546 10455 10598 10464
rect 10546 10421 10555 10455
rect 10555 10421 10589 10455
rect 10589 10421 10598 10455
rect 10546 10412 10598 10421
rect 9916 10310 9968 10362
rect 9980 10310 10032 10362
rect 10044 10310 10096 10362
rect 10108 10310 10160 10362
rect 19916 10310 19968 10362
rect 19980 10310 20032 10362
rect 20044 10310 20096 10362
rect 20108 10310 20160 10362
rect 22966 10251 23018 10260
rect 22966 10217 22975 10251
rect 22975 10217 23009 10251
rect 23009 10217 23018 10251
rect 22966 10208 23018 10217
rect 4916 9766 4968 9818
rect 4980 9766 5032 9818
rect 5044 9766 5096 9818
rect 5108 9766 5160 9818
rect 14916 9766 14968 9818
rect 14980 9766 15032 9818
rect 15044 9766 15096 9818
rect 15108 9766 15160 9818
rect 24916 9766 24968 9818
rect 24980 9766 25032 9818
rect 25044 9766 25096 9818
rect 25108 9766 25160 9818
rect 9916 9222 9968 9274
rect 9980 9222 10032 9274
rect 10044 9222 10096 9274
rect 10108 9222 10160 9274
rect 19916 9222 19968 9274
rect 19980 9222 20032 9274
rect 20044 9222 20096 9274
rect 20108 9222 20160 9274
rect 4916 8678 4968 8730
rect 4980 8678 5032 8730
rect 5044 8678 5096 8730
rect 5108 8678 5160 8730
rect 14916 8678 14968 8730
rect 14980 8678 15032 8730
rect 15044 8678 15096 8730
rect 15108 8678 15160 8730
rect 24916 8678 24968 8730
rect 24980 8678 25032 8730
rect 25044 8678 25096 8730
rect 25108 8678 25160 8730
rect 9916 8134 9968 8186
rect 9980 8134 10032 8186
rect 10044 8134 10096 8186
rect 10108 8134 10160 8186
rect 19916 8134 19968 8186
rect 19980 8134 20032 8186
rect 20044 8134 20096 8186
rect 20108 8134 20160 8186
rect 4916 7590 4968 7642
rect 4980 7590 5032 7642
rect 5044 7590 5096 7642
rect 5108 7590 5160 7642
rect 14916 7590 14968 7642
rect 14980 7590 15032 7642
rect 15044 7590 15096 7642
rect 15108 7590 15160 7642
rect 24916 7590 24968 7642
rect 24980 7590 25032 7642
rect 25044 7590 25096 7642
rect 25108 7590 25160 7642
rect 9916 7046 9968 7098
rect 9980 7046 10032 7098
rect 10044 7046 10096 7098
rect 10108 7046 10160 7098
rect 19916 7046 19968 7098
rect 19980 7046 20032 7098
rect 20044 7046 20096 7098
rect 20108 7046 20160 7098
rect 4916 6502 4968 6554
rect 4980 6502 5032 6554
rect 5044 6502 5096 6554
rect 5108 6502 5160 6554
rect 14916 6502 14968 6554
rect 14980 6502 15032 6554
rect 15044 6502 15096 6554
rect 15108 6502 15160 6554
rect 24916 6502 24968 6554
rect 24980 6502 25032 6554
rect 25044 6502 25096 6554
rect 25108 6502 25160 6554
rect 9916 5958 9968 6010
rect 9980 5958 10032 6010
rect 10044 5958 10096 6010
rect 10108 5958 10160 6010
rect 19916 5958 19968 6010
rect 19980 5958 20032 6010
rect 20044 5958 20096 6010
rect 20108 5958 20160 6010
rect 4916 5414 4968 5466
rect 4980 5414 5032 5466
rect 5044 5414 5096 5466
rect 5108 5414 5160 5466
rect 14916 5414 14968 5466
rect 14980 5414 15032 5466
rect 15044 5414 15096 5466
rect 15108 5414 15160 5466
rect 24916 5414 24968 5466
rect 24980 5414 25032 5466
rect 25044 5414 25096 5466
rect 25108 5414 25160 5466
rect 9916 4870 9968 4922
rect 9980 4870 10032 4922
rect 10044 4870 10096 4922
rect 10108 4870 10160 4922
rect 19916 4870 19968 4922
rect 19980 4870 20032 4922
rect 20044 4870 20096 4922
rect 20108 4870 20160 4922
rect 4916 4326 4968 4378
rect 4980 4326 5032 4378
rect 5044 4326 5096 4378
rect 5108 4326 5160 4378
rect 14916 4326 14968 4378
rect 14980 4326 15032 4378
rect 15044 4326 15096 4378
rect 15108 4326 15160 4378
rect 24916 4326 24968 4378
rect 24980 4326 25032 4378
rect 25044 4326 25096 4378
rect 25108 4326 25160 4378
rect 9916 3782 9968 3834
rect 9980 3782 10032 3834
rect 10044 3782 10096 3834
rect 10108 3782 10160 3834
rect 19916 3782 19968 3834
rect 19980 3782 20032 3834
rect 20044 3782 20096 3834
rect 20108 3782 20160 3834
rect 4916 3238 4968 3290
rect 4980 3238 5032 3290
rect 5044 3238 5096 3290
rect 5108 3238 5160 3290
rect 14916 3238 14968 3290
rect 14980 3238 15032 3290
rect 15044 3238 15096 3290
rect 15108 3238 15160 3290
rect 24916 3238 24968 3290
rect 24980 3238 25032 3290
rect 25044 3238 25096 3290
rect 25108 3238 25160 3290
rect 9916 2694 9968 2746
rect 9980 2694 10032 2746
rect 10044 2694 10096 2746
rect 10108 2694 10160 2746
rect 19916 2694 19968 2746
rect 19980 2694 20032 2746
rect 20044 2694 20096 2746
rect 20108 2694 20160 2746
rect 20482 2635 20534 2644
rect 20482 2601 20491 2635
rect 20491 2601 20525 2635
rect 20525 2601 20534 2635
rect 20482 2592 20534 2601
rect 22046 2635 22098 2644
rect 22046 2601 22055 2635
rect 22055 2601 22089 2635
rect 22089 2601 22098 2635
rect 22046 2592 22098 2601
rect 23886 2320 23938 2372
rect 4916 2150 4968 2202
rect 4980 2150 5032 2202
rect 5044 2150 5096 2202
rect 5108 2150 5160 2202
rect 14916 2150 14968 2202
rect 14980 2150 15032 2202
rect 15044 2150 15096 2202
rect 15108 2150 15160 2202
rect 24916 2150 24968 2202
rect 24980 2150 25032 2202
rect 25044 2150 25096 2202
rect 25108 2150 25160 2202
<< metal2 >>
rect 2632 23520 2688 24000
rect 10084 23520 10140 24000
rect 17628 23520 17684 24000
rect 25080 23520 25136 24000
rect 2646 23474 2674 23520
rect 2646 23446 3042 23474
rect 3014 10577 3042 23446
rect 4890 21788 5186 21808
rect 4946 21786 4970 21788
rect 5026 21786 5050 21788
rect 5106 21786 5130 21788
rect 4968 21734 4970 21786
rect 5032 21734 5044 21786
rect 5106 21734 5108 21786
rect 4946 21732 4970 21734
rect 5026 21732 5050 21734
rect 5106 21732 5130 21734
rect 4890 21712 5186 21732
rect 10098 21434 10126 23520
rect 14890 21788 15186 21808
rect 14946 21786 14970 21788
rect 15026 21786 15050 21788
rect 15106 21786 15130 21788
rect 14968 21734 14970 21786
rect 15032 21734 15044 21786
rect 15106 21734 15108 21786
rect 14946 21732 14970 21734
rect 15026 21732 15050 21734
rect 15106 21732 15130 21734
rect 14890 21712 15186 21732
rect 10098 21406 10310 21434
rect 9890 21244 10186 21264
rect 9946 21242 9970 21244
rect 10026 21242 10050 21244
rect 10106 21242 10130 21244
rect 9968 21190 9970 21242
rect 10032 21190 10044 21242
rect 10106 21190 10108 21242
rect 9946 21188 9970 21190
rect 10026 21188 10050 21190
rect 10106 21188 10130 21190
rect 9890 21168 10186 21188
rect 4890 20700 5186 20720
rect 4946 20698 4970 20700
rect 5026 20698 5050 20700
rect 5106 20698 5130 20700
rect 4968 20646 4970 20698
rect 5032 20646 5044 20698
rect 5106 20646 5108 20698
rect 4946 20644 4970 20646
rect 5026 20644 5050 20646
rect 5106 20644 5130 20646
rect 4890 20624 5186 20644
rect 9890 20156 10186 20176
rect 9946 20154 9970 20156
rect 10026 20154 10050 20156
rect 10106 20154 10130 20156
rect 9968 20102 9970 20154
rect 10032 20102 10044 20154
rect 10106 20102 10108 20154
rect 9946 20100 9970 20102
rect 10026 20100 10050 20102
rect 10106 20100 10130 20102
rect 9890 20080 10186 20100
rect 4890 19612 5186 19632
rect 4946 19610 4970 19612
rect 5026 19610 5050 19612
rect 5106 19610 5130 19612
rect 4968 19558 4970 19610
rect 5032 19558 5044 19610
rect 5106 19558 5108 19610
rect 4946 19556 4970 19558
rect 5026 19556 5050 19558
rect 5106 19556 5130 19558
rect 4890 19536 5186 19556
rect 10282 19417 10310 21406
rect 14890 20700 15186 20720
rect 14946 20698 14970 20700
rect 15026 20698 15050 20700
rect 15106 20698 15130 20700
rect 14968 20646 14970 20698
rect 15032 20646 15044 20698
rect 15106 20646 15108 20698
rect 14946 20644 14970 20646
rect 15026 20644 15050 20646
rect 15106 20644 15130 20646
rect 14890 20624 15186 20644
rect 17642 20505 17670 23520
rect 25094 21962 25122 23520
rect 23794 21956 23846 21962
rect 23794 21898 23846 21904
rect 25082 21956 25134 21962
rect 25082 21898 25134 21904
rect 19890 21244 20186 21264
rect 19946 21242 19970 21244
rect 20026 21242 20050 21244
rect 20106 21242 20130 21244
rect 19968 21190 19970 21242
rect 20032 21190 20044 21242
rect 20106 21190 20108 21242
rect 19946 21188 19970 21190
rect 20026 21188 20050 21190
rect 20106 21188 20130 21190
rect 19890 21168 20186 21188
rect 15328 20496 15384 20505
rect 15328 20431 15384 20440
rect 17628 20496 17684 20505
rect 17628 20431 17684 20440
rect 14890 19612 15186 19632
rect 14946 19610 14970 19612
rect 15026 19610 15050 19612
rect 15106 19610 15130 19612
rect 14968 19558 14970 19610
rect 15032 19558 15044 19610
rect 15106 19558 15108 19610
rect 14946 19556 14970 19558
rect 15026 19556 15050 19558
rect 15106 19556 15130 19558
rect 14890 19536 15186 19556
rect 10268 19408 10324 19417
rect 10268 19343 10324 19352
rect 13396 19408 13452 19417
rect 13396 19343 13452 19352
rect 9890 19068 10186 19088
rect 9946 19066 9970 19068
rect 10026 19066 10050 19068
rect 10106 19066 10130 19068
rect 9968 19014 9970 19066
rect 10032 19014 10044 19066
rect 10106 19014 10108 19066
rect 9946 19012 9970 19014
rect 10026 19012 10050 19014
rect 10106 19012 10130 19014
rect 9890 18992 10186 19012
rect 4890 18524 5186 18544
rect 4946 18522 4970 18524
rect 5026 18522 5050 18524
rect 5106 18522 5130 18524
rect 4968 18470 4970 18522
rect 5032 18470 5044 18522
rect 5106 18470 5108 18522
rect 4946 18468 4970 18470
rect 5026 18468 5050 18470
rect 5106 18468 5130 18470
rect 4890 18448 5186 18468
rect 13410 18426 13438 19343
rect 15342 18970 15370 20431
rect 19890 20156 20186 20176
rect 19946 20154 19970 20156
rect 20026 20154 20050 20156
rect 20106 20154 20130 20156
rect 19968 20102 19970 20154
rect 20032 20102 20044 20154
rect 20106 20102 20108 20154
rect 19946 20100 19970 20102
rect 20026 20100 20050 20102
rect 20106 20100 20130 20102
rect 19890 20080 20186 20100
rect 19890 19068 20186 19088
rect 19946 19066 19970 19068
rect 20026 19066 20050 19068
rect 20106 19066 20130 19068
rect 19968 19014 19970 19066
rect 20032 19014 20044 19066
rect 20106 19014 20108 19066
rect 19946 19012 19970 19014
rect 20026 19012 20050 19014
rect 20106 19012 20130 19014
rect 19890 18992 20186 19012
rect 15330 18964 15382 18970
rect 15330 18906 15382 18912
rect 15144 18864 15200 18873
rect 15144 18799 15146 18808
rect 15198 18799 15200 18808
rect 15146 18770 15198 18776
rect 15158 18714 15186 18770
rect 15158 18686 15278 18714
rect 14890 18524 15186 18544
rect 14946 18522 14970 18524
rect 15026 18522 15050 18524
rect 15106 18522 15130 18524
rect 14968 18470 14970 18522
rect 15032 18470 15044 18522
rect 15106 18470 15108 18522
rect 14946 18468 14970 18470
rect 15026 18468 15050 18470
rect 15106 18468 15130 18470
rect 14890 18448 15186 18468
rect 15250 18426 15278 18686
rect 13398 18420 13450 18426
rect 13398 18362 13450 18368
rect 15238 18420 15290 18426
rect 15238 18362 15290 18368
rect 9890 17980 10186 18000
rect 9946 17978 9970 17980
rect 10026 17978 10050 17980
rect 10106 17978 10130 17980
rect 9968 17926 9970 17978
rect 10032 17926 10044 17978
rect 10106 17926 10108 17978
rect 9946 17924 9970 17926
rect 10026 17924 10050 17926
rect 10106 17924 10130 17926
rect 9890 17904 10186 17924
rect 19890 17980 20186 18000
rect 19946 17978 19970 17980
rect 20026 17978 20050 17980
rect 20106 17978 20130 17980
rect 19968 17926 19970 17978
rect 20032 17926 20044 17978
rect 20106 17926 20108 17978
rect 19946 17924 19970 17926
rect 20026 17924 20050 17926
rect 20106 17924 20130 17926
rect 19890 17904 20186 17924
rect 4890 17436 5186 17456
rect 4946 17434 4970 17436
rect 5026 17434 5050 17436
rect 5106 17434 5130 17436
rect 4968 17382 4970 17434
rect 5032 17382 5044 17434
rect 5106 17382 5108 17434
rect 4946 17380 4970 17382
rect 5026 17380 5050 17382
rect 5106 17380 5130 17382
rect 4890 17360 5186 17380
rect 14890 17436 15186 17456
rect 14946 17434 14970 17436
rect 15026 17434 15050 17436
rect 15106 17434 15130 17436
rect 14968 17382 14970 17434
rect 15032 17382 15044 17434
rect 15106 17382 15108 17434
rect 14946 17380 14970 17382
rect 15026 17380 15050 17382
rect 15106 17380 15130 17382
rect 14890 17360 15186 17380
rect 9890 16892 10186 16912
rect 9946 16890 9970 16892
rect 10026 16890 10050 16892
rect 10106 16890 10130 16892
rect 9968 16838 9970 16890
rect 10032 16838 10044 16890
rect 10106 16838 10108 16890
rect 9946 16836 9970 16838
rect 10026 16836 10050 16838
rect 10106 16836 10130 16838
rect 9890 16816 10186 16836
rect 19890 16892 20186 16912
rect 19946 16890 19970 16892
rect 20026 16890 20050 16892
rect 20106 16890 20130 16892
rect 19968 16838 19970 16890
rect 20032 16838 20044 16890
rect 20106 16838 20108 16890
rect 19946 16836 19970 16838
rect 20026 16836 20050 16838
rect 20106 16836 20130 16838
rect 19890 16816 20186 16836
rect 4890 16348 5186 16368
rect 4946 16346 4970 16348
rect 5026 16346 5050 16348
rect 5106 16346 5130 16348
rect 4968 16294 4970 16346
rect 5032 16294 5044 16346
rect 5106 16294 5108 16346
rect 4946 16292 4970 16294
rect 5026 16292 5050 16294
rect 5106 16292 5130 16294
rect 4890 16272 5186 16292
rect 14890 16348 15186 16368
rect 14946 16346 14970 16348
rect 15026 16346 15050 16348
rect 15106 16346 15130 16348
rect 14968 16294 14970 16346
rect 15032 16294 15044 16346
rect 15106 16294 15108 16346
rect 14946 16292 14970 16294
rect 15026 16292 15050 16294
rect 15106 16292 15130 16294
rect 14890 16272 15186 16292
rect 9890 15804 10186 15824
rect 9946 15802 9970 15804
rect 10026 15802 10050 15804
rect 10106 15802 10130 15804
rect 9968 15750 9970 15802
rect 10032 15750 10044 15802
rect 10106 15750 10108 15802
rect 9946 15748 9970 15750
rect 10026 15748 10050 15750
rect 10106 15748 10130 15750
rect 9890 15728 10186 15748
rect 19890 15804 20186 15824
rect 19946 15802 19970 15804
rect 20026 15802 20050 15804
rect 20106 15802 20130 15804
rect 19968 15750 19970 15802
rect 20032 15750 20044 15802
rect 20106 15750 20108 15802
rect 19946 15748 19970 15750
rect 20026 15748 20050 15750
rect 20106 15748 20130 15750
rect 19890 15728 20186 15748
rect 4890 15260 5186 15280
rect 4946 15258 4970 15260
rect 5026 15258 5050 15260
rect 5106 15258 5130 15260
rect 4968 15206 4970 15258
rect 5032 15206 5044 15258
rect 5106 15206 5108 15258
rect 4946 15204 4970 15206
rect 5026 15204 5050 15206
rect 5106 15204 5130 15206
rect 4890 15184 5186 15204
rect 14890 15260 15186 15280
rect 14946 15258 14970 15260
rect 15026 15258 15050 15260
rect 15106 15258 15130 15260
rect 14968 15206 14970 15258
rect 15032 15206 15044 15258
rect 15106 15206 15108 15258
rect 14946 15204 14970 15206
rect 15026 15204 15050 15206
rect 15106 15204 15130 15206
rect 14890 15184 15186 15204
rect 9890 14716 10186 14736
rect 9946 14714 9970 14716
rect 10026 14714 10050 14716
rect 10106 14714 10130 14716
rect 9968 14662 9970 14714
rect 10032 14662 10044 14714
rect 10106 14662 10108 14714
rect 9946 14660 9970 14662
rect 10026 14660 10050 14662
rect 10106 14660 10130 14662
rect 9890 14640 10186 14660
rect 19890 14716 20186 14736
rect 19946 14714 19970 14716
rect 20026 14714 20050 14716
rect 20106 14714 20130 14716
rect 19968 14662 19970 14714
rect 20032 14662 20044 14714
rect 20106 14662 20108 14714
rect 19946 14660 19970 14662
rect 20026 14660 20050 14662
rect 20106 14660 20130 14662
rect 19890 14640 20186 14660
rect 4890 14172 5186 14192
rect 4946 14170 4970 14172
rect 5026 14170 5050 14172
rect 5106 14170 5130 14172
rect 4968 14118 4970 14170
rect 5032 14118 5044 14170
rect 5106 14118 5108 14170
rect 4946 14116 4970 14118
rect 5026 14116 5050 14118
rect 5106 14116 5130 14118
rect 4890 14096 5186 14116
rect 14890 14172 15186 14192
rect 14946 14170 14970 14172
rect 15026 14170 15050 14172
rect 15106 14170 15130 14172
rect 14968 14118 14970 14170
rect 15032 14118 15044 14170
rect 15106 14118 15108 14170
rect 14946 14116 14970 14118
rect 15026 14116 15050 14118
rect 15106 14116 15130 14118
rect 14890 14096 15186 14116
rect 9890 13628 10186 13648
rect 9946 13626 9970 13628
rect 10026 13626 10050 13628
rect 10106 13626 10130 13628
rect 9968 13574 9970 13626
rect 10032 13574 10044 13626
rect 10106 13574 10108 13626
rect 9946 13572 9970 13574
rect 10026 13572 10050 13574
rect 10106 13572 10130 13574
rect 9890 13552 10186 13572
rect 19890 13628 20186 13648
rect 19946 13626 19970 13628
rect 20026 13626 20050 13628
rect 20106 13626 20130 13628
rect 19968 13574 19970 13626
rect 20032 13574 20044 13626
rect 20106 13574 20108 13626
rect 19946 13572 19970 13574
rect 20026 13572 20050 13574
rect 20106 13572 20130 13574
rect 19890 13552 20186 13572
rect 4890 13084 5186 13104
rect 4946 13082 4970 13084
rect 5026 13082 5050 13084
rect 5106 13082 5130 13084
rect 4968 13030 4970 13082
rect 5032 13030 5044 13082
rect 5106 13030 5108 13082
rect 4946 13028 4970 13030
rect 5026 13028 5050 13030
rect 5106 13028 5130 13030
rect 4890 13008 5186 13028
rect 14890 13084 15186 13104
rect 14946 13082 14970 13084
rect 15026 13082 15050 13084
rect 15106 13082 15130 13084
rect 14968 13030 14970 13082
rect 15032 13030 15044 13082
rect 15106 13030 15108 13082
rect 14946 13028 14970 13030
rect 15026 13028 15050 13030
rect 15106 13028 15130 13030
rect 14890 13008 15186 13028
rect 9890 12540 10186 12560
rect 9946 12538 9970 12540
rect 10026 12538 10050 12540
rect 10106 12538 10130 12540
rect 9968 12486 9970 12538
rect 10032 12486 10044 12538
rect 10106 12486 10108 12538
rect 9946 12484 9970 12486
rect 10026 12484 10050 12486
rect 10106 12484 10130 12486
rect 9890 12464 10186 12484
rect 19890 12540 20186 12560
rect 19946 12538 19970 12540
rect 20026 12538 20050 12540
rect 20106 12538 20130 12540
rect 19968 12486 19970 12538
rect 20032 12486 20044 12538
rect 20106 12486 20108 12538
rect 19946 12484 19970 12486
rect 20026 12484 20050 12486
rect 20106 12484 20130 12486
rect 19890 12464 20186 12484
rect 4890 11996 5186 12016
rect 4946 11994 4970 11996
rect 5026 11994 5050 11996
rect 5106 11994 5130 11996
rect 4968 11942 4970 11994
rect 5032 11942 5044 11994
rect 5106 11942 5108 11994
rect 4946 11940 4970 11942
rect 5026 11940 5050 11942
rect 5106 11940 5130 11942
rect 4890 11920 5186 11940
rect 14890 11996 15186 12016
rect 14946 11994 14970 11996
rect 15026 11994 15050 11996
rect 15106 11994 15130 11996
rect 14968 11942 14970 11994
rect 15032 11942 15044 11994
rect 15106 11942 15108 11994
rect 14946 11940 14970 11942
rect 15026 11940 15050 11942
rect 15106 11940 15130 11942
rect 14890 11920 15186 11940
rect 9890 11452 10186 11472
rect 9946 11450 9970 11452
rect 10026 11450 10050 11452
rect 10106 11450 10130 11452
rect 9968 11398 9970 11450
rect 10032 11398 10044 11450
rect 10106 11398 10108 11450
rect 9946 11396 9970 11398
rect 10026 11396 10050 11398
rect 10106 11396 10130 11398
rect 9890 11376 10186 11396
rect 19890 11452 20186 11472
rect 19946 11450 19970 11452
rect 20026 11450 20050 11452
rect 20106 11450 20130 11452
rect 19968 11398 19970 11450
rect 20032 11398 20044 11450
rect 20106 11398 20108 11450
rect 19946 11396 19970 11398
rect 20026 11396 20050 11398
rect 20106 11396 20130 11398
rect 19890 11376 20186 11396
rect 22874 11008 22926 11014
rect 22874 10950 22926 10956
rect 4890 10908 5186 10928
rect 4946 10906 4970 10908
rect 5026 10906 5050 10908
rect 5106 10906 5130 10908
rect 4968 10854 4970 10906
rect 5032 10854 5044 10906
rect 5106 10854 5108 10906
rect 4946 10852 4970 10854
rect 5026 10852 5050 10854
rect 5106 10852 5130 10854
rect 4890 10832 5186 10852
rect 14890 10908 15186 10928
rect 14946 10906 14970 10908
rect 15026 10906 15050 10908
rect 15106 10906 15130 10908
rect 14968 10854 14970 10906
rect 15032 10854 15044 10906
rect 15106 10854 15108 10906
rect 14946 10852 14970 10854
rect 15026 10852 15050 10854
rect 15106 10852 15130 10854
rect 14890 10832 15186 10852
rect 10178 10736 10230 10742
rect 10178 10678 10230 10684
rect 10190 10577 10218 10678
rect 22886 10606 22914 10950
rect 22874 10600 22926 10606
rect 3000 10568 3056 10577
rect 3000 10503 3056 10512
rect 10176 10568 10232 10577
rect 22874 10542 22926 10548
rect 22966 10600 23018 10606
rect 22966 10542 23018 10548
rect 10176 10503 10232 10512
rect 10546 10464 10598 10470
rect 10546 10406 10598 10412
rect 9890 10364 10186 10384
rect 9946 10362 9970 10364
rect 10026 10362 10050 10364
rect 10106 10362 10130 10364
rect 9968 10310 9970 10362
rect 10032 10310 10044 10362
rect 10106 10310 10108 10362
rect 9946 10308 9970 10310
rect 10026 10308 10050 10310
rect 10106 10308 10130 10310
rect 9890 10288 10186 10308
rect 4890 9820 5186 9840
rect 4946 9818 4970 9820
rect 5026 9818 5050 9820
rect 5106 9818 5130 9820
rect 4968 9766 4970 9818
rect 5032 9766 5044 9818
rect 5106 9766 5108 9818
rect 4946 9764 4970 9766
rect 5026 9764 5050 9766
rect 5106 9764 5130 9766
rect 4890 9744 5186 9764
rect 9890 9276 10186 9296
rect 9946 9274 9970 9276
rect 10026 9274 10050 9276
rect 10106 9274 10130 9276
rect 9968 9222 9970 9274
rect 10032 9222 10044 9274
rect 10106 9222 10108 9274
rect 9946 9220 9970 9222
rect 10026 9220 10050 9222
rect 10106 9220 10130 9222
rect 9890 9200 10186 9220
rect 4890 8732 5186 8752
rect 4946 8730 4970 8732
rect 5026 8730 5050 8732
rect 5106 8730 5130 8732
rect 4968 8678 4970 8730
rect 5032 8678 5044 8730
rect 5106 8678 5108 8730
rect 4946 8676 4970 8678
rect 5026 8676 5050 8678
rect 5106 8676 5130 8678
rect 4890 8656 5186 8676
rect 9890 8188 10186 8208
rect 9946 8186 9970 8188
rect 10026 8186 10050 8188
rect 10106 8186 10130 8188
rect 9968 8134 9970 8186
rect 10032 8134 10044 8186
rect 10106 8134 10108 8186
rect 9946 8132 9970 8134
rect 10026 8132 10050 8134
rect 10106 8132 10130 8134
rect 9890 8112 10186 8132
rect 4890 7644 5186 7664
rect 4946 7642 4970 7644
rect 5026 7642 5050 7644
rect 5106 7642 5130 7644
rect 4968 7590 4970 7642
rect 5032 7590 5044 7642
rect 5106 7590 5108 7642
rect 4946 7588 4970 7590
rect 5026 7588 5050 7590
rect 5106 7588 5130 7590
rect 4890 7568 5186 7588
rect 9890 7100 10186 7120
rect 9946 7098 9970 7100
rect 10026 7098 10050 7100
rect 10106 7098 10130 7100
rect 9968 7046 9970 7098
rect 10032 7046 10044 7098
rect 10106 7046 10108 7098
rect 9946 7044 9970 7046
rect 10026 7044 10050 7046
rect 10106 7044 10130 7046
rect 9890 7024 10186 7044
rect 4890 6556 5186 6576
rect 4946 6554 4970 6556
rect 5026 6554 5050 6556
rect 5106 6554 5130 6556
rect 4968 6502 4970 6554
rect 5032 6502 5044 6554
rect 5106 6502 5108 6554
rect 4946 6500 4970 6502
rect 5026 6500 5050 6502
rect 5106 6500 5130 6502
rect 4890 6480 5186 6500
rect 9890 6012 10186 6032
rect 9946 6010 9970 6012
rect 10026 6010 10050 6012
rect 10106 6010 10130 6012
rect 9968 5958 9970 6010
rect 10032 5958 10044 6010
rect 10106 5958 10108 6010
rect 9946 5956 9970 5958
rect 10026 5956 10050 5958
rect 10106 5956 10130 5958
rect 9890 5936 10186 5956
rect 10558 5681 10586 10406
rect 19890 10364 20186 10384
rect 19946 10362 19970 10364
rect 20026 10362 20050 10364
rect 20106 10362 20130 10364
rect 19968 10310 19970 10362
rect 20032 10310 20044 10362
rect 20106 10310 20108 10362
rect 19946 10308 19970 10310
rect 20026 10308 20050 10310
rect 20106 10308 20130 10310
rect 19890 10288 20186 10308
rect 14890 9820 15186 9840
rect 14946 9818 14970 9820
rect 15026 9818 15050 9820
rect 15106 9818 15130 9820
rect 14968 9766 14970 9818
rect 15032 9766 15044 9818
rect 15106 9766 15108 9818
rect 14946 9764 14970 9766
rect 15026 9764 15050 9766
rect 15106 9764 15130 9766
rect 14890 9744 15186 9764
rect 19890 9276 20186 9296
rect 19946 9274 19970 9276
rect 20026 9274 20050 9276
rect 20106 9274 20130 9276
rect 19968 9222 19970 9274
rect 20032 9222 20044 9274
rect 20106 9222 20108 9274
rect 19946 9220 19970 9222
rect 20026 9220 20050 9222
rect 20106 9220 20130 9222
rect 19890 9200 20186 9220
rect 14890 8732 15186 8752
rect 14946 8730 14970 8732
rect 15026 8730 15050 8732
rect 15106 8730 15130 8732
rect 14968 8678 14970 8730
rect 15032 8678 15044 8730
rect 15106 8678 15108 8730
rect 14946 8676 14970 8678
rect 15026 8676 15050 8678
rect 15106 8676 15130 8678
rect 14890 8656 15186 8676
rect 19890 8188 20186 8208
rect 19946 8186 19970 8188
rect 20026 8186 20050 8188
rect 20106 8186 20130 8188
rect 19968 8134 19970 8186
rect 20032 8134 20044 8186
rect 20106 8134 20108 8186
rect 19946 8132 19970 8134
rect 20026 8132 20050 8134
rect 20106 8132 20130 8134
rect 19890 8112 20186 8132
rect 14890 7644 15186 7664
rect 14946 7642 14970 7644
rect 15026 7642 15050 7644
rect 15106 7642 15130 7644
rect 14968 7590 14970 7642
rect 15032 7590 15044 7642
rect 15106 7590 15108 7642
rect 14946 7588 14970 7590
rect 15026 7588 15050 7590
rect 15106 7588 15130 7590
rect 14890 7568 15186 7588
rect 19890 7100 20186 7120
rect 19946 7098 19970 7100
rect 20026 7098 20050 7100
rect 20106 7098 20130 7100
rect 19968 7046 19970 7098
rect 20032 7046 20044 7098
rect 20106 7046 20108 7098
rect 19946 7044 19970 7046
rect 20026 7044 20050 7046
rect 20106 7044 20130 7046
rect 19890 7024 20186 7044
rect 14890 6556 15186 6576
rect 14946 6554 14970 6556
rect 15026 6554 15050 6556
rect 15106 6554 15130 6556
rect 14968 6502 14970 6554
rect 15032 6502 15044 6554
rect 15106 6502 15108 6554
rect 14946 6500 14970 6502
rect 15026 6500 15050 6502
rect 15106 6500 15130 6502
rect 14890 6480 15186 6500
rect 19890 6012 20186 6032
rect 19946 6010 19970 6012
rect 20026 6010 20050 6012
rect 20106 6010 20130 6012
rect 19968 5958 19970 6010
rect 20032 5958 20044 6010
rect 20106 5958 20108 6010
rect 19946 5956 19970 5958
rect 20026 5956 20050 5958
rect 20106 5956 20130 5958
rect 19890 5936 20186 5956
rect 10544 5672 10600 5681
rect 10544 5607 10600 5616
rect 13856 5672 13912 5681
rect 13856 5607 13912 5616
rect 4890 5468 5186 5488
rect 4946 5466 4970 5468
rect 5026 5466 5050 5468
rect 5106 5466 5130 5468
rect 4968 5414 4970 5466
rect 5032 5414 5044 5466
rect 5106 5414 5108 5466
rect 4946 5412 4970 5414
rect 5026 5412 5050 5414
rect 5106 5412 5130 5414
rect 4890 5392 5186 5412
rect 9890 4924 10186 4944
rect 9946 4922 9970 4924
rect 10026 4922 10050 4924
rect 10106 4922 10130 4924
rect 9968 4870 9970 4922
rect 10032 4870 10044 4922
rect 10106 4870 10108 4922
rect 9946 4868 9970 4870
rect 10026 4868 10050 4870
rect 10106 4868 10130 4870
rect 9890 4848 10186 4868
rect 4890 4380 5186 4400
rect 4946 4378 4970 4380
rect 5026 4378 5050 4380
rect 5106 4378 5130 4380
rect 4968 4326 4970 4378
rect 5032 4326 5044 4378
rect 5106 4326 5108 4378
rect 4946 4324 4970 4326
rect 5026 4324 5050 4326
rect 5106 4324 5130 4326
rect 4890 4304 5186 4324
rect 9890 3836 10186 3856
rect 9946 3834 9970 3836
rect 10026 3834 10050 3836
rect 10106 3834 10130 3836
rect 9968 3782 9970 3834
rect 10032 3782 10044 3834
rect 10106 3782 10108 3834
rect 9946 3780 9970 3782
rect 10026 3780 10050 3782
rect 10106 3780 10130 3782
rect 9890 3760 10186 3780
rect 4890 3292 5186 3312
rect 4946 3290 4970 3292
rect 5026 3290 5050 3292
rect 5106 3290 5130 3292
rect 4968 3238 4970 3290
rect 5032 3238 5044 3290
rect 5106 3238 5108 3290
rect 4946 3236 4970 3238
rect 5026 3236 5050 3238
rect 5106 3236 5130 3238
rect 4890 3216 5186 3236
rect 3920 2952 3976 2961
rect 3920 2887 3976 2896
rect 3934 480 3962 2887
rect 9890 2748 10186 2768
rect 9946 2746 9970 2748
rect 10026 2746 10050 2748
rect 10106 2746 10130 2748
rect 9968 2694 9970 2746
rect 10032 2694 10044 2746
rect 10106 2694 10108 2746
rect 9946 2692 9970 2694
rect 10026 2692 10050 2694
rect 10106 2692 10130 2694
rect 9890 2672 10186 2692
rect 4890 2204 5186 2224
rect 4946 2202 4970 2204
rect 5026 2202 5050 2204
rect 5106 2202 5130 2204
rect 4968 2150 4970 2202
rect 5032 2150 5044 2202
rect 5106 2150 5108 2202
rect 4946 2148 4970 2150
rect 5026 2148 5050 2150
rect 5106 2148 5130 2150
rect 4890 2128 5186 2148
rect 13870 480 13898 5607
rect 14890 5468 15186 5488
rect 14946 5466 14970 5468
rect 15026 5466 15050 5468
rect 15106 5466 15130 5468
rect 14968 5414 14970 5466
rect 15032 5414 15044 5466
rect 15106 5414 15108 5466
rect 14946 5412 14970 5414
rect 15026 5412 15050 5414
rect 15106 5412 15130 5414
rect 14890 5392 15186 5412
rect 19890 4924 20186 4944
rect 19946 4922 19970 4924
rect 20026 4922 20050 4924
rect 20106 4922 20130 4924
rect 19968 4870 19970 4922
rect 20032 4870 20044 4922
rect 20106 4870 20108 4922
rect 19946 4868 19970 4870
rect 20026 4868 20050 4870
rect 20106 4868 20130 4870
rect 19890 4848 20186 4868
rect 14890 4380 15186 4400
rect 14946 4378 14970 4380
rect 15026 4378 15050 4380
rect 15106 4378 15130 4380
rect 14968 4326 14970 4378
rect 15032 4326 15044 4378
rect 15106 4326 15108 4378
rect 14946 4324 14970 4326
rect 15026 4324 15050 4326
rect 15106 4324 15130 4326
rect 14890 4304 15186 4324
rect 22886 4049 22914 10542
rect 22978 10266 23006 10542
rect 22966 10260 23018 10266
rect 22966 10202 23018 10208
rect 22872 4040 22928 4049
rect 22872 3975 22928 3984
rect 19890 3836 20186 3856
rect 19946 3834 19970 3836
rect 20026 3834 20050 3836
rect 20106 3834 20130 3836
rect 19968 3782 19970 3834
rect 20032 3782 20044 3834
rect 20106 3782 20108 3834
rect 19946 3780 19970 3782
rect 20026 3780 20050 3782
rect 20106 3780 20130 3782
rect 19890 3760 20186 3780
rect 14890 3292 15186 3312
rect 14946 3290 14970 3292
rect 15026 3290 15050 3292
rect 15106 3290 15130 3292
rect 14968 3238 14970 3290
rect 15032 3238 15044 3290
rect 15106 3238 15108 3290
rect 14946 3236 14970 3238
rect 15026 3236 15050 3238
rect 15106 3236 15130 3238
rect 14890 3216 15186 3236
rect 20480 2952 20536 2961
rect 20480 2887 20536 2896
rect 19890 2748 20186 2768
rect 19946 2746 19970 2748
rect 20026 2746 20050 2748
rect 20106 2746 20130 2748
rect 19968 2694 19970 2746
rect 20032 2694 20044 2746
rect 20106 2694 20108 2746
rect 19946 2692 19970 2694
rect 20026 2692 20050 2694
rect 20106 2692 20130 2694
rect 19890 2672 20186 2692
rect 20494 2650 20522 2887
rect 23806 2689 23834 21898
rect 24890 21788 25186 21808
rect 24946 21786 24970 21788
rect 25026 21786 25050 21788
rect 25106 21786 25130 21788
rect 24968 21734 24970 21786
rect 25032 21734 25044 21786
rect 25106 21734 25108 21786
rect 24946 21732 24970 21734
rect 25026 21732 25050 21734
rect 25106 21732 25130 21734
rect 24890 21712 25186 21732
rect 24890 20700 25186 20720
rect 24946 20698 24970 20700
rect 25026 20698 25050 20700
rect 25106 20698 25130 20700
rect 24968 20646 24970 20698
rect 25032 20646 25044 20698
rect 25106 20646 25108 20698
rect 24946 20644 24970 20646
rect 25026 20644 25050 20646
rect 25106 20644 25130 20646
rect 24890 20624 25186 20644
rect 24436 19952 24492 19961
rect 24436 19887 24492 19896
rect 24450 18873 24478 19887
rect 24890 19612 25186 19632
rect 24946 19610 24970 19612
rect 25026 19610 25050 19612
rect 25106 19610 25130 19612
rect 24968 19558 24970 19610
rect 25032 19558 25044 19610
rect 25106 19558 25108 19610
rect 24946 19556 24970 19558
rect 25026 19556 25050 19558
rect 25106 19556 25130 19558
rect 24890 19536 25186 19556
rect 24436 18864 24492 18873
rect 24436 18799 24492 18808
rect 23884 11792 23940 11801
rect 23884 11727 23940 11736
rect 23898 10606 23926 11727
rect 24450 10810 24478 18799
rect 24890 18524 25186 18544
rect 24946 18522 24970 18524
rect 25026 18522 25050 18524
rect 25106 18522 25130 18524
rect 24968 18470 24970 18522
rect 25032 18470 25044 18522
rect 25106 18470 25108 18522
rect 24946 18468 24970 18470
rect 25026 18468 25050 18470
rect 25106 18468 25130 18470
rect 24890 18448 25186 18468
rect 24890 17436 25186 17456
rect 24946 17434 24970 17436
rect 25026 17434 25050 17436
rect 25106 17434 25130 17436
rect 24968 17382 24970 17434
rect 25032 17382 25044 17434
rect 25106 17382 25108 17434
rect 24946 17380 24970 17382
rect 25026 17380 25050 17382
rect 25106 17380 25130 17382
rect 24890 17360 25186 17380
rect 24890 16348 25186 16368
rect 24946 16346 24970 16348
rect 25026 16346 25050 16348
rect 25106 16346 25130 16348
rect 24968 16294 24970 16346
rect 25032 16294 25044 16346
rect 25106 16294 25108 16346
rect 24946 16292 24970 16294
rect 25026 16292 25050 16294
rect 25106 16292 25130 16294
rect 24890 16272 25186 16292
rect 24890 15260 25186 15280
rect 24946 15258 24970 15260
rect 25026 15258 25050 15260
rect 25106 15258 25130 15260
rect 24968 15206 24970 15258
rect 25032 15206 25044 15258
rect 25106 15206 25108 15258
rect 24946 15204 24970 15206
rect 25026 15204 25050 15206
rect 25106 15204 25130 15206
rect 24890 15184 25186 15204
rect 24890 14172 25186 14192
rect 24946 14170 24970 14172
rect 25026 14170 25050 14172
rect 25106 14170 25130 14172
rect 24968 14118 24970 14170
rect 25032 14118 25044 14170
rect 25106 14118 25108 14170
rect 24946 14116 24970 14118
rect 25026 14116 25050 14118
rect 25106 14116 25130 14118
rect 24890 14096 25186 14116
rect 24890 13084 25186 13104
rect 24946 13082 24970 13084
rect 25026 13082 25050 13084
rect 25106 13082 25130 13084
rect 24968 13030 24970 13082
rect 25032 13030 25044 13082
rect 25106 13030 25108 13082
rect 24946 13028 24970 13030
rect 25026 13028 25050 13030
rect 25106 13028 25130 13030
rect 24890 13008 25186 13028
rect 24890 11996 25186 12016
rect 24946 11994 24970 11996
rect 25026 11994 25050 11996
rect 25106 11994 25130 11996
rect 24968 11942 24970 11994
rect 25032 11942 25044 11994
rect 25106 11942 25108 11994
rect 24946 11940 24970 11942
rect 25026 11940 25050 11942
rect 25106 11940 25130 11942
rect 24890 11920 25186 11940
rect 24890 10908 25186 10928
rect 24946 10906 24970 10908
rect 25026 10906 25050 10908
rect 25106 10906 25130 10908
rect 24968 10854 24970 10906
rect 25032 10854 25044 10906
rect 25106 10854 25108 10906
rect 24946 10852 24970 10854
rect 25026 10852 25050 10854
rect 25106 10852 25130 10854
rect 24890 10832 25186 10852
rect 24438 10804 24490 10810
rect 24438 10746 24490 10752
rect 23886 10600 23938 10606
rect 23886 10542 23938 10548
rect 24890 9820 25186 9840
rect 24946 9818 24970 9820
rect 25026 9818 25050 9820
rect 25106 9818 25130 9820
rect 24968 9766 24970 9818
rect 25032 9766 25044 9818
rect 25106 9766 25108 9818
rect 24946 9764 24970 9766
rect 25026 9764 25050 9766
rect 25106 9764 25130 9766
rect 24890 9744 25186 9764
rect 24890 8732 25186 8752
rect 24946 8730 24970 8732
rect 25026 8730 25050 8732
rect 25106 8730 25130 8732
rect 24968 8678 24970 8730
rect 25032 8678 25044 8730
rect 25106 8678 25108 8730
rect 24946 8676 24970 8678
rect 25026 8676 25050 8678
rect 25106 8676 25130 8678
rect 24890 8656 25186 8676
rect 24890 7644 25186 7664
rect 24946 7642 24970 7644
rect 25026 7642 25050 7644
rect 25106 7642 25130 7644
rect 24968 7590 24970 7642
rect 25032 7590 25044 7642
rect 25106 7590 25108 7642
rect 24946 7588 24970 7590
rect 25026 7588 25050 7590
rect 25106 7588 25130 7590
rect 24890 7568 25186 7588
rect 24890 6556 25186 6576
rect 24946 6554 24970 6556
rect 25026 6554 25050 6556
rect 25106 6554 25130 6556
rect 24968 6502 24970 6554
rect 25032 6502 25044 6554
rect 25106 6502 25108 6554
rect 24946 6500 24970 6502
rect 25026 6500 25050 6502
rect 25106 6500 25130 6502
rect 24890 6480 25186 6500
rect 24890 5468 25186 5488
rect 24946 5466 24970 5468
rect 25026 5466 25050 5468
rect 25106 5466 25130 5468
rect 24968 5414 24970 5466
rect 25032 5414 25044 5466
rect 25106 5414 25108 5466
rect 24946 5412 24970 5414
rect 25026 5412 25050 5414
rect 25106 5412 25130 5414
rect 24890 5392 25186 5412
rect 24890 4380 25186 4400
rect 24946 4378 24970 4380
rect 25026 4378 25050 4380
rect 25106 4378 25130 4380
rect 24968 4326 24970 4378
rect 25032 4326 25044 4378
rect 25106 4326 25108 4378
rect 24946 4324 24970 4326
rect 25026 4324 25050 4326
rect 25106 4324 25130 4326
rect 24890 4304 25186 4324
rect 24890 3292 25186 3312
rect 24946 3290 24970 3292
rect 25026 3290 25050 3292
rect 25106 3290 25130 3292
rect 24968 3238 24970 3290
rect 25032 3238 25044 3290
rect 25106 3238 25108 3290
rect 24946 3236 24970 3238
rect 25026 3236 25050 3238
rect 25106 3236 25130 3238
rect 24890 3216 25186 3236
rect 22044 2680 22100 2689
rect 20482 2644 20534 2650
rect 22044 2615 22046 2624
rect 20482 2586 20534 2592
rect 22098 2615 22100 2624
rect 23792 2680 23848 2689
rect 23792 2615 23848 2624
rect 22046 2586 22098 2592
rect 23886 2372 23938 2378
rect 23886 2314 23938 2320
rect 14890 2204 15186 2224
rect 14946 2202 14970 2204
rect 15026 2202 15050 2204
rect 15106 2202 15130 2204
rect 14968 2150 14970 2202
rect 15032 2150 15044 2202
rect 15106 2150 15108 2202
rect 14946 2148 14970 2150
rect 15026 2148 15050 2150
rect 15106 2148 15130 2150
rect 14890 2128 15186 2148
rect 23898 480 23926 2314
rect 24890 2204 25186 2224
rect 24946 2202 24970 2204
rect 25026 2202 25050 2204
rect 25106 2202 25130 2204
rect 24968 2150 24970 2202
rect 25032 2150 25044 2202
rect 25106 2150 25108 2202
rect 24946 2148 24970 2150
rect 25026 2148 25050 2150
rect 25106 2148 25130 2150
rect 24890 2128 25186 2148
rect 3920 0 3976 480
rect 13856 0 13912 480
rect 23884 0 23940 480
<< via2 >>
rect 4890 21786 4946 21788
rect 4970 21786 5026 21788
rect 5050 21786 5106 21788
rect 5130 21786 5186 21788
rect 4890 21734 4916 21786
rect 4916 21734 4946 21786
rect 4970 21734 4980 21786
rect 4980 21734 5026 21786
rect 5050 21734 5096 21786
rect 5096 21734 5106 21786
rect 5130 21734 5160 21786
rect 5160 21734 5186 21786
rect 4890 21732 4946 21734
rect 4970 21732 5026 21734
rect 5050 21732 5106 21734
rect 5130 21732 5186 21734
rect 14890 21786 14946 21788
rect 14970 21786 15026 21788
rect 15050 21786 15106 21788
rect 15130 21786 15186 21788
rect 14890 21734 14916 21786
rect 14916 21734 14946 21786
rect 14970 21734 14980 21786
rect 14980 21734 15026 21786
rect 15050 21734 15096 21786
rect 15096 21734 15106 21786
rect 15130 21734 15160 21786
rect 15160 21734 15186 21786
rect 14890 21732 14946 21734
rect 14970 21732 15026 21734
rect 15050 21732 15106 21734
rect 15130 21732 15186 21734
rect 9890 21242 9946 21244
rect 9970 21242 10026 21244
rect 10050 21242 10106 21244
rect 10130 21242 10186 21244
rect 9890 21190 9916 21242
rect 9916 21190 9946 21242
rect 9970 21190 9980 21242
rect 9980 21190 10026 21242
rect 10050 21190 10096 21242
rect 10096 21190 10106 21242
rect 10130 21190 10160 21242
rect 10160 21190 10186 21242
rect 9890 21188 9946 21190
rect 9970 21188 10026 21190
rect 10050 21188 10106 21190
rect 10130 21188 10186 21190
rect 4890 20698 4946 20700
rect 4970 20698 5026 20700
rect 5050 20698 5106 20700
rect 5130 20698 5186 20700
rect 4890 20646 4916 20698
rect 4916 20646 4946 20698
rect 4970 20646 4980 20698
rect 4980 20646 5026 20698
rect 5050 20646 5096 20698
rect 5096 20646 5106 20698
rect 5130 20646 5160 20698
rect 5160 20646 5186 20698
rect 4890 20644 4946 20646
rect 4970 20644 5026 20646
rect 5050 20644 5106 20646
rect 5130 20644 5186 20646
rect 9890 20154 9946 20156
rect 9970 20154 10026 20156
rect 10050 20154 10106 20156
rect 10130 20154 10186 20156
rect 9890 20102 9916 20154
rect 9916 20102 9946 20154
rect 9970 20102 9980 20154
rect 9980 20102 10026 20154
rect 10050 20102 10096 20154
rect 10096 20102 10106 20154
rect 10130 20102 10160 20154
rect 10160 20102 10186 20154
rect 9890 20100 9946 20102
rect 9970 20100 10026 20102
rect 10050 20100 10106 20102
rect 10130 20100 10186 20102
rect 4890 19610 4946 19612
rect 4970 19610 5026 19612
rect 5050 19610 5106 19612
rect 5130 19610 5186 19612
rect 4890 19558 4916 19610
rect 4916 19558 4946 19610
rect 4970 19558 4980 19610
rect 4980 19558 5026 19610
rect 5050 19558 5096 19610
rect 5096 19558 5106 19610
rect 5130 19558 5160 19610
rect 5160 19558 5186 19610
rect 4890 19556 4946 19558
rect 4970 19556 5026 19558
rect 5050 19556 5106 19558
rect 5130 19556 5186 19558
rect 14890 20698 14946 20700
rect 14970 20698 15026 20700
rect 15050 20698 15106 20700
rect 15130 20698 15186 20700
rect 14890 20646 14916 20698
rect 14916 20646 14946 20698
rect 14970 20646 14980 20698
rect 14980 20646 15026 20698
rect 15050 20646 15096 20698
rect 15096 20646 15106 20698
rect 15130 20646 15160 20698
rect 15160 20646 15186 20698
rect 14890 20644 14946 20646
rect 14970 20644 15026 20646
rect 15050 20644 15106 20646
rect 15130 20644 15186 20646
rect 19890 21242 19946 21244
rect 19970 21242 20026 21244
rect 20050 21242 20106 21244
rect 20130 21242 20186 21244
rect 19890 21190 19916 21242
rect 19916 21190 19946 21242
rect 19970 21190 19980 21242
rect 19980 21190 20026 21242
rect 20050 21190 20096 21242
rect 20096 21190 20106 21242
rect 20130 21190 20160 21242
rect 20160 21190 20186 21242
rect 19890 21188 19946 21190
rect 19970 21188 20026 21190
rect 20050 21188 20106 21190
rect 20130 21188 20186 21190
rect 15328 20440 15384 20496
rect 17628 20440 17684 20496
rect 14890 19610 14946 19612
rect 14970 19610 15026 19612
rect 15050 19610 15106 19612
rect 15130 19610 15186 19612
rect 14890 19558 14916 19610
rect 14916 19558 14946 19610
rect 14970 19558 14980 19610
rect 14980 19558 15026 19610
rect 15050 19558 15096 19610
rect 15096 19558 15106 19610
rect 15130 19558 15160 19610
rect 15160 19558 15186 19610
rect 14890 19556 14946 19558
rect 14970 19556 15026 19558
rect 15050 19556 15106 19558
rect 15130 19556 15186 19558
rect 10268 19352 10324 19408
rect 13396 19352 13452 19408
rect 9890 19066 9946 19068
rect 9970 19066 10026 19068
rect 10050 19066 10106 19068
rect 10130 19066 10186 19068
rect 9890 19014 9916 19066
rect 9916 19014 9946 19066
rect 9970 19014 9980 19066
rect 9980 19014 10026 19066
rect 10050 19014 10096 19066
rect 10096 19014 10106 19066
rect 10130 19014 10160 19066
rect 10160 19014 10186 19066
rect 9890 19012 9946 19014
rect 9970 19012 10026 19014
rect 10050 19012 10106 19014
rect 10130 19012 10186 19014
rect 4890 18522 4946 18524
rect 4970 18522 5026 18524
rect 5050 18522 5106 18524
rect 5130 18522 5186 18524
rect 4890 18470 4916 18522
rect 4916 18470 4946 18522
rect 4970 18470 4980 18522
rect 4980 18470 5026 18522
rect 5050 18470 5096 18522
rect 5096 18470 5106 18522
rect 5130 18470 5160 18522
rect 5160 18470 5186 18522
rect 4890 18468 4946 18470
rect 4970 18468 5026 18470
rect 5050 18468 5106 18470
rect 5130 18468 5186 18470
rect 19890 20154 19946 20156
rect 19970 20154 20026 20156
rect 20050 20154 20106 20156
rect 20130 20154 20186 20156
rect 19890 20102 19916 20154
rect 19916 20102 19946 20154
rect 19970 20102 19980 20154
rect 19980 20102 20026 20154
rect 20050 20102 20096 20154
rect 20096 20102 20106 20154
rect 20130 20102 20160 20154
rect 20160 20102 20186 20154
rect 19890 20100 19946 20102
rect 19970 20100 20026 20102
rect 20050 20100 20106 20102
rect 20130 20100 20186 20102
rect 19890 19066 19946 19068
rect 19970 19066 20026 19068
rect 20050 19066 20106 19068
rect 20130 19066 20186 19068
rect 19890 19014 19916 19066
rect 19916 19014 19946 19066
rect 19970 19014 19980 19066
rect 19980 19014 20026 19066
rect 20050 19014 20096 19066
rect 20096 19014 20106 19066
rect 20130 19014 20160 19066
rect 20160 19014 20186 19066
rect 19890 19012 19946 19014
rect 19970 19012 20026 19014
rect 20050 19012 20106 19014
rect 20130 19012 20186 19014
rect 15144 18828 15200 18864
rect 15144 18808 15146 18828
rect 15146 18808 15198 18828
rect 15198 18808 15200 18828
rect 14890 18522 14946 18524
rect 14970 18522 15026 18524
rect 15050 18522 15106 18524
rect 15130 18522 15186 18524
rect 14890 18470 14916 18522
rect 14916 18470 14946 18522
rect 14970 18470 14980 18522
rect 14980 18470 15026 18522
rect 15050 18470 15096 18522
rect 15096 18470 15106 18522
rect 15130 18470 15160 18522
rect 15160 18470 15186 18522
rect 14890 18468 14946 18470
rect 14970 18468 15026 18470
rect 15050 18468 15106 18470
rect 15130 18468 15186 18470
rect 9890 17978 9946 17980
rect 9970 17978 10026 17980
rect 10050 17978 10106 17980
rect 10130 17978 10186 17980
rect 9890 17926 9916 17978
rect 9916 17926 9946 17978
rect 9970 17926 9980 17978
rect 9980 17926 10026 17978
rect 10050 17926 10096 17978
rect 10096 17926 10106 17978
rect 10130 17926 10160 17978
rect 10160 17926 10186 17978
rect 9890 17924 9946 17926
rect 9970 17924 10026 17926
rect 10050 17924 10106 17926
rect 10130 17924 10186 17926
rect 19890 17978 19946 17980
rect 19970 17978 20026 17980
rect 20050 17978 20106 17980
rect 20130 17978 20186 17980
rect 19890 17926 19916 17978
rect 19916 17926 19946 17978
rect 19970 17926 19980 17978
rect 19980 17926 20026 17978
rect 20050 17926 20096 17978
rect 20096 17926 20106 17978
rect 20130 17926 20160 17978
rect 20160 17926 20186 17978
rect 19890 17924 19946 17926
rect 19970 17924 20026 17926
rect 20050 17924 20106 17926
rect 20130 17924 20186 17926
rect 4890 17434 4946 17436
rect 4970 17434 5026 17436
rect 5050 17434 5106 17436
rect 5130 17434 5186 17436
rect 4890 17382 4916 17434
rect 4916 17382 4946 17434
rect 4970 17382 4980 17434
rect 4980 17382 5026 17434
rect 5050 17382 5096 17434
rect 5096 17382 5106 17434
rect 5130 17382 5160 17434
rect 5160 17382 5186 17434
rect 4890 17380 4946 17382
rect 4970 17380 5026 17382
rect 5050 17380 5106 17382
rect 5130 17380 5186 17382
rect 14890 17434 14946 17436
rect 14970 17434 15026 17436
rect 15050 17434 15106 17436
rect 15130 17434 15186 17436
rect 14890 17382 14916 17434
rect 14916 17382 14946 17434
rect 14970 17382 14980 17434
rect 14980 17382 15026 17434
rect 15050 17382 15096 17434
rect 15096 17382 15106 17434
rect 15130 17382 15160 17434
rect 15160 17382 15186 17434
rect 14890 17380 14946 17382
rect 14970 17380 15026 17382
rect 15050 17380 15106 17382
rect 15130 17380 15186 17382
rect 9890 16890 9946 16892
rect 9970 16890 10026 16892
rect 10050 16890 10106 16892
rect 10130 16890 10186 16892
rect 9890 16838 9916 16890
rect 9916 16838 9946 16890
rect 9970 16838 9980 16890
rect 9980 16838 10026 16890
rect 10050 16838 10096 16890
rect 10096 16838 10106 16890
rect 10130 16838 10160 16890
rect 10160 16838 10186 16890
rect 9890 16836 9946 16838
rect 9970 16836 10026 16838
rect 10050 16836 10106 16838
rect 10130 16836 10186 16838
rect 19890 16890 19946 16892
rect 19970 16890 20026 16892
rect 20050 16890 20106 16892
rect 20130 16890 20186 16892
rect 19890 16838 19916 16890
rect 19916 16838 19946 16890
rect 19970 16838 19980 16890
rect 19980 16838 20026 16890
rect 20050 16838 20096 16890
rect 20096 16838 20106 16890
rect 20130 16838 20160 16890
rect 20160 16838 20186 16890
rect 19890 16836 19946 16838
rect 19970 16836 20026 16838
rect 20050 16836 20106 16838
rect 20130 16836 20186 16838
rect 4890 16346 4946 16348
rect 4970 16346 5026 16348
rect 5050 16346 5106 16348
rect 5130 16346 5186 16348
rect 4890 16294 4916 16346
rect 4916 16294 4946 16346
rect 4970 16294 4980 16346
rect 4980 16294 5026 16346
rect 5050 16294 5096 16346
rect 5096 16294 5106 16346
rect 5130 16294 5160 16346
rect 5160 16294 5186 16346
rect 4890 16292 4946 16294
rect 4970 16292 5026 16294
rect 5050 16292 5106 16294
rect 5130 16292 5186 16294
rect 14890 16346 14946 16348
rect 14970 16346 15026 16348
rect 15050 16346 15106 16348
rect 15130 16346 15186 16348
rect 14890 16294 14916 16346
rect 14916 16294 14946 16346
rect 14970 16294 14980 16346
rect 14980 16294 15026 16346
rect 15050 16294 15096 16346
rect 15096 16294 15106 16346
rect 15130 16294 15160 16346
rect 15160 16294 15186 16346
rect 14890 16292 14946 16294
rect 14970 16292 15026 16294
rect 15050 16292 15106 16294
rect 15130 16292 15186 16294
rect 9890 15802 9946 15804
rect 9970 15802 10026 15804
rect 10050 15802 10106 15804
rect 10130 15802 10186 15804
rect 9890 15750 9916 15802
rect 9916 15750 9946 15802
rect 9970 15750 9980 15802
rect 9980 15750 10026 15802
rect 10050 15750 10096 15802
rect 10096 15750 10106 15802
rect 10130 15750 10160 15802
rect 10160 15750 10186 15802
rect 9890 15748 9946 15750
rect 9970 15748 10026 15750
rect 10050 15748 10106 15750
rect 10130 15748 10186 15750
rect 19890 15802 19946 15804
rect 19970 15802 20026 15804
rect 20050 15802 20106 15804
rect 20130 15802 20186 15804
rect 19890 15750 19916 15802
rect 19916 15750 19946 15802
rect 19970 15750 19980 15802
rect 19980 15750 20026 15802
rect 20050 15750 20096 15802
rect 20096 15750 20106 15802
rect 20130 15750 20160 15802
rect 20160 15750 20186 15802
rect 19890 15748 19946 15750
rect 19970 15748 20026 15750
rect 20050 15748 20106 15750
rect 20130 15748 20186 15750
rect 4890 15258 4946 15260
rect 4970 15258 5026 15260
rect 5050 15258 5106 15260
rect 5130 15258 5186 15260
rect 4890 15206 4916 15258
rect 4916 15206 4946 15258
rect 4970 15206 4980 15258
rect 4980 15206 5026 15258
rect 5050 15206 5096 15258
rect 5096 15206 5106 15258
rect 5130 15206 5160 15258
rect 5160 15206 5186 15258
rect 4890 15204 4946 15206
rect 4970 15204 5026 15206
rect 5050 15204 5106 15206
rect 5130 15204 5186 15206
rect 14890 15258 14946 15260
rect 14970 15258 15026 15260
rect 15050 15258 15106 15260
rect 15130 15258 15186 15260
rect 14890 15206 14916 15258
rect 14916 15206 14946 15258
rect 14970 15206 14980 15258
rect 14980 15206 15026 15258
rect 15050 15206 15096 15258
rect 15096 15206 15106 15258
rect 15130 15206 15160 15258
rect 15160 15206 15186 15258
rect 14890 15204 14946 15206
rect 14970 15204 15026 15206
rect 15050 15204 15106 15206
rect 15130 15204 15186 15206
rect 9890 14714 9946 14716
rect 9970 14714 10026 14716
rect 10050 14714 10106 14716
rect 10130 14714 10186 14716
rect 9890 14662 9916 14714
rect 9916 14662 9946 14714
rect 9970 14662 9980 14714
rect 9980 14662 10026 14714
rect 10050 14662 10096 14714
rect 10096 14662 10106 14714
rect 10130 14662 10160 14714
rect 10160 14662 10186 14714
rect 9890 14660 9946 14662
rect 9970 14660 10026 14662
rect 10050 14660 10106 14662
rect 10130 14660 10186 14662
rect 19890 14714 19946 14716
rect 19970 14714 20026 14716
rect 20050 14714 20106 14716
rect 20130 14714 20186 14716
rect 19890 14662 19916 14714
rect 19916 14662 19946 14714
rect 19970 14662 19980 14714
rect 19980 14662 20026 14714
rect 20050 14662 20096 14714
rect 20096 14662 20106 14714
rect 20130 14662 20160 14714
rect 20160 14662 20186 14714
rect 19890 14660 19946 14662
rect 19970 14660 20026 14662
rect 20050 14660 20106 14662
rect 20130 14660 20186 14662
rect 4890 14170 4946 14172
rect 4970 14170 5026 14172
rect 5050 14170 5106 14172
rect 5130 14170 5186 14172
rect 4890 14118 4916 14170
rect 4916 14118 4946 14170
rect 4970 14118 4980 14170
rect 4980 14118 5026 14170
rect 5050 14118 5096 14170
rect 5096 14118 5106 14170
rect 5130 14118 5160 14170
rect 5160 14118 5186 14170
rect 4890 14116 4946 14118
rect 4970 14116 5026 14118
rect 5050 14116 5106 14118
rect 5130 14116 5186 14118
rect 14890 14170 14946 14172
rect 14970 14170 15026 14172
rect 15050 14170 15106 14172
rect 15130 14170 15186 14172
rect 14890 14118 14916 14170
rect 14916 14118 14946 14170
rect 14970 14118 14980 14170
rect 14980 14118 15026 14170
rect 15050 14118 15096 14170
rect 15096 14118 15106 14170
rect 15130 14118 15160 14170
rect 15160 14118 15186 14170
rect 14890 14116 14946 14118
rect 14970 14116 15026 14118
rect 15050 14116 15106 14118
rect 15130 14116 15186 14118
rect 9890 13626 9946 13628
rect 9970 13626 10026 13628
rect 10050 13626 10106 13628
rect 10130 13626 10186 13628
rect 9890 13574 9916 13626
rect 9916 13574 9946 13626
rect 9970 13574 9980 13626
rect 9980 13574 10026 13626
rect 10050 13574 10096 13626
rect 10096 13574 10106 13626
rect 10130 13574 10160 13626
rect 10160 13574 10186 13626
rect 9890 13572 9946 13574
rect 9970 13572 10026 13574
rect 10050 13572 10106 13574
rect 10130 13572 10186 13574
rect 19890 13626 19946 13628
rect 19970 13626 20026 13628
rect 20050 13626 20106 13628
rect 20130 13626 20186 13628
rect 19890 13574 19916 13626
rect 19916 13574 19946 13626
rect 19970 13574 19980 13626
rect 19980 13574 20026 13626
rect 20050 13574 20096 13626
rect 20096 13574 20106 13626
rect 20130 13574 20160 13626
rect 20160 13574 20186 13626
rect 19890 13572 19946 13574
rect 19970 13572 20026 13574
rect 20050 13572 20106 13574
rect 20130 13572 20186 13574
rect 4890 13082 4946 13084
rect 4970 13082 5026 13084
rect 5050 13082 5106 13084
rect 5130 13082 5186 13084
rect 4890 13030 4916 13082
rect 4916 13030 4946 13082
rect 4970 13030 4980 13082
rect 4980 13030 5026 13082
rect 5050 13030 5096 13082
rect 5096 13030 5106 13082
rect 5130 13030 5160 13082
rect 5160 13030 5186 13082
rect 4890 13028 4946 13030
rect 4970 13028 5026 13030
rect 5050 13028 5106 13030
rect 5130 13028 5186 13030
rect 14890 13082 14946 13084
rect 14970 13082 15026 13084
rect 15050 13082 15106 13084
rect 15130 13082 15186 13084
rect 14890 13030 14916 13082
rect 14916 13030 14946 13082
rect 14970 13030 14980 13082
rect 14980 13030 15026 13082
rect 15050 13030 15096 13082
rect 15096 13030 15106 13082
rect 15130 13030 15160 13082
rect 15160 13030 15186 13082
rect 14890 13028 14946 13030
rect 14970 13028 15026 13030
rect 15050 13028 15106 13030
rect 15130 13028 15186 13030
rect 9890 12538 9946 12540
rect 9970 12538 10026 12540
rect 10050 12538 10106 12540
rect 10130 12538 10186 12540
rect 9890 12486 9916 12538
rect 9916 12486 9946 12538
rect 9970 12486 9980 12538
rect 9980 12486 10026 12538
rect 10050 12486 10096 12538
rect 10096 12486 10106 12538
rect 10130 12486 10160 12538
rect 10160 12486 10186 12538
rect 9890 12484 9946 12486
rect 9970 12484 10026 12486
rect 10050 12484 10106 12486
rect 10130 12484 10186 12486
rect 19890 12538 19946 12540
rect 19970 12538 20026 12540
rect 20050 12538 20106 12540
rect 20130 12538 20186 12540
rect 19890 12486 19916 12538
rect 19916 12486 19946 12538
rect 19970 12486 19980 12538
rect 19980 12486 20026 12538
rect 20050 12486 20096 12538
rect 20096 12486 20106 12538
rect 20130 12486 20160 12538
rect 20160 12486 20186 12538
rect 19890 12484 19946 12486
rect 19970 12484 20026 12486
rect 20050 12484 20106 12486
rect 20130 12484 20186 12486
rect 4890 11994 4946 11996
rect 4970 11994 5026 11996
rect 5050 11994 5106 11996
rect 5130 11994 5186 11996
rect 4890 11942 4916 11994
rect 4916 11942 4946 11994
rect 4970 11942 4980 11994
rect 4980 11942 5026 11994
rect 5050 11942 5096 11994
rect 5096 11942 5106 11994
rect 5130 11942 5160 11994
rect 5160 11942 5186 11994
rect 4890 11940 4946 11942
rect 4970 11940 5026 11942
rect 5050 11940 5106 11942
rect 5130 11940 5186 11942
rect 14890 11994 14946 11996
rect 14970 11994 15026 11996
rect 15050 11994 15106 11996
rect 15130 11994 15186 11996
rect 14890 11942 14916 11994
rect 14916 11942 14946 11994
rect 14970 11942 14980 11994
rect 14980 11942 15026 11994
rect 15050 11942 15096 11994
rect 15096 11942 15106 11994
rect 15130 11942 15160 11994
rect 15160 11942 15186 11994
rect 14890 11940 14946 11942
rect 14970 11940 15026 11942
rect 15050 11940 15106 11942
rect 15130 11940 15186 11942
rect 9890 11450 9946 11452
rect 9970 11450 10026 11452
rect 10050 11450 10106 11452
rect 10130 11450 10186 11452
rect 9890 11398 9916 11450
rect 9916 11398 9946 11450
rect 9970 11398 9980 11450
rect 9980 11398 10026 11450
rect 10050 11398 10096 11450
rect 10096 11398 10106 11450
rect 10130 11398 10160 11450
rect 10160 11398 10186 11450
rect 9890 11396 9946 11398
rect 9970 11396 10026 11398
rect 10050 11396 10106 11398
rect 10130 11396 10186 11398
rect 19890 11450 19946 11452
rect 19970 11450 20026 11452
rect 20050 11450 20106 11452
rect 20130 11450 20186 11452
rect 19890 11398 19916 11450
rect 19916 11398 19946 11450
rect 19970 11398 19980 11450
rect 19980 11398 20026 11450
rect 20050 11398 20096 11450
rect 20096 11398 20106 11450
rect 20130 11398 20160 11450
rect 20160 11398 20186 11450
rect 19890 11396 19946 11398
rect 19970 11396 20026 11398
rect 20050 11396 20106 11398
rect 20130 11396 20186 11398
rect 4890 10906 4946 10908
rect 4970 10906 5026 10908
rect 5050 10906 5106 10908
rect 5130 10906 5186 10908
rect 4890 10854 4916 10906
rect 4916 10854 4946 10906
rect 4970 10854 4980 10906
rect 4980 10854 5026 10906
rect 5050 10854 5096 10906
rect 5096 10854 5106 10906
rect 5130 10854 5160 10906
rect 5160 10854 5186 10906
rect 4890 10852 4946 10854
rect 4970 10852 5026 10854
rect 5050 10852 5106 10854
rect 5130 10852 5186 10854
rect 14890 10906 14946 10908
rect 14970 10906 15026 10908
rect 15050 10906 15106 10908
rect 15130 10906 15186 10908
rect 14890 10854 14916 10906
rect 14916 10854 14946 10906
rect 14970 10854 14980 10906
rect 14980 10854 15026 10906
rect 15050 10854 15096 10906
rect 15096 10854 15106 10906
rect 15130 10854 15160 10906
rect 15160 10854 15186 10906
rect 14890 10852 14946 10854
rect 14970 10852 15026 10854
rect 15050 10852 15106 10854
rect 15130 10852 15186 10854
rect 3000 10512 3056 10568
rect 10176 10512 10232 10568
rect 9890 10362 9946 10364
rect 9970 10362 10026 10364
rect 10050 10362 10106 10364
rect 10130 10362 10186 10364
rect 9890 10310 9916 10362
rect 9916 10310 9946 10362
rect 9970 10310 9980 10362
rect 9980 10310 10026 10362
rect 10050 10310 10096 10362
rect 10096 10310 10106 10362
rect 10130 10310 10160 10362
rect 10160 10310 10186 10362
rect 9890 10308 9946 10310
rect 9970 10308 10026 10310
rect 10050 10308 10106 10310
rect 10130 10308 10186 10310
rect 4890 9818 4946 9820
rect 4970 9818 5026 9820
rect 5050 9818 5106 9820
rect 5130 9818 5186 9820
rect 4890 9766 4916 9818
rect 4916 9766 4946 9818
rect 4970 9766 4980 9818
rect 4980 9766 5026 9818
rect 5050 9766 5096 9818
rect 5096 9766 5106 9818
rect 5130 9766 5160 9818
rect 5160 9766 5186 9818
rect 4890 9764 4946 9766
rect 4970 9764 5026 9766
rect 5050 9764 5106 9766
rect 5130 9764 5186 9766
rect 9890 9274 9946 9276
rect 9970 9274 10026 9276
rect 10050 9274 10106 9276
rect 10130 9274 10186 9276
rect 9890 9222 9916 9274
rect 9916 9222 9946 9274
rect 9970 9222 9980 9274
rect 9980 9222 10026 9274
rect 10050 9222 10096 9274
rect 10096 9222 10106 9274
rect 10130 9222 10160 9274
rect 10160 9222 10186 9274
rect 9890 9220 9946 9222
rect 9970 9220 10026 9222
rect 10050 9220 10106 9222
rect 10130 9220 10186 9222
rect 4890 8730 4946 8732
rect 4970 8730 5026 8732
rect 5050 8730 5106 8732
rect 5130 8730 5186 8732
rect 4890 8678 4916 8730
rect 4916 8678 4946 8730
rect 4970 8678 4980 8730
rect 4980 8678 5026 8730
rect 5050 8678 5096 8730
rect 5096 8678 5106 8730
rect 5130 8678 5160 8730
rect 5160 8678 5186 8730
rect 4890 8676 4946 8678
rect 4970 8676 5026 8678
rect 5050 8676 5106 8678
rect 5130 8676 5186 8678
rect 9890 8186 9946 8188
rect 9970 8186 10026 8188
rect 10050 8186 10106 8188
rect 10130 8186 10186 8188
rect 9890 8134 9916 8186
rect 9916 8134 9946 8186
rect 9970 8134 9980 8186
rect 9980 8134 10026 8186
rect 10050 8134 10096 8186
rect 10096 8134 10106 8186
rect 10130 8134 10160 8186
rect 10160 8134 10186 8186
rect 9890 8132 9946 8134
rect 9970 8132 10026 8134
rect 10050 8132 10106 8134
rect 10130 8132 10186 8134
rect 4890 7642 4946 7644
rect 4970 7642 5026 7644
rect 5050 7642 5106 7644
rect 5130 7642 5186 7644
rect 4890 7590 4916 7642
rect 4916 7590 4946 7642
rect 4970 7590 4980 7642
rect 4980 7590 5026 7642
rect 5050 7590 5096 7642
rect 5096 7590 5106 7642
rect 5130 7590 5160 7642
rect 5160 7590 5186 7642
rect 4890 7588 4946 7590
rect 4970 7588 5026 7590
rect 5050 7588 5106 7590
rect 5130 7588 5186 7590
rect 9890 7098 9946 7100
rect 9970 7098 10026 7100
rect 10050 7098 10106 7100
rect 10130 7098 10186 7100
rect 9890 7046 9916 7098
rect 9916 7046 9946 7098
rect 9970 7046 9980 7098
rect 9980 7046 10026 7098
rect 10050 7046 10096 7098
rect 10096 7046 10106 7098
rect 10130 7046 10160 7098
rect 10160 7046 10186 7098
rect 9890 7044 9946 7046
rect 9970 7044 10026 7046
rect 10050 7044 10106 7046
rect 10130 7044 10186 7046
rect 4890 6554 4946 6556
rect 4970 6554 5026 6556
rect 5050 6554 5106 6556
rect 5130 6554 5186 6556
rect 4890 6502 4916 6554
rect 4916 6502 4946 6554
rect 4970 6502 4980 6554
rect 4980 6502 5026 6554
rect 5050 6502 5096 6554
rect 5096 6502 5106 6554
rect 5130 6502 5160 6554
rect 5160 6502 5186 6554
rect 4890 6500 4946 6502
rect 4970 6500 5026 6502
rect 5050 6500 5106 6502
rect 5130 6500 5186 6502
rect 9890 6010 9946 6012
rect 9970 6010 10026 6012
rect 10050 6010 10106 6012
rect 10130 6010 10186 6012
rect 9890 5958 9916 6010
rect 9916 5958 9946 6010
rect 9970 5958 9980 6010
rect 9980 5958 10026 6010
rect 10050 5958 10096 6010
rect 10096 5958 10106 6010
rect 10130 5958 10160 6010
rect 10160 5958 10186 6010
rect 9890 5956 9946 5958
rect 9970 5956 10026 5958
rect 10050 5956 10106 5958
rect 10130 5956 10186 5958
rect 19890 10362 19946 10364
rect 19970 10362 20026 10364
rect 20050 10362 20106 10364
rect 20130 10362 20186 10364
rect 19890 10310 19916 10362
rect 19916 10310 19946 10362
rect 19970 10310 19980 10362
rect 19980 10310 20026 10362
rect 20050 10310 20096 10362
rect 20096 10310 20106 10362
rect 20130 10310 20160 10362
rect 20160 10310 20186 10362
rect 19890 10308 19946 10310
rect 19970 10308 20026 10310
rect 20050 10308 20106 10310
rect 20130 10308 20186 10310
rect 14890 9818 14946 9820
rect 14970 9818 15026 9820
rect 15050 9818 15106 9820
rect 15130 9818 15186 9820
rect 14890 9766 14916 9818
rect 14916 9766 14946 9818
rect 14970 9766 14980 9818
rect 14980 9766 15026 9818
rect 15050 9766 15096 9818
rect 15096 9766 15106 9818
rect 15130 9766 15160 9818
rect 15160 9766 15186 9818
rect 14890 9764 14946 9766
rect 14970 9764 15026 9766
rect 15050 9764 15106 9766
rect 15130 9764 15186 9766
rect 19890 9274 19946 9276
rect 19970 9274 20026 9276
rect 20050 9274 20106 9276
rect 20130 9274 20186 9276
rect 19890 9222 19916 9274
rect 19916 9222 19946 9274
rect 19970 9222 19980 9274
rect 19980 9222 20026 9274
rect 20050 9222 20096 9274
rect 20096 9222 20106 9274
rect 20130 9222 20160 9274
rect 20160 9222 20186 9274
rect 19890 9220 19946 9222
rect 19970 9220 20026 9222
rect 20050 9220 20106 9222
rect 20130 9220 20186 9222
rect 14890 8730 14946 8732
rect 14970 8730 15026 8732
rect 15050 8730 15106 8732
rect 15130 8730 15186 8732
rect 14890 8678 14916 8730
rect 14916 8678 14946 8730
rect 14970 8678 14980 8730
rect 14980 8678 15026 8730
rect 15050 8678 15096 8730
rect 15096 8678 15106 8730
rect 15130 8678 15160 8730
rect 15160 8678 15186 8730
rect 14890 8676 14946 8678
rect 14970 8676 15026 8678
rect 15050 8676 15106 8678
rect 15130 8676 15186 8678
rect 19890 8186 19946 8188
rect 19970 8186 20026 8188
rect 20050 8186 20106 8188
rect 20130 8186 20186 8188
rect 19890 8134 19916 8186
rect 19916 8134 19946 8186
rect 19970 8134 19980 8186
rect 19980 8134 20026 8186
rect 20050 8134 20096 8186
rect 20096 8134 20106 8186
rect 20130 8134 20160 8186
rect 20160 8134 20186 8186
rect 19890 8132 19946 8134
rect 19970 8132 20026 8134
rect 20050 8132 20106 8134
rect 20130 8132 20186 8134
rect 14890 7642 14946 7644
rect 14970 7642 15026 7644
rect 15050 7642 15106 7644
rect 15130 7642 15186 7644
rect 14890 7590 14916 7642
rect 14916 7590 14946 7642
rect 14970 7590 14980 7642
rect 14980 7590 15026 7642
rect 15050 7590 15096 7642
rect 15096 7590 15106 7642
rect 15130 7590 15160 7642
rect 15160 7590 15186 7642
rect 14890 7588 14946 7590
rect 14970 7588 15026 7590
rect 15050 7588 15106 7590
rect 15130 7588 15186 7590
rect 19890 7098 19946 7100
rect 19970 7098 20026 7100
rect 20050 7098 20106 7100
rect 20130 7098 20186 7100
rect 19890 7046 19916 7098
rect 19916 7046 19946 7098
rect 19970 7046 19980 7098
rect 19980 7046 20026 7098
rect 20050 7046 20096 7098
rect 20096 7046 20106 7098
rect 20130 7046 20160 7098
rect 20160 7046 20186 7098
rect 19890 7044 19946 7046
rect 19970 7044 20026 7046
rect 20050 7044 20106 7046
rect 20130 7044 20186 7046
rect 14890 6554 14946 6556
rect 14970 6554 15026 6556
rect 15050 6554 15106 6556
rect 15130 6554 15186 6556
rect 14890 6502 14916 6554
rect 14916 6502 14946 6554
rect 14970 6502 14980 6554
rect 14980 6502 15026 6554
rect 15050 6502 15096 6554
rect 15096 6502 15106 6554
rect 15130 6502 15160 6554
rect 15160 6502 15186 6554
rect 14890 6500 14946 6502
rect 14970 6500 15026 6502
rect 15050 6500 15106 6502
rect 15130 6500 15186 6502
rect 19890 6010 19946 6012
rect 19970 6010 20026 6012
rect 20050 6010 20106 6012
rect 20130 6010 20186 6012
rect 19890 5958 19916 6010
rect 19916 5958 19946 6010
rect 19970 5958 19980 6010
rect 19980 5958 20026 6010
rect 20050 5958 20096 6010
rect 20096 5958 20106 6010
rect 20130 5958 20160 6010
rect 20160 5958 20186 6010
rect 19890 5956 19946 5958
rect 19970 5956 20026 5958
rect 20050 5956 20106 5958
rect 20130 5956 20186 5958
rect 10544 5616 10600 5672
rect 13856 5616 13912 5672
rect 4890 5466 4946 5468
rect 4970 5466 5026 5468
rect 5050 5466 5106 5468
rect 5130 5466 5186 5468
rect 4890 5414 4916 5466
rect 4916 5414 4946 5466
rect 4970 5414 4980 5466
rect 4980 5414 5026 5466
rect 5050 5414 5096 5466
rect 5096 5414 5106 5466
rect 5130 5414 5160 5466
rect 5160 5414 5186 5466
rect 4890 5412 4946 5414
rect 4970 5412 5026 5414
rect 5050 5412 5106 5414
rect 5130 5412 5186 5414
rect 9890 4922 9946 4924
rect 9970 4922 10026 4924
rect 10050 4922 10106 4924
rect 10130 4922 10186 4924
rect 9890 4870 9916 4922
rect 9916 4870 9946 4922
rect 9970 4870 9980 4922
rect 9980 4870 10026 4922
rect 10050 4870 10096 4922
rect 10096 4870 10106 4922
rect 10130 4870 10160 4922
rect 10160 4870 10186 4922
rect 9890 4868 9946 4870
rect 9970 4868 10026 4870
rect 10050 4868 10106 4870
rect 10130 4868 10186 4870
rect 4890 4378 4946 4380
rect 4970 4378 5026 4380
rect 5050 4378 5106 4380
rect 5130 4378 5186 4380
rect 4890 4326 4916 4378
rect 4916 4326 4946 4378
rect 4970 4326 4980 4378
rect 4980 4326 5026 4378
rect 5050 4326 5096 4378
rect 5096 4326 5106 4378
rect 5130 4326 5160 4378
rect 5160 4326 5186 4378
rect 4890 4324 4946 4326
rect 4970 4324 5026 4326
rect 5050 4324 5106 4326
rect 5130 4324 5186 4326
rect 9890 3834 9946 3836
rect 9970 3834 10026 3836
rect 10050 3834 10106 3836
rect 10130 3834 10186 3836
rect 9890 3782 9916 3834
rect 9916 3782 9946 3834
rect 9970 3782 9980 3834
rect 9980 3782 10026 3834
rect 10050 3782 10096 3834
rect 10096 3782 10106 3834
rect 10130 3782 10160 3834
rect 10160 3782 10186 3834
rect 9890 3780 9946 3782
rect 9970 3780 10026 3782
rect 10050 3780 10106 3782
rect 10130 3780 10186 3782
rect 4890 3290 4946 3292
rect 4970 3290 5026 3292
rect 5050 3290 5106 3292
rect 5130 3290 5186 3292
rect 4890 3238 4916 3290
rect 4916 3238 4946 3290
rect 4970 3238 4980 3290
rect 4980 3238 5026 3290
rect 5050 3238 5096 3290
rect 5096 3238 5106 3290
rect 5130 3238 5160 3290
rect 5160 3238 5186 3290
rect 4890 3236 4946 3238
rect 4970 3236 5026 3238
rect 5050 3236 5106 3238
rect 5130 3236 5186 3238
rect 3920 2896 3976 2952
rect 9890 2746 9946 2748
rect 9970 2746 10026 2748
rect 10050 2746 10106 2748
rect 10130 2746 10186 2748
rect 9890 2694 9916 2746
rect 9916 2694 9946 2746
rect 9970 2694 9980 2746
rect 9980 2694 10026 2746
rect 10050 2694 10096 2746
rect 10096 2694 10106 2746
rect 10130 2694 10160 2746
rect 10160 2694 10186 2746
rect 9890 2692 9946 2694
rect 9970 2692 10026 2694
rect 10050 2692 10106 2694
rect 10130 2692 10186 2694
rect 4890 2202 4946 2204
rect 4970 2202 5026 2204
rect 5050 2202 5106 2204
rect 5130 2202 5186 2204
rect 4890 2150 4916 2202
rect 4916 2150 4946 2202
rect 4970 2150 4980 2202
rect 4980 2150 5026 2202
rect 5050 2150 5096 2202
rect 5096 2150 5106 2202
rect 5130 2150 5160 2202
rect 5160 2150 5186 2202
rect 4890 2148 4946 2150
rect 4970 2148 5026 2150
rect 5050 2148 5106 2150
rect 5130 2148 5186 2150
rect 14890 5466 14946 5468
rect 14970 5466 15026 5468
rect 15050 5466 15106 5468
rect 15130 5466 15186 5468
rect 14890 5414 14916 5466
rect 14916 5414 14946 5466
rect 14970 5414 14980 5466
rect 14980 5414 15026 5466
rect 15050 5414 15096 5466
rect 15096 5414 15106 5466
rect 15130 5414 15160 5466
rect 15160 5414 15186 5466
rect 14890 5412 14946 5414
rect 14970 5412 15026 5414
rect 15050 5412 15106 5414
rect 15130 5412 15186 5414
rect 19890 4922 19946 4924
rect 19970 4922 20026 4924
rect 20050 4922 20106 4924
rect 20130 4922 20186 4924
rect 19890 4870 19916 4922
rect 19916 4870 19946 4922
rect 19970 4870 19980 4922
rect 19980 4870 20026 4922
rect 20050 4870 20096 4922
rect 20096 4870 20106 4922
rect 20130 4870 20160 4922
rect 20160 4870 20186 4922
rect 19890 4868 19946 4870
rect 19970 4868 20026 4870
rect 20050 4868 20106 4870
rect 20130 4868 20186 4870
rect 14890 4378 14946 4380
rect 14970 4378 15026 4380
rect 15050 4378 15106 4380
rect 15130 4378 15186 4380
rect 14890 4326 14916 4378
rect 14916 4326 14946 4378
rect 14970 4326 14980 4378
rect 14980 4326 15026 4378
rect 15050 4326 15096 4378
rect 15096 4326 15106 4378
rect 15130 4326 15160 4378
rect 15160 4326 15186 4378
rect 14890 4324 14946 4326
rect 14970 4324 15026 4326
rect 15050 4324 15106 4326
rect 15130 4324 15186 4326
rect 22872 3984 22928 4040
rect 19890 3834 19946 3836
rect 19970 3834 20026 3836
rect 20050 3834 20106 3836
rect 20130 3834 20186 3836
rect 19890 3782 19916 3834
rect 19916 3782 19946 3834
rect 19970 3782 19980 3834
rect 19980 3782 20026 3834
rect 20050 3782 20096 3834
rect 20096 3782 20106 3834
rect 20130 3782 20160 3834
rect 20160 3782 20186 3834
rect 19890 3780 19946 3782
rect 19970 3780 20026 3782
rect 20050 3780 20106 3782
rect 20130 3780 20186 3782
rect 14890 3290 14946 3292
rect 14970 3290 15026 3292
rect 15050 3290 15106 3292
rect 15130 3290 15186 3292
rect 14890 3238 14916 3290
rect 14916 3238 14946 3290
rect 14970 3238 14980 3290
rect 14980 3238 15026 3290
rect 15050 3238 15096 3290
rect 15096 3238 15106 3290
rect 15130 3238 15160 3290
rect 15160 3238 15186 3290
rect 14890 3236 14946 3238
rect 14970 3236 15026 3238
rect 15050 3236 15106 3238
rect 15130 3236 15186 3238
rect 20480 2896 20536 2952
rect 19890 2746 19946 2748
rect 19970 2746 20026 2748
rect 20050 2746 20106 2748
rect 20130 2746 20186 2748
rect 19890 2694 19916 2746
rect 19916 2694 19946 2746
rect 19970 2694 19980 2746
rect 19980 2694 20026 2746
rect 20050 2694 20096 2746
rect 20096 2694 20106 2746
rect 20130 2694 20160 2746
rect 20160 2694 20186 2746
rect 19890 2692 19946 2694
rect 19970 2692 20026 2694
rect 20050 2692 20106 2694
rect 20130 2692 20186 2694
rect 24890 21786 24946 21788
rect 24970 21786 25026 21788
rect 25050 21786 25106 21788
rect 25130 21786 25186 21788
rect 24890 21734 24916 21786
rect 24916 21734 24946 21786
rect 24970 21734 24980 21786
rect 24980 21734 25026 21786
rect 25050 21734 25096 21786
rect 25096 21734 25106 21786
rect 25130 21734 25160 21786
rect 25160 21734 25186 21786
rect 24890 21732 24946 21734
rect 24970 21732 25026 21734
rect 25050 21732 25106 21734
rect 25130 21732 25186 21734
rect 24890 20698 24946 20700
rect 24970 20698 25026 20700
rect 25050 20698 25106 20700
rect 25130 20698 25186 20700
rect 24890 20646 24916 20698
rect 24916 20646 24946 20698
rect 24970 20646 24980 20698
rect 24980 20646 25026 20698
rect 25050 20646 25096 20698
rect 25096 20646 25106 20698
rect 25130 20646 25160 20698
rect 25160 20646 25186 20698
rect 24890 20644 24946 20646
rect 24970 20644 25026 20646
rect 25050 20644 25106 20646
rect 25130 20644 25186 20646
rect 24436 19896 24492 19952
rect 24890 19610 24946 19612
rect 24970 19610 25026 19612
rect 25050 19610 25106 19612
rect 25130 19610 25186 19612
rect 24890 19558 24916 19610
rect 24916 19558 24946 19610
rect 24970 19558 24980 19610
rect 24980 19558 25026 19610
rect 25050 19558 25096 19610
rect 25096 19558 25106 19610
rect 25130 19558 25160 19610
rect 25160 19558 25186 19610
rect 24890 19556 24946 19558
rect 24970 19556 25026 19558
rect 25050 19556 25106 19558
rect 25130 19556 25186 19558
rect 24436 18808 24492 18864
rect 23884 11736 23940 11792
rect 24890 18522 24946 18524
rect 24970 18522 25026 18524
rect 25050 18522 25106 18524
rect 25130 18522 25186 18524
rect 24890 18470 24916 18522
rect 24916 18470 24946 18522
rect 24970 18470 24980 18522
rect 24980 18470 25026 18522
rect 25050 18470 25096 18522
rect 25096 18470 25106 18522
rect 25130 18470 25160 18522
rect 25160 18470 25186 18522
rect 24890 18468 24946 18470
rect 24970 18468 25026 18470
rect 25050 18468 25106 18470
rect 25130 18468 25186 18470
rect 24890 17434 24946 17436
rect 24970 17434 25026 17436
rect 25050 17434 25106 17436
rect 25130 17434 25186 17436
rect 24890 17382 24916 17434
rect 24916 17382 24946 17434
rect 24970 17382 24980 17434
rect 24980 17382 25026 17434
rect 25050 17382 25096 17434
rect 25096 17382 25106 17434
rect 25130 17382 25160 17434
rect 25160 17382 25186 17434
rect 24890 17380 24946 17382
rect 24970 17380 25026 17382
rect 25050 17380 25106 17382
rect 25130 17380 25186 17382
rect 24890 16346 24946 16348
rect 24970 16346 25026 16348
rect 25050 16346 25106 16348
rect 25130 16346 25186 16348
rect 24890 16294 24916 16346
rect 24916 16294 24946 16346
rect 24970 16294 24980 16346
rect 24980 16294 25026 16346
rect 25050 16294 25096 16346
rect 25096 16294 25106 16346
rect 25130 16294 25160 16346
rect 25160 16294 25186 16346
rect 24890 16292 24946 16294
rect 24970 16292 25026 16294
rect 25050 16292 25106 16294
rect 25130 16292 25186 16294
rect 24890 15258 24946 15260
rect 24970 15258 25026 15260
rect 25050 15258 25106 15260
rect 25130 15258 25186 15260
rect 24890 15206 24916 15258
rect 24916 15206 24946 15258
rect 24970 15206 24980 15258
rect 24980 15206 25026 15258
rect 25050 15206 25096 15258
rect 25096 15206 25106 15258
rect 25130 15206 25160 15258
rect 25160 15206 25186 15258
rect 24890 15204 24946 15206
rect 24970 15204 25026 15206
rect 25050 15204 25106 15206
rect 25130 15204 25186 15206
rect 24890 14170 24946 14172
rect 24970 14170 25026 14172
rect 25050 14170 25106 14172
rect 25130 14170 25186 14172
rect 24890 14118 24916 14170
rect 24916 14118 24946 14170
rect 24970 14118 24980 14170
rect 24980 14118 25026 14170
rect 25050 14118 25096 14170
rect 25096 14118 25106 14170
rect 25130 14118 25160 14170
rect 25160 14118 25186 14170
rect 24890 14116 24946 14118
rect 24970 14116 25026 14118
rect 25050 14116 25106 14118
rect 25130 14116 25186 14118
rect 24890 13082 24946 13084
rect 24970 13082 25026 13084
rect 25050 13082 25106 13084
rect 25130 13082 25186 13084
rect 24890 13030 24916 13082
rect 24916 13030 24946 13082
rect 24970 13030 24980 13082
rect 24980 13030 25026 13082
rect 25050 13030 25096 13082
rect 25096 13030 25106 13082
rect 25130 13030 25160 13082
rect 25160 13030 25186 13082
rect 24890 13028 24946 13030
rect 24970 13028 25026 13030
rect 25050 13028 25106 13030
rect 25130 13028 25186 13030
rect 24890 11994 24946 11996
rect 24970 11994 25026 11996
rect 25050 11994 25106 11996
rect 25130 11994 25186 11996
rect 24890 11942 24916 11994
rect 24916 11942 24946 11994
rect 24970 11942 24980 11994
rect 24980 11942 25026 11994
rect 25050 11942 25096 11994
rect 25096 11942 25106 11994
rect 25130 11942 25160 11994
rect 25160 11942 25186 11994
rect 24890 11940 24946 11942
rect 24970 11940 25026 11942
rect 25050 11940 25106 11942
rect 25130 11940 25186 11942
rect 24890 10906 24946 10908
rect 24970 10906 25026 10908
rect 25050 10906 25106 10908
rect 25130 10906 25186 10908
rect 24890 10854 24916 10906
rect 24916 10854 24946 10906
rect 24970 10854 24980 10906
rect 24980 10854 25026 10906
rect 25050 10854 25096 10906
rect 25096 10854 25106 10906
rect 25130 10854 25160 10906
rect 25160 10854 25186 10906
rect 24890 10852 24946 10854
rect 24970 10852 25026 10854
rect 25050 10852 25106 10854
rect 25130 10852 25186 10854
rect 24890 9818 24946 9820
rect 24970 9818 25026 9820
rect 25050 9818 25106 9820
rect 25130 9818 25186 9820
rect 24890 9766 24916 9818
rect 24916 9766 24946 9818
rect 24970 9766 24980 9818
rect 24980 9766 25026 9818
rect 25050 9766 25096 9818
rect 25096 9766 25106 9818
rect 25130 9766 25160 9818
rect 25160 9766 25186 9818
rect 24890 9764 24946 9766
rect 24970 9764 25026 9766
rect 25050 9764 25106 9766
rect 25130 9764 25186 9766
rect 24890 8730 24946 8732
rect 24970 8730 25026 8732
rect 25050 8730 25106 8732
rect 25130 8730 25186 8732
rect 24890 8678 24916 8730
rect 24916 8678 24946 8730
rect 24970 8678 24980 8730
rect 24980 8678 25026 8730
rect 25050 8678 25096 8730
rect 25096 8678 25106 8730
rect 25130 8678 25160 8730
rect 25160 8678 25186 8730
rect 24890 8676 24946 8678
rect 24970 8676 25026 8678
rect 25050 8676 25106 8678
rect 25130 8676 25186 8678
rect 24890 7642 24946 7644
rect 24970 7642 25026 7644
rect 25050 7642 25106 7644
rect 25130 7642 25186 7644
rect 24890 7590 24916 7642
rect 24916 7590 24946 7642
rect 24970 7590 24980 7642
rect 24980 7590 25026 7642
rect 25050 7590 25096 7642
rect 25096 7590 25106 7642
rect 25130 7590 25160 7642
rect 25160 7590 25186 7642
rect 24890 7588 24946 7590
rect 24970 7588 25026 7590
rect 25050 7588 25106 7590
rect 25130 7588 25186 7590
rect 24890 6554 24946 6556
rect 24970 6554 25026 6556
rect 25050 6554 25106 6556
rect 25130 6554 25186 6556
rect 24890 6502 24916 6554
rect 24916 6502 24946 6554
rect 24970 6502 24980 6554
rect 24980 6502 25026 6554
rect 25050 6502 25096 6554
rect 25096 6502 25106 6554
rect 25130 6502 25160 6554
rect 25160 6502 25186 6554
rect 24890 6500 24946 6502
rect 24970 6500 25026 6502
rect 25050 6500 25106 6502
rect 25130 6500 25186 6502
rect 24890 5466 24946 5468
rect 24970 5466 25026 5468
rect 25050 5466 25106 5468
rect 25130 5466 25186 5468
rect 24890 5414 24916 5466
rect 24916 5414 24946 5466
rect 24970 5414 24980 5466
rect 24980 5414 25026 5466
rect 25050 5414 25096 5466
rect 25096 5414 25106 5466
rect 25130 5414 25160 5466
rect 25160 5414 25186 5466
rect 24890 5412 24946 5414
rect 24970 5412 25026 5414
rect 25050 5412 25106 5414
rect 25130 5412 25186 5414
rect 24890 4378 24946 4380
rect 24970 4378 25026 4380
rect 25050 4378 25106 4380
rect 25130 4378 25186 4380
rect 24890 4326 24916 4378
rect 24916 4326 24946 4378
rect 24970 4326 24980 4378
rect 24980 4326 25026 4378
rect 25050 4326 25096 4378
rect 25096 4326 25106 4378
rect 25130 4326 25160 4378
rect 25160 4326 25186 4378
rect 24890 4324 24946 4326
rect 24970 4324 25026 4326
rect 25050 4324 25106 4326
rect 25130 4324 25186 4326
rect 24890 3290 24946 3292
rect 24970 3290 25026 3292
rect 25050 3290 25106 3292
rect 25130 3290 25186 3292
rect 24890 3238 24916 3290
rect 24916 3238 24946 3290
rect 24970 3238 24980 3290
rect 24980 3238 25026 3290
rect 25050 3238 25096 3290
rect 25096 3238 25106 3290
rect 25130 3238 25160 3290
rect 25160 3238 25186 3290
rect 24890 3236 24946 3238
rect 24970 3236 25026 3238
rect 25050 3236 25106 3238
rect 25130 3236 25186 3238
rect 22044 2644 22100 2680
rect 22044 2624 22046 2644
rect 22046 2624 22098 2644
rect 22098 2624 22100 2644
rect 23792 2624 23848 2680
rect 14890 2202 14946 2204
rect 14970 2202 15026 2204
rect 15050 2202 15106 2204
rect 15130 2202 15186 2204
rect 14890 2150 14916 2202
rect 14916 2150 14946 2202
rect 14970 2150 14980 2202
rect 14980 2150 15026 2202
rect 15050 2150 15096 2202
rect 15096 2150 15106 2202
rect 15130 2150 15160 2202
rect 15160 2150 15186 2202
rect 14890 2148 14946 2150
rect 14970 2148 15026 2150
rect 15050 2148 15106 2150
rect 15130 2148 15186 2150
rect 24890 2202 24946 2204
rect 24970 2202 25026 2204
rect 25050 2202 25106 2204
rect 25130 2202 25186 2204
rect 24890 2150 24916 2202
rect 24916 2150 24946 2202
rect 24970 2150 24980 2202
rect 24980 2150 25026 2202
rect 25050 2150 25096 2202
rect 25096 2150 25106 2202
rect 25130 2150 25160 2202
rect 25160 2150 25186 2202
rect 24890 2148 24946 2150
rect 24970 2148 25026 2150
rect 25050 2148 25106 2150
rect 25130 2148 25186 2150
<< metal3 >>
rect 4878 21792 5198 21793
rect 4878 21728 4886 21792
rect 4950 21728 4966 21792
rect 5030 21728 5046 21792
rect 5110 21728 5126 21792
rect 5190 21728 5198 21792
rect 4878 21727 5198 21728
rect 14878 21792 15198 21793
rect 14878 21728 14886 21792
rect 14950 21728 14966 21792
rect 15030 21728 15046 21792
rect 15110 21728 15126 21792
rect 15190 21728 15198 21792
rect 14878 21727 15198 21728
rect 24878 21792 25198 21793
rect 24878 21728 24886 21792
rect 24950 21728 24966 21792
rect 25030 21728 25046 21792
rect 25110 21728 25126 21792
rect 25190 21728 25198 21792
rect 24878 21727 25198 21728
rect 9878 21248 10198 21249
rect 9878 21184 9886 21248
rect 9950 21184 9966 21248
rect 10030 21184 10046 21248
rect 10110 21184 10126 21248
rect 10190 21184 10198 21248
rect 9878 21183 10198 21184
rect 19878 21248 20198 21249
rect 19878 21184 19886 21248
rect 19950 21184 19966 21248
rect 20030 21184 20046 21248
rect 20110 21184 20126 21248
rect 20190 21184 20198 21248
rect 19878 21183 20198 21184
rect 4878 20704 5198 20705
rect 4878 20640 4886 20704
rect 4950 20640 4966 20704
rect 5030 20640 5046 20704
rect 5110 20640 5126 20704
rect 5190 20640 5198 20704
rect 4878 20639 5198 20640
rect 14878 20704 15198 20705
rect 14878 20640 14886 20704
rect 14950 20640 14966 20704
rect 15030 20640 15046 20704
rect 15110 20640 15126 20704
rect 15190 20640 15198 20704
rect 14878 20639 15198 20640
rect 24878 20704 25198 20705
rect 24878 20640 24886 20704
rect 24950 20640 24966 20704
rect 25030 20640 25046 20704
rect 25110 20640 25126 20704
rect 25190 20640 25198 20704
rect 24878 20639 25198 20640
rect 15323 20498 15389 20501
rect 17623 20498 17689 20501
rect 15323 20496 17689 20498
rect 15323 20440 15328 20496
rect 15384 20440 17628 20496
rect 17684 20440 17689 20496
rect 15323 20438 17689 20440
rect 15323 20435 15389 20438
rect 17623 20435 17689 20438
rect 9878 20160 10198 20161
rect 9878 20096 9886 20160
rect 9950 20096 9966 20160
rect 10030 20096 10046 20160
rect 10110 20096 10126 20160
rect 10190 20096 10198 20160
rect 9878 20095 10198 20096
rect 19878 20160 20198 20161
rect 19878 20096 19886 20160
rect 19950 20096 19966 20160
rect 20030 20096 20046 20160
rect 20110 20096 20126 20160
rect 20190 20096 20198 20160
rect 19878 20095 20198 20096
rect 24431 19954 24497 19957
rect 28454 19954 28934 19984
rect 24431 19952 28934 19954
rect 24431 19896 24436 19952
rect 24492 19896 28934 19952
rect 24431 19894 28934 19896
rect 24431 19891 24497 19894
rect 28454 19864 28934 19894
rect 4878 19616 5198 19617
rect 4878 19552 4886 19616
rect 4950 19552 4966 19616
rect 5030 19552 5046 19616
rect 5110 19552 5126 19616
rect 5190 19552 5198 19616
rect 4878 19551 5198 19552
rect 14878 19616 15198 19617
rect 14878 19552 14886 19616
rect 14950 19552 14966 19616
rect 15030 19552 15046 19616
rect 15110 19552 15126 19616
rect 15190 19552 15198 19616
rect 14878 19551 15198 19552
rect 24878 19616 25198 19617
rect 24878 19552 24886 19616
rect 24950 19552 24966 19616
rect 25030 19552 25046 19616
rect 25110 19552 25126 19616
rect 25190 19552 25198 19616
rect 24878 19551 25198 19552
rect 10263 19410 10329 19413
rect 13391 19410 13457 19413
rect 10263 19408 13457 19410
rect 10263 19352 10268 19408
rect 10324 19352 13396 19408
rect 13452 19352 13457 19408
rect 10263 19350 13457 19352
rect 10263 19347 10329 19350
rect 13391 19347 13457 19350
rect 9878 19072 10198 19073
rect 9878 19008 9886 19072
rect 9950 19008 9966 19072
rect 10030 19008 10046 19072
rect 10110 19008 10126 19072
rect 10190 19008 10198 19072
rect 9878 19007 10198 19008
rect 19878 19072 20198 19073
rect 19878 19008 19886 19072
rect 19950 19008 19966 19072
rect 20030 19008 20046 19072
rect 20110 19008 20126 19072
rect 20190 19008 20198 19072
rect 19878 19007 20198 19008
rect 15139 18866 15205 18869
rect 24431 18866 24497 18869
rect 15139 18864 24497 18866
rect 15139 18808 15144 18864
rect 15200 18808 24436 18864
rect 24492 18808 24497 18864
rect 15139 18806 24497 18808
rect 15139 18803 15205 18806
rect 24431 18803 24497 18806
rect 4878 18528 5198 18529
rect 4878 18464 4886 18528
rect 4950 18464 4966 18528
rect 5030 18464 5046 18528
rect 5110 18464 5126 18528
rect 5190 18464 5198 18528
rect 4878 18463 5198 18464
rect 14878 18528 15198 18529
rect 14878 18464 14886 18528
rect 14950 18464 14966 18528
rect 15030 18464 15046 18528
rect 15110 18464 15126 18528
rect 15190 18464 15198 18528
rect 14878 18463 15198 18464
rect 24878 18528 25198 18529
rect 24878 18464 24886 18528
rect 24950 18464 24966 18528
rect 25030 18464 25046 18528
rect 25110 18464 25126 18528
rect 25190 18464 25198 18528
rect 24878 18463 25198 18464
rect 9878 17984 10198 17985
rect 9878 17920 9886 17984
rect 9950 17920 9966 17984
rect 10030 17920 10046 17984
rect 10110 17920 10126 17984
rect 10190 17920 10198 17984
rect 9878 17919 10198 17920
rect 19878 17984 20198 17985
rect 19878 17920 19886 17984
rect 19950 17920 19966 17984
rect 20030 17920 20046 17984
rect 20110 17920 20126 17984
rect 20190 17920 20198 17984
rect 19878 17919 20198 17920
rect 4878 17440 5198 17441
rect 4878 17376 4886 17440
rect 4950 17376 4966 17440
rect 5030 17376 5046 17440
rect 5110 17376 5126 17440
rect 5190 17376 5198 17440
rect 4878 17375 5198 17376
rect 14878 17440 15198 17441
rect 14878 17376 14886 17440
rect 14950 17376 14966 17440
rect 15030 17376 15046 17440
rect 15110 17376 15126 17440
rect 15190 17376 15198 17440
rect 14878 17375 15198 17376
rect 24878 17440 25198 17441
rect 24878 17376 24886 17440
rect 24950 17376 24966 17440
rect 25030 17376 25046 17440
rect 25110 17376 25126 17440
rect 25190 17376 25198 17440
rect 24878 17375 25198 17376
rect 9878 16896 10198 16897
rect 9878 16832 9886 16896
rect 9950 16832 9966 16896
rect 10030 16832 10046 16896
rect 10110 16832 10126 16896
rect 10190 16832 10198 16896
rect 9878 16831 10198 16832
rect 19878 16896 20198 16897
rect 19878 16832 19886 16896
rect 19950 16832 19966 16896
rect 20030 16832 20046 16896
rect 20110 16832 20126 16896
rect 20190 16832 20198 16896
rect 19878 16831 20198 16832
rect 4878 16352 5198 16353
rect 4878 16288 4886 16352
rect 4950 16288 4966 16352
rect 5030 16288 5046 16352
rect 5110 16288 5126 16352
rect 5190 16288 5198 16352
rect 4878 16287 5198 16288
rect 14878 16352 15198 16353
rect 14878 16288 14886 16352
rect 14950 16288 14966 16352
rect 15030 16288 15046 16352
rect 15110 16288 15126 16352
rect 15190 16288 15198 16352
rect 14878 16287 15198 16288
rect 24878 16352 25198 16353
rect 24878 16288 24886 16352
rect 24950 16288 24966 16352
rect 25030 16288 25046 16352
rect 25110 16288 25126 16352
rect 25190 16288 25198 16352
rect 24878 16287 25198 16288
rect 9878 15808 10198 15809
rect 9878 15744 9886 15808
rect 9950 15744 9966 15808
rect 10030 15744 10046 15808
rect 10110 15744 10126 15808
rect 10190 15744 10198 15808
rect 9878 15743 10198 15744
rect 19878 15808 20198 15809
rect 19878 15744 19886 15808
rect 19950 15744 19966 15808
rect 20030 15744 20046 15808
rect 20110 15744 20126 15808
rect 20190 15744 20198 15808
rect 19878 15743 20198 15744
rect 4878 15264 5198 15265
rect 4878 15200 4886 15264
rect 4950 15200 4966 15264
rect 5030 15200 5046 15264
rect 5110 15200 5126 15264
rect 5190 15200 5198 15264
rect 4878 15199 5198 15200
rect 14878 15264 15198 15265
rect 14878 15200 14886 15264
rect 14950 15200 14966 15264
rect 15030 15200 15046 15264
rect 15110 15200 15126 15264
rect 15190 15200 15198 15264
rect 14878 15199 15198 15200
rect 24878 15264 25198 15265
rect 24878 15200 24886 15264
rect 24950 15200 24966 15264
rect 25030 15200 25046 15264
rect 25110 15200 25126 15264
rect 25190 15200 25198 15264
rect 24878 15199 25198 15200
rect 9878 14720 10198 14721
rect 9878 14656 9886 14720
rect 9950 14656 9966 14720
rect 10030 14656 10046 14720
rect 10110 14656 10126 14720
rect 10190 14656 10198 14720
rect 9878 14655 10198 14656
rect 19878 14720 20198 14721
rect 19878 14656 19886 14720
rect 19950 14656 19966 14720
rect 20030 14656 20046 14720
rect 20110 14656 20126 14720
rect 20190 14656 20198 14720
rect 19878 14655 20198 14656
rect 4878 14176 5198 14177
rect 4878 14112 4886 14176
rect 4950 14112 4966 14176
rect 5030 14112 5046 14176
rect 5110 14112 5126 14176
rect 5190 14112 5198 14176
rect 4878 14111 5198 14112
rect 14878 14176 15198 14177
rect 14878 14112 14886 14176
rect 14950 14112 14966 14176
rect 15030 14112 15046 14176
rect 15110 14112 15126 14176
rect 15190 14112 15198 14176
rect 14878 14111 15198 14112
rect 24878 14176 25198 14177
rect 24878 14112 24886 14176
rect 24950 14112 24966 14176
rect 25030 14112 25046 14176
rect 25110 14112 25126 14176
rect 25190 14112 25198 14176
rect 24878 14111 25198 14112
rect 9878 13632 10198 13633
rect 9878 13568 9886 13632
rect 9950 13568 9966 13632
rect 10030 13568 10046 13632
rect 10110 13568 10126 13632
rect 10190 13568 10198 13632
rect 9878 13567 10198 13568
rect 19878 13632 20198 13633
rect 19878 13568 19886 13632
rect 19950 13568 19966 13632
rect 20030 13568 20046 13632
rect 20110 13568 20126 13632
rect 20190 13568 20198 13632
rect 19878 13567 20198 13568
rect 4878 13088 5198 13089
rect 4878 13024 4886 13088
rect 4950 13024 4966 13088
rect 5030 13024 5046 13088
rect 5110 13024 5126 13088
rect 5190 13024 5198 13088
rect 4878 13023 5198 13024
rect 14878 13088 15198 13089
rect 14878 13024 14886 13088
rect 14950 13024 14966 13088
rect 15030 13024 15046 13088
rect 15110 13024 15126 13088
rect 15190 13024 15198 13088
rect 14878 13023 15198 13024
rect 24878 13088 25198 13089
rect 24878 13024 24886 13088
rect 24950 13024 24966 13088
rect 25030 13024 25046 13088
rect 25110 13024 25126 13088
rect 25190 13024 25198 13088
rect 24878 13023 25198 13024
rect 9878 12544 10198 12545
rect 9878 12480 9886 12544
rect 9950 12480 9966 12544
rect 10030 12480 10046 12544
rect 10110 12480 10126 12544
rect 10190 12480 10198 12544
rect 9878 12479 10198 12480
rect 19878 12544 20198 12545
rect 19878 12480 19886 12544
rect 19950 12480 19966 12544
rect 20030 12480 20046 12544
rect 20110 12480 20126 12544
rect 20190 12480 20198 12544
rect 19878 12479 20198 12480
rect 4878 12000 5198 12001
rect 4878 11936 4886 12000
rect 4950 11936 4966 12000
rect 5030 11936 5046 12000
rect 5110 11936 5126 12000
rect 5190 11936 5198 12000
rect 4878 11935 5198 11936
rect 14878 12000 15198 12001
rect 14878 11936 14886 12000
rect 14950 11936 14966 12000
rect 15030 11936 15046 12000
rect 15110 11936 15126 12000
rect 15190 11936 15198 12000
rect 14878 11935 15198 11936
rect 24878 12000 25198 12001
rect 24878 11936 24886 12000
rect 24950 11936 24966 12000
rect 25030 11936 25046 12000
rect 25110 11936 25126 12000
rect 25190 11936 25198 12000
rect 24878 11935 25198 11936
rect 28454 11930 28934 11960
rect 26780 11870 28934 11930
rect 23879 11794 23945 11797
rect 26780 11794 26840 11870
rect 28454 11840 28934 11870
rect 23879 11792 26840 11794
rect 23879 11736 23884 11792
rect 23940 11736 26840 11792
rect 23879 11734 26840 11736
rect 23879 11731 23945 11734
rect 9878 11456 10198 11457
rect 9878 11392 9886 11456
rect 9950 11392 9966 11456
rect 10030 11392 10046 11456
rect 10110 11392 10126 11456
rect 10190 11392 10198 11456
rect 9878 11391 10198 11392
rect 19878 11456 20198 11457
rect 19878 11392 19886 11456
rect 19950 11392 19966 11456
rect 20030 11392 20046 11456
rect 20110 11392 20126 11456
rect 20190 11392 20198 11456
rect 19878 11391 20198 11392
rect 4878 10912 5198 10913
rect 4878 10848 4886 10912
rect 4950 10848 4966 10912
rect 5030 10848 5046 10912
rect 5110 10848 5126 10912
rect 5190 10848 5198 10912
rect 4878 10847 5198 10848
rect 14878 10912 15198 10913
rect 14878 10848 14886 10912
rect 14950 10848 14966 10912
rect 15030 10848 15046 10912
rect 15110 10848 15126 10912
rect 15190 10848 15198 10912
rect 14878 10847 15198 10848
rect 24878 10912 25198 10913
rect 24878 10848 24886 10912
rect 24950 10848 24966 10912
rect 25030 10848 25046 10912
rect 25110 10848 25126 10912
rect 25190 10848 25198 10912
rect 24878 10847 25198 10848
rect 2995 10570 3061 10573
rect 10171 10570 10237 10573
rect 2995 10568 10237 10570
rect 2995 10512 3000 10568
rect 3056 10512 10176 10568
rect 10232 10512 10237 10568
rect 2995 10510 10237 10512
rect 2995 10507 3061 10510
rect 10171 10507 10237 10510
rect 9878 10368 10198 10369
rect 9878 10304 9886 10368
rect 9950 10304 9966 10368
rect 10030 10304 10046 10368
rect 10110 10304 10126 10368
rect 10190 10304 10198 10368
rect 9878 10303 10198 10304
rect 19878 10368 20198 10369
rect 19878 10304 19886 10368
rect 19950 10304 19966 10368
rect 20030 10304 20046 10368
rect 20110 10304 20126 10368
rect 20190 10304 20198 10368
rect 19878 10303 20198 10304
rect 4878 9824 5198 9825
rect 4878 9760 4886 9824
rect 4950 9760 4966 9824
rect 5030 9760 5046 9824
rect 5110 9760 5126 9824
rect 5190 9760 5198 9824
rect 4878 9759 5198 9760
rect 14878 9824 15198 9825
rect 14878 9760 14886 9824
rect 14950 9760 14966 9824
rect 15030 9760 15046 9824
rect 15110 9760 15126 9824
rect 15190 9760 15198 9824
rect 14878 9759 15198 9760
rect 24878 9824 25198 9825
rect 24878 9760 24886 9824
rect 24950 9760 24966 9824
rect 25030 9760 25046 9824
rect 25110 9760 25126 9824
rect 25190 9760 25198 9824
rect 24878 9759 25198 9760
rect 9878 9280 10198 9281
rect 9878 9216 9886 9280
rect 9950 9216 9966 9280
rect 10030 9216 10046 9280
rect 10110 9216 10126 9280
rect 10190 9216 10198 9280
rect 9878 9215 10198 9216
rect 19878 9280 20198 9281
rect 19878 9216 19886 9280
rect 19950 9216 19966 9280
rect 20030 9216 20046 9280
rect 20110 9216 20126 9280
rect 20190 9216 20198 9280
rect 19878 9215 20198 9216
rect 4878 8736 5198 8737
rect 4878 8672 4886 8736
rect 4950 8672 4966 8736
rect 5030 8672 5046 8736
rect 5110 8672 5126 8736
rect 5190 8672 5198 8736
rect 4878 8671 5198 8672
rect 14878 8736 15198 8737
rect 14878 8672 14886 8736
rect 14950 8672 14966 8736
rect 15030 8672 15046 8736
rect 15110 8672 15126 8736
rect 15190 8672 15198 8736
rect 14878 8671 15198 8672
rect 24878 8736 25198 8737
rect 24878 8672 24886 8736
rect 24950 8672 24966 8736
rect 25030 8672 25046 8736
rect 25110 8672 25126 8736
rect 25190 8672 25198 8736
rect 24878 8671 25198 8672
rect 9878 8192 10198 8193
rect 9878 8128 9886 8192
rect 9950 8128 9966 8192
rect 10030 8128 10046 8192
rect 10110 8128 10126 8192
rect 10190 8128 10198 8192
rect 9878 8127 10198 8128
rect 19878 8192 20198 8193
rect 19878 8128 19886 8192
rect 19950 8128 19966 8192
rect 20030 8128 20046 8192
rect 20110 8128 20126 8192
rect 20190 8128 20198 8192
rect 19878 8127 20198 8128
rect 4878 7648 5198 7649
rect 4878 7584 4886 7648
rect 4950 7584 4966 7648
rect 5030 7584 5046 7648
rect 5110 7584 5126 7648
rect 5190 7584 5198 7648
rect 4878 7583 5198 7584
rect 14878 7648 15198 7649
rect 14878 7584 14886 7648
rect 14950 7584 14966 7648
rect 15030 7584 15046 7648
rect 15110 7584 15126 7648
rect 15190 7584 15198 7648
rect 14878 7583 15198 7584
rect 24878 7648 25198 7649
rect 24878 7584 24886 7648
rect 24950 7584 24966 7648
rect 25030 7584 25046 7648
rect 25110 7584 25126 7648
rect 25190 7584 25198 7648
rect 24878 7583 25198 7584
rect 9878 7104 10198 7105
rect 9878 7040 9886 7104
rect 9950 7040 9966 7104
rect 10030 7040 10046 7104
rect 10110 7040 10126 7104
rect 10190 7040 10198 7104
rect 9878 7039 10198 7040
rect 19878 7104 20198 7105
rect 19878 7040 19886 7104
rect 19950 7040 19966 7104
rect 20030 7040 20046 7104
rect 20110 7040 20126 7104
rect 20190 7040 20198 7104
rect 19878 7039 20198 7040
rect 4878 6560 5198 6561
rect 4878 6496 4886 6560
rect 4950 6496 4966 6560
rect 5030 6496 5046 6560
rect 5110 6496 5126 6560
rect 5190 6496 5198 6560
rect 4878 6495 5198 6496
rect 14878 6560 15198 6561
rect 14878 6496 14886 6560
rect 14950 6496 14966 6560
rect 15030 6496 15046 6560
rect 15110 6496 15126 6560
rect 15190 6496 15198 6560
rect 14878 6495 15198 6496
rect 24878 6560 25198 6561
rect 24878 6496 24886 6560
rect 24950 6496 24966 6560
rect 25030 6496 25046 6560
rect 25110 6496 25126 6560
rect 25190 6496 25198 6560
rect 24878 6495 25198 6496
rect 9878 6016 10198 6017
rect 9878 5952 9886 6016
rect 9950 5952 9966 6016
rect 10030 5952 10046 6016
rect 10110 5952 10126 6016
rect 10190 5952 10198 6016
rect 9878 5951 10198 5952
rect 19878 6016 20198 6017
rect 19878 5952 19886 6016
rect 19950 5952 19966 6016
rect 20030 5952 20046 6016
rect 20110 5952 20126 6016
rect 20190 5952 20198 6016
rect 19878 5951 20198 5952
rect 10539 5674 10605 5677
rect 13851 5674 13917 5677
rect 10539 5672 13917 5674
rect 10539 5616 10544 5672
rect 10600 5616 13856 5672
rect 13912 5616 13917 5672
rect 10539 5614 13917 5616
rect 10539 5611 10605 5614
rect 13851 5611 13917 5614
rect 4878 5472 5198 5473
rect 4878 5408 4886 5472
rect 4950 5408 4966 5472
rect 5030 5408 5046 5472
rect 5110 5408 5126 5472
rect 5190 5408 5198 5472
rect 4878 5407 5198 5408
rect 14878 5472 15198 5473
rect 14878 5408 14886 5472
rect 14950 5408 14966 5472
rect 15030 5408 15046 5472
rect 15110 5408 15126 5472
rect 15190 5408 15198 5472
rect 14878 5407 15198 5408
rect 24878 5472 25198 5473
rect 24878 5408 24886 5472
rect 24950 5408 24966 5472
rect 25030 5408 25046 5472
rect 25110 5408 25126 5472
rect 25190 5408 25198 5472
rect 24878 5407 25198 5408
rect 9878 4928 10198 4929
rect 9878 4864 9886 4928
rect 9950 4864 9966 4928
rect 10030 4864 10046 4928
rect 10110 4864 10126 4928
rect 10190 4864 10198 4928
rect 9878 4863 10198 4864
rect 19878 4928 20198 4929
rect 19878 4864 19886 4928
rect 19950 4864 19966 4928
rect 20030 4864 20046 4928
rect 20110 4864 20126 4928
rect 20190 4864 20198 4928
rect 19878 4863 20198 4864
rect 4878 4384 5198 4385
rect 4878 4320 4886 4384
rect 4950 4320 4966 4384
rect 5030 4320 5046 4384
rect 5110 4320 5126 4384
rect 5190 4320 5198 4384
rect 4878 4319 5198 4320
rect 14878 4384 15198 4385
rect 14878 4320 14886 4384
rect 14950 4320 14966 4384
rect 15030 4320 15046 4384
rect 15110 4320 15126 4384
rect 15190 4320 15198 4384
rect 14878 4319 15198 4320
rect 24878 4384 25198 4385
rect 24878 4320 24886 4384
rect 24950 4320 24966 4384
rect 25030 4320 25046 4384
rect 25110 4320 25126 4384
rect 25190 4320 25198 4384
rect 24878 4319 25198 4320
rect 22867 4042 22933 4045
rect 28454 4042 28934 4072
rect 22867 4040 28934 4042
rect 22867 3984 22872 4040
rect 22928 3984 28934 4040
rect 22867 3982 28934 3984
rect 22867 3979 22933 3982
rect 28454 3952 28934 3982
rect 9878 3840 10198 3841
rect 9878 3776 9886 3840
rect 9950 3776 9966 3840
rect 10030 3776 10046 3840
rect 10110 3776 10126 3840
rect 10190 3776 10198 3840
rect 9878 3775 10198 3776
rect 19878 3840 20198 3841
rect 19878 3776 19886 3840
rect 19950 3776 19966 3840
rect 20030 3776 20046 3840
rect 20110 3776 20126 3840
rect 20190 3776 20198 3840
rect 19878 3775 20198 3776
rect 4878 3296 5198 3297
rect 4878 3232 4886 3296
rect 4950 3232 4966 3296
rect 5030 3232 5046 3296
rect 5110 3232 5126 3296
rect 5190 3232 5198 3296
rect 4878 3231 5198 3232
rect 14878 3296 15198 3297
rect 14878 3232 14886 3296
rect 14950 3232 14966 3296
rect 15030 3232 15046 3296
rect 15110 3232 15126 3296
rect 15190 3232 15198 3296
rect 14878 3231 15198 3232
rect 24878 3296 25198 3297
rect 24878 3232 24886 3296
rect 24950 3232 24966 3296
rect 25030 3232 25046 3296
rect 25110 3232 25126 3296
rect 25190 3232 25198 3296
rect 24878 3231 25198 3232
rect 3915 2954 3981 2957
rect 20475 2954 20541 2957
rect 3915 2952 20541 2954
rect 3915 2896 3920 2952
rect 3976 2896 20480 2952
rect 20536 2896 20541 2952
rect 3915 2894 20541 2896
rect 3915 2891 3981 2894
rect 20475 2891 20541 2894
rect 9878 2752 10198 2753
rect 9878 2688 9886 2752
rect 9950 2688 9966 2752
rect 10030 2688 10046 2752
rect 10110 2688 10126 2752
rect 10190 2688 10198 2752
rect 9878 2687 10198 2688
rect 19878 2752 20198 2753
rect 19878 2688 19886 2752
rect 19950 2688 19966 2752
rect 20030 2688 20046 2752
rect 20110 2688 20126 2752
rect 20190 2688 20198 2752
rect 19878 2687 20198 2688
rect 22039 2682 22105 2685
rect 23787 2682 23853 2685
rect 22039 2680 23853 2682
rect 22039 2624 22044 2680
rect 22100 2624 23792 2680
rect 23848 2624 23853 2680
rect 22039 2622 23853 2624
rect 22039 2619 22105 2622
rect 23787 2619 23853 2622
rect 4878 2208 5198 2209
rect 4878 2144 4886 2208
rect 4950 2144 4966 2208
rect 5030 2144 5046 2208
rect 5110 2144 5126 2208
rect 5190 2144 5198 2208
rect 4878 2143 5198 2144
rect 14878 2208 15198 2209
rect 14878 2144 14886 2208
rect 14950 2144 14966 2208
rect 15030 2144 15046 2208
rect 15110 2144 15126 2208
rect 15190 2144 15198 2208
rect 14878 2143 15198 2144
rect 24878 2208 25198 2209
rect 24878 2144 24886 2208
rect 24950 2144 24966 2208
rect 25030 2144 25046 2208
rect 25110 2144 25126 2208
rect 25190 2144 25198 2208
rect 24878 2143 25198 2144
<< via3 >>
rect 4886 21788 4950 21792
rect 4886 21732 4890 21788
rect 4890 21732 4946 21788
rect 4946 21732 4950 21788
rect 4886 21728 4950 21732
rect 4966 21788 5030 21792
rect 4966 21732 4970 21788
rect 4970 21732 5026 21788
rect 5026 21732 5030 21788
rect 4966 21728 5030 21732
rect 5046 21788 5110 21792
rect 5046 21732 5050 21788
rect 5050 21732 5106 21788
rect 5106 21732 5110 21788
rect 5046 21728 5110 21732
rect 5126 21788 5190 21792
rect 5126 21732 5130 21788
rect 5130 21732 5186 21788
rect 5186 21732 5190 21788
rect 5126 21728 5190 21732
rect 14886 21788 14950 21792
rect 14886 21732 14890 21788
rect 14890 21732 14946 21788
rect 14946 21732 14950 21788
rect 14886 21728 14950 21732
rect 14966 21788 15030 21792
rect 14966 21732 14970 21788
rect 14970 21732 15026 21788
rect 15026 21732 15030 21788
rect 14966 21728 15030 21732
rect 15046 21788 15110 21792
rect 15046 21732 15050 21788
rect 15050 21732 15106 21788
rect 15106 21732 15110 21788
rect 15046 21728 15110 21732
rect 15126 21788 15190 21792
rect 15126 21732 15130 21788
rect 15130 21732 15186 21788
rect 15186 21732 15190 21788
rect 15126 21728 15190 21732
rect 24886 21788 24950 21792
rect 24886 21732 24890 21788
rect 24890 21732 24946 21788
rect 24946 21732 24950 21788
rect 24886 21728 24950 21732
rect 24966 21788 25030 21792
rect 24966 21732 24970 21788
rect 24970 21732 25026 21788
rect 25026 21732 25030 21788
rect 24966 21728 25030 21732
rect 25046 21788 25110 21792
rect 25046 21732 25050 21788
rect 25050 21732 25106 21788
rect 25106 21732 25110 21788
rect 25046 21728 25110 21732
rect 25126 21788 25190 21792
rect 25126 21732 25130 21788
rect 25130 21732 25186 21788
rect 25186 21732 25190 21788
rect 25126 21728 25190 21732
rect 9886 21244 9950 21248
rect 9886 21188 9890 21244
rect 9890 21188 9946 21244
rect 9946 21188 9950 21244
rect 9886 21184 9950 21188
rect 9966 21244 10030 21248
rect 9966 21188 9970 21244
rect 9970 21188 10026 21244
rect 10026 21188 10030 21244
rect 9966 21184 10030 21188
rect 10046 21244 10110 21248
rect 10046 21188 10050 21244
rect 10050 21188 10106 21244
rect 10106 21188 10110 21244
rect 10046 21184 10110 21188
rect 10126 21244 10190 21248
rect 10126 21188 10130 21244
rect 10130 21188 10186 21244
rect 10186 21188 10190 21244
rect 10126 21184 10190 21188
rect 19886 21244 19950 21248
rect 19886 21188 19890 21244
rect 19890 21188 19946 21244
rect 19946 21188 19950 21244
rect 19886 21184 19950 21188
rect 19966 21244 20030 21248
rect 19966 21188 19970 21244
rect 19970 21188 20026 21244
rect 20026 21188 20030 21244
rect 19966 21184 20030 21188
rect 20046 21244 20110 21248
rect 20046 21188 20050 21244
rect 20050 21188 20106 21244
rect 20106 21188 20110 21244
rect 20046 21184 20110 21188
rect 20126 21244 20190 21248
rect 20126 21188 20130 21244
rect 20130 21188 20186 21244
rect 20186 21188 20190 21244
rect 20126 21184 20190 21188
rect 4886 20700 4950 20704
rect 4886 20644 4890 20700
rect 4890 20644 4946 20700
rect 4946 20644 4950 20700
rect 4886 20640 4950 20644
rect 4966 20700 5030 20704
rect 4966 20644 4970 20700
rect 4970 20644 5026 20700
rect 5026 20644 5030 20700
rect 4966 20640 5030 20644
rect 5046 20700 5110 20704
rect 5046 20644 5050 20700
rect 5050 20644 5106 20700
rect 5106 20644 5110 20700
rect 5046 20640 5110 20644
rect 5126 20700 5190 20704
rect 5126 20644 5130 20700
rect 5130 20644 5186 20700
rect 5186 20644 5190 20700
rect 5126 20640 5190 20644
rect 14886 20700 14950 20704
rect 14886 20644 14890 20700
rect 14890 20644 14946 20700
rect 14946 20644 14950 20700
rect 14886 20640 14950 20644
rect 14966 20700 15030 20704
rect 14966 20644 14970 20700
rect 14970 20644 15026 20700
rect 15026 20644 15030 20700
rect 14966 20640 15030 20644
rect 15046 20700 15110 20704
rect 15046 20644 15050 20700
rect 15050 20644 15106 20700
rect 15106 20644 15110 20700
rect 15046 20640 15110 20644
rect 15126 20700 15190 20704
rect 15126 20644 15130 20700
rect 15130 20644 15186 20700
rect 15186 20644 15190 20700
rect 15126 20640 15190 20644
rect 24886 20700 24950 20704
rect 24886 20644 24890 20700
rect 24890 20644 24946 20700
rect 24946 20644 24950 20700
rect 24886 20640 24950 20644
rect 24966 20700 25030 20704
rect 24966 20644 24970 20700
rect 24970 20644 25026 20700
rect 25026 20644 25030 20700
rect 24966 20640 25030 20644
rect 25046 20700 25110 20704
rect 25046 20644 25050 20700
rect 25050 20644 25106 20700
rect 25106 20644 25110 20700
rect 25046 20640 25110 20644
rect 25126 20700 25190 20704
rect 25126 20644 25130 20700
rect 25130 20644 25186 20700
rect 25186 20644 25190 20700
rect 25126 20640 25190 20644
rect 9886 20156 9950 20160
rect 9886 20100 9890 20156
rect 9890 20100 9946 20156
rect 9946 20100 9950 20156
rect 9886 20096 9950 20100
rect 9966 20156 10030 20160
rect 9966 20100 9970 20156
rect 9970 20100 10026 20156
rect 10026 20100 10030 20156
rect 9966 20096 10030 20100
rect 10046 20156 10110 20160
rect 10046 20100 10050 20156
rect 10050 20100 10106 20156
rect 10106 20100 10110 20156
rect 10046 20096 10110 20100
rect 10126 20156 10190 20160
rect 10126 20100 10130 20156
rect 10130 20100 10186 20156
rect 10186 20100 10190 20156
rect 10126 20096 10190 20100
rect 19886 20156 19950 20160
rect 19886 20100 19890 20156
rect 19890 20100 19946 20156
rect 19946 20100 19950 20156
rect 19886 20096 19950 20100
rect 19966 20156 20030 20160
rect 19966 20100 19970 20156
rect 19970 20100 20026 20156
rect 20026 20100 20030 20156
rect 19966 20096 20030 20100
rect 20046 20156 20110 20160
rect 20046 20100 20050 20156
rect 20050 20100 20106 20156
rect 20106 20100 20110 20156
rect 20046 20096 20110 20100
rect 20126 20156 20190 20160
rect 20126 20100 20130 20156
rect 20130 20100 20186 20156
rect 20186 20100 20190 20156
rect 20126 20096 20190 20100
rect 4886 19612 4950 19616
rect 4886 19556 4890 19612
rect 4890 19556 4946 19612
rect 4946 19556 4950 19612
rect 4886 19552 4950 19556
rect 4966 19612 5030 19616
rect 4966 19556 4970 19612
rect 4970 19556 5026 19612
rect 5026 19556 5030 19612
rect 4966 19552 5030 19556
rect 5046 19612 5110 19616
rect 5046 19556 5050 19612
rect 5050 19556 5106 19612
rect 5106 19556 5110 19612
rect 5046 19552 5110 19556
rect 5126 19612 5190 19616
rect 5126 19556 5130 19612
rect 5130 19556 5186 19612
rect 5186 19556 5190 19612
rect 5126 19552 5190 19556
rect 14886 19612 14950 19616
rect 14886 19556 14890 19612
rect 14890 19556 14946 19612
rect 14946 19556 14950 19612
rect 14886 19552 14950 19556
rect 14966 19612 15030 19616
rect 14966 19556 14970 19612
rect 14970 19556 15026 19612
rect 15026 19556 15030 19612
rect 14966 19552 15030 19556
rect 15046 19612 15110 19616
rect 15046 19556 15050 19612
rect 15050 19556 15106 19612
rect 15106 19556 15110 19612
rect 15046 19552 15110 19556
rect 15126 19612 15190 19616
rect 15126 19556 15130 19612
rect 15130 19556 15186 19612
rect 15186 19556 15190 19612
rect 15126 19552 15190 19556
rect 24886 19612 24950 19616
rect 24886 19556 24890 19612
rect 24890 19556 24946 19612
rect 24946 19556 24950 19612
rect 24886 19552 24950 19556
rect 24966 19612 25030 19616
rect 24966 19556 24970 19612
rect 24970 19556 25026 19612
rect 25026 19556 25030 19612
rect 24966 19552 25030 19556
rect 25046 19612 25110 19616
rect 25046 19556 25050 19612
rect 25050 19556 25106 19612
rect 25106 19556 25110 19612
rect 25046 19552 25110 19556
rect 25126 19612 25190 19616
rect 25126 19556 25130 19612
rect 25130 19556 25186 19612
rect 25186 19556 25190 19612
rect 25126 19552 25190 19556
rect 9886 19068 9950 19072
rect 9886 19012 9890 19068
rect 9890 19012 9946 19068
rect 9946 19012 9950 19068
rect 9886 19008 9950 19012
rect 9966 19068 10030 19072
rect 9966 19012 9970 19068
rect 9970 19012 10026 19068
rect 10026 19012 10030 19068
rect 9966 19008 10030 19012
rect 10046 19068 10110 19072
rect 10046 19012 10050 19068
rect 10050 19012 10106 19068
rect 10106 19012 10110 19068
rect 10046 19008 10110 19012
rect 10126 19068 10190 19072
rect 10126 19012 10130 19068
rect 10130 19012 10186 19068
rect 10186 19012 10190 19068
rect 10126 19008 10190 19012
rect 19886 19068 19950 19072
rect 19886 19012 19890 19068
rect 19890 19012 19946 19068
rect 19946 19012 19950 19068
rect 19886 19008 19950 19012
rect 19966 19068 20030 19072
rect 19966 19012 19970 19068
rect 19970 19012 20026 19068
rect 20026 19012 20030 19068
rect 19966 19008 20030 19012
rect 20046 19068 20110 19072
rect 20046 19012 20050 19068
rect 20050 19012 20106 19068
rect 20106 19012 20110 19068
rect 20046 19008 20110 19012
rect 20126 19068 20190 19072
rect 20126 19012 20130 19068
rect 20130 19012 20186 19068
rect 20186 19012 20190 19068
rect 20126 19008 20190 19012
rect 4886 18524 4950 18528
rect 4886 18468 4890 18524
rect 4890 18468 4946 18524
rect 4946 18468 4950 18524
rect 4886 18464 4950 18468
rect 4966 18524 5030 18528
rect 4966 18468 4970 18524
rect 4970 18468 5026 18524
rect 5026 18468 5030 18524
rect 4966 18464 5030 18468
rect 5046 18524 5110 18528
rect 5046 18468 5050 18524
rect 5050 18468 5106 18524
rect 5106 18468 5110 18524
rect 5046 18464 5110 18468
rect 5126 18524 5190 18528
rect 5126 18468 5130 18524
rect 5130 18468 5186 18524
rect 5186 18468 5190 18524
rect 5126 18464 5190 18468
rect 14886 18524 14950 18528
rect 14886 18468 14890 18524
rect 14890 18468 14946 18524
rect 14946 18468 14950 18524
rect 14886 18464 14950 18468
rect 14966 18524 15030 18528
rect 14966 18468 14970 18524
rect 14970 18468 15026 18524
rect 15026 18468 15030 18524
rect 14966 18464 15030 18468
rect 15046 18524 15110 18528
rect 15046 18468 15050 18524
rect 15050 18468 15106 18524
rect 15106 18468 15110 18524
rect 15046 18464 15110 18468
rect 15126 18524 15190 18528
rect 15126 18468 15130 18524
rect 15130 18468 15186 18524
rect 15186 18468 15190 18524
rect 15126 18464 15190 18468
rect 24886 18524 24950 18528
rect 24886 18468 24890 18524
rect 24890 18468 24946 18524
rect 24946 18468 24950 18524
rect 24886 18464 24950 18468
rect 24966 18524 25030 18528
rect 24966 18468 24970 18524
rect 24970 18468 25026 18524
rect 25026 18468 25030 18524
rect 24966 18464 25030 18468
rect 25046 18524 25110 18528
rect 25046 18468 25050 18524
rect 25050 18468 25106 18524
rect 25106 18468 25110 18524
rect 25046 18464 25110 18468
rect 25126 18524 25190 18528
rect 25126 18468 25130 18524
rect 25130 18468 25186 18524
rect 25186 18468 25190 18524
rect 25126 18464 25190 18468
rect 9886 17980 9950 17984
rect 9886 17924 9890 17980
rect 9890 17924 9946 17980
rect 9946 17924 9950 17980
rect 9886 17920 9950 17924
rect 9966 17980 10030 17984
rect 9966 17924 9970 17980
rect 9970 17924 10026 17980
rect 10026 17924 10030 17980
rect 9966 17920 10030 17924
rect 10046 17980 10110 17984
rect 10046 17924 10050 17980
rect 10050 17924 10106 17980
rect 10106 17924 10110 17980
rect 10046 17920 10110 17924
rect 10126 17980 10190 17984
rect 10126 17924 10130 17980
rect 10130 17924 10186 17980
rect 10186 17924 10190 17980
rect 10126 17920 10190 17924
rect 19886 17980 19950 17984
rect 19886 17924 19890 17980
rect 19890 17924 19946 17980
rect 19946 17924 19950 17980
rect 19886 17920 19950 17924
rect 19966 17980 20030 17984
rect 19966 17924 19970 17980
rect 19970 17924 20026 17980
rect 20026 17924 20030 17980
rect 19966 17920 20030 17924
rect 20046 17980 20110 17984
rect 20046 17924 20050 17980
rect 20050 17924 20106 17980
rect 20106 17924 20110 17980
rect 20046 17920 20110 17924
rect 20126 17980 20190 17984
rect 20126 17924 20130 17980
rect 20130 17924 20186 17980
rect 20186 17924 20190 17980
rect 20126 17920 20190 17924
rect 4886 17436 4950 17440
rect 4886 17380 4890 17436
rect 4890 17380 4946 17436
rect 4946 17380 4950 17436
rect 4886 17376 4950 17380
rect 4966 17436 5030 17440
rect 4966 17380 4970 17436
rect 4970 17380 5026 17436
rect 5026 17380 5030 17436
rect 4966 17376 5030 17380
rect 5046 17436 5110 17440
rect 5046 17380 5050 17436
rect 5050 17380 5106 17436
rect 5106 17380 5110 17436
rect 5046 17376 5110 17380
rect 5126 17436 5190 17440
rect 5126 17380 5130 17436
rect 5130 17380 5186 17436
rect 5186 17380 5190 17436
rect 5126 17376 5190 17380
rect 14886 17436 14950 17440
rect 14886 17380 14890 17436
rect 14890 17380 14946 17436
rect 14946 17380 14950 17436
rect 14886 17376 14950 17380
rect 14966 17436 15030 17440
rect 14966 17380 14970 17436
rect 14970 17380 15026 17436
rect 15026 17380 15030 17436
rect 14966 17376 15030 17380
rect 15046 17436 15110 17440
rect 15046 17380 15050 17436
rect 15050 17380 15106 17436
rect 15106 17380 15110 17436
rect 15046 17376 15110 17380
rect 15126 17436 15190 17440
rect 15126 17380 15130 17436
rect 15130 17380 15186 17436
rect 15186 17380 15190 17436
rect 15126 17376 15190 17380
rect 24886 17436 24950 17440
rect 24886 17380 24890 17436
rect 24890 17380 24946 17436
rect 24946 17380 24950 17436
rect 24886 17376 24950 17380
rect 24966 17436 25030 17440
rect 24966 17380 24970 17436
rect 24970 17380 25026 17436
rect 25026 17380 25030 17436
rect 24966 17376 25030 17380
rect 25046 17436 25110 17440
rect 25046 17380 25050 17436
rect 25050 17380 25106 17436
rect 25106 17380 25110 17436
rect 25046 17376 25110 17380
rect 25126 17436 25190 17440
rect 25126 17380 25130 17436
rect 25130 17380 25186 17436
rect 25186 17380 25190 17436
rect 25126 17376 25190 17380
rect 9886 16892 9950 16896
rect 9886 16836 9890 16892
rect 9890 16836 9946 16892
rect 9946 16836 9950 16892
rect 9886 16832 9950 16836
rect 9966 16892 10030 16896
rect 9966 16836 9970 16892
rect 9970 16836 10026 16892
rect 10026 16836 10030 16892
rect 9966 16832 10030 16836
rect 10046 16892 10110 16896
rect 10046 16836 10050 16892
rect 10050 16836 10106 16892
rect 10106 16836 10110 16892
rect 10046 16832 10110 16836
rect 10126 16892 10190 16896
rect 10126 16836 10130 16892
rect 10130 16836 10186 16892
rect 10186 16836 10190 16892
rect 10126 16832 10190 16836
rect 19886 16892 19950 16896
rect 19886 16836 19890 16892
rect 19890 16836 19946 16892
rect 19946 16836 19950 16892
rect 19886 16832 19950 16836
rect 19966 16892 20030 16896
rect 19966 16836 19970 16892
rect 19970 16836 20026 16892
rect 20026 16836 20030 16892
rect 19966 16832 20030 16836
rect 20046 16892 20110 16896
rect 20046 16836 20050 16892
rect 20050 16836 20106 16892
rect 20106 16836 20110 16892
rect 20046 16832 20110 16836
rect 20126 16892 20190 16896
rect 20126 16836 20130 16892
rect 20130 16836 20186 16892
rect 20186 16836 20190 16892
rect 20126 16832 20190 16836
rect 4886 16348 4950 16352
rect 4886 16292 4890 16348
rect 4890 16292 4946 16348
rect 4946 16292 4950 16348
rect 4886 16288 4950 16292
rect 4966 16348 5030 16352
rect 4966 16292 4970 16348
rect 4970 16292 5026 16348
rect 5026 16292 5030 16348
rect 4966 16288 5030 16292
rect 5046 16348 5110 16352
rect 5046 16292 5050 16348
rect 5050 16292 5106 16348
rect 5106 16292 5110 16348
rect 5046 16288 5110 16292
rect 5126 16348 5190 16352
rect 5126 16292 5130 16348
rect 5130 16292 5186 16348
rect 5186 16292 5190 16348
rect 5126 16288 5190 16292
rect 14886 16348 14950 16352
rect 14886 16292 14890 16348
rect 14890 16292 14946 16348
rect 14946 16292 14950 16348
rect 14886 16288 14950 16292
rect 14966 16348 15030 16352
rect 14966 16292 14970 16348
rect 14970 16292 15026 16348
rect 15026 16292 15030 16348
rect 14966 16288 15030 16292
rect 15046 16348 15110 16352
rect 15046 16292 15050 16348
rect 15050 16292 15106 16348
rect 15106 16292 15110 16348
rect 15046 16288 15110 16292
rect 15126 16348 15190 16352
rect 15126 16292 15130 16348
rect 15130 16292 15186 16348
rect 15186 16292 15190 16348
rect 15126 16288 15190 16292
rect 24886 16348 24950 16352
rect 24886 16292 24890 16348
rect 24890 16292 24946 16348
rect 24946 16292 24950 16348
rect 24886 16288 24950 16292
rect 24966 16348 25030 16352
rect 24966 16292 24970 16348
rect 24970 16292 25026 16348
rect 25026 16292 25030 16348
rect 24966 16288 25030 16292
rect 25046 16348 25110 16352
rect 25046 16292 25050 16348
rect 25050 16292 25106 16348
rect 25106 16292 25110 16348
rect 25046 16288 25110 16292
rect 25126 16348 25190 16352
rect 25126 16292 25130 16348
rect 25130 16292 25186 16348
rect 25186 16292 25190 16348
rect 25126 16288 25190 16292
rect 9886 15804 9950 15808
rect 9886 15748 9890 15804
rect 9890 15748 9946 15804
rect 9946 15748 9950 15804
rect 9886 15744 9950 15748
rect 9966 15804 10030 15808
rect 9966 15748 9970 15804
rect 9970 15748 10026 15804
rect 10026 15748 10030 15804
rect 9966 15744 10030 15748
rect 10046 15804 10110 15808
rect 10046 15748 10050 15804
rect 10050 15748 10106 15804
rect 10106 15748 10110 15804
rect 10046 15744 10110 15748
rect 10126 15804 10190 15808
rect 10126 15748 10130 15804
rect 10130 15748 10186 15804
rect 10186 15748 10190 15804
rect 10126 15744 10190 15748
rect 19886 15804 19950 15808
rect 19886 15748 19890 15804
rect 19890 15748 19946 15804
rect 19946 15748 19950 15804
rect 19886 15744 19950 15748
rect 19966 15804 20030 15808
rect 19966 15748 19970 15804
rect 19970 15748 20026 15804
rect 20026 15748 20030 15804
rect 19966 15744 20030 15748
rect 20046 15804 20110 15808
rect 20046 15748 20050 15804
rect 20050 15748 20106 15804
rect 20106 15748 20110 15804
rect 20046 15744 20110 15748
rect 20126 15804 20190 15808
rect 20126 15748 20130 15804
rect 20130 15748 20186 15804
rect 20186 15748 20190 15804
rect 20126 15744 20190 15748
rect 4886 15260 4950 15264
rect 4886 15204 4890 15260
rect 4890 15204 4946 15260
rect 4946 15204 4950 15260
rect 4886 15200 4950 15204
rect 4966 15260 5030 15264
rect 4966 15204 4970 15260
rect 4970 15204 5026 15260
rect 5026 15204 5030 15260
rect 4966 15200 5030 15204
rect 5046 15260 5110 15264
rect 5046 15204 5050 15260
rect 5050 15204 5106 15260
rect 5106 15204 5110 15260
rect 5046 15200 5110 15204
rect 5126 15260 5190 15264
rect 5126 15204 5130 15260
rect 5130 15204 5186 15260
rect 5186 15204 5190 15260
rect 5126 15200 5190 15204
rect 14886 15260 14950 15264
rect 14886 15204 14890 15260
rect 14890 15204 14946 15260
rect 14946 15204 14950 15260
rect 14886 15200 14950 15204
rect 14966 15260 15030 15264
rect 14966 15204 14970 15260
rect 14970 15204 15026 15260
rect 15026 15204 15030 15260
rect 14966 15200 15030 15204
rect 15046 15260 15110 15264
rect 15046 15204 15050 15260
rect 15050 15204 15106 15260
rect 15106 15204 15110 15260
rect 15046 15200 15110 15204
rect 15126 15260 15190 15264
rect 15126 15204 15130 15260
rect 15130 15204 15186 15260
rect 15186 15204 15190 15260
rect 15126 15200 15190 15204
rect 24886 15260 24950 15264
rect 24886 15204 24890 15260
rect 24890 15204 24946 15260
rect 24946 15204 24950 15260
rect 24886 15200 24950 15204
rect 24966 15260 25030 15264
rect 24966 15204 24970 15260
rect 24970 15204 25026 15260
rect 25026 15204 25030 15260
rect 24966 15200 25030 15204
rect 25046 15260 25110 15264
rect 25046 15204 25050 15260
rect 25050 15204 25106 15260
rect 25106 15204 25110 15260
rect 25046 15200 25110 15204
rect 25126 15260 25190 15264
rect 25126 15204 25130 15260
rect 25130 15204 25186 15260
rect 25186 15204 25190 15260
rect 25126 15200 25190 15204
rect 9886 14716 9950 14720
rect 9886 14660 9890 14716
rect 9890 14660 9946 14716
rect 9946 14660 9950 14716
rect 9886 14656 9950 14660
rect 9966 14716 10030 14720
rect 9966 14660 9970 14716
rect 9970 14660 10026 14716
rect 10026 14660 10030 14716
rect 9966 14656 10030 14660
rect 10046 14716 10110 14720
rect 10046 14660 10050 14716
rect 10050 14660 10106 14716
rect 10106 14660 10110 14716
rect 10046 14656 10110 14660
rect 10126 14716 10190 14720
rect 10126 14660 10130 14716
rect 10130 14660 10186 14716
rect 10186 14660 10190 14716
rect 10126 14656 10190 14660
rect 19886 14716 19950 14720
rect 19886 14660 19890 14716
rect 19890 14660 19946 14716
rect 19946 14660 19950 14716
rect 19886 14656 19950 14660
rect 19966 14716 20030 14720
rect 19966 14660 19970 14716
rect 19970 14660 20026 14716
rect 20026 14660 20030 14716
rect 19966 14656 20030 14660
rect 20046 14716 20110 14720
rect 20046 14660 20050 14716
rect 20050 14660 20106 14716
rect 20106 14660 20110 14716
rect 20046 14656 20110 14660
rect 20126 14716 20190 14720
rect 20126 14660 20130 14716
rect 20130 14660 20186 14716
rect 20186 14660 20190 14716
rect 20126 14656 20190 14660
rect 4886 14172 4950 14176
rect 4886 14116 4890 14172
rect 4890 14116 4946 14172
rect 4946 14116 4950 14172
rect 4886 14112 4950 14116
rect 4966 14172 5030 14176
rect 4966 14116 4970 14172
rect 4970 14116 5026 14172
rect 5026 14116 5030 14172
rect 4966 14112 5030 14116
rect 5046 14172 5110 14176
rect 5046 14116 5050 14172
rect 5050 14116 5106 14172
rect 5106 14116 5110 14172
rect 5046 14112 5110 14116
rect 5126 14172 5190 14176
rect 5126 14116 5130 14172
rect 5130 14116 5186 14172
rect 5186 14116 5190 14172
rect 5126 14112 5190 14116
rect 14886 14172 14950 14176
rect 14886 14116 14890 14172
rect 14890 14116 14946 14172
rect 14946 14116 14950 14172
rect 14886 14112 14950 14116
rect 14966 14172 15030 14176
rect 14966 14116 14970 14172
rect 14970 14116 15026 14172
rect 15026 14116 15030 14172
rect 14966 14112 15030 14116
rect 15046 14172 15110 14176
rect 15046 14116 15050 14172
rect 15050 14116 15106 14172
rect 15106 14116 15110 14172
rect 15046 14112 15110 14116
rect 15126 14172 15190 14176
rect 15126 14116 15130 14172
rect 15130 14116 15186 14172
rect 15186 14116 15190 14172
rect 15126 14112 15190 14116
rect 24886 14172 24950 14176
rect 24886 14116 24890 14172
rect 24890 14116 24946 14172
rect 24946 14116 24950 14172
rect 24886 14112 24950 14116
rect 24966 14172 25030 14176
rect 24966 14116 24970 14172
rect 24970 14116 25026 14172
rect 25026 14116 25030 14172
rect 24966 14112 25030 14116
rect 25046 14172 25110 14176
rect 25046 14116 25050 14172
rect 25050 14116 25106 14172
rect 25106 14116 25110 14172
rect 25046 14112 25110 14116
rect 25126 14172 25190 14176
rect 25126 14116 25130 14172
rect 25130 14116 25186 14172
rect 25186 14116 25190 14172
rect 25126 14112 25190 14116
rect 9886 13628 9950 13632
rect 9886 13572 9890 13628
rect 9890 13572 9946 13628
rect 9946 13572 9950 13628
rect 9886 13568 9950 13572
rect 9966 13628 10030 13632
rect 9966 13572 9970 13628
rect 9970 13572 10026 13628
rect 10026 13572 10030 13628
rect 9966 13568 10030 13572
rect 10046 13628 10110 13632
rect 10046 13572 10050 13628
rect 10050 13572 10106 13628
rect 10106 13572 10110 13628
rect 10046 13568 10110 13572
rect 10126 13628 10190 13632
rect 10126 13572 10130 13628
rect 10130 13572 10186 13628
rect 10186 13572 10190 13628
rect 10126 13568 10190 13572
rect 19886 13628 19950 13632
rect 19886 13572 19890 13628
rect 19890 13572 19946 13628
rect 19946 13572 19950 13628
rect 19886 13568 19950 13572
rect 19966 13628 20030 13632
rect 19966 13572 19970 13628
rect 19970 13572 20026 13628
rect 20026 13572 20030 13628
rect 19966 13568 20030 13572
rect 20046 13628 20110 13632
rect 20046 13572 20050 13628
rect 20050 13572 20106 13628
rect 20106 13572 20110 13628
rect 20046 13568 20110 13572
rect 20126 13628 20190 13632
rect 20126 13572 20130 13628
rect 20130 13572 20186 13628
rect 20186 13572 20190 13628
rect 20126 13568 20190 13572
rect 4886 13084 4950 13088
rect 4886 13028 4890 13084
rect 4890 13028 4946 13084
rect 4946 13028 4950 13084
rect 4886 13024 4950 13028
rect 4966 13084 5030 13088
rect 4966 13028 4970 13084
rect 4970 13028 5026 13084
rect 5026 13028 5030 13084
rect 4966 13024 5030 13028
rect 5046 13084 5110 13088
rect 5046 13028 5050 13084
rect 5050 13028 5106 13084
rect 5106 13028 5110 13084
rect 5046 13024 5110 13028
rect 5126 13084 5190 13088
rect 5126 13028 5130 13084
rect 5130 13028 5186 13084
rect 5186 13028 5190 13084
rect 5126 13024 5190 13028
rect 14886 13084 14950 13088
rect 14886 13028 14890 13084
rect 14890 13028 14946 13084
rect 14946 13028 14950 13084
rect 14886 13024 14950 13028
rect 14966 13084 15030 13088
rect 14966 13028 14970 13084
rect 14970 13028 15026 13084
rect 15026 13028 15030 13084
rect 14966 13024 15030 13028
rect 15046 13084 15110 13088
rect 15046 13028 15050 13084
rect 15050 13028 15106 13084
rect 15106 13028 15110 13084
rect 15046 13024 15110 13028
rect 15126 13084 15190 13088
rect 15126 13028 15130 13084
rect 15130 13028 15186 13084
rect 15186 13028 15190 13084
rect 15126 13024 15190 13028
rect 24886 13084 24950 13088
rect 24886 13028 24890 13084
rect 24890 13028 24946 13084
rect 24946 13028 24950 13084
rect 24886 13024 24950 13028
rect 24966 13084 25030 13088
rect 24966 13028 24970 13084
rect 24970 13028 25026 13084
rect 25026 13028 25030 13084
rect 24966 13024 25030 13028
rect 25046 13084 25110 13088
rect 25046 13028 25050 13084
rect 25050 13028 25106 13084
rect 25106 13028 25110 13084
rect 25046 13024 25110 13028
rect 25126 13084 25190 13088
rect 25126 13028 25130 13084
rect 25130 13028 25186 13084
rect 25186 13028 25190 13084
rect 25126 13024 25190 13028
rect 9886 12540 9950 12544
rect 9886 12484 9890 12540
rect 9890 12484 9946 12540
rect 9946 12484 9950 12540
rect 9886 12480 9950 12484
rect 9966 12540 10030 12544
rect 9966 12484 9970 12540
rect 9970 12484 10026 12540
rect 10026 12484 10030 12540
rect 9966 12480 10030 12484
rect 10046 12540 10110 12544
rect 10046 12484 10050 12540
rect 10050 12484 10106 12540
rect 10106 12484 10110 12540
rect 10046 12480 10110 12484
rect 10126 12540 10190 12544
rect 10126 12484 10130 12540
rect 10130 12484 10186 12540
rect 10186 12484 10190 12540
rect 10126 12480 10190 12484
rect 19886 12540 19950 12544
rect 19886 12484 19890 12540
rect 19890 12484 19946 12540
rect 19946 12484 19950 12540
rect 19886 12480 19950 12484
rect 19966 12540 20030 12544
rect 19966 12484 19970 12540
rect 19970 12484 20026 12540
rect 20026 12484 20030 12540
rect 19966 12480 20030 12484
rect 20046 12540 20110 12544
rect 20046 12484 20050 12540
rect 20050 12484 20106 12540
rect 20106 12484 20110 12540
rect 20046 12480 20110 12484
rect 20126 12540 20190 12544
rect 20126 12484 20130 12540
rect 20130 12484 20186 12540
rect 20186 12484 20190 12540
rect 20126 12480 20190 12484
rect 4886 11996 4950 12000
rect 4886 11940 4890 11996
rect 4890 11940 4946 11996
rect 4946 11940 4950 11996
rect 4886 11936 4950 11940
rect 4966 11996 5030 12000
rect 4966 11940 4970 11996
rect 4970 11940 5026 11996
rect 5026 11940 5030 11996
rect 4966 11936 5030 11940
rect 5046 11996 5110 12000
rect 5046 11940 5050 11996
rect 5050 11940 5106 11996
rect 5106 11940 5110 11996
rect 5046 11936 5110 11940
rect 5126 11996 5190 12000
rect 5126 11940 5130 11996
rect 5130 11940 5186 11996
rect 5186 11940 5190 11996
rect 5126 11936 5190 11940
rect 14886 11996 14950 12000
rect 14886 11940 14890 11996
rect 14890 11940 14946 11996
rect 14946 11940 14950 11996
rect 14886 11936 14950 11940
rect 14966 11996 15030 12000
rect 14966 11940 14970 11996
rect 14970 11940 15026 11996
rect 15026 11940 15030 11996
rect 14966 11936 15030 11940
rect 15046 11996 15110 12000
rect 15046 11940 15050 11996
rect 15050 11940 15106 11996
rect 15106 11940 15110 11996
rect 15046 11936 15110 11940
rect 15126 11996 15190 12000
rect 15126 11940 15130 11996
rect 15130 11940 15186 11996
rect 15186 11940 15190 11996
rect 15126 11936 15190 11940
rect 24886 11996 24950 12000
rect 24886 11940 24890 11996
rect 24890 11940 24946 11996
rect 24946 11940 24950 11996
rect 24886 11936 24950 11940
rect 24966 11996 25030 12000
rect 24966 11940 24970 11996
rect 24970 11940 25026 11996
rect 25026 11940 25030 11996
rect 24966 11936 25030 11940
rect 25046 11996 25110 12000
rect 25046 11940 25050 11996
rect 25050 11940 25106 11996
rect 25106 11940 25110 11996
rect 25046 11936 25110 11940
rect 25126 11996 25190 12000
rect 25126 11940 25130 11996
rect 25130 11940 25186 11996
rect 25186 11940 25190 11996
rect 25126 11936 25190 11940
rect 9886 11452 9950 11456
rect 9886 11396 9890 11452
rect 9890 11396 9946 11452
rect 9946 11396 9950 11452
rect 9886 11392 9950 11396
rect 9966 11452 10030 11456
rect 9966 11396 9970 11452
rect 9970 11396 10026 11452
rect 10026 11396 10030 11452
rect 9966 11392 10030 11396
rect 10046 11452 10110 11456
rect 10046 11396 10050 11452
rect 10050 11396 10106 11452
rect 10106 11396 10110 11452
rect 10046 11392 10110 11396
rect 10126 11452 10190 11456
rect 10126 11396 10130 11452
rect 10130 11396 10186 11452
rect 10186 11396 10190 11452
rect 10126 11392 10190 11396
rect 19886 11452 19950 11456
rect 19886 11396 19890 11452
rect 19890 11396 19946 11452
rect 19946 11396 19950 11452
rect 19886 11392 19950 11396
rect 19966 11452 20030 11456
rect 19966 11396 19970 11452
rect 19970 11396 20026 11452
rect 20026 11396 20030 11452
rect 19966 11392 20030 11396
rect 20046 11452 20110 11456
rect 20046 11396 20050 11452
rect 20050 11396 20106 11452
rect 20106 11396 20110 11452
rect 20046 11392 20110 11396
rect 20126 11452 20190 11456
rect 20126 11396 20130 11452
rect 20130 11396 20186 11452
rect 20186 11396 20190 11452
rect 20126 11392 20190 11396
rect 4886 10908 4950 10912
rect 4886 10852 4890 10908
rect 4890 10852 4946 10908
rect 4946 10852 4950 10908
rect 4886 10848 4950 10852
rect 4966 10908 5030 10912
rect 4966 10852 4970 10908
rect 4970 10852 5026 10908
rect 5026 10852 5030 10908
rect 4966 10848 5030 10852
rect 5046 10908 5110 10912
rect 5046 10852 5050 10908
rect 5050 10852 5106 10908
rect 5106 10852 5110 10908
rect 5046 10848 5110 10852
rect 5126 10908 5190 10912
rect 5126 10852 5130 10908
rect 5130 10852 5186 10908
rect 5186 10852 5190 10908
rect 5126 10848 5190 10852
rect 14886 10908 14950 10912
rect 14886 10852 14890 10908
rect 14890 10852 14946 10908
rect 14946 10852 14950 10908
rect 14886 10848 14950 10852
rect 14966 10908 15030 10912
rect 14966 10852 14970 10908
rect 14970 10852 15026 10908
rect 15026 10852 15030 10908
rect 14966 10848 15030 10852
rect 15046 10908 15110 10912
rect 15046 10852 15050 10908
rect 15050 10852 15106 10908
rect 15106 10852 15110 10908
rect 15046 10848 15110 10852
rect 15126 10908 15190 10912
rect 15126 10852 15130 10908
rect 15130 10852 15186 10908
rect 15186 10852 15190 10908
rect 15126 10848 15190 10852
rect 24886 10908 24950 10912
rect 24886 10852 24890 10908
rect 24890 10852 24946 10908
rect 24946 10852 24950 10908
rect 24886 10848 24950 10852
rect 24966 10908 25030 10912
rect 24966 10852 24970 10908
rect 24970 10852 25026 10908
rect 25026 10852 25030 10908
rect 24966 10848 25030 10852
rect 25046 10908 25110 10912
rect 25046 10852 25050 10908
rect 25050 10852 25106 10908
rect 25106 10852 25110 10908
rect 25046 10848 25110 10852
rect 25126 10908 25190 10912
rect 25126 10852 25130 10908
rect 25130 10852 25186 10908
rect 25186 10852 25190 10908
rect 25126 10848 25190 10852
rect 9886 10364 9950 10368
rect 9886 10308 9890 10364
rect 9890 10308 9946 10364
rect 9946 10308 9950 10364
rect 9886 10304 9950 10308
rect 9966 10364 10030 10368
rect 9966 10308 9970 10364
rect 9970 10308 10026 10364
rect 10026 10308 10030 10364
rect 9966 10304 10030 10308
rect 10046 10364 10110 10368
rect 10046 10308 10050 10364
rect 10050 10308 10106 10364
rect 10106 10308 10110 10364
rect 10046 10304 10110 10308
rect 10126 10364 10190 10368
rect 10126 10308 10130 10364
rect 10130 10308 10186 10364
rect 10186 10308 10190 10364
rect 10126 10304 10190 10308
rect 19886 10364 19950 10368
rect 19886 10308 19890 10364
rect 19890 10308 19946 10364
rect 19946 10308 19950 10364
rect 19886 10304 19950 10308
rect 19966 10364 20030 10368
rect 19966 10308 19970 10364
rect 19970 10308 20026 10364
rect 20026 10308 20030 10364
rect 19966 10304 20030 10308
rect 20046 10364 20110 10368
rect 20046 10308 20050 10364
rect 20050 10308 20106 10364
rect 20106 10308 20110 10364
rect 20046 10304 20110 10308
rect 20126 10364 20190 10368
rect 20126 10308 20130 10364
rect 20130 10308 20186 10364
rect 20186 10308 20190 10364
rect 20126 10304 20190 10308
rect 4886 9820 4950 9824
rect 4886 9764 4890 9820
rect 4890 9764 4946 9820
rect 4946 9764 4950 9820
rect 4886 9760 4950 9764
rect 4966 9820 5030 9824
rect 4966 9764 4970 9820
rect 4970 9764 5026 9820
rect 5026 9764 5030 9820
rect 4966 9760 5030 9764
rect 5046 9820 5110 9824
rect 5046 9764 5050 9820
rect 5050 9764 5106 9820
rect 5106 9764 5110 9820
rect 5046 9760 5110 9764
rect 5126 9820 5190 9824
rect 5126 9764 5130 9820
rect 5130 9764 5186 9820
rect 5186 9764 5190 9820
rect 5126 9760 5190 9764
rect 14886 9820 14950 9824
rect 14886 9764 14890 9820
rect 14890 9764 14946 9820
rect 14946 9764 14950 9820
rect 14886 9760 14950 9764
rect 14966 9820 15030 9824
rect 14966 9764 14970 9820
rect 14970 9764 15026 9820
rect 15026 9764 15030 9820
rect 14966 9760 15030 9764
rect 15046 9820 15110 9824
rect 15046 9764 15050 9820
rect 15050 9764 15106 9820
rect 15106 9764 15110 9820
rect 15046 9760 15110 9764
rect 15126 9820 15190 9824
rect 15126 9764 15130 9820
rect 15130 9764 15186 9820
rect 15186 9764 15190 9820
rect 15126 9760 15190 9764
rect 24886 9820 24950 9824
rect 24886 9764 24890 9820
rect 24890 9764 24946 9820
rect 24946 9764 24950 9820
rect 24886 9760 24950 9764
rect 24966 9820 25030 9824
rect 24966 9764 24970 9820
rect 24970 9764 25026 9820
rect 25026 9764 25030 9820
rect 24966 9760 25030 9764
rect 25046 9820 25110 9824
rect 25046 9764 25050 9820
rect 25050 9764 25106 9820
rect 25106 9764 25110 9820
rect 25046 9760 25110 9764
rect 25126 9820 25190 9824
rect 25126 9764 25130 9820
rect 25130 9764 25186 9820
rect 25186 9764 25190 9820
rect 25126 9760 25190 9764
rect 9886 9276 9950 9280
rect 9886 9220 9890 9276
rect 9890 9220 9946 9276
rect 9946 9220 9950 9276
rect 9886 9216 9950 9220
rect 9966 9276 10030 9280
rect 9966 9220 9970 9276
rect 9970 9220 10026 9276
rect 10026 9220 10030 9276
rect 9966 9216 10030 9220
rect 10046 9276 10110 9280
rect 10046 9220 10050 9276
rect 10050 9220 10106 9276
rect 10106 9220 10110 9276
rect 10046 9216 10110 9220
rect 10126 9276 10190 9280
rect 10126 9220 10130 9276
rect 10130 9220 10186 9276
rect 10186 9220 10190 9276
rect 10126 9216 10190 9220
rect 19886 9276 19950 9280
rect 19886 9220 19890 9276
rect 19890 9220 19946 9276
rect 19946 9220 19950 9276
rect 19886 9216 19950 9220
rect 19966 9276 20030 9280
rect 19966 9220 19970 9276
rect 19970 9220 20026 9276
rect 20026 9220 20030 9276
rect 19966 9216 20030 9220
rect 20046 9276 20110 9280
rect 20046 9220 20050 9276
rect 20050 9220 20106 9276
rect 20106 9220 20110 9276
rect 20046 9216 20110 9220
rect 20126 9276 20190 9280
rect 20126 9220 20130 9276
rect 20130 9220 20186 9276
rect 20186 9220 20190 9276
rect 20126 9216 20190 9220
rect 4886 8732 4950 8736
rect 4886 8676 4890 8732
rect 4890 8676 4946 8732
rect 4946 8676 4950 8732
rect 4886 8672 4950 8676
rect 4966 8732 5030 8736
rect 4966 8676 4970 8732
rect 4970 8676 5026 8732
rect 5026 8676 5030 8732
rect 4966 8672 5030 8676
rect 5046 8732 5110 8736
rect 5046 8676 5050 8732
rect 5050 8676 5106 8732
rect 5106 8676 5110 8732
rect 5046 8672 5110 8676
rect 5126 8732 5190 8736
rect 5126 8676 5130 8732
rect 5130 8676 5186 8732
rect 5186 8676 5190 8732
rect 5126 8672 5190 8676
rect 14886 8732 14950 8736
rect 14886 8676 14890 8732
rect 14890 8676 14946 8732
rect 14946 8676 14950 8732
rect 14886 8672 14950 8676
rect 14966 8732 15030 8736
rect 14966 8676 14970 8732
rect 14970 8676 15026 8732
rect 15026 8676 15030 8732
rect 14966 8672 15030 8676
rect 15046 8732 15110 8736
rect 15046 8676 15050 8732
rect 15050 8676 15106 8732
rect 15106 8676 15110 8732
rect 15046 8672 15110 8676
rect 15126 8732 15190 8736
rect 15126 8676 15130 8732
rect 15130 8676 15186 8732
rect 15186 8676 15190 8732
rect 15126 8672 15190 8676
rect 24886 8732 24950 8736
rect 24886 8676 24890 8732
rect 24890 8676 24946 8732
rect 24946 8676 24950 8732
rect 24886 8672 24950 8676
rect 24966 8732 25030 8736
rect 24966 8676 24970 8732
rect 24970 8676 25026 8732
rect 25026 8676 25030 8732
rect 24966 8672 25030 8676
rect 25046 8732 25110 8736
rect 25046 8676 25050 8732
rect 25050 8676 25106 8732
rect 25106 8676 25110 8732
rect 25046 8672 25110 8676
rect 25126 8732 25190 8736
rect 25126 8676 25130 8732
rect 25130 8676 25186 8732
rect 25186 8676 25190 8732
rect 25126 8672 25190 8676
rect 9886 8188 9950 8192
rect 9886 8132 9890 8188
rect 9890 8132 9946 8188
rect 9946 8132 9950 8188
rect 9886 8128 9950 8132
rect 9966 8188 10030 8192
rect 9966 8132 9970 8188
rect 9970 8132 10026 8188
rect 10026 8132 10030 8188
rect 9966 8128 10030 8132
rect 10046 8188 10110 8192
rect 10046 8132 10050 8188
rect 10050 8132 10106 8188
rect 10106 8132 10110 8188
rect 10046 8128 10110 8132
rect 10126 8188 10190 8192
rect 10126 8132 10130 8188
rect 10130 8132 10186 8188
rect 10186 8132 10190 8188
rect 10126 8128 10190 8132
rect 19886 8188 19950 8192
rect 19886 8132 19890 8188
rect 19890 8132 19946 8188
rect 19946 8132 19950 8188
rect 19886 8128 19950 8132
rect 19966 8188 20030 8192
rect 19966 8132 19970 8188
rect 19970 8132 20026 8188
rect 20026 8132 20030 8188
rect 19966 8128 20030 8132
rect 20046 8188 20110 8192
rect 20046 8132 20050 8188
rect 20050 8132 20106 8188
rect 20106 8132 20110 8188
rect 20046 8128 20110 8132
rect 20126 8188 20190 8192
rect 20126 8132 20130 8188
rect 20130 8132 20186 8188
rect 20186 8132 20190 8188
rect 20126 8128 20190 8132
rect 4886 7644 4950 7648
rect 4886 7588 4890 7644
rect 4890 7588 4946 7644
rect 4946 7588 4950 7644
rect 4886 7584 4950 7588
rect 4966 7644 5030 7648
rect 4966 7588 4970 7644
rect 4970 7588 5026 7644
rect 5026 7588 5030 7644
rect 4966 7584 5030 7588
rect 5046 7644 5110 7648
rect 5046 7588 5050 7644
rect 5050 7588 5106 7644
rect 5106 7588 5110 7644
rect 5046 7584 5110 7588
rect 5126 7644 5190 7648
rect 5126 7588 5130 7644
rect 5130 7588 5186 7644
rect 5186 7588 5190 7644
rect 5126 7584 5190 7588
rect 14886 7644 14950 7648
rect 14886 7588 14890 7644
rect 14890 7588 14946 7644
rect 14946 7588 14950 7644
rect 14886 7584 14950 7588
rect 14966 7644 15030 7648
rect 14966 7588 14970 7644
rect 14970 7588 15026 7644
rect 15026 7588 15030 7644
rect 14966 7584 15030 7588
rect 15046 7644 15110 7648
rect 15046 7588 15050 7644
rect 15050 7588 15106 7644
rect 15106 7588 15110 7644
rect 15046 7584 15110 7588
rect 15126 7644 15190 7648
rect 15126 7588 15130 7644
rect 15130 7588 15186 7644
rect 15186 7588 15190 7644
rect 15126 7584 15190 7588
rect 24886 7644 24950 7648
rect 24886 7588 24890 7644
rect 24890 7588 24946 7644
rect 24946 7588 24950 7644
rect 24886 7584 24950 7588
rect 24966 7644 25030 7648
rect 24966 7588 24970 7644
rect 24970 7588 25026 7644
rect 25026 7588 25030 7644
rect 24966 7584 25030 7588
rect 25046 7644 25110 7648
rect 25046 7588 25050 7644
rect 25050 7588 25106 7644
rect 25106 7588 25110 7644
rect 25046 7584 25110 7588
rect 25126 7644 25190 7648
rect 25126 7588 25130 7644
rect 25130 7588 25186 7644
rect 25186 7588 25190 7644
rect 25126 7584 25190 7588
rect 9886 7100 9950 7104
rect 9886 7044 9890 7100
rect 9890 7044 9946 7100
rect 9946 7044 9950 7100
rect 9886 7040 9950 7044
rect 9966 7100 10030 7104
rect 9966 7044 9970 7100
rect 9970 7044 10026 7100
rect 10026 7044 10030 7100
rect 9966 7040 10030 7044
rect 10046 7100 10110 7104
rect 10046 7044 10050 7100
rect 10050 7044 10106 7100
rect 10106 7044 10110 7100
rect 10046 7040 10110 7044
rect 10126 7100 10190 7104
rect 10126 7044 10130 7100
rect 10130 7044 10186 7100
rect 10186 7044 10190 7100
rect 10126 7040 10190 7044
rect 19886 7100 19950 7104
rect 19886 7044 19890 7100
rect 19890 7044 19946 7100
rect 19946 7044 19950 7100
rect 19886 7040 19950 7044
rect 19966 7100 20030 7104
rect 19966 7044 19970 7100
rect 19970 7044 20026 7100
rect 20026 7044 20030 7100
rect 19966 7040 20030 7044
rect 20046 7100 20110 7104
rect 20046 7044 20050 7100
rect 20050 7044 20106 7100
rect 20106 7044 20110 7100
rect 20046 7040 20110 7044
rect 20126 7100 20190 7104
rect 20126 7044 20130 7100
rect 20130 7044 20186 7100
rect 20186 7044 20190 7100
rect 20126 7040 20190 7044
rect 4886 6556 4950 6560
rect 4886 6500 4890 6556
rect 4890 6500 4946 6556
rect 4946 6500 4950 6556
rect 4886 6496 4950 6500
rect 4966 6556 5030 6560
rect 4966 6500 4970 6556
rect 4970 6500 5026 6556
rect 5026 6500 5030 6556
rect 4966 6496 5030 6500
rect 5046 6556 5110 6560
rect 5046 6500 5050 6556
rect 5050 6500 5106 6556
rect 5106 6500 5110 6556
rect 5046 6496 5110 6500
rect 5126 6556 5190 6560
rect 5126 6500 5130 6556
rect 5130 6500 5186 6556
rect 5186 6500 5190 6556
rect 5126 6496 5190 6500
rect 14886 6556 14950 6560
rect 14886 6500 14890 6556
rect 14890 6500 14946 6556
rect 14946 6500 14950 6556
rect 14886 6496 14950 6500
rect 14966 6556 15030 6560
rect 14966 6500 14970 6556
rect 14970 6500 15026 6556
rect 15026 6500 15030 6556
rect 14966 6496 15030 6500
rect 15046 6556 15110 6560
rect 15046 6500 15050 6556
rect 15050 6500 15106 6556
rect 15106 6500 15110 6556
rect 15046 6496 15110 6500
rect 15126 6556 15190 6560
rect 15126 6500 15130 6556
rect 15130 6500 15186 6556
rect 15186 6500 15190 6556
rect 15126 6496 15190 6500
rect 24886 6556 24950 6560
rect 24886 6500 24890 6556
rect 24890 6500 24946 6556
rect 24946 6500 24950 6556
rect 24886 6496 24950 6500
rect 24966 6556 25030 6560
rect 24966 6500 24970 6556
rect 24970 6500 25026 6556
rect 25026 6500 25030 6556
rect 24966 6496 25030 6500
rect 25046 6556 25110 6560
rect 25046 6500 25050 6556
rect 25050 6500 25106 6556
rect 25106 6500 25110 6556
rect 25046 6496 25110 6500
rect 25126 6556 25190 6560
rect 25126 6500 25130 6556
rect 25130 6500 25186 6556
rect 25186 6500 25190 6556
rect 25126 6496 25190 6500
rect 9886 6012 9950 6016
rect 9886 5956 9890 6012
rect 9890 5956 9946 6012
rect 9946 5956 9950 6012
rect 9886 5952 9950 5956
rect 9966 6012 10030 6016
rect 9966 5956 9970 6012
rect 9970 5956 10026 6012
rect 10026 5956 10030 6012
rect 9966 5952 10030 5956
rect 10046 6012 10110 6016
rect 10046 5956 10050 6012
rect 10050 5956 10106 6012
rect 10106 5956 10110 6012
rect 10046 5952 10110 5956
rect 10126 6012 10190 6016
rect 10126 5956 10130 6012
rect 10130 5956 10186 6012
rect 10186 5956 10190 6012
rect 10126 5952 10190 5956
rect 19886 6012 19950 6016
rect 19886 5956 19890 6012
rect 19890 5956 19946 6012
rect 19946 5956 19950 6012
rect 19886 5952 19950 5956
rect 19966 6012 20030 6016
rect 19966 5956 19970 6012
rect 19970 5956 20026 6012
rect 20026 5956 20030 6012
rect 19966 5952 20030 5956
rect 20046 6012 20110 6016
rect 20046 5956 20050 6012
rect 20050 5956 20106 6012
rect 20106 5956 20110 6012
rect 20046 5952 20110 5956
rect 20126 6012 20190 6016
rect 20126 5956 20130 6012
rect 20130 5956 20186 6012
rect 20186 5956 20190 6012
rect 20126 5952 20190 5956
rect 4886 5468 4950 5472
rect 4886 5412 4890 5468
rect 4890 5412 4946 5468
rect 4946 5412 4950 5468
rect 4886 5408 4950 5412
rect 4966 5468 5030 5472
rect 4966 5412 4970 5468
rect 4970 5412 5026 5468
rect 5026 5412 5030 5468
rect 4966 5408 5030 5412
rect 5046 5468 5110 5472
rect 5046 5412 5050 5468
rect 5050 5412 5106 5468
rect 5106 5412 5110 5468
rect 5046 5408 5110 5412
rect 5126 5468 5190 5472
rect 5126 5412 5130 5468
rect 5130 5412 5186 5468
rect 5186 5412 5190 5468
rect 5126 5408 5190 5412
rect 14886 5468 14950 5472
rect 14886 5412 14890 5468
rect 14890 5412 14946 5468
rect 14946 5412 14950 5468
rect 14886 5408 14950 5412
rect 14966 5468 15030 5472
rect 14966 5412 14970 5468
rect 14970 5412 15026 5468
rect 15026 5412 15030 5468
rect 14966 5408 15030 5412
rect 15046 5468 15110 5472
rect 15046 5412 15050 5468
rect 15050 5412 15106 5468
rect 15106 5412 15110 5468
rect 15046 5408 15110 5412
rect 15126 5468 15190 5472
rect 15126 5412 15130 5468
rect 15130 5412 15186 5468
rect 15186 5412 15190 5468
rect 15126 5408 15190 5412
rect 24886 5468 24950 5472
rect 24886 5412 24890 5468
rect 24890 5412 24946 5468
rect 24946 5412 24950 5468
rect 24886 5408 24950 5412
rect 24966 5468 25030 5472
rect 24966 5412 24970 5468
rect 24970 5412 25026 5468
rect 25026 5412 25030 5468
rect 24966 5408 25030 5412
rect 25046 5468 25110 5472
rect 25046 5412 25050 5468
rect 25050 5412 25106 5468
rect 25106 5412 25110 5468
rect 25046 5408 25110 5412
rect 25126 5468 25190 5472
rect 25126 5412 25130 5468
rect 25130 5412 25186 5468
rect 25186 5412 25190 5468
rect 25126 5408 25190 5412
rect 9886 4924 9950 4928
rect 9886 4868 9890 4924
rect 9890 4868 9946 4924
rect 9946 4868 9950 4924
rect 9886 4864 9950 4868
rect 9966 4924 10030 4928
rect 9966 4868 9970 4924
rect 9970 4868 10026 4924
rect 10026 4868 10030 4924
rect 9966 4864 10030 4868
rect 10046 4924 10110 4928
rect 10046 4868 10050 4924
rect 10050 4868 10106 4924
rect 10106 4868 10110 4924
rect 10046 4864 10110 4868
rect 10126 4924 10190 4928
rect 10126 4868 10130 4924
rect 10130 4868 10186 4924
rect 10186 4868 10190 4924
rect 10126 4864 10190 4868
rect 19886 4924 19950 4928
rect 19886 4868 19890 4924
rect 19890 4868 19946 4924
rect 19946 4868 19950 4924
rect 19886 4864 19950 4868
rect 19966 4924 20030 4928
rect 19966 4868 19970 4924
rect 19970 4868 20026 4924
rect 20026 4868 20030 4924
rect 19966 4864 20030 4868
rect 20046 4924 20110 4928
rect 20046 4868 20050 4924
rect 20050 4868 20106 4924
rect 20106 4868 20110 4924
rect 20046 4864 20110 4868
rect 20126 4924 20190 4928
rect 20126 4868 20130 4924
rect 20130 4868 20186 4924
rect 20186 4868 20190 4924
rect 20126 4864 20190 4868
rect 4886 4380 4950 4384
rect 4886 4324 4890 4380
rect 4890 4324 4946 4380
rect 4946 4324 4950 4380
rect 4886 4320 4950 4324
rect 4966 4380 5030 4384
rect 4966 4324 4970 4380
rect 4970 4324 5026 4380
rect 5026 4324 5030 4380
rect 4966 4320 5030 4324
rect 5046 4380 5110 4384
rect 5046 4324 5050 4380
rect 5050 4324 5106 4380
rect 5106 4324 5110 4380
rect 5046 4320 5110 4324
rect 5126 4380 5190 4384
rect 5126 4324 5130 4380
rect 5130 4324 5186 4380
rect 5186 4324 5190 4380
rect 5126 4320 5190 4324
rect 14886 4380 14950 4384
rect 14886 4324 14890 4380
rect 14890 4324 14946 4380
rect 14946 4324 14950 4380
rect 14886 4320 14950 4324
rect 14966 4380 15030 4384
rect 14966 4324 14970 4380
rect 14970 4324 15026 4380
rect 15026 4324 15030 4380
rect 14966 4320 15030 4324
rect 15046 4380 15110 4384
rect 15046 4324 15050 4380
rect 15050 4324 15106 4380
rect 15106 4324 15110 4380
rect 15046 4320 15110 4324
rect 15126 4380 15190 4384
rect 15126 4324 15130 4380
rect 15130 4324 15186 4380
rect 15186 4324 15190 4380
rect 15126 4320 15190 4324
rect 24886 4380 24950 4384
rect 24886 4324 24890 4380
rect 24890 4324 24946 4380
rect 24946 4324 24950 4380
rect 24886 4320 24950 4324
rect 24966 4380 25030 4384
rect 24966 4324 24970 4380
rect 24970 4324 25026 4380
rect 25026 4324 25030 4380
rect 24966 4320 25030 4324
rect 25046 4380 25110 4384
rect 25046 4324 25050 4380
rect 25050 4324 25106 4380
rect 25106 4324 25110 4380
rect 25046 4320 25110 4324
rect 25126 4380 25190 4384
rect 25126 4324 25130 4380
rect 25130 4324 25186 4380
rect 25186 4324 25190 4380
rect 25126 4320 25190 4324
rect 9886 3836 9950 3840
rect 9886 3780 9890 3836
rect 9890 3780 9946 3836
rect 9946 3780 9950 3836
rect 9886 3776 9950 3780
rect 9966 3836 10030 3840
rect 9966 3780 9970 3836
rect 9970 3780 10026 3836
rect 10026 3780 10030 3836
rect 9966 3776 10030 3780
rect 10046 3836 10110 3840
rect 10046 3780 10050 3836
rect 10050 3780 10106 3836
rect 10106 3780 10110 3836
rect 10046 3776 10110 3780
rect 10126 3836 10190 3840
rect 10126 3780 10130 3836
rect 10130 3780 10186 3836
rect 10186 3780 10190 3836
rect 10126 3776 10190 3780
rect 19886 3836 19950 3840
rect 19886 3780 19890 3836
rect 19890 3780 19946 3836
rect 19946 3780 19950 3836
rect 19886 3776 19950 3780
rect 19966 3836 20030 3840
rect 19966 3780 19970 3836
rect 19970 3780 20026 3836
rect 20026 3780 20030 3836
rect 19966 3776 20030 3780
rect 20046 3836 20110 3840
rect 20046 3780 20050 3836
rect 20050 3780 20106 3836
rect 20106 3780 20110 3836
rect 20046 3776 20110 3780
rect 20126 3836 20190 3840
rect 20126 3780 20130 3836
rect 20130 3780 20186 3836
rect 20186 3780 20190 3836
rect 20126 3776 20190 3780
rect 4886 3292 4950 3296
rect 4886 3236 4890 3292
rect 4890 3236 4946 3292
rect 4946 3236 4950 3292
rect 4886 3232 4950 3236
rect 4966 3292 5030 3296
rect 4966 3236 4970 3292
rect 4970 3236 5026 3292
rect 5026 3236 5030 3292
rect 4966 3232 5030 3236
rect 5046 3292 5110 3296
rect 5046 3236 5050 3292
rect 5050 3236 5106 3292
rect 5106 3236 5110 3292
rect 5046 3232 5110 3236
rect 5126 3292 5190 3296
rect 5126 3236 5130 3292
rect 5130 3236 5186 3292
rect 5186 3236 5190 3292
rect 5126 3232 5190 3236
rect 14886 3292 14950 3296
rect 14886 3236 14890 3292
rect 14890 3236 14946 3292
rect 14946 3236 14950 3292
rect 14886 3232 14950 3236
rect 14966 3292 15030 3296
rect 14966 3236 14970 3292
rect 14970 3236 15026 3292
rect 15026 3236 15030 3292
rect 14966 3232 15030 3236
rect 15046 3292 15110 3296
rect 15046 3236 15050 3292
rect 15050 3236 15106 3292
rect 15106 3236 15110 3292
rect 15046 3232 15110 3236
rect 15126 3292 15190 3296
rect 15126 3236 15130 3292
rect 15130 3236 15186 3292
rect 15186 3236 15190 3292
rect 15126 3232 15190 3236
rect 24886 3292 24950 3296
rect 24886 3236 24890 3292
rect 24890 3236 24946 3292
rect 24946 3236 24950 3292
rect 24886 3232 24950 3236
rect 24966 3292 25030 3296
rect 24966 3236 24970 3292
rect 24970 3236 25026 3292
rect 25026 3236 25030 3292
rect 24966 3232 25030 3236
rect 25046 3292 25110 3296
rect 25046 3236 25050 3292
rect 25050 3236 25106 3292
rect 25106 3236 25110 3292
rect 25046 3232 25110 3236
rect 25126 3292 25190 3296
rect 25126 3236 25130 3292
rect 25130 3236 25186 3292
rect 25186 3236 25190 3292
rect 25126 3232 25190 3236
rect 9886 2748 9950 2752
rect 9886 2692 9890 2748
rect 9890 2692 9946 2748
rect 9946 2692 9950 2748
rect 9886 2688 9950 2692
rect 9966 2748 10030 2752
rect 9966 2692 9970 2748
rect 9970 2692 10026 2748
rect 10026 2692 10030 2748
rect 9966 2688 10030 2692
rect 10046 2748 10110 2752
rect 10046 2692 10050 2748
rect 10050 2692 10106 2748
rect 10106 2692 10110 2748
rect 10046 2688 10110 2692
rect 10126 2748 10190 2752
rect 10126 2692 10130 2748
rect 10130 2692 10186 2748
rect 10186 2692 10190 2748
rect 10126 2688 10190 2692
rect 19886 2748 19950 2752
rect 19886 2692 19890 2748
rect 19890 2692 19946 2748
rect 19946 2692 19950 2748
rect 19886 2688 19950 2692
rect 19966 2748 20030 2752
rect 19966 2692 19970 2748
rect 19970 2692 20026 2748
rect 20026 2692 20030 2748
rect 19966 2688 20030 2692
rect 20046 2748 20110 2752
rect 20046 2692 20050 2748
rect 20050 2692 20106 2748
rect 20106 2692 20110 2748
rect 20046 2688 20110 2692
rect 20126 2748 20190 2752
rect 20126 2692 20130 2748
rect 20130 2692 20186 2748
rect 20186 2692 20190 2748
rect 20126 2688 20190 2692
rect 4886 2204 4950 2208
rect 4886 2148 4890 2204
rect 4890 2148 4946 2204
rect 4946 2148 4950 2204
rect 4886 2144 4950 2148
rect 4966 2204 5030 2208
rect 4966 2148 4970 2204
rect 4970 2148 5026 2204
rect 5026 2148 5030 2204
rect 4966 2144 5030 2148
rect 5046 2204 5110 2208
rect 5046 2148 5050 2204
rect 5050 2148 5106 2204
rect 5106 2148 5110 2204
rect 5046 2144 5110 2148
rect 5126 2204 5190 2208
rect 5126 2148 5130 2204
rect 5130 2148 5186 2204
rect 5186 2148 5190 2204
rect 5126 2144 5190 2148
rect 14886 2204 14950 2208
rect 14886 2148 14890 2204
rect 14890 2148 14946 2204
rect 14946 2148 14950 2204
rect 14886 2144 14950 2148
rect 14966 2204 15030 2208
rect 14966 2148 14970 2204
rect 14970 2148 15026 2204
rect 15026 2148 15030 2204
rect 14966 2144 15030 2148
rect 15046 2204 15110 2208
rect 15046 2148 15050 2204
rect 15050 2148 15106 2204
rect 15106 2148 15110 2204
rect 15046 2144 15110 2148
rect 15126 2204 15190 2208
rect 15126 2148 15130 2204
rect 15130 2148 15186 2204
rect 15186 2148 15190 2204
rect 15126 2144 15190 2148
rect 24886 2204 24950 2208
rect 24886 2148 24890 2204
rect 24890 2148 24946 2204
rect 24946 2148 24950 2204
rect 24886 2144 24950 2148
rect 24966 2204 25030 2208
rect 24966 2148 24970 2204
rect 24970 2148 25026 2204
rect 25026 2148 25030 2204
rect 24966 2144 25030 2148
rect 25046 2204 25110 2208
rect 25046 2148 25050 2204
rect 25050 2148 25106 2204
rect 25106 2148 25110 2204
rect 25046 2144 25110 2148
rect 25126 2204 25190 2208
rect 25126 2148 25130 2204
rect 25130 2148 25186 2204
rect 25186 2148 25190 2204
rect 25126 2144 25190 2148
<< metal4 >>
rect 4878 21792 5198 21808
rect 4878 21728 4886 21792
rect 4950 21728 4966 21792
rect 5030 21728 5046 21792
rect 5110 21728 5126 21792
rect 5190 21728 5198 21792
rect 4878 20704 5198 21728
rect 4878 20640 4886 20704
rect 4950 20640 4966 20704
rect 5030 20640 5046 20704
rect 5110 20640 5126 20704
rect 5190 20640 5198 20704
rect 4878 19616 5198 20640
rect 4878 19552 4886 19616
rect 4950 19552 4966 19616
rect 5030 19552 5046 19616
rect 5110 19552 5126 19616
rect 5190 19552 5198 19616
rect 4878 18528 5198 19552
rect 4878 18464 4886 18528
rect 4950 18464 4966 18528
rect 5030 18464 5046 18528
rect 5110 18464 5126 18528
rect 5190 18464 5198 18528
rect 4878 17440 5198 18464
rect 4878 17376 4886 17440
rect 4950 17376 4966 17440
rect 5030 17376 5046 17440
rect 5110 17376 5126 17440
rect 5190 17376 5198 17440
rect 4878 16352 5198 17376
rect 4878 16288 4886 16352
rect 4950 16288 4966 16352
rect 5030 16288 5046 16352
rect 5110 16288 5126 16352
rect 5190 16288 5198 16352
rect 4878 15264 5198 16288
rect 4878 15200 4886 15264
rect 4950 15200 4966 15264
rect 5030 15200 5046 15264
rect 5110 15200 5126 15264
rect 5190 15200 5198 15264
rect 4878 14176 5198 15200
rect 4878 14112 4886 14176
rect 4950 14112 4966 14176
rect 5030 14112 5046 14176
rect 5110 14112 5126 14176
rect 5190 14112 5198 14176
rect 4878 13088 5198 14112
rect 4878 13024 4886 13088
rect 4950 13024 4966 13088
rect 5030 13024 5046 13088
rect 5110 13024 5126 13088
rect 5190 13024 5198 13088
rect 4878 12000 5198 13024
rect 4878 11936 4886 12000
rect 4950 11936 4966 12000
rect 5030 11936 5046 12000
rect 5110 11936 5126 12000
rect 5190 11936 5198 12000
rect 4878 10912 5198 11936
rect 4878 10848 4886 10912
rect 4950 10848 4966 10912
rect 5030 10848 5046 10912
rect 5110 10848 5126 10912
rect 5190 10848 5198 10912
rect 4878 9824 5198 10848
rect 4878 9760 4886 9824
rect 4950 9760 4966 9824
rect 5030 9760 5046 9824
rect 5110 9760 5126 9824
rect 5190 9760 5198 9824
rect 4878 8736 5198 9760
rect 4878 8672 4886 8736
rect 4950 8672 4966 8736
rect 5030 8672 5046 8736
rect 5110 8672 5126 8736
rect 5190 8672 5198 8736
rect 4878 7648 5198 8672
rect 4878 7584 4886 7648
rect 4950 7584 4966 7648
rect 5030 7584 5046 7648
rect 5110 7584 5126 7648
rect 5190 7584 5198 7648
rect 4878 6560 5198 7584
rect 4878 6496 4886 6560
rect 4950 6496 4966 6560
rect 5030 6496 5046 6560
rect 5110 6496 5126 6560
rect 5190 6496 5198 6560
rect 4878 5472 5198 6496
rect 4878 5408 4886 5472
rect 4950 5408 4966 5472
rect 5030 5408 5046 5472
rect 5110 5408 5126 5472
rect 5190 5408 5198 5472
rect 4878 4384 5198 5408
rect 4878 4320 4886 4384
rect 4950 4320 4966 4384
rect 5030 4320 5046 4384
rect 5110 4320 5126 4384
rect 5190 4320 5198 4384
rect 4878 3296 5198 4320
rect 4878 3232 4886 3296
rect 4950 3232 4966 3296
rect 5030 3232 5046 3296
rect 5110 3232 5126 3296
rect 5190 3232 5198 3296
rect 4878 2208 5198 3232
rect 4878 2144 4886 2208
rect 4950 2144 4966 2208
rect 5030 2144 5046 2208
rect 5110 2144 5126 2208
rect 5190 2144 5198 2208
rect 4878 2128 5198 2144
rect 9878 21248 10198 21808
rect 9878 21184 9886 21248
rect 9950 21184 9966 21248
rect 10030 21184 10046 21248
rect 10110 21184 10126 21248
rect 10190 21184 10198 21248
rect 9878 20160 10198 21184
rect 9878 20096 9886 20160
rect 9950 20096 9966 20160
rect 10030 20096 10046 20160
rect 10110 20096 10126 20160
rect 10190 20096 10198 20160
rect 9878 19072 10198 20096
rect 9878 19008 9886 19072
rect 9950 19008 9966 19072
rect 10030 19008 10046 19072
rect 10110 19008 10126 19072
rect 10190 19008 10198 19072
rect 9878 17984 10198 19008
rect 9878 17920 9886 17984
rect 9950 17920 9966 17984
rect 10030 17920 10046 17984
rect 10110 17920 10126 17984
rect 10190 17920 10198 17984
rect 9878 16896 10198 17920
rect 9878 16832 9886 16896
rect 9950 16832 9966 16896
rect 10030 16832 10046 16896
rect 10110 16832 10126 16896
rect 10190 16832 10198 16896
rect 9878 15808 10198 16832
rect 9878 15744 9886 15808
rect 9950 15744 9966 15808
rect 10030 15744 10046 15808
rect 10110 15744 10126 15808
rect 10190 15744 10198 15808
rect 9878 14720 10198 15744
rect 9878 14656 9886 14720
rect 9950 14656 9966 14720
rect 10030 14656 10046 14720
rect 10110 14656 10126 14720
rect 10190 14656 10198 14720
rect 9878 13632 10198 14656
rect 9878 13568 9886 13632
rect 9950 13568 9966 13632
rect 10030 13568 10046 13632
rect 10110 13568 10126 13632
rect 10190 13568 10198 13632
rect 9878 12544 10198 13568
rect 9878 12480 9886 12544
rect 9950 12480 9966 12544
rect 10030 12480 10046 12544
rect 10110 12480 10126 12544
rect 10190 12480 10198 12544
rect 9878 11456 10198 12480
rect 9878 11392 9886 11456
rect 9950 11392 9966 11456
rect 10030 11392 10046 11456
rect 10110 11392 10126 11456
rect 10190 11392 10198 11456
rect 9878 10368 10198 11392
rect 9878 10304 9886 10368
rect 9950 10304 9966 10368
rect 10030 10304 10046 10368
rect 10110 10304 10126 10368
rect 10190 10304 10198 10368
rect 9878 9280 10198 10304
rect 9878 9216 9886 9280
rect 9950 9216 9966 9280
rect 10030 9216 10046 9280
rect 10110 9216 10126 9280
rect 10190 9216 10198 9280
rect 9878 8192 10198 9216
rect 9878 8128 9886 8192
rect 9950 8128 9966 8192
rect 10030 8128 10046 8192
rect 10110 8128 10126 8192
rect 10190 8128 10198 8192
rect 9878 7104 10198 8128
rect 9878 7040 9886 7104
rect 9950 7040 9966 7104
rect 10030 7040 10046 7104
rect 10110 7040 10126 7104
rect 10190 7040 10198 7104
rect 9878 6016 10198 7040
rect 9878 5952 9886 6016
rect 9950 5952 9966 6016
rect 10030 5952 10046 6016
rect 10110 5952 10126 6016
rect 10190 5952 10198 6016
rect 9878 4928 10198 5952
rect 9878 4864 9886 4928
rect 9950 4864 9966 4928
rect 10030 4864 10046 4928
rect 10110 4864 10126 4928
rect 10190 4864 10198 4928
rect 9878 3840 10198 4864
rect 9878 3776 9886 3840
rect 9950 3776 9966 3840
rect 10030 3776 10046 3840
rect 10110 3776 10126 3840
rect 10190 3776 10198 3840
rect 9878 2752 10198 3776
rect 9878 2688 9886 2752
rect 9950 2688 9966 2752
rect 10030 2688 10046 2752
rect 10110 2688 10126 2752
rect 10190 2688 10198 2752
rect 9878 2128 10198 2688
rect 14878 21792 15198 21808
rect 14878 21728 14886 21792
rect 14950 21728 14966 21792
rect 15030 21728 15046 21792
rect 15110 21728 15126 21792
rect 15190 21728 15198 21792
rect 14878 20704 15198 21728
rect 14878 20640 14886 20704
rect 14950 20640 14966 20704
rect 15030 20640 15046 20704
rect 15110 20640 15126 20704
rect 15190 20640 15198 20704
rect 14878 19616 15198 20640
rect 14878 19552 14886 19616
rect 14950 19552 14966 19616
rect 15030 19552 15046 19616
rect 15110 19552 15126 19616
rect 15190 19552 15198 19616
rect 14878 18528 15198 19552
rect 14878 18464 14886 18528
rect 14950 18464 14966 18528
rect 15030 18464 15046 18528
rect 15110 18464 15126 18528
rect 15190 18464 15198 18528
rect 14878 17440 15198 18464
rect 14878 17376 14886 17440
rect 14950 17376 14966 17440
rect 15030 17376 15046 17440
rect 15110 17376 15126 17440
rect 15190 17376 15198 17440
rect 14878 16352 15198 17376
rect 14878 16288 14886 16352
rect 14950 16288 14966 16352
rect 15030 16288 15046 16352
rect 15110 16288 15126 16352
rect 15190 16288 15198 16352
rect 14878 15264 15198 16288
rect 14878 15200 14886 15264
rect 14950 15200 14966 15264
rect 15030 15200 15046 15264
rect 15110 15200 15126 15264
rect 15190 15200 15198 15264
rect 14878 14176 15198 15200
rect 14878 14112 14886 14176
rect 14950 14112 14966 14176
rect 15030 14112 15046 14176
rect 15110 14112 15126 14176
rect 15190 14112 15198 14176
rect 14878 13088 15198 14112
rect 14878 13024 14886 13088
rect 14950 13024 14966 13088
rect 15030 13024 15046 13088
rect 15110 13024 15126 13088
rect 15190 13024 15198 13088
rect 14878 12000 15198 13024
rect 14878 11936 14886 12000
rect 14950 11936 14966 12000
rect 15030 11936 15046 12000
rect 15110 11936 15126 12000
rect 15190 11936 15198 12000
rect 14878 10912 15198 11936
rect 14878 10848 14886 10912
rect 14950 10848 14966 10912
rect 15030 10848 15046 10912
rect 15110 10848 15126 10912
rect 15190 10848 15198 10912
rect 14878 9824 15198 10848
rect 14878 9760 14886 9824
rect 14950 9760 14966 9824
rect 15030 9760 15046 9824
rect 15110 9760 15126 9824
rect 15190 9760 15198 9824
rect 14878 8736 15198 9760
rect 14878 8672 14886 8736
rect 14950 8672 14966 8736
rect 15030 8672 15046 8736
rect 15110 8672 15126 8736
rect 15190 8672 15198 8736
rect 14878 7648 15198 8672
rect 14878 7584 14886 7648
rect 14950 7584 14966 7648
rect 15030 7584 15046 7648
rect 15110 7584 15126 7648
rect 15190 7584 15198 7648
rect 14878 6560 15198 7584
rect 14878 6496 14886 6560
rect 14950 6496 14966 6560
rect 15030 6496 15046 6560
rect 15110 6496 15126 6560
rect 15190 6496 15198 6560
rect 14878 5472 15198 6496
rect 14878 5408 14886 5472
rect 14950 5408 14966 5472
rect 15030 5408 15046 5472
rect 15110 5408 15126 5472
rect 15190 5408 15198 5472
rect 14878 4384 15198 5408
rect 14878 4320 14886 4384
rect 14950 4320 14966 4384
rect 15030 4320 15046 4384
rect 15110 4320 15126 4384
rect 15190 4320 15198 4384
rect 14878 3296 15198 4320
rect 14878 3232 14886 3296
rect 14950 3232 14966 3296
rect 15030 3232 15046 3296
rect 15110 3232 15126 3296
rect 15190 3232 15198 3296
rect 14878 2208 15198 3232
rect 14878 2144 14886 2208
rect 14950 2144 14966 2208
rect 15030 2144 15046 2208
rect 15110 2144 15126 2208
rect 15190 2144 15198 2208
rect 14878 2128 15198 2144
rect 19878 21248 20198 21808
rect 19878 21184 19886 21248
rect 19950 21184 19966 21248
rect 20030 21184 20046 21248
rect 20110 21184 20126 21248
rect 20190 21184 20198 21248
rect 19878 20160 20198 21184
rect 19878 20096 19886 20160
rect 19950 20096 19966 20160
rect 20030 20096 20046 20160
rect 20110 20096 20126 20160
rect 20190 20096 20198 20160
rect 19878 19072 20198 20096
rect 19878 19008 19886 19072
rect 19950 19008 19966 19072
rect 20030 19008 20046 19072
rect 20110 19008 20126 19072
rect 20190 19008 20198 19072
rect 19878 17984 20198 19008
rect 19878 17920 19886 17984
rect 19950 17920 19966 17984
rect 20030 17920 20046 17984
rect 20110 17920 20126 17984
rect 20190 17920 20198 17984
rect 19878 16896 20198 17920
rect 19878 16832 19886 16896
rect 19950 16832 19966 16896
rect 20030 16832 20046 16896
rect 20110 16832 20126 16896
rect 20190 16832 20198 16896
rect 19878 15808 20198 16832
rect 19878 15744 19886 15808
rect 19950 15744 19966 15808
rect 20030 15744 20046 15808
rect 20110 15744 20126 15808
rect 20190 15744 20198 15808
rect 19878 14720 20198 15744
rect 19878 14656 19886 14720
rect 19950 14656 19966 14720
rect 20030 14656 20046 14720
rect 20110 14656 20126 14720
rect 20190 14656 20198 14720
rect 19878 13632 20198 14656
rect 19878 13568 19886 13632
rect 19950 13568 19966 13632
rect 20030 13568 20046 13632
rect 20110 13568 20126 13632
rect 20190 13568 20198 13632
rect 19878 12544 20198 13568
rect 19878 12480 19886 12544
rect 19950 12480 19966 12544
rect 20030 12480 20046 12544
rect 20110 12480 20126 12544
rect 20190 12480 20198 12544
rect 19878 11456 20198 12480
rect 19878 11392 19886 11456
rect 19950 11392 19966 11456
rect 20030 11392 20046 11456
rect 20110 11392 20126 11456
rect 20190 11392 20198 11456
rect 19878 10368 20198 11392
rect 19878 10304 19886 10368
rect 19950 10304 19966 10368
rect 20030 10304 20046 10368
rect 20110 10304 20126 10368
rect 20190 10304 20198 10368
rect 19878 9280 20198 10304
rect 19878 9216 19886 9280
rect 19950 9216 19966 9280
rect 20030 9216 20046 9280
rect 20110 9216 20126 9280
rect 20190 9216 20198 9280
rect 19878 8192 20198 9216
rect 19878 8128 19886 8192
rect 19950 8128 19966 8192
rect 20030 8128 20046 8192
rect 20110 8128 20126 8192
rect 20190 8128 20198 8192
rect 19878 7104 20198 8128
rect 19878 7040 19886 7104
rect 19950 7040 19966 7104
rect 20030 7040 20046 7104
rect 20110 7040 20126 7104
rect 20190 7040 20198 7104
rect 19878 6016 20198 7040
rect 19878 5952 19886 6016
rect 19950 5952 19966 6016
rect 20030 5952 20046 6016
rect 20110 5952 20126 6016
rect 20190 5952 20198 6016
rect 19878 4928 20198 5952
rect 19878 4864 19886 4928
rect 19950 4864 19966 4928
rect 20030 4864 20046 4928
rect 20110 4864 20126 4928
rect 20190 4864 20198 4928
rect 19878 3840 20198 4864
rect 19878 3776 19886 3840
rect 19950 3776 19966 3840
rect 20030 3776 20046 3840
rect 20110 3776 20126 3840
rect 20190 3776 20198 3840
rect 19878 2752 20198 3776
rect 19878 2688 19886 2752
rect 19950 2688 19966 2752
rect 20030 2688 20046 2752
rect 20110 2688 20126 2752
rect 20190 2688 20198 2752
rect 19878 2128 20198 2688
rect 24878 21792 25198 21808
rect 24878 21728 24886 21792
rect 24950 21728 24966 21792
rect 25030 21728 25046 21792
rect 25110 21728 25126 21792
rect 25190 21728 25198 21792
rect 24878 20704 25198 21728
rect 24878 20640 24886 20704
rect 24950 20640 24966 20704
rect 25030 20640 25046 20704
rect 25110 20640 25126 20704
rect 25190 20640 25198 20704
rect 24878 19616 25198 20640
rect 24878 19552 24886 19616
rect 24950 19552 24966 19616
rect 25030 19552 25046 19616
rect 25110 19552 25126 19616
rect 25190 19552 25198 19616
rect 24878 18528 25198 19552
rect 24878 18464 24886 18528
rect 24950 18464 24966 18528
rect 25030 18464 25046 18528
rect 25110 18464 25126 18528
rect 25190 18464 25198 18528
rect 24878 17440 25198 18464
rect 24878 17376 24886 17440
rect 24950 17376 24966 17440
rect 25030 17376 25046 17440
rect 25110 17376 25126 17440
rect 25190 17376 25198 17440
rect 24878 16352 25198 17376
rect 24878 16288 24886 16352
rect 24950 16288 24966 16352
rect 25030 16288 25046 16352
rect 25110 16288 25126 16352
rect 25190 16288 25198 16352
rect 24878 15264 25198 16288
rect 24878 15200 24886 15264
rect 24950 15200 24966 15264
rect 25030 15200 25046 15264
rect 25110 15200 25126 15264
rect 25190 15200 25198 15264
rect 24878 14176 25198 15200
rect 24878 14112 24886 14176
rect 24950 14112 24966 14176
rect 25030 14112 25046 14176
rect 25110 14112 25126 14176
rect 25190 14112 25198 14176
rect 24878 13088 25198 14112
rect 24878 13024 24886 13088
rect 24950 13024 24966 13088
rect 25030 13024 25046 13088
rect 25110 13024 25126 13088
rect 25190 13024 25198 13088
rect 24878 12000 25198 13024
rect 24878 11936 24886 12000
rect 24950 11936 24966 12000
rect 25030 11936 25046 12000
rect 25110 11936 25126 12000
rect 25190 11936 25198 12000
rect 24878 10912 25198 11936
rect 24878 10848 24886 10912
rect 24950 10848 24966 10912
rect 25030 10848 25046 10912
rect 25110 10848 25126 10912
rect 25190 10848 25198 10912
rect 24878 9824 25198 10848
rect 24878 9760 24886 9824
rect 24950 9760 24966 9824
rect 25030 9760 25046 9824
rect 25110 9760 25126 9824
rect 25190 9760 25198 9824
rect 24878 8736 25198 9760
rect 24878 8672 24886 8736
rect 24950 8672 24966 8736
rect 25030 8672 25046 8736
rect 25110 8672 25126 8736
rect 25190 8672 25198 8736
rect 24878 7648 25198 8672
rect 24878 7584 24886 7648
rect 24950 7584 24966 7648
rect 25030 7584 25046 7648
rect 25110 7584 25126 7648
rect 25190 7584 25198 7648
rect 24878 6560 25198 7584
rect 24878 6496 24886 6560
rect 24950 6496 24966 6560
rect 25030 6496 25046 6560
rect 25110 6496 25126 6560
rect 25190 6496 25198 6560
rect 24878 5472 25198 6496
rect 24878 5408 24886 5472
rect 24950 5408 24966 5472
rect 25030 5408 25046 5472
rect 25110 5408 25126 5472
rect 25190 5408 25198 5472
rect 24878 4384 25198 5408
rect 24878 4320 24886 4384
rect 24950 4320 24966 4384
rect 25030 4320 25046 4384
rect 25110 4320 25126 4384
rect 25190 4320 25198 4384
rect 24878 3296 25198 4320
rect 24878 3232 24886 3296
rect 24950 3232 24966 3296
rect 25030 3232 25046 3296
rect 25110 3232 25126 3296
rect 25190 3232 25198 3296
rect 24878 2208 25198 3232
rect 24878 2144 24886 2208
rect 24950 2144 24966 2208
rect 25030 2144 25046 2208
rect 25110 2144 25126 2208
rect 25190 2144 25198 2208
rect 24878 2128 25198 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 38 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 38 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 314 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 1418 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 314 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 1418 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_72 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2890 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2522 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 2982 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 2522 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 3626 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 4086 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5190 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4730 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5466 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 5742 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 5650 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 5834 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 6938 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 5742 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 6846 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 8594 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 8042 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 8686 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 7950 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 9054 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 9790 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 10894 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 10158 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 11446 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 11262 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 11538 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 12642 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 11354 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 12458 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 14298 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 13746 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 14390 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 13562 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 15494 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 14666 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 15770 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 17150 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 16874 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 16598 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 17242 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 16966 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 18070 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 20002 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 18346 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 19450 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_218
timestamp 1586364061
transform 1 0 20094 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 19174 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21382 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _1_
timestamp 1586364061
transform 1 0 20278 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__1__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20830 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__0__A
timestamp 1586364061
transform 1 0 21934 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_224
timestamp 1586364061
transform 1 0 20646 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_228
timestamp 1586364061
transform 1 0 21014 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_236
timestamp 1586364061
transform 1 0 21750 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 20278 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 21382 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 22854 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 22486 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_240
timestamp 1586364061
transform 1 0 22118 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 22946 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 22578 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 23682 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 24050 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_273
timestamp 1586364061
transform 1 0 25154 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_269
timestamp 1586364061
transform 1 0 24786 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 25706 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_280
timestamp 1586364061
transform 1 0 25798 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_292
timestamp 1586364061
transform 1 0 26902 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_281
timestamp 1586364061
transform 1 0 25890 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_293
timestamp 1586364061
transform 1 0 26994 0 1 2720
box -38 -48 590 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 27822 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 27822 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_298 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 27454 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 38 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 314 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 1418 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 2890 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 2522 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 2982 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 4086 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 5190 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 6294 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 8502 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 7398 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 8594 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 9698 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 10802 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 11906 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 14114 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 13010 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 14206 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 15310 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 16414 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 17518 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 19726 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 18622 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 19818 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 20922 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 22026 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 23130 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 25338 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 24234 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_276
timestamp 1586364061
transform 1 0 25430 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_288
timestamp 1586364061
transform 1 0 26534 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_296
timestamp 1586364061
transform 1 0 27270 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 27822 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 38 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 314 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 1418 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 2522 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 3626 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 4730 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 5466 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 5650 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 5742 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 6846 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 7950 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 9054 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 10158 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 11262 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 11354 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 12458 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 13562 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 14666 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 15770 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 16874 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 16966 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 18070 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 19174 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 20278 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 21382 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 22486 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 22578 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 23682 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_269
timestamp 1586364061
transform 1 0 24786 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_281
timestamp 1586364061
transform 1 0 25890 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_3_293
timestamp 1586364061
transform 1 0 26994 0 1 3808
box -38 -48 590 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 27822 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 38 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 314 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 1418 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 2890 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 2522 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 2982 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 4086 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 5190 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 6294 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 8502 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 7398 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 8594 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 9698 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 10802 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 11906 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 14114 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 13010 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 14206 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 15310 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 16414 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 17518 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 19726 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 18622 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 19818 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 20922 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 22026 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 23130 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 25338 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 24234 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_276
timestamp 1586364061
transform 1 0 25430 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_288
timestamp 1586364061
transform 1 0 26534 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_4_296
timestamp 1586364061
transform 1 0 27270 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 27822 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 38 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 314 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 1418 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 2522 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 3626 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 4730 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 5466 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 5650 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 5742 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 6846 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 7950 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 9054 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 10158 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 11262 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 11354 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 12458 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 13562 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 14666 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 15770 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 16874 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 16966 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 18070 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 19174 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 20278 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 21382 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 22486 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 22578 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 23682 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_269
timestamp 1586364061
transform 1 0 24786 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_281
timestamp 1586364061
transform 1 0 25890 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_5_293
timestamp 1586364061
transform 1 0 26994 0 1 4896
box -38 -48 590 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 27822 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 38 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 38 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 314 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 1418 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 314 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 1418 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 2890 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 2522 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 2982 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 2522 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 3626 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 4086 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 5190 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 4730 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 5466 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 5650 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 6294 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 5742 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 6846 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 8502 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 7398 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 8594 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 7950 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 9054 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 9698 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 10802 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 10158 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 11262 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 11906 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 11354 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 12458 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 14114 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 13010 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 14206 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_147
timestamp 1586364061
transform 1 0 13562 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 15310 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 16414 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_159
timestamp 1586364061
transform 1 0 14666 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_171
timestamp 1586364061
transform 1 0 15770 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 16874 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 17518 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 16966 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 18070 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 19726 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 18622 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 19818 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 19174 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 20922 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 20278 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 21382 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 22486 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 22026 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 23130 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 22578 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 23682 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 25338 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 24234 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_276
timestamp 1586364061
transform 1 0 25430 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_269
timestamp 1586364061
transform 1 0 24786 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_288
timestamp 1586364061
transform 1 0 26534 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_296
timestamp 1586364061
transform 1 0 27270 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_281
timestamp 1586364061
transform 1 0 25890 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_293
timestamp 1586364061
transform 1 0 26994 0 1 5984
box -38 -48 590 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 27822 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 27822 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 38 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 314 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 1418 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 2890 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 2522 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 2982 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 4086 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 5190 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 6294 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 8502 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 7398 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 8594 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 9698 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 10802 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 11906 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 14114 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 13010 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 14206 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 15310 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 16414 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 17518 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 19726 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 18622 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 19818 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 20922 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 22026 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 23130 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 25338 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 24234 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_276
timestamp 1586364061
transform 1 0 25430 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_288
timestamp 1586364061
transform 1 0 26534 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_296
timestamp 1586364061
transform 1 0 27270 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 27822 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 38 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 314 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 1418 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 2522 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 3626 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 4730 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 5466 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 5650 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 5742 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 6846 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 7950 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 9054 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_110
timestamp 1586364061
transform 1 0 10158 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 11262 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 11354 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 12458 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 13562 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 14666 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_171
timestamp 1586364061
transform 1 0 15770 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 16874 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 16966 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 18070 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 19174 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 20278 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 21382 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 22486 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 22578 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 23682 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_269
timestamp 1586364061
transform 1 0 24786 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_281
timestamp 1586364061
transform 1 0 25890 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_293
timestamp 1586364061
transform 1 0 26994 0 1 7072
box -38 -48 590 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 27822 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 38 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 314 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 1418 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 2890 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 2522 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 2982 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 4086 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 5190 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 6294 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 8502 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 7398 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 8594 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 9698 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 10802 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 11906 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 14114 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 13010 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 14206 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 15310 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 16414 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_190
timestamp 1586364061
transform 1 0 17518 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 19726 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_202
timestamp 1586364061
transform 1 0 18622 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 19818 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 20922 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 22026 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 23130 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 25338 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 24234 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_276
timestamp 1586364061
transform 1 0 25430 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_288
timestamp 1586364061
transform 1 0 26534 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_296
timestamp 1586364061
transform 1 0 27270 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 27822 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 38 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 314 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 1418 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 2522 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 3626 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 4730 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 5466 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 5650 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 5742 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 6846 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 7950 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 9054 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 10158 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 11262 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 11354 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 12458 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 13562 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_159
timestamp 1586364061
transform 1 0 14666 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_171
timestamp 1586364061
transform 1 0 15770 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 16874 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 16966 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 18070 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 19174 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 20278 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 21382 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 22486 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 22578 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 23682 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_269
timestamp 1586364061
transform 1 0 24786 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_281
timestamp 1586364061
transform 1 0 25890 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_11_293
timestamp 1586364061
transform 1 0 26994 0 1 8160
box -38 -48 590 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 27822 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 38 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 314 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 1418 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 2890 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 2522 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 2982 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 4086 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 5190 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 6294 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 8502 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 7398 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 8594 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 9698 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 10802 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 11906 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 14114 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 13010 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 14206 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 15310 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 16414 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_190
timestamp 1586364061
transform 1 0 17518 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 19726 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_202
timestamp 1586364061
transform 1 0 18622 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 19818 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 20922 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 22026 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 23130 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 25338 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 24234 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_276
timestamp 1586364061
transform 1 0 25430 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_288
timestamp 1586364061
transform 1 0 26534 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_296
timestamp 1586364061
transform 1 0 27270 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 27822 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 38 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 38 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 314 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 1418 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 314 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 1418 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 2890 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 2522 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 3626 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 2522 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 2982 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 4730 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 5466 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 4086 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 5190 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 5650 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 5742 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 6846 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 6294 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 8502 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 7950 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 9054 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 7398 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 8594 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 10158 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 9698 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 10802 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 11262 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 11354 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 12458 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 11906 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 14114 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_147
timestamp 1586364061
transform 1 0 13562 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 13010 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 14206 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_159
timestamp 1586364061
transform 1 0 14666 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_171
timestamp 1586364061
transform 1 0 15770 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 15310 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 16414 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 16874 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 16966 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 18070 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 17518 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 19726 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 19174 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 18622 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 19818 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 20278 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 21382 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 20922 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 22486 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_scs8hd_dfxbp_1_mem.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 22854 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 22578 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 23682 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_239
timestamp 1586364061
transform 1 0 22026 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_247
timestamp 1586364061
transform 1 0 22762 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_250
timestamp 1586364061
transform 1 0 23038 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 25338 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_269
timestamp 1586364061
transform 1 0 24786 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_262
timestamp 1586364061
transform 1 0 24142 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_274
timestamp 1586364061
transform 1 0 25246 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_276
timestamp 1586364061
transform 1 0 25430 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_281
timestamp 1586364061
transform 1 0 25890 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_13_293
timestamp 1586364061
transform 1 0 26994 0 1 9248
box -38 -48 590 592
use scs8hd_decap_8  FILLER_14_288
timestamp 1586364061
transform 1 0 26534 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_296
timestamp 1586364061
transform 1 0 27270 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 27822 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 27822 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 38 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 314 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 1418 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 2522 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 3626 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 4730 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 5466 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 5650 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 5742 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 6846 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 7950 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_98
timestamp 1586364061
transform 1 0 9054 0 1 10336
box -38 -48 774 592
use scs8hd_buf_2  _2_
timestamp 1586364061
transform 1 0 9974 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__2__A
timestamp 1586364061
transform 1 0 10526 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_106
timestamp 1586364061
transform 1 0 9790 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_112
timestamp 1586364061
transform 1 0 10342 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_116
timestamp 1586364061
transform 1 0 10710 0 1 10336
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 11262 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 11354 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 12458 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 13562 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_159
timestamp 1586364061
transform 1 0 14666 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_171
timestamp 1586364061
transform 1 0 15770 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 16874 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 16966 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 18070 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 19174 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 20278 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 21382 0 1 10336
box -38 -48 1142 592
use scs8hd_dfxbp_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_scs8hd_dfxbp_1_mem.scs8hd_dfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 22854 0 1 10336
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 22486 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_245
timestamp 1586364061
transform 1 0 22578 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_267
timestamp 1586364061
transform 1 0 24602 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_279
timestamp 1586364061
transform 1 0 25706 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_291
timestamp 1586364061
transform 1 0 26810 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 27822 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 38 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 314 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 1418 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 2890 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 2522 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 2982 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 4086 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 5190 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 6294 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 8502 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 7398 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 8594 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 9698 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 10802 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 11906 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 14114 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 13010 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 14206 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 15310 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 16414 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 17518 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 19726 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 18622 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 19818 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 20922 0 -1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_scs8hd_dfxbp_1_mem.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 22854 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_239
timestamp 1586364061
transform 1 0 22026 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_247
timestamp 1586364061
transform 1 0 22762 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_250
timestamp 1586364061
transform 1 0 23038 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 25338 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_262
timestamp 1586364061
transform 1 0 24142 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 25246 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_276
timestamp 1586364061
transform 1 0 25430 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_288
timestamp 1586364061
transform 1 0 26534 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_296
timestamp 1586364061
transform 1 0 27270 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 27822 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 38 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 314 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 1418 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 2522 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 3626 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 4730 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 5466 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 5650 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 5742 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 6846 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 7950 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 9054 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 10158 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 11262 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 11354 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 12458 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_147
timestamp 1586364061
transform 1 0 13562 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_159
timestamp 1586364061
transform 1 0 14666 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_171
timestamp 1586364061
transform 1 0 15770 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 16874 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 16966 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 18070 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 19174 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 20278 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 21382 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 22486 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 22578 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 23682 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_269
timestamp 1586364061
transform 1 0 24786 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_281
timestamp 1586364061
transform 1 0 25890 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_17_293
timestamp 1586364061
transform 1 0 26994 0 1 11424
box -38 -48 590 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 27822 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 38 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 314 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 1418 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 2890 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 2522 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 2982 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 4086 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 5190 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 6294 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 8502 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 7398 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 8594 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 9698 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 10802 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_129
timestamp 1586364061
transform 1 0 11906 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 14114 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 13010 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 14206 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 15310 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 16414 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 17518 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 19726 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 18622 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 19818 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 20922 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 22026 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 23130 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 25338 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 24234 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_276
timestamp 1586364061
transform 1 0 25430 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_288
timestamp 1586364061
transform 1 0 26534 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_296
timestamp 1586364061
transform 1 0 27270 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 27822 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 38 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 38 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 314 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 1418 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 314 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 1418 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 2890 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 2522 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 3626 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 2522 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 2982 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 4730 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 5466 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 4086 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 5190 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 5650 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 5742 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 6846 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 6294 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 8502 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 7950 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 9054 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 7398 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 8594 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 10158 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 9698 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_117
timestamp 1586364061
transform 1 0 10802 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 11262 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 11354 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 12458 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_129
timestamp 1586364061
transform 1 0 11906 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 14114 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 13562 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_141
timestamp 1586364061
transform 1 0 13010 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_154
timestamp 1586364061
transform 1 0 14206 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 14666 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 15770 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_166
timestamp 1586364061
transform 1 0 15310 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_178
timestamp 1586364061
transform 1 0 16414 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 16874 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 16966 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 18070 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_190
timestamp 1586364061
transform 1 0 17518 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 19726 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 19174 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_202
timestamp 1586364061
transform 1 0 18622 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 19818 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 20278 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 21382 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 20922 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 22486 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 22578 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 23682 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 22026 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_251
timestamp 1586364061
transform 1 0 23130 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 25338 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_269
timestamp 1586364061
transform 1 0 24786 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 24234 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_276
timestamp 1586364061
transform 1 0 25430 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_281
timestamp 1586364061
transform 1 0 25890 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_19_293
timestamp 1586364061
transform 1 0 26994 0 1 12512
box -38 -48 590 592
use scs8hd_decap_8  FILLER_20_288
timestamp 1586364061
transform 1 0 26534 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_20_296
timestamp 1586364061
transform 1 0 27270 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 27822 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 27822 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 38 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 314 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 1418 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 2522 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 3626 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 4730 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 5466 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 5650 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 5742 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 6846 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_86
timestamp 1586364061
transform 1 0 7950 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_98
timestamp 1586364061
transform 1 0 9054 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_110
timestamp 1586364061
transform 1 0 10158 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 11262 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 11354 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_135
timestamp 1586364061
transform 1 0 12458 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_147
timestamp 1586364061
transform 1 0 13562 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_159
timestamp 1586364061
transform 1 0 14666 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 15770 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 16874 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 16966 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 18070 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 19174 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 20278 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 21382 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 22486 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 22578 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 23682 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_269
timestamp 1586364061
transform 1 0 24786 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_281
timestamp 1586364061
transform 1 0 25890 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_21_293
timestamp 1586364061
transform 1 0 26994 0 1 13600
box -38 -48 590 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 27822 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 38 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 314 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 1418 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 2890 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 2522 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 2982 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 4086 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 5190 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 6294 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 8502 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 7398 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 8594 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 9698 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_117
timestamp 1586364061
transform 1 0 10802 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_129
timestamp 1586364061
transform 1 0 11906 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 14114 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_141
timestamp 1586364061
transform 1 0 13010 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_154
timestamp 1586364061
transform 1 0 14206 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_166
timestamp 1586364061
transform 1 0 15310 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_178
timestamp 1586364061
transform 1 0 16414 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_190
timestamp 1586364061
transform 1 0 17518 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 19726 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_202
timestamp 1586364061
transform 1 0 18622 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 19818 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 20922 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 22026 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 23130 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 25338 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 24234 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_276
timestamp 1586364061
transform 1 0 25430 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_288
timestamp 1586364061
transform 1 0 26534 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_296
timestamp 1586364061
transform 1 0 27270 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 27822 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 38 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 314 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 1418 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 2522 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 3626 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 4730 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 5466 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 5650 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 5742 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 6846 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 7950 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 9054 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_110
timestamp 1586364061
transform 1 0 10158 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 11262 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 11354 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_135
timestamp 1586364061
transform 1 0 12458 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_147
timestamp 1586364061
transform 1 0 13562 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_159
timestamp 1586364061
transform 1 0 14666 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_171
timestamp 1586364061
transform 1 0 15770 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 16874 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 16966 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 18070 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 19174 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 20278 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_232
timestamp 1586364061
transform 1 0 21382 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 22486 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 22578 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 23682 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_269
timestamp 1586364061
transform 1 0 24786 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_281
timestamp 1586364061
transform 1 0 25890 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_23_293
timestamp 1586364061
transform 1 0 26994 0 1 14688
box -38 -48 590 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 27822 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 38 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 314 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 1418 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 2890 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 2522 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 2982 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 4086 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 5190 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 6294 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 8502 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 7398 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 8594 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 9698 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 10802 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 11906 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 14114 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_141
timestamp 1586364061
transform 1 0 13010 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 14206 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 15310 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 16414 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_190
timestamp 1586364061
transform 1 0 17518 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 19726 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 18622 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 19818 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 20922 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 22026 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 23130 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 25338 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 24234 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_276
timestamp 1586364061
transform 1 0 25430 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_288
timestamp 1586364061
transform 1 0 26534 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_24_296
timestamp 1586364061
transform 1 0 27270 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 27822 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 38 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 314 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 1418 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 2522 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 3626 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 4730 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 5466 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 5650 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 5742 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 6846 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_86
timestamp 1586364061
transform 1 0 7950 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_98
timestamp 1586364061
transform 1 0 9054 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_110
timestamp 1586364061
transform 1 0 10158 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 11262 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 11354 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 12458 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_147
timestamp 1586364061
transform 1 0 13562 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_159
timestamp 1586364061
transform 1 0 14666 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_171
timestamp 1586364061
transform 1 0 15770 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 16874 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 16966 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 18070 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 19174 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 20278 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_232
timestamp 1586364061
transform 1 0 21382 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 22486 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 22578 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 23682 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_269
timestamp 1586364061
transform 1 0 24786 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_281
timestamp 1586364061
transform 1 0 25890 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_25_293
timestamp 1586364061
transform 1 0 26994 0 1 15776
box -38 -48 590 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 27822 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 38 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 38 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 314 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 1418 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 314 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 1418 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 2890 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 2522 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 2982 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 2522 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 3626 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 4086 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 5190 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 4730 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 5466 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 5650 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 6294 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 5742 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 6846 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 8502 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 7398 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 8594 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 7950 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 9054 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 9698 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 10802 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_110
timestamp 1586364061
transform 1 0 10158 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 11262 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 11906 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 11354 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 12458 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 14114 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 13010 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 14206 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 13562 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 15310 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 16414 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 14666 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 15770 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 16874 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 17518 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 16966 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 18070 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 19726 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 18622 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 19818 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 19174 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 20922 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 20278 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 21382 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 22486 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 22026 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 23130 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 22578 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 23682 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 25338 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 24234 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_276
timestamp 1586364061
transform 1 0 25430 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_269
timestamp 1586364061
transform 1 0 24786 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_26_288
timestamp 1586364061
transform 1 0 26534 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_296
timestamp 1586364061
transform 1 0 27270 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_281
timestamp 1586364061
transform 1 0 25890 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_27_293
timestamp 1586364061
transform 1 0 26994 0 1 16864
box -38 -48 590 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 27822 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 27822 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 38 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 314 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 1418 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 2890 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 2522 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 2982 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 4086 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 5190 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 6294 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 8502 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 7398 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 8594 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 9698 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 10802 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 11906 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 14114 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 13010 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 14206 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 15310 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 16414 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 17518 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 19726 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 18622 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 19818 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 20922 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 22026 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 23130 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 25338 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 24234 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_276
timestamp 1586364061
transform 1 0 25430 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_28_288
timestamp 1586364061
transform 1 0 26534 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_296
timestamp 1586364061
transform 1 0 27270 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 27822 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 38 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 314 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 1418 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 2522 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 3626 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 4730 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 5466 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 5650 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 5742 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 6846 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 7950 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 9054 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 10158 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 11262 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 11354 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_135
timestamp 1586364061
transform 1 0 12458 0 1 17952
box -38 -48 774 592
use scs8hd_buf_2  _3_
timestamp 1586364061
transform 1 0 13194 0 1 17952
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__3__A
timestamp 1586364061
transform 1 0 13746 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_147
timestamp 1586364061
transform 1 0 13562 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_151
timestamp 1586364061
transform 1 0 13930 0 1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.ie_oe_inv_A
timestamp 1586364061
transform 1 0 15034 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_165
timestamp 1586364061
transform 1 0 15218 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_29_177
timestamp 1586364061
transform 1 0 16322 0 1 17952
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 16874 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 16966 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 18070 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 19174 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 20278 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 21382 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 22486 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 22578 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 23682 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_269
timestamp 1586364061
transform 1 0 24786 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_281
timestamp 1586364061
transform 1 0 25890 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_29_293
timestamp 1586364061
transform 1 0 26994 0 1 17952
box -38 -48 590 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 27822 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 38 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 314 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 1418 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 2890 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 2522 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 2982 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 4086 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 5190 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 6294 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 8502 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 7398 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 8594 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 9698 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 10802 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 11906 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 14114 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 13010 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_154
timestamp 1586364061
transform 1 0 14206 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.ie_oe_inv tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15034 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_1  FILLER_30_162
timestamp 1586364061
transform 1 0 14942 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 15310 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 16414 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 17518 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 19726 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 18622 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 19818 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 20922 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 22026 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 23130 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 25338 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 24234 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_276
timestamp 1586364061
transform 1 0 25430 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_288
timestamp 1586364061
transform 1 0 26534 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_30_296
timestamp 1586364061
transform 1 0 27270 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 27822 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 38 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 314 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 1418 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 2522 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 3626 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 4730 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 5466 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 5650 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 5742 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 6846 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 7950 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 9054 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 10158 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 11262 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 11354 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 12458 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 13562 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 14666 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 15770 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 16874 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 16966 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 18070 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 19174 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 20278 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 21382 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 22486 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 22578 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 23682 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_269
timestamp 1586364061
transform 1 0 24786 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_281
timestamp 1586364061
transform 1 0 25890 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_31_293
timestamp 1586364061
transform 1 0 26994 0 1 19040
box -38 -48 590 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 27822 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 38 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 314 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 1418 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 2890 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 2522 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 2982 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 4086 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 5190 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 6294 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 8502 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 7398 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 8594 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 9698 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 10802 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 11906 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 14114 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 13010 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 14206 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 15310 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 16414 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 17518 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 19726 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 18622 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 19818 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 20922 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 22026 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 23130 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 25338 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 24234 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_276
timestamp 1586364061
transform 1 0 25430 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_288
timestamp 1586364061
transform 1 0 26534 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_32_296
timestamp 1586364061
transform 1 0 27270 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 27822 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 38 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 38 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 314 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 1418 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 314 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 1418 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 2890 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 2522 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 3626 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 2522 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 2982 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 4730 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 5466 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 4086 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 5190 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 5650 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 5742 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 6846 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 6294 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 8502 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 7950 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 9054 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 7398 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 8594 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 10158 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 9698 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 10802 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 11262 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 11354 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 12458 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 11906 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 14114 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 13562 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 13010 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 14206 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 14666 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 15770 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 15310 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 16414 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 16874 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 16966 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 18070 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 17518 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 19726 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 19174 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 18622 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 19818 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 20278 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 21382 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 20922 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 22486 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 22578 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 23682 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 22026 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 23130 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 25338 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_269
timestamp 1586364061
transform 1 0 24786 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 24234 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_276
timestamp 1586364061
transform 1 0 25430 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_281
timestamp 1586364061
transform 1 0 25890 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_33_293
timestamp 1586364061
transform 1 0 26994 0 1 20128
box -38 -48 590 592
use scs8hd_decap_8  FILLER_34_288
timestamp 1586364061
transform 1 0 26534 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  FILLER_34_296
timestamp 1586364061
transform 1 0 27270 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 27822 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 27822 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 38 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 314 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 1418 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 2890 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_27
timestamp 1586364061
transform 1 0 2522 0 1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_35_32
timestamp 1586364061
transform 1 0 2982 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_44
timestamp 1586364061
transform 1 0 4086 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_56
timestamp 1586364061
transform 1 0 5190 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 5742 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_63
timestamp 1586364061
transform 1 0 5834 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_75
timestamp 1586364061
transform 1 0 6938 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 8594 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_87
timestamp 1586364061
transform 1 0 8042 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_94
timestamp 1586364061
transform 1 0 8686 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_106
timestamp 1586364061
transform 1 0 9790 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_118
timestamp 1586364061
transform 1 0 10894 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 11446 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_125
timestamp 1586364061
transform 1 0 11538 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_137
timestamp 1586364061
transform 1 0 12642 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 14298 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_149
timestamp 1586364061
transform 1 0 13746 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_156
timestamp 1586364061
transform 1 0 14390 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_168
timestamp 1586364061
transform 1 0 15494 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 17150 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_180
timestamp 1586364061
transform 1 0 16598 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_187
timestamp 1586364061
transform 1 0 17242 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 20002 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_199
timestamp 1586364061
transform 1 0 18346 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_211
timestamp 1586364061
transform 1 0 19450 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_218
timestamp 1586364061
transform 1 0 20094 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_230
timestamp 1586364061
transform 1 0 21198 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 22854 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_242
timestamp 1586364061
transform 1 0 22302 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_249
timestamp 1586364061
transform 1 0 22946 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_261
timestamp 1586364061
transform 1 0 24050 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_273
timestamp 1586364061
transform 1 0 25154 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 25706 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_280
timestamp 1586364061
transform 1 0 25798 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_292
timestamp 1586364061
transform 1 0 26902 0 1 21216
box -38 -48 590 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 27822 0 1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_35_298
timestamp 1586364061
transform 1 0 27454 0 1 21216
box -38 -48 130 592
<< labels >>
rlabel metal2 s 13856 0 13912 480 6 bottom_width_0_height_0__pin_0_
port 0 nsew default input
rlabel metal2 s 23884 0 23940 480 6 bottom_width_0_height_0__pin_1_lower
port 1 nsew default tristate
rlabel metal2 s 3920 0 3976 480 6 bottom_width_0_height_0__pin_1_upper
port 2 nsew default tristate
rlabel metal3 s 28454 11840 28934 11960 6 ccff_head
port 3 nsew default input
rlabel metal3 s 28454 19864 28934 19984 6 ccff_tail
port 4 nsew default tristate
rlabel metal2 s 2632 23520 2688 24000 6 gfpga_pad_GPIO_A
port 5 nsew default tristate
rlabel metal2 s 10084 23520 10140 24000 6 gfpga_pad_GPIO_IE
port 6 nsew default tristate
rlabel metal2 s 17628 23520 17684 24000 6 gfpga_pad_GPIO_OE
port 7 nsew default tristate
rlabel metal2 s 25080 23520 25136 24000 6 gfpga_pad_GPIO_Y
port 8 nsew default bidirectional
rlabel metal3 s 28454 3952 28934 4072 6 prog_clk
port 9 nsew default input
rlabel metal4 s 4878 2128 5198 21808 6 vpwr
port 10 nsew default input
rlabel metal4 s 9878 2128 10198 21808 6 vgnd
port 11 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28934 24000
<< end >>
