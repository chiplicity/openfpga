VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_2__1_
  CLASS BLOCK ;
  FOREIGN sb_2__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 115.000 BY 115.000 ;
  PIN bottom_left_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 2.400 ;
    END
  END bottom_left_grid_pin_42_
  PIN bottom_left_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 2.400 ;
    END
  END bottom_left_grid_pin_43_
  PIN bottom_left_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 2.400 ;
    END
  END bottom_left_grid_pin_44_
  PIN bottom_left_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 2.400 ;
    END
  END bottom_left_grid_pin_45_
  PIN bottom_left_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 2.400 ;
    END
  END bottom_left_grid_pin_46_
  PIN bottom_left_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 2.400 ;
    END
  END bottom_left_grid_pin_47_
  PIN bottom_left_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 2.400 ;
    END
  END bottom_left_grid_pin_48_
  PIN bottom_left_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 2.400 ;
    END
  END bottom_left_grid_pin_49_
  PIN bottom_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 2.400 ;
    END
  END bottom_right_grid_pin_1_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 57.160 115.000 57.760 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 112.600 95.240 115.000 95.840 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 2.400 20.360 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 2.400 44.160 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 2.400 46.200 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 2.400 48.920 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 2.400 50.960 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 2.400 53.680 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 2.400 55.720 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 2.400 58.440 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 2.400 61.160 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 2.400 63.200 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 2.400 65.920 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 2.400 22.400 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 2.400 25.120 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 2.400 27.160 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 2.400 29.880 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 2.400 31.920 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 2.400 34.640 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 2.400 36.680 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 2.400 39.400 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.400 41.440 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 2.400 67.960 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 2.400 91.760 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 2.400 94.480 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 2.400 96.520 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 2.400 99.240 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 2.400 101.280 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 2.400 104.000 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 2.400 106.040 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 2.400 108.760 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 2.400 110.800 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 2.400 113.520 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 2.400 70.680 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 2.400 72.720 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 2.400 75.440 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 2.400 77.480 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.400 80.200 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 2.400 82.240 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 2.400 84.960 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 2.400 87.000 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 2.400 89.720 ;
    END
  END chanx_left_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 2.400 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 2.400 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 2.400 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 2.400 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 2.400 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 2.400 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 2.400 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 2.400 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 2.400 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 2.400 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 2.400 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 2.400 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 2.400 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 2.400 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 2.400 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 2.400 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 2.400 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 2.400 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 2.400 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 2.400 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 2.400 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 2.400 ;
    END
  END chany_bottom_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 112.600 19.690 115.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.870 112.600 43.150 115.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 112.600 45.450 115.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.930 112.600 48.210 115.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 112.600 50.510 115.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 112.600 52.810 115.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.830 112.600 55.110 115.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.130 112.600 57.410 115.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.430 112.600 59.710 115.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.730 112.600 62.010 115.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.030 112.600 64.310 115.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 112.600 21.990 115.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.470 112.600 24.750 115.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 112.600 27.050 115.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.070 112.600 29.350 115.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.370 112.600 31.650 115.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.670 112.600 33.950 115.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.970 112.600 36.250 115.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 112.600 38.550 115.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.570 112.600 40.850 115.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 66.330 112.600 66.610 115.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 112.600 90.070 115.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.090 112.600 92.370 115.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.850 112.600 95.130 115.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.150 112.600 97.430 115.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 99.450 112.600 99.730 115.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.750 112.600 102.030 115.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.050 112.600 104.330 115.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.350 112.600 106.630 115.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.650 112.600 108.930 115.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.950 112.600 111.230 115.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.630 112.600 68.910 115.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.390 112.600 71.670 115.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 112.600 73.970 115.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.990 112.600 76.270 115.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.290 112.600 78.570 115.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.590 112.600 80.870 115.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.890 112.600 83.170 115.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.190 112.600 85.470 115.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.490 112.600 87.770 115.000 ;
    END
  END chany_top_out[9]
  PIN left_bottom_grid_pin_34_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 2.400 1.320 ;
    END
  END left_bottom_grid_pin_34_
  PIN left_bottom_grid_pin_35_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 2.400 3.360 ;
    END
  END left_bottom_grid_pin_35_
  PIN left_bottom_grid_pin_36_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 2.400 6.080 ;
    END
  END left_bottom_grid_pin_36_
  PIN left_bottom_grid_pin_37_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 2.400 8.120 ;
    END
  END left_bottom_grid_pin_37_
  PIN left_bottom_grid_pin_38_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 2.400 10.840 ;
    END
  END left_bottom_grid_pin_38_
  PIN left_bottom_grid_pin_39_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END left_bottom_grid_pin_39_
  PIN left_bottom_grid_pin_40_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 2.400 15.600 ;
    END
  END left_bottom_grid_pin_40_
  PIN left_bottom_grid_pin_41_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 2.400 17.640 ;
    END
  END left_bottom_grid_pin_41_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 112.600 19.080 115.000 19.680 ;
    END
  END prog_clk
  PIN top_left_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 112.600 1.290 115.000 ;
    END
  END top_left_grid_pin_42_
  PIN top_left_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 112.600 3.590 115.000 ;
    END
  END top_left_grid_pin_43_
  PIN top_left_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 112.600 5.890 115.000 ;
    END
  END top_left_grid_pin_44_
  PIN top_left_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.910 112.600 8.190 115.000 ;
    END
  END top_left_grid_pin_45_
  PIN top_left_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 112.600 10.490 115.000 ;
    END
  END top_left_grid_pin_46_
  PIN top_left_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 112.600 12.790 115.000 ;
    END
  END top_left_grid_pin_47_
  PIN top_left_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.810 112.600 15.090 115.000 ;
    END
  END top_left_grid_pin_48_
  PIN top_left_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 112.600 17.390 115.000 ;
    END
  END top_left_grid_pin_49_
  PIN top_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.250 112.600 113.530 115.000 ;
    END
  END top_right_grid_pin_1_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.045 10.640 23.645 103.600 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.375 10.640 40.975 103.600 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 109.480 103.445 ;
      LAYER met1 ;
        RECT 0.990 2.760 113.550 104.000 ;
      LAYER met2 ;
        RECT 1.570 112.320 3.030 113.405 ;
        RECT 3.870 112.320 5.330 113.405 ;
        RECT 6.170 112.320 7.630 113.405 ;
        RECT 8.470 112.320 9.930 113.405 ;
        RECT 10.770 112.320 12.230 113.405 ;
        RECT 13.070 112.320 14.530 113.405 ;
        RECT 15.370 112.320 16.830 113.405 ;
        RECT 17.670 112.320 19.130 113.405 ;
        RECT 19.970 112.320 21.430 113.405 ;
        RECT 22.270 112.320 24.190 113.405 ;
        RECT 25.030 112.320 26.490 113.405 ;
        RECT 27.330 112.320 28.790 113.405 ;
        RECT 29.630 112.320 31.090 113.405 ;
        RECT 31.930 112.320 33.390 113.405 ;
        RECT 34.230 112.320 35.690 113.405 ;
        RECT 36.530 112.320 37.990 113.405 ;
        RECT 38.830 112.320 40.290 113.405 ;
        RECT 41.130 112.320 42.590 113.405 ;
        RECT 43.430 112.320 44.890 113.405 ;
        RECT 45.730 112.320 47.650 113.405 ;
        RECT 48.490 112.320 49.950 113.405 ;
        RECT 50.790 112.320 52.250 113.405 ;
        RECT 53.090 112.320 54.550 113.405 ;
        RECT 55.390 112.320 56.850 113.405 ;
        RECT 57.690 112.320 59.150 113.405 ;
        RECT 59.990 112.320 61.450 113.405 ;
        RECT 62.290 112.320 63.750 113.405 ;
        RECT 64.590 112.320 66.050 113.405 ;
        RECT 66.890 112.320 68.350 113.405 ;
        RECT 69.190 112.320 71.110 113.405 ;
        RECT 71.950 112.320 73.410 113.405 ;
        RECT 74.250 112.320 75.710 113.405 ;
        RECT 76.550 112.320 78.010 113.405 ;
        RECT 78.850 112.320 80.310 113.405 ;
        RECT 81.150 112.320 82.610 113.405 ;
        RECT 83.450 112.320 84.910 113.405 ;
        RECT 85.750 112.320 87.210 113.405 ;
        RECT 88.050 112.320 89.510 113.405 ;
        RECT 90.350 112.320 91.810 113.405 ;
        RECT 92.650 112.320 94.570 113.405 ;
        RECT 95.410 112.320 96.870 113.405 ;
        RECT 97.710 112.320 99.170 113.405 ;
        RECT 100.010 112.320 101.470 113.405 ;
        RECT 102.310 112.320 103.770 113.405 ;
        RECT 104.610 112.320 106.070 113.405 ;
        RECT 106.910 112.320 108.370 113.405 ;
        RECT 109.210 112.320 110.670 113.405 ;
        RECT 111.510 112.320 112.970 113.405 ;
        RECT 1.020 2.680 113.520 112.320 ;
        RECT 1.570 2.400 3.030 2.680 ;
        RECT 3.870 2.400 5.330 2.680 ;
        RECT 6.170 2.400 7.630 2.680 ;
        RECT 8.470 2.400 9.930 2.680 ;
        RECT 10.770 2.400 12.230 2.680 ;
        RECT 13.070 2.400 14.530 2.680 ;
        RECT 15.370 2.400 16.830 2.680 ;
        RECT 17.670 2.400 19.130 2.680 ;
        RECT 19.970 2.400 21.430 2.680 ;
        RECT 22.270 2.400 24.190 2.680 ;
        RECT 25.030 2.400 26.490 2.680 ;
        RECT 27.330 2.400 28.790 2.680 ;
        RECT 29.630 2.400 31.090 2.680 ;
        RECT 31.930 2.400 33.390 2.680 ;
        RECT 34.230 2.400 35.690 2.680 ;
        RECT 36.530 2.400 37.990 2.680 ;
        RECT 38.830 2.400 40.290 2.680 ;
        RECT 41.130 2.400 42.590 2.680 ;
        RECT 43.430 2.400 44.890 2.680 ;
        RECT 45.730 2.400 47.650 2.680 ;
        RECT 48.490 2.400 49.950 2.680 ;
        RECT 50.790 2.400 52.250 2.680 ;
        RECT 53.090 2.400 54.550 2.680 ;
        RECT 55.390 2.400 56.850 2.680 ;
        RECT 57.690 2.400 59.150 2.680 ;
        RECT 59.990 2.400 61.450 2.680 ;
        RECT 62.290 2.400 63.750 2.680 ;
        RECT 64.590 2.400 66.050 2.680 ;
        RECT 66.890 2.400 68.350 2.680 ;
        RECT 69.190 2.400 71.110 2.680 ;
        RECT 71.950 2.400 73.410 2.680 ;
        RECT 74.250 2.400 75.710 2.680 ;
        RECT 76.550 2.400 78.010 2.680 ;
        RECT 78.850 2.400 80.310 2.680 ;
        RECT 81.150 2.400 82.610 2.680 ;
        RECT 83.450 2.400 84.910 2.680 ;
        RECT 85.750 2.400 87.210 2.680 ;
        RECT 88.050 2.400 89.510 2.680 ;
        RECT 90.350 2.400 91.810 2.680 ;
        RECT 92.650 2.400 94.570 2.680 ;
        RECT 95.410 2.400 96.870 2.680 ;
        RECT 97.710 2.400 99.170 2.680 ;
        RECT 100.010 2.400 101.470 2.680 ;
        RECT 102.310 2.400 103.770 2.680 ;
        RECT 104.610 2.400 106.070 2.680 ;
        RECT 106.910 2.400 108.370 2.680 ;
        RECT 109.210 2.400 110.670 2.680 ;
        RECT 111.510 2.400 112.970 2.680 ;
      LAYER met3 ;
        RECT 2.800 112.520 112.600 113.385 ;
        RECT 2.400 111.200 112.600 112.520 ;
        RECT 2.800 109.800 112.600 111.200 ;
        RECT 2.400 109.160 112.600 109.800 ;
        RECT 2.800 107.760 112.600 109.160 ;
        RECT 2.400 106.440 112.600 107.760 ;
        RECT 2.800 105.040 112.600 106.440 ;
        RECT 2.400 104.400 112.600 105.040 ;
        RECT 2.800 103.000 112.600 104.400 ;
        RECT 2.400 101.680 112.600 103.000 ;
        RECT 2.800 100.280 112.600 101.680 ;
        RECT 2.400 99.640 112.600 100.280 ;
        RECT 2.800 98.240 112.600 99.640 ;
        RECT 2.400 96.920 112.600 98.240 ;
        RECT 2.800 96.240 112.600 96.920 ;
        RECT 2.800 95.520 112.200 96.240 ;
        RECT 2.400 94.880 112.200 95.520 ;
        RECT 2.800 94.840 112.200 94.880 ;
        RECT 2.800 93.480 112.600 94.840 ;
        RECT 2.400 92.160 112.600 93.480 ;
        RECT 2.800 90.760 112.600 92.160 ;
        RECT 2.400 90.120 112.600 90.760 ;
        RECT 2.800 88.720 112.600 90.120 ;
        RECT 2.400 87.400 112.600 88.720 ;
        RECT 2.800 86.000 112.600 87.400 ;
        RECT 2.400 85.360 112.600 86.000 ;
        RECT 2.800 83.960 112.600 85.360 ;
        RECT 2.400 82.640 112.600 83.960 ;
        RECT 2.800 81.240 112.600 82.640 ;
        RECT 2.400 80.600 112.600 81.240 ;
        RECT 2.800 79.200 112.600 80.600 ;
        RECT 2.400 77.880 112.600 79.200 ;
        RECT 2.800 76.480 112.600 77.880 ;
        RECT 2.400 75.840 112.600 76.480 ;
        RECT 2.800 74.440 112.600 75.840 ;
        RECT 2.400 73.120 112.600 74.440 ;
        RECT 2.800 71.720 112.600 73.120 ;
        RECT 2.400 71.080 112.600 71.720 ;
        RECT 2.800 69.680 112.600 71.080 ;
        RECT 2.400 68.360 112.600 69.680 ;
        RECT 2.800 66.960 112.600 68.360 ;
        RECT 2.400 66.320 112.600 66.960 ;
        RECT 2.800 64.920 112.600 66.320 ;
        RECT 2.400 63.600 112.600 64.920 ;
        RECT 2.800 62.200 112.600 63.600 ;
        RECT 2.400 61.560 112.600 62.200 ;
        RECT 2.800 60.160 112.600 61.560 ;
        RECT 2.400 58.840 112.600 60.160 ;
        RECT 2.800 58.160 112.600 58.840 ;
        RECT 2.800 57.440 112.200 58.160 ;
        RECT 2.400 56.760 112.200 57.440 ;
        RECT 2.400 56.120 112.600 56.760 ;
        RECT 2.800 54.720 112.600 56.120 ;
        RECT 2.400 54.080 112.600 54.720 ;
        RECT 2.800 52.680 112.600 54.080 ;
        RECT 2.400 51.360 112.600 52.680 ;
        RECT 2.800 49.960 112.600 51.360 ;
        RECT 2.400 49.320 112.600 49.960 ;
        RECT 2.800 47.920 112.600 49.320 ;
        RECT 2.400 46.600 112.600 47.920 ;
        RECT 2.800 45.200 112.600 46.600 ;
        RECT 2.400 44.560 112.600 45.200 ;
        RECT 2.800 43.160 112.600 44.560 ;
        RECT 2.400 41.840 112.600 43.160 ;
        RECT 2.800 40.440 112.600 41.840 ;
        RECT 2.400 39.800 112.600 40.440 ;
        RECT 2.800 38.400 112.600 39.800 ;
        RECT 2.400 37.080 112.600 38.400 ;
        RECT 2.800 35.680 112.600 37.080 ;
        RECT 2.400 35.040 112.600 35.680 ;
        RECT 2.800 33.640 112.600 35.040 ;
        RECT 2.400 32.320 112.600 33.640 ;
        RECT 2.800 30.920 112.600 32.320 ;
        RECT 2.400 30.280 112.600 30.920 ;
        RECT 2.800 28.880 112.600 30.280 ;
        RECT 2.400 27.560 112.600 28.880 ;
        RECT 2.800 26.160 112.600 27.560 ;
        RECT 2.400 25.520 112.600 26.160 ;
        RECT 2.800 24.120 112.600 25.520 ;
        RECT 2.400 22.800 112.600 24.120 ;
        RECT 2.800 21.400 112.600 22.800 ;
        RECT 2.400 20.760 112.600 21.400 ;
        RECT 2.800 20.080 112.600 20.760 ;
        RECT 2.800 19.360 112.200 20.080 ;
        RECT 2.400 18.680 112.200 19.360 ;
        RECT 2.400 18.040 112.600 18.680 ;
        RECT 2.800 16.640 112.600 18.040 ;
        RECT 2.400 16.000 112.600 16.640 ;
        RECT 2.800 14.600 112.600 16.000 ;
        RECT 2.400 13.280 112.600 14.600 ;
        RECT 2.800 11.880 112.600 13.280 ;
        RECT 2.400 11.240 112.600 11.880 ;
        RECT 2.800 9.840 112.600 11.240 ;
        RECT 2.400 8.520 112.600 9.840 ;
        RECT 2.800 7.120 112.600 8.520 ;
        RECT 2.400 6.480 112.600 7.120 ;
        RECT 2.800 5.080 112.600 6.480 ;
        RECT 2.400 3.760 112.600 5.080 ;
        RECT 2.800 2.360 112.600 3.760 ;
        RECT 2.400 1.720 112.600 2.360 ;
        RECT 2.800 0.860 112.600 1.720 ;
      LAYER met4 ;
        RECT 7.655 10.240 21.645 103.600 ;
        RECT 24.045 10.240 38.975 103.600 ;
        RECT 41.375 10.240 96.305 103.600 ;
        RECT 7.655 0.855 96.305 10.240 ;
      LAYER met5 ;
        RECT 15.300 45.100 46.340 46.700 ;
  END
END sb_2__1_
END LIBRARY

