VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_3__1_
  CLASS BLOCK ;
  FOREIGN sb_3__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 137.930 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.830 137.600 78.110 140.000 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.510 137.600 81.790 140.000 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.650 137.600 85.930 140.000 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.790 137.600 90.070 140.000 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.470 137.600 93.750 140.000 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.610 137.600 97.890 140.000 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.750 137.600 102.030 140.000 ;
    END
  END address[6]
  PIN bottom_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 2.400 ;
    END
  END bottom_left_grid_pin_13_
  PIN bottom_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 2.400 ;
    END
  END bottom_right_grid_pin_11_
  PIN bottom_right_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 2.400 ;
    END
  END bottom_right_grid_pin_13_
  PIN bottom_right_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 2.400 ;
    END
  END bottom_right_grid_pin_15_
  PIN bottom_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 2.400 ;
    END
  END bottom_right_grid_pin_1_
  PIN bottom_right_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 2.400 ;
    END
  END bottom_right_grid_pin_3_
  PIN bottom_right_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 2.400 ;
    END
  END bottom_right_grid_pin_5_
  PIN bottom_right_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 2.400 ;
    END
  END bottom_right_grid_pin_7_
  PIN bottom_right_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 2.400 ;
    END
  END bottom_right_grid_pin_9_
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 2.400 4.040 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 2.400 10.840 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 2.400 17.640 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 2.400 24.440 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 2.400 31.920 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 2.400 38.720 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 2.400 45.520 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 2.400 53.000 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 2.400 59.800 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 2.400 80.880 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 2.400 87.680 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 2.400 94.480 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 2.400 101.960 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 2.400 108.760 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 2.400 115.560 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 2.400 123.040 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 2.400 129.840 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 2.400 136.640 ;
    END
  END chanx_left_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.930 137.600 2.210 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 137.600 5.890 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 137.600 10.030 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 137.600 14.170 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 137.600 17.850 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 137.600 21.990 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.850 137.600 26.130 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 137.600 29.810 140.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.670 137.600 33.950 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.430 137.600 105.710 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.570 137.600 109.850 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.710 137.600 113.990 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.390 137.600 117.670 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.530 137.600 121.810 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 125.670 137.600 125.950 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.350 137.600 129.630 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 133.490 137.600 133.770 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.630 137.600 137.910 140.000 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.690 137.600 73.970 140.000 ;
    END
  END enable
  PIN left_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 2.400 74.080 ;
    END
  END left_bottom_grid_pin_12_
  PIN left_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 2.400 66.600 ;
    END
  END left_top_grid_pin_10_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.810 137.600 38.090 140.000 ;
    END
  END top_left_grid_pin_13_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.730 137.600 62.010 140.000 ;
    END
  END top_right_grid_pin_11_
  PIN top_right_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.410 137.600 65.690 140.000 ;
    END
  END top_right_grid_pin_13_
  PIN top_right_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 137.600 69.830 140.000 ;
    END
  END top_right_grid_pin_15_
  PIN top_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.490 137.600 41.770 140.000 ;
    END
  END top_right_grid_pin_1_
  PIN top_right_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 137.600 45.910 140.000 ;
    END
  END top_right_grid_pin_3_
  PIN top_right_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 137.600 50.050 140.000 ;
    END
  END top_right_grid_pin_5_
  PIN top_right_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.450 137.600 53.730 140.000 ;
    END
  END top_right_grid_pin_7_
  PIN top_right_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.590 137.600 57.870 140.000 ;
    END
  END top_right_grid_pin_9_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 0.070 4.120 137.930 128.080 ;
      LAYER met2 ;
        RECT 0.100 137.320 1.650 137.770 ;
        RECT 2.490 137.320 5.330 137.770 ;
        RECT 6.170 137.320 9.470 137.770 ;
        RECT 10.310 137.320 13.610 137.770 ;
        RECT 14.450 137.320 17.290 137.770 ;
        RECT 18.130 137.320 21.430 137.770 ;
        RECT 22.270 137.320 25.570 137.770 ;
        RECT 26.410 137.320 29.250 137.770 ;
        RECT 30.090 137.320 33.390 137.770 ;
        RECT 34.230 137.320 37.530 137.770 ;
        RECT 38.370 137.320 41.210 137.770 ;
        RECT 42.050 137.320 45.350 137.770 ;
        RECT 46.190 137.320 49.490 137.770 ;
        RECT 50.330 137.320 53.170 137.770 ;
        RECT 54.010 137.320 57.310 137.770 ;
        RECT 58.150 137.320 61.450 137.770 ;
        RECT 62.290 137.320 65.130 137.770 ;
        RECT 65.970 137.320 69.270 137.770 ;
        RECT 70.110 137.320 73.410 137.770 ;
        RECT 74.250 137.320 77.550 137.770 ;
        RECT 78.390 137.320 81.230 137.770 ;
        RECT 82.070 137.320 85.370 137.770 ;
        RECT 86.210 137.320 89.510 137.770 ;
        RECT 90.350 137.320 93.190 137.770 ;
        RECT 94.030 137.320 97.330 137.770 ;
        RECT 98.170 137.320 101.470 137.770 ;
        RECT 102.310 137.320 105.150 137.770 ;
        RECT 105.990 137.320 109.290 137.770 ;
        RECT 110.130 137.320 113.430 137.770 ;
        RECT 114.270 137.320 117.110 137.770 ;
        RECT 117.950 137.320 121.250 137.770 ;
        RECT 122.090 137.320 125.390 137.770 ;
        RECT 126.230 137.320 129.070 137.770 ;
        RECT 129.910 137.320 133.210 137.770 ;
        RECT 134.050 137.320 137.350 137.770 ;
        RECT 0.100 2.680 137.900 137.320 ;
        RECT 0.100 0.270 2.110 2.680 ;
        RECT 2.950 0.270 6.710 2.680 ;
        RECT 7.550 0.270 11.770 2.680 ;
        RECT 12.610 0.270 16.830 2.680 ;
        RECT 17.670 0.270 21.890 2.680 ;
        RECT 22.730 0.270 26.950 2.680 ;
        RECT 27.790 0.270 32.010 2.680 ;
        RECT 32.850 0.270 37.070 2.680 ;
        RECT 37.910 0.270 41.670 2.680 ;
        RECT 42.510 0.270 46.730 2.680 ;
        RECT 47.570 0.270 51.790 2.680 ;
        RECT 52.630 0.270 56.850 2.680 ;
        RECT 57.690 0.270 61.910 2.680 ;
        RECT 62.750 0.270 66.970 2.680 ;
        RECT 67.810 0.270 72.030 2.680 ;
        RECT 72.870 0.270 76.630 2.680 ;
        RECT 77.470 0.270 81.690 2.680 ;
        RECT 82.530 0.270 86.750 2.680 ;
        RECT 87.590 0.270 91.810 2.680 ;
        RECT 92.650 0.270 96.870 2.680 ;
        RECT 97.710 0.270 101.930 2.680 ;
        RECT 102.770 0.270 106.990 2.680 ;
        RECT 107.830 0.270 111.590 2.680 ;
        RECT 112.430 0.270 116.650 2.680 ;
        RECT 117.490 0.270 121.710 2.680 ;
        RECT 122.550 0.270 126.770 2.680 ;
        RECT 127.610 0.270 131.830 2.680 ;
        RECT 132.670 0.270 136.890 2.680 ;
        RECT 137.730 0.270 137.900 2.680 ;
      LAYER met3 ;
        RECT 2.800 135.640 133.795 136.040 ;
        RECT 0.270 130.240 133.795 135.640 ;
        RECT 2.800 128.840 133.795 130.240 ;
        RECT 0.270 123.440 133.795 128.840 ;
        RECT 2.800 122.040 133.795 123.440 ;
        RECT 0.270 115.960 133.795 122.040 ;
        RECT 2.800 114.560 133.795 115.960 ;
        RECT 0.270 109.160 133.795 114.560 ;
        RECT 2.800 107.760 133.795 109.160 ;
        RECT 0.270 102.360 133.795 107.760 ;
        RECT 2.800 100.960 133.795 102.360 ;
        RECT 0.270 94.880 133.795 100.960 ;
        RECT 2.800 93.480 133.795 94.880 ;
        RECT 0.270 88.080 133.795 93.480 ;
        RECT 2.800 86.680 133.795 88.080 ;
        RECT 0.270 81.280 133.795 86.680 ;
        RECT 2.800 79.880 133.795 81.280 ;
        RECT 0.270 74.480 133.795 79.880 ;
        RECT 2.800 73.080 133.795 74.480 ;
        RECT 0.270 67.000 133.795 73.080 ;
        RECT 2.800 65.600 133.795 67.000 ;
        RECT 0.270 60.200 133.795 65.600 ;
        RECT 2.800 58.800 133.795 60.200 ;
        RECT 0.270 53.400 133.795 58.800 ;
        RECT 2.800 52.000 133.795 53.400 ;
        RECT 0.270 45.920 133.795 52.000 ;
        RECT 2.800 44.520 133.795 45.920 ;
        RECT 0.270 39.120 133.795 44.520 ;
        RECT 2.800 37.720 133.795 39.120 ;
        RECT 0.270 32.320 133.795 37.720 ;
        RECT 2.800 30.920 133.795 32.320 ;
        RECT 0.270 24.840 133.795 30.920 ;
        RECT 2.800 23.440 133.795 24.840 ;
        RECT 0.270 18.040 133.795 23.440 ;
        RECT 2.800 16.640 133.795 18.040 ;
        RECT 0.270 11.240 133.795 16.640 ;
        RECT 2.800 9.840 133.795 11.240 ;
        RECT 0.270 4.440 133.795 9.840 ;
        RECT 2.800 4.040 133.795 4.440 ;
      LAYER met4 ;
        RECT 0.295 10.640 27.655 128.080 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 122.985 128.080 ;
  END
END sb_3__1_
END LIBRARY

