magic
tech sky130A
magscale 1 2
timestamp 1604669221
<< locali >>
rect 9873 18207 9907 18309
rect 9137 16983 9171 17153
rect 3341 5083 3375 5321
rect 4905 5015 4939 5253
<< viali >>
rect 1409 25313 1443 25347
rect 2513 25313 2547 25347
rect 1593 25177 1627 25211
rect 2237 25109 2271 25143
rect 2697 25109 2731 25143
rect 3157 25109 3191 25143
rect 3525 25109 3559 25143
rect 4353 25109 4387 25143
rect 2421 24905 2455 24939
rect 2053 24769 2087 24803
rect 3249 24769 3283 24803
rect 4813 24769 4847 24803
rect 1409 24701 1443 24735
rect 2973 24701 3007 24735
rect 3709 24701 3743 24735
rect 4629 24701 4663 24735
rect 16037 24701 16071 24735
rect 16589 24701 16623 24735
rect 4077 24633 4111 24667
rect 4537 24633 4571 24667
rect 1593 24565 1627 24599
rect 2605 24565 2639 24599
rect 3065 24565 3099 24599
rect 4169 24565 4203 24599
rect 7205 24565 7239 24599
rect 7481 24565 7515 24599
rect 7849 24565 7883 24599
rect 16221 24565 16255 24599
rect 1869 24361 1903 24395
rect 2421 24361 2455 24395
rect 3433 24361 3467 24395
rect 6377 24361 6411 24395
rect 10793 24361 10827 24395
rect 14289 24361 14323 24395
rect 15485 24361 15519 24395
rect 16681 24361 16715 24395
rect 18981 24361 19015 24395
rect 21097 24361 21131 24395
rect 2881 24293 2915 24327
rect 6285 24293 6319 24327
rect 1409 24225 1443 24259
rect 2789 24225 2823 24259
rect 4537 24225 4571 24259
rect 7849 24225 7883 24259
rect 10609 24225 10643 24259
rect 12081 24225 12115 24259
rect 14105 24225 14139 24259
rect 15301 24225 15335 24259
rect 16497 24225 16531 24259
rect 17601 24225 17635 24259
rect 18797 24225 18831 24259
rect 20913 24225 20947 24259
rect 3065 24157 3099 24191
rect 4629 24157 4663 24191
rect 4813 24157 4847 24191
rect 6561 24157 6595 24191
rect 7941 24157 7975 24191
rect 8125 24157 8159 24191
rect 3893 24089 3927 24123
rect 5917 24089 5951 24123
rect 12265 24089 12299 24123
rect 17785 24089 17819 24123
rect 2329 24021 2363 24055
rect 4169 24021 4203 24055
rect 5273 24021 5307 24055
rect 7113 24021 7147 24055
rect 7481 24021 7515 24055
rect 2053 23817 2087 23851
rect 3157 23817 3191 23851
rect 3709 23817 3743 23851
rect 5641 23817 5675 23851
rect 6193 23817 6227 23851
rect 13093 23817 13127 23851
rect 13737 23817 13771 23851
rect 14473 23817 14507 23851
rect 18337 23817 18371 23851
rect 19533 23817 19567 23851
rect 21281 23817 21315 23851
rect 23857 23817 23891 23851
rect 4169 23749 4203 23783
rect 6561 23749 6595 23783
rect 15209 23749 15243 23783
rect 16957 23749 16991 23783
rect 2605 23681 2639 23715
rect 2697 23681 2731 23715
rect 2513 23613 2547 23647
rect 4261 23613 4295 23647
rect 7113 23613 7147 23647
rect 10609 23613 10643 23647
rect 11253 23613 11287 23647
rect 11805 23613 11839 23647
rect 12449 23613 12483 23647
rect 13829 23613 13863 23647
rect 15025 23613 15059 23647
rect 16773 23613 16807 23647
rect 17325 23613 17359 23647
rect 18153 23613 18187 23647
rect 19349 23613 19383 23647
rect 19901 23613 19935 23647
rect 21097 23613 21131 23647
rect 21649 23613 21683 23647
rect 23673 23613 23707 23647
rect 24225 23613 24259 23647
rect 1685 23545 1719 23579
rect 4528 23545 4562 23579
rect 7380 23545 7414 23579
rect 2145 23477 2179 23511
rect 8493 23477 8527 23511
rect 9045 23477 9079 23511
rect 11437 23477 11471 23511
rect 12173 23477 12207 23511
rect 12633 23477 12667 23511
rect 14013 23477 14047 23511
rect 14841 23477 14875 23511
rect 15577 23477 15611 23511
rect 16589 23477 16623 23511
rect 17693 23477 17727 23511
rect 18705 23477 18739 23511
rect 19073 23477 19107 23511
rect 20913 23477 20947 23511
rect 3157 23273 3191 23307
rect 6009 23273 6043 23307
rect 9873 23273 9907 23307
rect 14013 23273 14047 23307
rect 17233 23273 17267 23307
rect 18337 23273 18371 23307
rect 21097 23273 21131 23307
rect 22569 23273 22603 23307
rect 2881 23205 2915 23239
rect 5089 23205 5123 23239
rect 6552 23205 6586 23239
rect 2145 23137 2179 23171
rect 4353 23137 4387 23171
rect 9689 23137 9723 23171
rect 12725 23137 12759 23171
rect 13829 23137 13863 23171
rect 15301 23137 15335 23171
rect 17049 23137 17083 23171
rect 18153 23137 18187 23171
rect 20913 23137 20947 23171
rect 22385 23137 22419 23171
rect 2237 23069 2271 23103
rect 2421 23069 2455 23103
rect 5181 23069 5215 23103
rect 5365 23069 5399 23103
rect 6285 23069 6319 23103
rect 1685 23001 1719 23035
rect 3893 23001 3927 23035
rect 12909 23001 12943 23035
rect 1777 22933 1811 22967
rect 4721 22933 4755 22967
rect 7665 22933 7699 22967
rect 8493 22933 8527 22967
rect 13645 22933 13679 22967
rect 14289 22933 14323 22967
rect 15485 22933 15519 22967
rect 2053 22729 2087 22763
rect 2605 22729 2639 22763
rect 4813 22729 4847 22763
rect 6193 22729 6227 22763
rect 6561 22729 6595 22763
rect 15669 22729 15703 22763
rect 16773 22729 16807 22763
rect 20913 22729 20947 22763
rect 6837 22661 6871 22695
rect 8401 22661 8435 22695
rect 2697 22593 2731 22627
rect 5641 22593 5675 22627
rect 5825 22593 5859 22627
rect 7297 22593 7331 22627
rect 7481 22593 7515 22627
rect 7941 22593 7975 22627
rect 8953 22593 8987 22627
rect 14197 22593 14231 22627
rect 1409 22525 1443 22559
rect 2964 22525 2998 22559
rect 5549 22525 5583 22559
rect 7205 22525 7239 22559
rect 8769 22525 8803 22559
rect 15485 22525 15519 22559
rect 16037 22525 16071 22559
rect 16589 22525 16623 22559
rect 13369 22457 13403 22491
rect 14013 22457 14047 22491
rect 15393 22457 15427 22491
rect 1593 22389 1627 22423
rect 4077 22389 4111 22423
rect 5181 22389 5215 22423
rect 8217 22389 8251 22423
rect 8861 22389 8895 22423
rect 9689 22389 9723 22423
rect 10885 22389 10919 22423
rect 12817 22389 12851 22423
rect 13553 22389 13587 22423
rect 13921 22389 13955 22423
rect 14657 22389 14691 22423
rect 17049 22389 17083 22423
rect 17509 22389 17543 22423
rect 18245 22389 18279 22423
rect 22385 22389 22419 22423
rect 5641 22185 5675 22219
rect 6009 22185 6043 22219
rect 8033 22185 8067 22219
rect 10885 22185 10919 22219
rect 13277 22185 13311 22219
rect 13737 22185 13771 22219
rect 4445 22117 4479 22151
rect 12357 22117 12391 22151
rect 1676 22049 1710 22083
rect 3893 22049 3927 22083
rect 5273 22049 5307 22083
rect 6837 22049 6871 22083
rect 15557 22049 15591 22083
rect 1409 21981 1443 22015
rect 3525 21981 3559 22015
rect 4537 21981 4571 22015
rect 4629 21981 4663 22015
rect 6929 21981 6963 22015
rect 7113 21981 7147 22015
rect 10977 21981 11011 22015
rect 11069 21981 11103 22015
rect 13829 21981 13863 22015
rect 13921 21981 13955 22015
rect 15301 21981 15335 22015
rect 2789 21913 2823 21947
rect 4077 21913 4111 21947
rect 6469 21913 6503 21947
rect 7573 21913 7607 21947
rect 10517 21913 10551 21947
rect 16681 21913 16715 21947
rect 6377 21845 6411 21879
rect 7849 21845 7883 21879
rect 9045 21845 9079 21879
rect 10333 21845 10367 21879
rect 11529 21845 11563 21879
rect 13369 21845 13403 21879
rect 14473 21845 14507 21879
rect 1685 21641 1719 21675
rect 2145 21641 2179 21675
rect 4721 21641 4755 21675
rect 10609 21641 10643 21675
rect 13553 21641 13587 21675
rect 15577 21641 15611 21675
rect 2237 21505 2271 21539
rect 5365 21505 5399 21539
rect 5457 21505 5491 21539
rect 7665 21505 7699 21539
rect 8033 21505 8067 21539
rect 9505 21505 9539 21539
rect 11345 21505 11379 21539
rect 13001 21505 13035 21539
rect 6101 21437 6135 21471
rect 11161 21437 11195 21471
rect 12265 21437 12299 21471
rect 12817 21437 12851 21471
rect 14197 21437 14231 21471
rect 2482 21369 2516 21403
rect 4445 21369 4479 21403
rect 7389 21369 7423 21403
rect 8401 21369 8435 21403
rect 8861 21369 8895 21403
rect 9413 21369 9447 21403
rect 10241 21369 10275 21403
rect 11897 21369 11931 21403
rect 14442 21369 14476 21403
rect 3617 21301 3651 21335
rect 4905 21301 4939 21335
rect 5273 21301 5307 21335
rect 6561 21301 6595 21335
rect 7021 21301 7055 21335
rect 7481 21301 7515 21335
rect 8953 21301 8987 21335
rect 9321 21301 9355 21335
rect 10793 21301 10827 21335
rect 11253 21301 11287 21335
rect 12449 21301 12483 21335
rect 12909 21301 12943 21335
rect 14105 21301 14139 21335
rect 16129 21301 16163 21335
rect 1685 21097 1719 21131
rect 2329 21097 2363 21131
rect 2605 21097 2639 21131
rect 3525 21097 3559 21131
rect 5733 21097 5767 21131
rect 6285 21097 6319 21131
rect 7481 21097 7515 21131
rect 9045 21097 9079 21131
rect 13461 21097 13495 21131
rect 13645 21097 13679 21131
rect 15577 21097 15611 21131
rect 9956 21029 9990 21063
rect 13093 21029 13127 21063
rect 4721 20961 4755 20995
rect 7849 20961 7883 20995
rect 9689 20961 9723 20995
rect 12165 20961 12199 20995
rect 14013 20961 14047 20995
rect 14105 20961 14139 20995
rect 3801 20893 3835 20927
rect 4813 20893 4847 20927
rect 4905 20893 4939 20927
rect 6377 20893 6411 20927
rect 6469 20893 6503 20927
rect 7941 20893 7975 20927
rect 8125 20893 8159 20927
rect 12633 20893 12667 20927
rect 14289 20893 14323 20927
rect 5917 20825 5951 20859
rect 7297 20825 7331 20859
rect 4353 20757 4387 20791
rect 5365 20757 5399 20791
rect 7021 20757 7055 20791
rect 8493 20757 8527 20791
rect 11069 20757 11103 20791
rect 11621 20757 11655 20791
rect 12357 20757 12391 20791
rect 2329 20553 2363 20587
rect 4813 20553 4847 20587
rect 5549 20553 5583 20587
rect 6285 20553 6319 20587
rect 7205 20553 7239 20587
rect 8769 20553 8803 20587
rect 9321 20553 9355 20587
rect 11253 20553 11287 20587
rect 11897 20553 11931 20587
rect 15209 20553 15243 20587
rect 3341 20417 3375 20451
rect 3433 20417 3467 20451
rect 1501 20349 1535 20383
rect 2973 20349 3007 20383
rect 7389 20349 7423 20383
rect 9873 20349 9907 20383
rect 10129 20349 10163 20383
rect 12265 20349 12299 20383
rect 12449 20349 12483 20383
rect 3678 20281 3712 20315
rect 7656 20281 7690 20315
rect 12694 20281 12728 20315
rect 14473 20281 14507 20315
rect 1685 20213 1719 20247
rect 2053 20213 2087 20247
rect 6009 20213 6043 20247
rect 9781 20213 9815 20247
rect 13829 20213 13863 20247
rect 14749 20213 14783 20247
rect 2973 20009 3007 20043
rect 3525 20009 3559 20043
rect 6929 20009 6963 20043
rect 7757 20009 7791 20043
rect 8033 20009 8067 20043
rect 8585 20009 8619 20043
rect 10241 20009 10275 20043
rect 11897 20009 11931 20043
rect 3893 19941 3927 19975
rect 4344 19941 4378 19975
rect 9229 19941 9263 19975
rect 10784 19941 10818 19975
rect 1409 19873 1443 19907
rect 4077 19873 4111 19907
rect 7021 19873 7055 19907
rect 13737 19873 13771 19907
rect 14749 19873 14783 19907
rect 7113 19805 7147 19839
rect 9965 19805 9999 19839
rect 10517 19805 10551 19839
rect 12725 19805 12759 19839
rect 13829 19805 13863 19839
rect 13921 19805 13955 19839
rect 2053 19737 2087 19771
rect 1593 19669 1627 19703
rect 5457 19669 5491 19703
rect 6561 19669 6595 19703
rect 8493 19669 8527 19703
rect 13093 19669 13127 19703
rect 13369 19669 13403 19703
rect 14381 19669 14415 19703
rect 3341 19465 3375 19499
rect 6193 19465 6227 19499
rect 7665 19465 7699 19499
rect 10609 19465 10643 19499
rect 9137 19397 9171 19431
rect 12633 19397 12667 19431
rect 4445 19329 4479 19363
rect 8125 19329 8159 19363
rect 8309 19329 8343 19363
rect 9873 19329 9907 19363
rect 11437 19329 11471 19363
rect 13185 19329 13219 19363
rect 1409 19261 1443 19295
rect 2421 19261 2455 19295
rect 2513 19261 2547 19295
rect 3709 19261 3743 19295
rect 4169 19261 4203 19295
rect 5181 19261 5215 19295
rect 5365 19261 5399 19295
rect 6653 19261 6687 19295
rect 9597 19261 9631 19295
rect 11161 19261 11195 19295
rect 13093 19261 13127 19295
rect 14197 19261 14231 19295
rect 14464 19261 14498 19295
rect 11897 19193 11931 19227
rect 13737 19193 13771 19227
rect 1593 19125 1627 19159
rect 2053 19125 2087 19159
rect 2697 19125 2731 19159
rect 3801 19125 3835 19159
rect 4261 19125 4295 19159
rect 4813 19125 4847 19159
rect 7021 19125 7055 19159
rect 7573 19125 7607 19159
rect 8033 19125 8067 19159
rect 8677 19125 8711 19159
rect 9229 19125 9263 19159
rect 9689 19125 9723 19159
rect 10793 19125 10827 19159
rect 11253 19125 11287 19159
rect 12265 19125 12299 19159
rect 13001 19125 13035 19159
rect 14013 19125 14047 19159
rect 15577 19125 15611 19159
rect 1961 18921 1995 18955
rect 2697 18921 2731 18955
rect 3157 18921 3191 18955
rect 3893 18921 3927 18955
rect 4537 18921 4571 18955
rect 4997 18921 5031 18955
rect 6101 18921 6135 18955
rect 7481 18921 7515 18955
rect 8125 18921 8159 18955
rect 9321 18921 9355 18955
rect 11253 18921 11287 18955
rect 11805 18921 11839 18955
rect 14657 18921 14691 18955
rect 3525 18853 3559 18887
rect 4353 18853 4387 18887
rect 4905 18853 4939 18887
rect 6469 18853 6503 18887
rect 10057 18853 10091 18887
rect 12081 18853 12115 18887
rect 12992 18853 13026 18887
rect 1409 18785 1443 18819
rect 2513 18785 2547 18819
rect 8033 18785 8067 18819
rect 11161 18785 11195 18819
rect 12725 18785 12759 18819
rect 5089 18717 5123 18751
rect 6561 18717 6595 18751
rect 6653 18717 6687 18751
rect 8217 18717 8251 18751
rect 10149 18717 10183 18751
rect 10333 18717 10367 18751
rect 15301 18717 15335 18751
rect 14105 18649 14139 18683
rect 1593 18581 1627 18615
rect 2421 18581 2455 18615
rect 7113 18581 7147 18615
rect 7665 18581 7699 18615
rect 9689 18581 9723 18615
rect 10701 18581 10735 18615
rect 12541 18581 12575 18615
rect 2513 18377 2547 18411
rect 3801 18377 3835 18411
rect 8493 18377 8527 18411
rect 10977 18377 11011 18411
rect 14013 18377 14047 18411
rect 9413 18309 9447 18343
rect 9873 18309 9907 18343
rect 13829 18309 13863 18343
rect 15025 18309 15059 18343
rect 2237 18241 2271 18275
rect 3157 18241 3191 18275
rect 3341 18241 3375 18275
rect 10517 18241 10551 18275
rect 12265 18241 12299 18275
rect 12909 18241 12943 18275
rect 13001 18241 13035 18275
rect 14565 18241 14599 18275
rect 1409 18173 1443 18207
rect 3065 18173 3099 18207
rect 4261 18173 4295 18207
rect 4517 18173 4551 18207
rect 7113 18173 7147 18207
rect 9873 18173 9907 18207
rect 10333 18173 10367 18207
rect 11897 18173 11931 18207
rect 14381 18173 14415 18207
rect 6285 18105 6319 18139
rect 7380 18105 7414 18139
rect 9781 18105 9815 18139
rect 1593 18037 1627 18071
rect 2697 18037 2731 18071
rect 4169 18037 4203 18071
rect 5641 18037 5675 18071
rect 6561 18037 6595 18071
rect 9965 18037 9999 18071
rect 10425 18037 10459 18071
rect 11345 18037 11379 18071
rect 12449 18037 12483 18071
rect 12817 18037 12851 18071
rect 13461 18037 13495 18071
rect 14473 18037 14507 18071
rect 2789 17833 2823 17867
rect 4077 17833 4111 17867
rect 4537 17833 4571 17867
rect 5181 17833 5215 17867
rect 6193 17833 6227 17867
rect 12357 17833 12391 17867
rect 13001 17833 13035 17867
rect 13921 17833 13955 17867
rect 14473 17833 14507 17867
rect 2237 17765 2271 17799
rect 3893 17765 3927 17799
rect 5641 17765 5675 17799
rect 11244 17765 11278 17799
rect 1409 17697 1443 17731
rect 4445 17697 4479 17731
rect 6920 17697 6954 17731
rect 9965 17697 9999 17731
rect 13829 17697 13863 17731
rect 2881 17629 2915 17663
rect 3065 17629 3099 17663
rect 3525 17629 3559 17663
rect 4721 17629 4755 17663
rect 6653 17629 6687 17663
rect 10977 17629 11011 17663
rect 14013 17629 14047 17663
rect 10149 17561 10183 17595
rect 1961 17493 1995 17527
rect 2421 17493 2455 17527
rect 5549 17493 5583 17527
rect 6469 17493 6503 17527
rect 8033 17493 8067 17527
rect 8677 17493 8711 17527
rect 10517 17493 10551 17527
rect 13277 17493 13311 17527
rect 13461 17493 13495 17527
rect 4905 17289 4939 17323
rect 5273 17289 5307 17323
rect 6285 17289 6319 17323
rect 7941 17289 7975 17323
rect 11345 17289 11379 17323
rect 14657 17289 14691 17323
rect 7389 17153 7423 17187
rect 8861 17153 8895 17187
rect 9137 17153 9171 17187
rect 9413 17153 9447 17187
rect 1409 17085 1443 17119
rect 2881 17085 2915 17119
rect 2973 17085 3007 17119
rect 3240 17085 3274 17119
rect 5457 17085 5491 17119
rect 7205 17085 7239 17119
rect 8401 17085 8435 17119
rect 2513 17017 2547 17051
rect 8309 17017 8343 17051
rect 13277 17085 13311 17119
rect 9658 17017 9692 17051
rect 12817 17017 12851 17051
rect 13544 17017 13578 17051
rect 1593 16949 1627 16983
rect 2145 16949 2179 16983
rect 4353 16949 4387 16983
rect 5641 16949 5675 16983
rect 6561 16949 6595 16983
rect 6837 16949 6871 16983
rect 7297 16949 7331 16983
rect 8585 16949 8619 16983
rect 9137 16949 9171 16983
rect 9229 16949 9263 16983
rect 10793 16949 10827 16983
rect 11713 16949 11747 16983
rect 13093 16949 13127 16983
rect 1593 16745 1627 16779
rect 2053 16745 2087 16779
rect 2421 16745 2455 16779
rect 2697 16745 2731 16779
rect 3157 16745 3191 16779
rect 4445 16745 4479 16779
rect 5641 16745 5675 16779
rect 6009 16745 6043 16779
rect 7205 16745 7239 16779
rect 8217 16745 8251 16779
rect 8677 16745 8711 16779
rect 9505 16745 9539 16779
rect 9689 16745 9723 16779
rect 10149 16745 10183 16779
rect 10793 16745 10827 16779
rect 13093 16745 13127 16779
rect 14013 16745 14047 16779
rect 4537 16677 4571 16711
rect 7665 16677 7699 16711
rect 13645 16677 13679 16711
rect 1409 16609 1443 16643
rect 2513 16609 2547 16643
rect 3433 16609 3467 16643
rect 5089 16609 5123 16643
rect 5549 16609 5583 16643
rect 6745 16609 6779 16643
rect 7573 16609 7607 16643
rect 10057 16609 10091 16643
rect 11980 16609 12014 16643
rect 4721 16541 4755 16575
rect 6101 16541 6135 16575
rect 6285 16541 6319 16575
rect 7849 16541 7883 16575
rect 10241 16541 10275 16575
rect 11713 16541 11747 16575
rect 3893 16473 3927 16507
rect 4077 16405 4111 16439
rect 7021 16405 7055 16439
rect 2053 16201 2087 16235
rect 4813 16201 4847 16235
rect 5273 16201 5307 16235
rect 5641 16201 5675 16235
rect 11161 16201 11195 16235
rect 12081 16201 12115 16235
rect 11713 16133 11747 16167
rect 2421 16065 2455 16099
rect 7113 16065 7147 16099
rect 9781 16065 9815 16099
rect 12449 16065 12483 16099
rect 1409 15997 1443 16031
rect 2881 15997 2915 16031
rect 3137 15997 3171 16031
rect 7369 15997 7403 16031
rect 9689 15997 9723 16031
rect 10048 15997 10082 16031
rect 13737 15997 13771 16031
rect 13982 15929 14016 15963
rect 1593 15861 1627 15895
rect 2789 15861 2823 15895
rect 4261 15861 4295 15895
rect 5733 15861 5767 15895
rect 6285 15861 6319 15895
rect 6653 15861 6687 15895
rect 8493 15861 8527 15895
rect 9229 15861 9263 15895
rect 13645 15861 13679 15895
rect 15117 15861 15151 15895
rect 1593 15657 1627 15691
rect 1869 15657 1903 15691
rect 2329 15657 2363 15691
rect 2789 15657 2823 15691
rect 2881 15657 2915 15691
rect 4261 15657 4295 15691
rect 4537 15657 4571 15691
rect 5273 15657 5307 15691
rect 7113 15657 7147 15691
rect 7757 15657 7791 15691
rect 8033 15657 8067 15691
rect 9505 15657 9539 15691
rect 10241 15657 10275 15691
rect 10793 15657 10827 15691
rect 11253 15657 11287 15691
rect 12357 15657 12391 15691
rect 13829 15657 13863 15691
rect 14381 15657 14415 15691
rect 3893 15589 3927 15623
rect 11161 15589 11195 15623
rect 12725 15589 12759 15623
rect 15117 15589 15151 15623
rect 15761 15589 15795 15623
rect 1409 15521 1443 15555
rect 4077 15521 4111 15555
rect 5733 15521 5767 15555
rect 6000 15521 6034 15555
rect 9965 15521 9999 15555
rect 14197 15521 14231 15555
rect 15669 15521 15703 15555
rect 3065 15453 3099 15487
rect 8585 15453 8619 15487
rect 11437 15453 11471 15487
rect 12817 15453 12851 15487
rect 13001 15453 13035 15487
rect 15945 15453 15979 15487
rect 3433 15385 3467 15419
rect 14657 15385 14691 15419
rect 2421 15317 2455 15351
rect 5641 15317 5675 15351
rect 8401 15317 8435 15351
rect 9045 15317 9079 15351
rect 15301 15317 15335 15351
rect 16497 15317 16531 15351
rect 2053 15113 2087 15147
rect 3525 15113 3559 15147
rect 5181 15113 5215 15147
rect 6653 15113 6687 15147
rect 8493 15113 8527 15147
rect 10057 15113 10091 15147
rect 10885 15113 10919 15147
rect 11253 15113 11287 15147
rect 11621 15113 11655 15147
rect 12265 15113 12299 15147
rect 13093 15113 13127 15147
rect 16405 15113 16439 15147
rect 2421 15045 2455 15079
rect 3801 15045 3835 15079
rect 4169 15045 4203 15079
rect 4721 14977 4755 15011
rect 5733 14977 5767 15011
rect 7389 14977 7423 15011
rect 8677 14977 8711 15011
rect 17049 14977 17083 15011
rect 1409 14909 1443 14943
rect 2513 14909 2547 14943
rect 3617 14909 3651 14943
rect 5549 14909 5583 14943
rect 7205 14909 7239 14943
rect 7297 14909 7331 14943
rect 13921 14909 13955 14943
rect 3157 14841 3191 14875
rect 5089 14841 5123 14875
rect 5641 14841 5675 14875
rect 8922 14841 8956 14875
rect 13461 14841 13495 14875
rect 14166 14841 14200 14875
rect 16865 14841 16899 14875
rect 1593 14773 1627 14807
rect 2697 14773 2731 14807
rect 6193 14773 6227 14807
rect 6837 14773 6871 14807
rect 7849 14773 7883 14807
rect 12725 14773 12759 14807
rect 13829 14773 13863 14807
rect 15301 14773 15335 14807
rect 15853 14773 15887 14807
rect 16221 14773 16255 14807
rect 16773 14773 16807 14807
rect 1593 14569 1627 14603
rect 3617 14569 3651 14603
rect 5457 14569 5491 14603
rect 6009 14569 6043 14603
rect 7941 14569 7975 14603
rect 9689 14569 9723 14603
rect 10149 14569 10183 14603
rect 14105 14569 14139 14603
rect 15761 14569 15795 14603
rect 16865 14569 16899 14603
rect 6806 14501 6840 14535
rect 1409 14433 1443 14467
rect 2789 14433 2823 14467
rect 4077 14433 4111 14467
rect 4344 14433 4378 14467
rect 9505 14433 9539 14467
rect 10057 14433 10091 14467
rect 12992 14433 13026 14467
rect 15025 14433 15059 14467
rect 15669 14433 15703 14467
rect 17233 14433 17267 14467
rect 2881 14365 2915 14399
rect 3065 14365 3099 14399
rect 6561 14365 6595 14399
rect 10333 14365 10367 14399
rect 12725 14365 12759 14399
rect 15853 14365 15887 14399
rect 16405 14365 16439 14399
rect 17325 14365 17359 14399
rect 17509 14365 17543 14399
rect 2329 14297 2363 14331
rect 1869 14229 1903 14263
rect 2421 14229 2455 14263
rect 6377 14229 6411 14263
rect 8769 14229 8803 14263
rect 9137 14229 9171 14263
rect 12541 14229 12575 14263
rect 14657 14229 14691 14263
rect 15301 14229 15335 14263
rect 4445 14025 4479 14059
rect 4997 14025 5031 14059
rect 5181 14025 5215 14059
rect 6193 14025 6227 14059
rect 6837 14025 6871 14059
rect 9413 14025 9447 14059
rect 9781 14025 9815 14059
rect 9965 14025 9999 14059
rect 11069 14025 11103 14059
rect 13277 14025 13311 14059
rect 1593 13957 1627 13991
rect 2881 13957 2915 13991
rect 8401 13957 8435 13991
rect 11345 13957 11379 13991
rect 12817 13957 12851 13991
rect 3341 13889 3375 13923
rect 3525 13889 3559 13923
rect 5641 13889 5675 13923
rect 5825 13889 5859 13923
rect 7389 13889 7423 13923
rect 7941 13889 7975 13923
rect 9045 13889 9079 13923
rect 10517 13889 10551 13923
rect 12265 13889 12299 13923
rect 13185 13889 13219 13923
rect 13921 13889 13955 13923
rect 1409 13821 1443 13855
rect 2421 13821 2455 13855
rect 4169 13821 4203 13855
rect 6653 13821 6687 13855
rect 7297 13821 7331 13855
rect 8309 13821 8343 13855
rect 8861 13821 8895 13855
rect 10425 13821 10459 13855
rect 14289 13821 14323 13855
rect 14749 13821 14783 13855
rect 14841 13821 14875 13855
rect 15108 13821 15142 13855
rect 16865 13821 16899 13855
rect 17233 13821 17267 13855
rect 3249 13753 3283 13787
rect 10333 13753 10367 13787
rect 2145 13685 2179 13719
rect 5549 13685 5583 13719
rect 7205 13685 7239 13719
rect 8769 13685 8803 13719
rect 13645 13685 13679 13719
rect 13737 13685 13771 13719
rect 16221 13685 16255 13719
rect 17693 13685 17727 13719
rect 1593 13481 1627 13515
rect 2237 13481 2271 13515
rect 2789 13481 2823 13515
rect 4077 13481 4111 13515
rect 4445 13481 4479 13515
rect 6009 13481 6043 13515
rect 6653 13481 6687 13515
rect 7205 13481 7239 13515
rect 7665 13481 7699 13515
rect 9413 13481 9447 13515
rect 10057 13481 10091 13515
rect 10701 13481 10735 13515
rect 11253 13481 11287 13515
rect 11713 13481 11747 13515
rect 13185 13481 13219 13515
rect 13553 13481 13587 13515
rect 14013 13481 14047 13515
rect 14933 13481 14967 13515
rect 16313 13481 16347 13515
rect 2881 13413 2915 13447
rect 3893 13413 3927 13447
rect 6101 13413 6135 13447
rect 18236 13413 18270 13447
rect 1409 13345 1443 13379
rect 1961 13345 1995 13379
rect 4537 13345 4571 13379
rect 7113 13345 7147 13379
rect 7573 13345 7607 13379
rect 11621 13345 11655 13379
rect 15669 13345 15703 13379
rect 17969 13345 18003 13379
rect 2973 13277 3007 13311
rect 4721 13277 4755 13311
rect 6285 13277 6319 13311
rect 7757 13277 7791 13311
rect 10149 13277 10183 13311
rect 10333 13277 10367 13311
rect 11897 13277 11931 13311
rect 14105 13277 14139 13311
rect 14289 13277 14323 13311
rect 15761 13277 15795 13311
rect 15945 13277 15979 13311
rect 16681 13277 16715 13311
rect 3525 13209 3559 13243
rect 5641 13209 5675 13243
rect 9137 13209 9171 13243
rect 13645 13209 13679 13243
rect 2421 13141 2455 13175
rect 5273 13141 5307 13175
rect 8401 13141 8435 13175
rect 9689 13141 9723 13175
rect 11069 13141 11103 13175
rect 12449 13141 12483 13175
rect 12817 13141 12851 13175
rect 15301 13141 15335 13175
rect 19349 13141 19383 13175
rect 1961 12937 1995 12971
rect 4997 12937 5031 12971
rect 5181 12937 5215 12971
rect 6193 12937 6227 12971
rect 6561 12937 6595 12971
rect 7849 12937 7883 12971
rect 8309 12937 8343 12971
rect 8953 12937 8987 12971
rect 11345 12937 11379 12971
rect 11989 12937 12023 12971
rect 12449 12937 12483 12971
rect 14013 12937 14047 12971
rect 15025 12937 15059 12971
rect 17417 12937 17451 12971
rect 18245 12937 18279 12971
rect 18613 12937 18647 12971
rect 4169 12869 4203 12903
rect 2053 12801 2087 12835
rect 5733 12801 5767 12835
rect 7481 12801 7515 12835
rect 9045 12801 9079 12835
rect 11621 12801 11655 12835
rect 13093 12801 13127 12835
rect 14473 12801 14507 12835
rect 2309 12733 2343 12767
rect 4445 12733 4479 12767
rect 7205 12733 7239 12767
rect 12817 12733 12851 12767
rect 13645 12733 13679 12767
rect 15393 12733 15427 12767
rect 15485 12733 15519 12767
rect 15752 12733 15786 12767
rect 9290 12665 9324 12699
rect 3433 12597 3467 12631
rect 5549 12597 5583 12631
rect 5641 12597 5675 12631
rect 6837 12597 6871 12631
rect 7297 12597 7331 12631
rect 10425 12597 10459 12631
rect 12909 12597 12943 12631
rect 16865 12597 16899 12631
rect 3709 12393 3743 12427
rect 5273 12393 5307 12427
rect 7389 12393 7423 12427
rect 7665 12393 7699 12427
rect 8309 12393 8343 12427
rect 9045 12393 9079 12427
rect 9413 12393 9447 12427
rect 9689 12393 9723 12427
rect 12541 12393 12575 12427
rect 13185 12393 13219 12427
rect 15577 12393 15611 12427
rect 16313 12393 16347 12427
rect 1676 12325 1710 12359
rect 10057 12325 10091 12359
rect 13277 12325 13311 12359
rect 14289 12325 14323 12359
rect 4077 12257 4111 12291
rect 5621 12257 5655 12291
rect 8217 12257 8251 12291
rect 10149 12257 10183 12291
rect 10701 12257 10735 12291
rect 11621 12257 11655 12291
rect 11713 12257 11747 12291
rect 15025 12257 15059 12291
rect 16221 12257 16255 12291
rect 17785 12257 17819 12291
rect 1409 12189 1443 12223
rect 5365 12189 5399 12223
rect 8401 12189 8435 12223
rect 10241 12189 10275 12223
rect 11897 12189 11931 12223
rect 13369 12189 13403 12223
rect 16405 12189 16439 12223
rect 17877 12189 17911 12223
rect 17969 12189 18003 12223
rect 18797 12189 18831 12223
rect 7849 12121 7883 12155
rect 11253 12121 11287 12155
rect 12817 12121 12851 12155
rect 16865 12121 16899 12155
rect 2789 12053 2823 12087
rect 3433 12053 3467 12087
rect 4261 12053 4295 12087
rect 4721 12053 4755 12087
rect 6745 12053 6779 12087
rect 11069 12053 11103 12087
rect 13829 12053 13863 12087
rect 14749 12053 14783 12087
rect 15853 12053 15887 12087
rect 17417 12053 17451 12087
rect 18429 12053 18463 12087
rect 1593 11849 1627 11883
rect 4813 11849 4847 11883
rect 5549 11849 5583 11883
rect 6193 11849 6227 11883
rect 8769 11849 8803 11883
rect 9137 11849 9171 11883
rect 9321 11849 9355 11883
rect 11253 11849 11287 11883
rect 13921 11849 13955 11883
rect 14473 11849 14507 11883
rect 16497 11849 16531 11883
rect 17785 11849 17819 11883
rect 19165 11849 19199 11883
rect 5825 11781 5859 11815
rect 10885 11781 10919 11815
rect 16037 11781 16071 11815
rect 2421 11713 2455 11747
rect 9873 11713 9907 11747
rect 15577 11713 15611 11747
rect 18521 11713 18555 11747
rect 18613 11713 18647 11747
rect 1409 11645 1443 11679
rect 2881 11645 2915 11679
rect 3148 11645 3182 11679
rect 5365 11645 5399 11679
rect 6561 11645 6595 11679
rect 6837 11645 6871 11679
rect 7093 11645 7127 11679
rect 9781 11645 9815 11679
rect 11805 11645 11839 11679
rect 12173 11645 12207 11679
rect 12541 11645 12575 11679
rect 17049 11645 17083 11679
rect 18429 11645 18463 11679
rect 12808 11577 12842 11611
rect 15393 11577 15427 11611
rect 2053 11509 2087 11543
rect 2697 11509 2731 11543
rect 4261 11509 4295 11543
rect 5273 11509 5307 11543
rect 8217 11509 8251 11543
rect 9689 11509 9723 11543
rect 10425 11509 10459 11543
rect 11345 11509 11379 11543
rect 14841 11509 14875 11543
rect 15025 11509 15059 11543
rect 15485 11509 15519 11543
rect 17509 11509 17543 11543
rect 18061 11509 18095 11543
rect 2421 11305 2455 11339
rect 3433 11305 3467 11339
rect 3893 11305 3927 11339
rect 4261 11305 4295 11339
rect 5273 11305 5307 11339
rect 6837 11305 6871 11339
rect 8309 11305 8343 11339
rect 8953 11305 8987 11339
rect 9413 11305 9447 11339
rect 9965 11305 9999 11339
rect 11805 11305 11839 11339
rect 12909 11305 12943 11339
rect 13369 11305 13403 11339
rect 17509 11305 17543 11339
rect 18061 11305 18095 11339
rect 5724 11237 5758 11271
rect 7481 11237 7515 11271
rect 7849 11237 7883 11271
rect 10670 11237 10704 11271
rect 13277 11237 13311 11271
rect 14657 11237 14691 11271
rect 18521 11237 18555 11271
rect 2789 11169 2823 11203
rect 4077 11169 4111 11203
rect 4537 11169 4571 11203
rect 5457 11169 5491 11203
rect 10425 11169 10459 11203
rect 15833 11169 15867 11203
rect 18429 11169 18463 11203
rect 1409 11101 1443 11135
rect 1869 11101 1903 11135
rect 2881 11101 2915 11135
rect 3065 11101 3099 11135
rect 8401 11101 8435 11135
rect 8493 11101 8527 11135
rect 13553 11101 13587 11135
rect 15025 11101 15059 11135
rect 15577 11101 15611 11135
rect 18705 11101 18739 11135
rect 7941 11033 7975 11067
rect 13921 11033 13955 11067
rect 14289 11033 14323 11067
rect 16957 11033 16991 11067
rect 2329 10965 2363 10999
rect 4997 10965 5031 10999
rect 10333 10965 10367 10999
rect 12541 10965 12575 10999
rect 1409 10761 1443 10795
rect 3157 10761 3191 10795
rect 3249 10761 3283 10795
rect 5181 10761 5215 10795
rect 6193 10761 6227 10795
rect 6653 10761 6687 10795
rect 9229 10761 9263 10795
rect 9781 10761 9815 10795
rect 11713 10761 11747 10795
rect 13461 10761 13495 10795
rect 14013 10761 14047 10795
rect 15117 10761 15151 10795
rect 16681 10761 16715 10795
rect 18061 10761 18095 10795
rect 7665 10693 7699 10727
rect 10333 10693 10367 10727
rect 13829 10693 13863 10727
rect 15485 10693 15519 10727
rect 16957 10693 16991 10727
rect 1869 10625 1903 10659
rect 2053 10625 2087 10659
rect 3709 10625 3743 10659
rect 3893 10625 3927 10659
rect 4721 10625 4755 10659
rect 5089 10625 5123 10659
rect 5825 10625 5859 10659
rect 7849 10625 7883 10659
rect 10885 10625 10919 10659
rect 13093 10625 13127 10659
rect 14473 10625 14507 10659
rect 14565 10625 14599 10659
rect 16037 10625 16071 10659
rect 16129 10625 16163 10659
rect 17509 10625 17543 10659
rect 18613 10625 18647 10659
rect 1777 10557 1811 10591
rect 2789 10557 2823 10591
rect 3617 10557 3651 10591
rect 5549 10557 5583 10591
rect 12173 10557 12207 10591
rect 12909 10557 12943 10591
rect 14381 10557 14415 10591
rect 15945 10557 15979 10591
rect 7297 10489 7331 10523
rect 8116 10489 8150 10523
rect 10793 10489 10827 10523
rect 11345 10489 11379 10523
rect 12817 10489 12851 10523
rect 18521 10489 18555 10523
rect 19073 10489 19107 10523
rect 4261 10421 4295 10455
rect 5641 10421 5675 10455
rect 10149 10421 10183 10455
rect 10701 10421 10735 10455
rect 12449 10421 12483 10455
rect 15577 10421 15611 10455
rect 17785 10421 17819 10455
rect 18429 10421 18463 10455
rect 1777 10217 1811 10251
rect 4261 10217 4295 10251
rect 4905 10217 4939 10251
rect 5457 10217 5491 10251
rect 7849 10217 7883 10251
rect 8493 10217 8527 10251
rect 9413 10217 9447 10251
rect 11069 10217 11103 10251
rect 12817 10217 12851 10251
rect 14013 10217 14047 10251
rect 14749 10217 14783 10251
rect 17417 10217 17451 10251
rect 18521 10217 18555 10251
rect 3525 10149 3559 10183
rect 5917 10149 5951 10183
rect 11621 10149 11655 10183
rect 12541 10149 12575 10183
rect 14381 10149 14415 10183
rect 16282 10149 16316 10183
rect 5825 10081 5859 10115
rect 8401 10081 8435 10115
rect 9945 10081 9979 10115
rect 13185 10081 13219 10115
rect 1869 10013 1903 10047
rect 2053 10013 2087 10047
rect 6009 10013 6043 10047
rect 7205 10013 7239 10047
rect 8677 10013 8711 10047
rect 9689 10013 9723 10047
rect 13277 10013 13311 10047
rect 13461 10013 13495 10047
rect 16037 10013 16071 10047
rect 1409 9945 1443 9979
rect 6561 9945 6595 9979
rect 8033 9945 8067 9979
rect 18153 9945 18187 9979
rect 2421 9877 2455 9911
rect 3065 9877 3099 9911
rect 3893 9877 3927 9911
rect 5273 9877 5307 9911
rect 6929 9877 6963 9911
rect 9045 9877 9079 9911
rect 11989 9877 12023 9911
rect 15669 9877 15703 9911
rect 18797 9877 18831 9911
rect 1409 9673 1443 9707
rect 6837 9673 6871 9707
rect 8493 9673 8527 9707
rect 9781 9673 9815 9707
rect 2421 9605 2455 9639
rect 5089 9605 5123 9639
rect 8125 9605 8159 9639
rect 8677 9605 8711 9639
rect 10609 9605 10643 9639
rect 12265 9605 12299 9639
rect 15209 9605 15243 9639
rect 16313 9605 16347 9639
rect 2053 9537 2087 9571
rect 3065 9537 3099 9571
rect 5457 9537 5491 9571
rect 5549 9537 5583 9571
rect 7389 9537 7423 9571
rect 9137 9537 9171 9571
rect 9321 9537 9355 9571
rect 10333 9537 10367 9571
rect 11345 9537 11379 9571
rect 16865 9537 16899 9571
rect 17325 9537 17359 9571
rect 1777 9469 1811 9503
rect 3332 9469 3366 9503
rect 9045 9469 9079 9503
rect 11253 9469 11287 9503
rect 13829 9469 13863 9503
rect 16681 9469 16715 9503
rect 18245 9469 18279 9503
rect 6653 9401 6687 9435
rect 7297 9401 7331 9435
rect 12909 9401 12943 9435
rect 14074 9401 14108 9435
rect 16773 9401 16807 9435
rect 1869 9333 1903 9367
rect 2789 9333 2823 9367
rect 4445 9333 4479 9367
rect 6009 9333 6043 9367
rect 7205 9333 7239 9367
rect 10793 9333 10827 9367
rect 11161 9333 11195 9367
rect 11805 9333 11839 9367
rect 13369 9333 13403 9367
rect 13737 9333 13771 9367
rect 16129 9333 16163 9367
rect 17693 9333 17727 9367
rect 2881 9129 2915 9163
rect 3525 9129 3559 9163
rect 4537 9129 4571 9163
rect 7757 9129 7791 9163
rect 8677 9129 8711 9163
rect 11253 9129 11287 9163
rect 16405 9129 16439 9163
rect 4445 9061 4479 9095
rect 10149 9061 10183 9095
rect 14933 9061 14967 9095
rect 16856 9061 16890 9095
rect 1768 8993 1802 9027
rect 6377 8993 6411 9027
rect 6644 8993 6678 9027
rect 10057 8993 10091 9027
rect 12061 8993 12095 9027
rect 16589 8993 16623 9027
rect 1501 8925 1535 8959
rect 3893 8925 3927 8959
rect 4629 8925 4663 8959
rect 5089 8925 5123 8959
rect 5549 8925 5583 8959
rect 10241 8925 10275 8959
rect 11805 8925 11839 8959
rect 15577 8925 15611 8959
rect 4077 8857 4111 8891
rect 9137 8857 9171 8891
rect 9505 8857 9539 8891
rect 5825 8789 5859 8823
rect 6285 8789 6319 8823
rect 8401 8789 8435 8823
rect 9689 8789 9723 8823
rect 10885 8789 10919 8823
rect 11621 8789 11655 8823
rect 13185 8789 13219 8823
rect 13921 8789 13955 8823
rect 14197 8789 14231 8823
rect 14565 8789 14599 8823
rect 16129 8789 16163 8823
rect 17969 8789 18003 8823
rect 2697 8585 2731 8619
rect 6837 8585 6871 8619
rect 7849 8585 7883 8619
rect 10057 8585 10091 8619
rect 10609 8585 10643 8619
rect 14381 8585 14415 8619
rect 15301 8585 15335 8619
rect 15577 8585 15611 8619
rect 15761 8585 15795 8619
rect 17233 8585 17267 8619
rect 1685 8449 1719 8483
rect 3341 8449 3375 8483
rect 7389 8449 7423 8483
rect 11345 8449 11379 8483
rect 16221 8449 16255 8483
rect 16405 8449 16439 8483
rect 4169 8381 4203 8415
rect 4261 8381 4295 8415
rect 6653 8381 6687 8415
rect 7205 8381 7239 8415
rect 8585 8381 8619 8415
rect 8677 8381 8711 8415
rect 13001 8381 13035 8415
rect 16129 8381 16163 8415
rect 2145 8313 2179 8347
rect 3065 8313 3099 8347
rect 3801 8313 3835 8347
rect 4506 8313 4540 8347
rect 8922 8313 8956 8347
rect 11069 8313 11103 8347
rect 11897 8313 11931 8347
rect 12909 8313 12943 8347
rect 13246 8313 13280 8347
rect 17509 8313 17543 8347
rect 2605 8245 2639 8279
rect 3157 8245 3191 8279
rect 5641 8245 5675 8279
rect 6285 8245 6319 8279
rect 7297 8245 7331 8279
rect 12265 8245 12299 8279
rect 16773 8245 16807 8279
rect 1777 8041 1811 8075
rect 2789 8041 2823 8075
rect 5917 8041 5951 8075
rect 9413 8041 9447 8075
rect 9689 8041 9723 8075
rect 11713 8041 11747 8075
rect 12081 8041 12115 8075
rect 13277 8041 13311 8075
rect 13645 8041 13679 8075
rect 16589 8041 16623 8075
rect 17693 8041 17727 8075
rect 4721 7973 4755 8007
rect 6377 7973 6411 8007
rect 9045 7973 9079 8007
rect 13737 7973 13771 8007
rect 14289 7973 14323 8007
rect 4813 7905 4847 7939
rect 6285 7905 6319 7939
rect 8401 7905 8435 7939
rect 8493 7905 8527 7939
rect 10057 7905 10091 7939
rect 16497 7905 16531 7939
rect 18061 7905 18095 7939
rect 1869 7837 1903 7871
rect 2053 7837 2087 7871
rect 3893 7837 3927 7871
rect 4905 7837 4939 7871
rect 6561 7837 6595 7871
rect 8585 7837 8619 7871
rect 10149 7837 10183 7871
rect 10241 7837 10275 7871
rect 12173 7837 12207 7871
rect 12265 7837 12299 7871
rect 13093 7837 13127 7871
rect 13921 7837 13955 7871
rect 16681 7837 16715 7871
rect 18153 7837 18187 7871
rect 18245 7837 18279 7871
rect 8033 7769 8067 7803
rect 14749 7769 14783 7803
rect 16129 7769 16163 7803
rect 17601 7769 17635 7803
rect 19717 7769 19751 7803
rect 1409 7701 1443 7735
rect 3157 7701 3191 7735
rect 3525 7701 3559 7735
rect 4353 7701 4387 7735
rect 5365 7701 5399 7735
rect 5825 7701 5859 7735
rect 6929 7701 6963 7735
rect 7297 7701 7331 7735
rect 7665 7701 7699 7735
rect 10885 7701 10919 7735
rect 11253 7701 11287 7735
rect 11529 7701 11563 7735
rect 15117 7701 15151 7735
rect 15761 7701 15795 7735
rect 17141 7701 17175 7735
rect 19993 7701 20027 7735
rect 1409 7497 1443 7531
rect 4997 7497 5031 7531
rect 5181 7497 5215 7531
rect 8217 7497 8251 7531
rect 8769 7497 8803 7531
rect 10793 7497 10827 7531
rect 11897 7497 11931 7531
rect 13645 7497 13679 7531
rect 15761 7497 15795 7531
rect 16773 7497 16807 7531
rect 3617 7429 3651 7463
rect 4721 7429 4755 7463
rect 9137 7429 9171 7463
rect 13185 7429 13219 7463
rect 17325 7429 17359 7463
rect 2053 7361 2087 7395
rect 4261 7361 4295 7395
rect 5825 7361 5859 7395
rect 11345 7361 11379 7395
rect 13553 7361 13587 7395
rect 14105 7361 14139 7395
rect 14289 7361 14323 7395
rect 16221 7361 16255 7395
rect 16405 7361 16439 7395
rect 18705 7361 18739 7395
rect 19533 7361 19567 7395
rect 20177 7361 20211 7395
rect 1869 7293 1903 7327
rect 5549 7293 5583 7327
rect 6837 7293 6871 7327
rect 10609 7293 10643 7327
rect 11161 7293 11195 7327
rect 14013 7293 14047 7327
rect 15577 7293 15611 7327
rect 16129 7293 16163 7327
rect 17693 7293 17727 7327
rect 18429 7293 18463 7327
rect 18521 7293 18555 7327
rect 19073 7293 19107 7327
rect 1777 7225 1811 7259
rect 2789 7225 2823 7259
rect 3985 7225 4019 7259
rect 7104 7225 7138 7259
rect 9321 7225 9355 7259
rect 10241 7225 10275 7259
rect 11253 7225 11287 7259
rect 19993 7225 20027 7259
rect 2421 7157 2455 7191
rect 3433 7157 3467 7191
rect 4077 7157 4111 7191
rect 5641 7157 5675 7191
rect 6285 7157 6319 7191
rect 6561 7157 6595 7191
rect 9873 7157 9907 7191
rect 12265 7157 12299 7191
rect 12449 7157 12483 7191
rect 14933 7157 14967 7191
rect 15301 7157 15335 7191
rect 18061 7157 18095 7191
rect 19625 7157 19659 7191
rect 20085 7157 20119 7191
rect 1409 6953 1443 6987
rect 1961 6953 1995 6987
rect 4445 6953 4479 6987
rect 9873 6953 9907 6987
rect 13737 6953 13771 6987
rect 15393 6953 15427 6987
rect 16221 6953 16255 6987
rect 18429 6953 18463 6987
rect 19257 6953 19291 6987
rect 2789 6885 2823 6919
rect 11437 6885 11471 6919
rect 6276 6817 6310 6851
rect 8125 6817 8159 6851
rect 8493 6817 8527 6851
rect 13001 6817 13035 6851
rect 14013 6817 14047 6851
rect 14197 6817 14231 6851
rect 16661 6817 16695 6851
rect 19349 6817 19383 6851
rect 22293 6817 22327 6851
rect 2881 6749 2915 6783
rect 3065 6749 3099 6783
rect 4537 6749 4571 6783
rect 4721 6749 4755 6783
rect 6009 6749 6043 6783
rect 11529 6749 11563 6783
rect 11621 6749 11655 6783
rect 12541 6749 12575 6783
rect 13093 6749 13127 6783
rect 13277 6749 13311 6783
rect 16405 6749 16439 6783
rect 19441 6749 19475 6783
rect 19901 6749 19935 6783
rect 5181 6681 5215 6715
rect 10793 6681 10827 6715
rect 12173 6681 12207 6715
rect 15025 6681 15059 6715
rect 18889 6681 18923 6715
rect 21189 6681 21223 6715
rect 2237 6613 2271 6647
rect 2421 6613 2455 6647
rect 3617 6613 3651 6647
rect 4077 6613 4111 6647
rect 5549 6613 5583 6647
rect 7389 6613 7423 6647
rect 8953 6613 8987 6647
rect 9321 6613 9355 6647
rect 10241 6613 10275 6647
rect 11069 6613 11103 6647
rect 12633 6613 12667 6647
rect 14381 6613 14415 6647
rect 14657 6613 14691 6647
rect 17785 6613 17819 6647
rect 18705 6613 18739 6647
rect 20269 6613 20303 6647
rect 21557 6613 21591 6647
rect 22477 6613 22511 6647
rect 1685 6409 1719 6443
rect 2145 6409 2179 6443
rect 4721 6409 4755 6443
rect 6101 6409 6135 6443
rect 6837 6409 6871 6443
rect 7849 6409 7883 6443
rect 8309 6409 8343 6443
rect 8585 6409 8619 6443
rect 9413 6409 9447 6443
rect 15669 6409 15703 6443
rect 17785 6409 17819 6443
rect 18061 6409 18095 6443
rect 19073 6409 19107 6443
rect 21189 6409 21223 6443
rect 22293 6409 22327 6443
rect 2237 6273 2271 6307
rect 5273 6273 5307 6307
rect 6377 6273 6411 6307
rect 7297 6273 7331 6307
rect 7481 6273 7515 6307
rect 9505 6273 9539 6307
rect 13093 6273 13127 6307
rect 18705 6273 18739 6307
rect 19533 6273 19567 6307
rect 20085 6273 20119 6307
rect 20177 6273 20211 6307
rect 20637 6273 20671 6307
rect 21649 6273 21683 6307
rect 21741 6273 21775 6307
rect 7205 6205 7239 6239
rect 11805 6205 11839 6239
rect 12265 6205 12299 6239
rect 12817 6205 12851 6239
rect 14197 6205 14231 6239
rect 14289 6205 14323 6239
rect 14556 6205 14590 6239
rect 16773 6205 16807 6239
rect 18429 6205 18463 6239
rect 19993 6205 20027 6239
rect 2504 6137 2538 6171
rect 4261 6137 4295 6171
rect 5089 6137 5123 6171
rect 9045 6137 9079 6171
rect 9772 6137 9806 6171
rect 17509 6137 17543 6171
rect 18521 6137 18555 6171
rect 21557 6137 21591 6171
rect 3617 6069 3651 6103
rect 4537 6069 4571 6103
rect 5181 6069 5215 6103
rect 10885 6069 10919 6103
rect 11529 6069 11563 6103
rect 12449 6069 12483 6103
rect 12909 6069 12943 6103
rect 13461 6069 13495 6103
rect 16497 6069 16531 6103
rect 16957 6069 16991 6103
rect 19625 6069 19659 6103
rect 21005 6069 21039 6103
rect 5457 5865 5491 5899
rect 6561 5865 6595 5899
rect 7665 5865 7699 5899
rect 8309 5865 8343 5899
rect 11069 5865 11103 5899
rect 11621 5865 11655 5899
rect 12081 5865 12115 5899
rect 14381 5865 14415 5899
rect 15761 5865 15795 5899
rect 16681 5865 16715 5899
rect 19993 5865 20027 5899
rect 20545 5865 20579 5899
rect 20913 5865 20947 5899
rect 21373 5865 21407 5899
rect 1676 5797 1710 5831
rect 6929 5797 6963 5831
rect 17132 5797 17166 5831
rect 1409 5729 1443 5763
rect 4077 5729 4111 5763
rect 4344 5729 4378 5763
rect 7021 5729 7055 5763
rect 8585 5729 8619 5763
rect 9689 5729 9723 5763
rect 9956 5729 9990 5763
rect 12173 5729 12207 5763
rect 12440 5729 12474 5763
rect 15669 5729 15703 5763
rect 16865 5729 16899 5763
rect 19349 5729 19383 5763
rect 21281 5729 21315 5763
rect 23305 5729 23339 5763
rect 7113 5661 7147 5695
rect 15945 5661 15979 5695
rect 21465 5661 21499 5695
rect 2789 5593 2823 5627
rect 9413 5593 9447 5627
rect 14657 5593 14691 5627
rect 15301 5593 15335 5627
rect 19533 5593 19567 5627
rect 3709 5525 3743 5559
rect 6101 5525 6135 5559
rect 6377 5525 6411 5559
rect 7941 5525 7975 5559
rect 13553 5525 13587 5559
rect 15025 5525 15059 5559
rect 16405 5525 16439 5559
rect 18245 5525 18279 5559
rect 18889 5525 18923 5559
rect 23489 5525 23523 5559
rect 3341 5321 3375 5355
rect 3617 5321 3651 5355
rect 4629 5321 4663 5355
rect 8861 5321 8895 5355
rect 10701 5321 10735 5355
rect 12173 5321 12207 5355
rect 13001 5321 13035 5355
rect 14933 5321 14967 5355
rect 15577 5321 15611 5355
rect 15945 5321 15979 5355
rect 16405 5321 16439 5355
rect 19441 5321 19475 5355
rect 21925 5321 21959 5355
rect 23305 5321 23339 5355
rect 1409 5253 1443 5287
rect 1869 5185 1903 5219
rect 2053 5185 2087 5219
rect 1777 5117 1811 5151
rect 2513 5117 2547 5151
rect 3157 5117 3191 5151
rect 4905 5253 4939 5287
rect 9229 5253 9263 5287
rect 13369 5253 13403 5287
rect 20085 5253 20119 5287
rect 22293 5253 22327 5287
rect 4261 5185 4295 5219
rect 3341 5049 3375 5083
rect 5733 5185 5767 5219
rect 9321 5185 9355 5219
rect 11253 5185 11287 5219
rect 13553 5185 13587 5219
rect 16313 5185 16347 5219
rect 16957 5185 16991 5219
rect 21097 5185 21131 5219
rect 6653 5117 6687 5151
rect 6837 5117 6871 5151
rect 9577 5117 9611 5151
rect 12541 5117 12575 5151
rect 16865 5117 16899 5151
rect 17417 5117 17451 5151
rect 18061 5117 18095 5151
rect 18317 5117 18351 5151
rect 21557 5117 21591 5151
rect 22109 5117 22143 5151
rect 22569 5117 22603 5151
rect 5641 5049 5675 5083
rect 6285 5049 6319 5083
rect 7082 5049 7116 5083
rect 11621 5049 11655 5083
rect 13798 5049 13832 5083
rect 16773 5049 16807 5083
rect 17877 5049 17911 5083
rect 3525 4981 3559 5015
rect 3985 4981 4019 5015
rect 4077 4981 4111 5015
rect 4905 4981 4939 5015
rect 4997 4981 5031 5015
rect 5181 4981 5215 5015
rect 5549 4981 5583 5015
rect 8217 4981 8251 5015
rect 12725 4981 12759 5015
rect 20361 4981 20395 5015
rect 20545 4981 20579 5015
rect 20913 4981 20947 5015
rect 21005 4981 21039 5015
rect 1685 4777 1719 4811
rect 2789 4777 2823 4811
rect 4445 4777 4479 4811
rect 6377 4777 6411 4811
rect 7113 4777 7147 4811
rect 7573 4777 7607 4811
rect 8033 4777 8067 4811
rect 8953 4777 8987 4811
rect 9321 4777 9355 4811
rect 10977 4777 11011 4811
rect 11437 4777 11471 4811
rect 13001 4777 13035 4811
rect 15485 4777 15519 4811
rect 16129 4777 16163 4811
rect 17877 4777 17911 4811
rect 21465 4777 21499 4811
rect 6469 4709 6503 4743
rect 10793 4709 10827 4743
rect 11345 4709 11379 4743
rect 12909 4709 12943 4743
rect 14657 4709 14691 4743
rect 15117 4709 15151 4743
rect 18429 4709 18463 4743
rect 19441 4709 19475 4743
rect 2881 4641 2915 4675
rect 4813 4641 4847 4675
rect 4905 4641 4939 4675
rect 5549 4641 5583 4675
rect 7941 4641 7975 4675
rect 9965 4641 9999 4675
rect 12449 4641 12483 4675
rect 13645 4641 13679 4675
rect 14105 4641 14139 4675
rect 15301 4641 15335 4675
rect 16865 4641 16899 4675
rect 17601 4641 17635 4675
rect 18521 4641 18555 4675
rect 19073 4641 19107 4675
rect 19625 4641 19659 4675
rect 20913 4641 20947 4675
rect 3065 4573 3099 4607
rect 5089 4573 5123 4607
rect 5917 4573 5951 4607
rect 6653 4573 6687 4607
rect 8125 4573 8159 4607
rect 10517 4573 10551 4607
rect 11621 4573 11655 4607
rect 13185 4573 13219 4607
rect 16957 4573 16991 4607
rect 17141 4573 17175 4607
rect 18613 4573 18647 4607
rect 20545 4573 20579 4607
rect 3709 4505 3743 4539
rect 6009 4505 6043 4539
rect 8677 4505 8711 4539
rect 12081 4505 12115 4539
rect 18061 4505 18095 4539
rect 21097 4505 21131 4539
rect 2329 4437 2363 4471
rect 2421 4437 2455 4471
rect 4353 4437 4387 4471
rect 7481 4437 7515 4471
rect 10149 4437 10183 4471
rect 12541 4437 12575 4471
rect 13921 4437 13955 4471
rect 14289 4437 14323 4471
rect 16497 4437 16531 4471
rect 19809 4437 19843 4471
rect 20177 4437 20211 4471
rect 21833 4437 21867 4471
rect 3801 4233 3835 4267
rect 6009 4233 6043 4267
rect 6377 4233 6411 4267
rect 7297 4233 7331 4267
rect 10701 4233 10735 4267
rect 11897 4233 11931 4267
rect 13921 4233 13955 4267
rect 15393 4233 15427 4267
rect 16129 4233 16163 4267
rect 18061 4233 18095 4267
rect 20913 4233 20947 4267
rect 11069 4165 11103 4199
rect 14013 4165 14047 4199
rect 1777 4097 1811 4131
rect 2789 4097 2823 4131
rect 2973 4097 3007 4131
rect 8309 4097 8343 4131
rect 8493 4097 8527 4131
rect 8953 4097 8987 4131
rect 10057 4097 10091 4131
rect 12909 4097 12943 4131
rect 13093 4097 13127 4131
rect 14565 4097 14599 4131
rect 16037 4097 16071 4131
rect 16681 4097 16715 4131
rect 18613 4097 18647 4131
rect 19165 4097 19199 4131
rect 20177 4097 20211 4131
rect 3433 4029 3467 4063
rect 3893 4029 3927 4063
rect 7573 4029 7607 4063
rect 9781 4029 9815 4063
rect 11253 4029 11287 4063
rect 12817 4029 12851 4063
rect 13461 4029 13495 4063
rect 14381 4029 14415 4063
rect 16589 4029 16623 4063
rect 19993 4029 20027 4063
rect 21189 4029 21223 4063
rect 21741 4029 21775 4063
rect 22293 4029 22327 4063
rect 22753 4029 22787 4063
rect 2145 3961 2179 3995
rect 4160 3961 4194 3995
rect 8217 3961 8251 3995
rect 9321 3961 9355 3995
rect 9873 3961 9907 3995
rect 12173 3961 12207 3995
rect 14473 3961 14507 3995
rect 18429 3961 18463 3995
rect 20085 3961 20119 3995
rect 2329 3893 2363 3927
rect 2697 3893 2731 3927
rect 5273 3893 5307 3927
rect 7849 3893 7883 3927
rect 9413 3893 9447 3927
rect 11437 3893 11471 3927
rect 12449 3893 12483 3927
rect 16497 3893 16531 3927
rect 17417 3893 17451 3927
rect 17785 3893 17819 3927
rect 18521 3893 18555 3927
rect 19441 3893 19475 3927
rect 19625 3893 19659 3927
rect 21373 3893 21407 3927
rect 22201 3893 22235 3927
rect 22477 3893 22511 3927
rect 1685 3689 1719 3723
rect 2053 3689 2087 3723
rect 2697 3689 2731 3723
rect 3893 3689 3927 3723
rect 5181 3689 5215 3723
rect 8401 3689 8435 3723
rect 9045 3689 9079 3723
rect 9413 3689 9447 3723
rect 9965 3689 9999 3723
rect 10609 3689 10643 3723
rect 11253 3689 11287 3723
rect 11621 3689 11655 3723
rect 14197 3689 14231 3723
rect 15025 3689 15059 3723
rect 15945 3689 15979 3723
rect 18061 3689 18095 3723
rect 18613 3689 18647 3723
rect 18981 3689 19015 3723
rect 19625 3689 19659 3723
rect 20177 3689 20211 3723
rect 3525 3621 3559 3655
rect 4905 3621 4939 3655
rect 5794 3621 5828 3655
rect 7573 3621 7607 3655
rect 10517 3621 10551 3655
rect 11958 3621 11992 3655
rect 14657 3621 14691 3655
rect 2145 3553 2179 3587
rect 5549 3553 5583 3587
rect 15301 3553 15335 3587
rect 16681 3553 16715 3587
rect 16948 3553 16982 3587
rect 19533 3553 19567 3587
rect 21097 3553 21131 3587
rect 21649 3553 21683 3587
rect 22201 3553 22235 3587
rect 2237 3485 2271 3519
rect 8493 3485 8527 3519
rect 8677 3485 8711 3519
rect 10793 3485 10827 3519
rect 11713 3485 11747 3519
rect 19809 3485 19843 3519
rect 6929 3417 6963 3451
rect 15485 3417 15519 3451
rect 20545 3417 20579 3451
rect 3157 3349 3191 3383
rect 4445 3349 4479 3383
rect 8033 3349 8067 3383
rect 10149 3349 10183 3383
rect 13093 3349 13127 3383
rect 13737 3349 13771 3383
rect 14105 3349 14139 3383
rect 16589 3349 16623 3383
rect 19165 3349 19199 3383
rect 21281 3349 21315 3383
rect 22385 3349 22419 3383
rect 4905 3145 4939 3179
rect 6009 3145 6043 3179
rect 6929 3145 6963 3179
rect 9873 3145 9907 3179
rect 10793 3145 10827 3179
rect 11897 3145 11931 3179
rect 12173 3145 12207 3179
rect 17141 3145 17175 3179
rect 17785 3145 17819 3179
rect 18061 3145 18095 3179
rect 19073 3145 19107 3179
rect 20637 3145 20671 3179
rect 21465 3145 21499 3179
rect 22569 3145 22603 3179
rect 23857 3145 23891 3179
rect 3433 3077 3467 3111
rect 8033 3077 8067 3111
rect 10425 3077 10459 3111
rect 16497 3077 16531 3111
rect 19625 3077 19659 3111
rect 21005 3077 21039 3111
rect 4445 3009 4479 3043
rect 5549 3009 5583 3043
rect 7573 3009 7607 3043
rect 12633 3009 12667 3043
rect 17509 3009 17543 3043
rect 18613 3009 18647 3043
rect 20177 3009 20211 3043
rect 2053 2941 2087 2975
rect 2320 2941 2354 2975
rect 4813 2941 4847 2975
rect 5273 2941 5307 2975
rect 7297 2941 7331 2975
rect 8493 2941 8527 2975
rect 8760 2941 8794 2975
rect 11253 2941 11287 2975
rect 14933 2941 14967 2975
rect 15117 2941 15151 2975
rect 18429 2941 18463 2975
rect 20085 2941 20119 2975
rect 21649 2941 21683 2975
rect 22201 2941 22235 2975
rect 23673 2941 23707 2975
rect 24225 2941 24259 2975
rect 4077 2873 4111 2907
rect 5365 2873 5399 2907
rect 6653 2873 6687 2907
rect 7389 2873 7423 2907
rect 12900 2873 12934 2907
rect 14657 2873 14691 2907
rect 15362 2873 15396 2907
rect 18521 2873 18555 2907
rect 19993 2873 20027 2907
rect 1685 2805 1719 2839
rect 11437 2805 11471 2839
rect 14013 2805 14047 2839
rect 19441 2805 19475 2839
rect 21833 2805 21867 2839
rect 2421 2601 2455 2635
rect 3801 2601 3835 2635
rect 6101 2601 6135 2635
rect 7205 2601 7239 2635
rect 8125 2601 8159 2635
rect 9597 2601 9631 2635
rect 10149 2601 10183 2635
rect 10793 2601 10827 2635
rect 11345 2601 11379 2635
rect 12633 2601 12667 2635
rect 13001 2601 13035 2635
rect 13093 2601 13127 2635
rect 14197 2601 14231 2635
rect 15485 2601 15519 2635
rect 16681 2601 16715 2635
rect 18153 2601 18187 2635
rect 18705 2601 18739 2635
rect 18797 2601 18831 2635
rect 1961 2533 1995 2567
rect 2789 2533 2823 2567
rect 7665 2533 7699 2567
rect 8585 2533 8619 2567
rect 10241 2533 10275 2567
rect 12449 2533 12483 2567
rect 4077 2465 4111 2499
rect 4344 2465 4378 2499
rect 8493 2465 8527 2499
rect 9137 2465 9171 2499
rect 11437 2465 11471 2499
rect 14289 2465 14323 2499
rect 14841 2465 14875 2499
rect 15853 2465 15887 2499
rect 17141 2465 17175 2499
rect 17693 2465 17727 2499
rect 19901 2465 19935 2499
rect 20453 2465 20487 2499
rect 21557 2465 21591 2499
rect 22753 2465 22787 2499
rect 23305 2465 23339 2499
rect 23673 2465 23707 2499
rect 24041 2465 24075 2499
rect 24593 2465 24627 2499
rect 1409 2397 1443 2431
rect 2329 2397 2363 2431
rect 2881 2397 2915 2431
rect 3065 2397 3099 2431
rect 3525 2397 3559 2431
rect 7941 2397 7975 2431
rect 8769 2397 8803 2431
rect 10425 2397 10459 2431
rect 11989 2397 12023 2431
rect 13277 2397 13311 2431
rect 13645 2397 13679 2431
rect 15945 2397 15979 2431
rect 16129 2397 16163 2431
rect 18889 2397 18923 2431
rect 21649 2397 21683 2431
rect 21741 2397 21775 2431
rect 9781 2329 9815 2363
rect 18337 2329 18371 2363
rect 22201 2329 22235 2363
rect 22937 2329 22971 2363
rect 5457 2261 5491 2295
rect 6469 2261 6503 2295
rect 11621 2261 11655 2295
rect 14473 2261 14507 2295
rect 15301 2261 15335 2295
rect 16957 2261 16991 2295
rect 17325 2261 17359 2295
rect 19625 2261 19659 2295
rect 20085 2261 20119 2295
rect 20913 2261 20947 2295
rect 21189 2261 21223 2295
rect 22569 2261 22603 2295
rect 24225 2261 24259 2295
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 1854 25344 1860 25356
rect 1443 25316 1860 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 1854 25304 1860 25316
rect 1912 25304 1918 25356
rect 2406 25304 2412 25356
rect 2464 25344 2470 25356
rect 2501 25347 2559 25353
rect 2501 25344 2513 25347
rect 2464 25316 2513 25344
rect 2464 25304 2470 25316
rect 2501 25313 2513 25316
rect 2547 25344 2559 25347
rect 5350 25344 5356 25356
rect 2547 25316 5356 25344
rect 2547 25313 2559 25316
rect 2501 25307 2559 25313
rect 5350 25304 5356 25316
rect 5408 25304 5414 25356
rect 1581 25211 1639 25217
rect 1581 25177 1593 25211
rect 1627 25208 1639 25211
rect 2958 25208 2964 25220
rect 1627 25180 2964 25208
rect 1627 25177 1639 25180
rect 1581 25171 1639 25177
rect 2958 25168 2964 25180
rect 3016 25168 3022 25220
rect 2222 25140 2228 25152
rect 2183 25112 2228 25140
rect 2222 25100 2228 25112
rect 2280 25100 2286 25152
rect 2685 25143 2743 25149
rect 2685 25109 2697 25143
rect 2731 25140 2743 25143
rect 2866 25140 2872 25152
rect 2731 25112 2872 25140
rect 2731 25109 2743 25112
rect 2685 25103 2743 25109
rect 2866 25100 2872 25112
rect 2924 25100 2930 25152
rect 3145 25143 3203 25149
rect 3145 25109 3157 25143
rect 3191 25140 3203 25143
rect 3234 25140 3240 25152
rect 3191 25112 3240 25140
rect 3191 25109 3203 25112
rect 3145 25103 3203 25109
rect 3234 25100 3240 25112
rect 3292 25100 3298 25152
rect 3513 25143 3571 25149
rect 3513 25109 3525 25143
rect 3559 25140 3571 25143
rect 4341 25143 4399 25149
rect 4341 25140 4353 25143
rect 3559 25112 4353 25140
rect 3559 25109 3571 25112
rect 3513 25103 3571 25109
rect 4341 25109 4353 25112
rect 4387 25140 4399 25143
rect 4890 25140 4896 25152
rect 4387 25112 4896 25140
rect 4387 25109 4399 25112
rect 4341 25103 4399 25109
rect 4890 25100 4896 25112
rect 4948 25100 4954 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 2406 24936 2412 24948
rect 2367 24908 2412 24936
rect 2406 24896 2412 24908
rect 2464 24896 2470 24948
rect 4062 24828 4068 24880
rect 4120 24868 4126 24880
rect 6086 24868 6092 24880
rect 4120 24840 6092 24868
rect 4120 24828 4126 24840
rect 6086 24828 6092 24840
rect 6144 24828 6150 24880
rect 2038 24800 2044 24812
rect 1412 24772 2044 24800
rect 1412 24741 1440 24772
rect 2038 24760 2044 24772
rect 2096 24760 2102 24812
rect 3237 24803 3295 24809
rect 3237 24769 3249 24803
rect 3283 24800 3295 24803
rect 4801 24803 4859 24809
rect 4801 24800 4813 24803
rect 3283 24772 4813 24800
rect 3283 24769 3295 24772
rect 3237 24763 3295 24769
rect 4801 24769 4813 24772
rect 4847 24800 4859 24803
rect 4890 24800 4896 24812
rect 4847 24772 4896 24800
rect 4847 24769 4859 24772
rect 4801 24763 4859 24769
rect 4890 24760 4896 24772
rect 4948 24760 4954 24812
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24701 1455 24735
rect 1397 24695 1455 24701
rect 2774 24692 2780 24744
rect 2832 24732 2838 24744
rect 2961 24735 3019 24741
rect 2961 24732 2973 24735
rect 2832 24704 2973 24732
rect 2832 24692 2838 24704
rect 2961 24701 2973 24704
rect 3007 24701 3019 24735
rect 2961 24695 3019 24701
rect 3697 24735 3755 24741
rect 3697 24701 3709 24735
rect 3743 24732 3755 24735
rect 4338 24732 4344 24744
rect 3743 24704 4344 24732
rect 3743 24701 3755 24704
rect 3697 24695 3755 24701
rect 4338 24692 4344 24704
rect 4396 24732 4402 24744
rect 4617 24735 4675 24741
rect 4617 24732 4629 24735
rect 4396 24704 4629 24732
rect 4396 24692 4402 24704
rect 4617 24701 4629 24704
rect 4663 24732 4675 24735
rect 7098 24732 7104 24744
rect 4663 24704 7104 24732
rect 4663 24701 4675 24704
rect 4617 24695 4675 24701
rect 7098 24692 7104 24704
rect 7156 24692 7162 24744
rect 16022 24732 16028 24744
rect 15983 24704 16028 24732
rect 16022 24692 16028 24704
rect 16080 24732 16086 24744
rect 16577 24735 16635 24741
rect 16577 24732 16589 24735
rect 16080 24704 16589 24732
rect 16080 24692 16086 24704
rect 16577 24701 16589 24704
rect 16623 24701 16635 24735
rect 16577 24695 16635 24701
rect 4065 24667 4123 24673
rect 4065 24633 4077 24667
rect 4111 24664 4123 24667
rect 4525 24667 4583 24673
rect 4525 24664 4537 24667
rect 4111 24636 4537 24664
rect 4111 24633 4123 24636
rect 4065 24627 4123 24633
rect 4525 24633 4537 24636
rect 4571 24664 4583 24667
rect 5074 24664 5080 24676
rect 4571 24636 5080 24664
rect 4571 24633 4583 24636
rect 4525 24627 4583 24633
rect 5074 24624 5080 24636
rect 5132 24624 5138 24676
rect 1578 24596 1584 24608
rect 1539 24568 1584 24596
rect 1578 24556 1584 24568
rect 1636 24556 1642 24608
rect 2590 24596 2596 24608
rect 2551 24568 2596 24596
rect 2590 24556 2596 24568
rect 2648 24556 2654 24608
rect 3053 24599 3111 24605
rect 3053 24565 3065 24599
rect 3099 24596 3111 24599
rect 3234 24596 3240 24608
rect 3099 24568 3240 24596
rect 3099 24565 3111 24568
rect 3053 24559 3111 24565
rect 3234 24556 3240 24568
rect 3292 24556 3298 24608
rect 4154 24596 4160 24608
rect 4115 24568 4160 24596
rect 4154 24556 4160 24568
rect 4212 24556 4218 24608
rect 7190 24596 7196 24608
rect 7151 24568 7196 24596
rect 7190 24556 7196 24568
rect 7248 24556 7254 24608
rect 7374 24556 7380 24608
rect 7432 24596 7438 24608
rect 7469 24599 7527 24605
rect 7469 24596 7481 24599
rect 7432 24568 7481 24596
rect 7432 24556 7438 24568
rect 7469 24565 7481 24568
rect 7515 24565 7527 24599
rect 7834 24596 7840 24608
rect 7795 24568 7840 24596
rect 7469 24559 7527 24565
rect 7834 24556 7840 24568
rect 7892 24556 7898 24608
rect 16206 24596 16212 24608
rect 16167 24568 16212 24596
rect 16206 24556 16212 24568
rect 16264 24556 16270 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1854 24392 1860 24404
rect 1815 24364 1860 24392
rect 1854 24352 1860 24364
rect 1912 24352 1918 24404
rect 2222 24352 2228 24404
rect 2280 24392 2286 24404
rect 2409 24395 2467 24401
rect 2409 24392 2421 24395
rect 2280 24364 2421 24392
rect 2280 24352 2286 24364
rect 2409 24361 2421 24364
rect 2455 24361 2467 24395
rect 2409 24355 2467 24361
rect 2774 24352 2780 24404
rect 2832 24392 2838 24404
rect 3421 24395 3479 24401
rect 3421 24392 3433 24395
rect 2832 24364 3433 24392
rect 2832 24352 2838 24364
rect 3421 24361 3433 24364
rect 3467 24392 3479 24395
rect 3510 24392 3516 24404
rect 3467 24364 3516 24392
rect 3467 24361 3479 24364
rect 3421 24355 3479 24361
rect 3510 24352 3516 24364
rect 3568 24352 3574 24404
rect 4798 24352 4804 24404
rect 4856 24392 4862 24404
rect 6178 24392 6184 24404
rect 4856 24364 6184 24392
rect 4856 24352 4862 24364
rect 6178 24352 6184 24364
rect 6236 24392 6242 24404
rect 6365 24395 6423 24401
rect 6365 24392 6377 24395
rect 6236 24364 6377 24392
rect 6236 24352 6242 24364
rect 6365 24361 6377 24364
rect 6411 24361 6423 24395
rect 10778 24392 10784 24404
rect 10739 24364 10784 24392
rect 6365 24355 6423 24361
rect 10778 24352 10784 24364
rect 10836 24352 10842 24404
rect 14274 24392 14280 24404
rect 14235 24364 14280 24392
rect 14274 24352 14280 24364
rect 14332 24352 14338 24404
rect 15473 24395 15531 24401
rect 15473 24361 15485 24395
rect 15519 24392 15531 24395
rect 16482 24392 16488 24404
rect 15519 24364 16488 24392
rect 15519 24361 15531 24364
rect 15473 24355 15531 24361
rect 16482 24352 16488 24364
rect 16540 24352 16546 24404
rect 16669 24395 16727 24401
rect 16669 24361 16681 24395
rect 16715 24392 16727 24395
rect 18506 24392 18512 24404
rect 16715 24364 18512 24392
rect 16715 24361 16727 24364
rect 16669 24355 16727 24361
rect 18506 24352 18512 24364
rect 18564 24352 18570 24404
rect 18966 24392 18972 24404
rect 18927 24364 18972 24392
rect 18966 24352 18972 24364
rect 19024 24352 19030 24404
rect 21085 24395 21143 24401
rect 21085 24361 21097 24395
rect 21131 24392 21143 24395
rect 22462 24392 22468 24404
rect 21131 24364 22468 24392
rect 21131 24361 21143 24364
rect 21085 24355 21143 24361
rect 22462 24352 22468 24364
rect 22520 24352 22526 24404
rect 2869 24327 2927 24333
rect 2869 24293 2881 24327
rect 2915 24324 2927 24327
rect 3050 24324 3056 24336
rect 2915 24296 3056 24324
rect 2915 24293 2927 24296
rect 2869 24287 2927 24293
rect 3050 24284 3056 24296
rect 3108 24284 3114 24336
rect 4246 24284 4252 24336
rect 4304 24324 4310 24336
rect 4706 24324 4712 24336
rect 4304 24296 4712 24324
rect 4304 24284 4310 24296
rect 4706 24284 4712 24296
rect 4764 24284 4770 24336
rect 5994 24284 6000 24336
rect 6052 24324 6058 24336
rect 6273 24327 6331 24333
rect 6273 24324 6285 24327
rect 6052 24296 6285 24324
rect 6052 24284 6058 24296
rect 6273 24293 6285 24296
rect 6319 24293 6331 24327
rect 6273 24287 6331 24293
rect 1397 24259 1455 24265
rect 1397 24225 1409 24259
rect 1443 24256 1455 24259
rect 2038 24256 2044 24268
rect 1443 24228 2044 24256
rect 1443 24225 1455 24228
rect 1397 24219 1455 24225
rect 2038 24216 2044 24228
rect 2096 24256 2102 24268
rect 2777 24259 2835 24265
rect 2777 24256 2789 24259
rect 2096 24228 2789 24256
rect 2096 24216 2102 24228
rect 2777 24225 2789 24228
rect 2823 24225 2835 24259
rect 2777 24219 2835 24225
rect 3694 24216 3700 24268
rect 3752 24256 3758 24268
rect 4525 24259 4583 24265
rect 4525 24256 4537 24259
rect 3752 24228 4537 24256
rect 3752 24216 3758 24228
rect 4525 24225 4537 24228
rect 4571 24225 4583 24259
rect 4525 24219 4583 24225
rect 6914 24216 6920 24268
rect 6972 24256 6978 24268
rect 7834 24256 7840 24268
rect 6972 24228 7840 24256
rect 6972 24216 6978 24228
rect 7834 24216 7840 24228
rect 7892 24216 7898 24268
rect 10594 24256 10600 24268
rect 10555 24228 10600 24256
rect 10594 24216 10600 24228
rect 10652 24216 10658 24268
rect 11974 24216 11980 24268
rect 12032 24256 12038 24268
rect 12069 24259 12127 24265
rect 12069 24256 12081 24259
rect 12032 24228 12081 24256
rect 12032 24216 12038 24228
rect 12069 24225 12081 24228
rect 12115 24225 12127 24259
rect 14090 24256 14096 24268
rect 14051 24228 14096 24256
rect 12069 24219 12127 24225
rect 14090 24216 14096 24228
rect 14148 24216 14154 24268
rect 15289 24259 15347 24265
rect 15289 24225 15301 24259
rect 15335 24256 15347 24259
rect 15470 24256 15476 24268
rect 15335 24228 15476 24256
rect 15335 24225 15347 24228
rect 15289 24219 15347 24225
rect 15470 24216 15476 24228
rect 15528 24216 15534 24268
rect 16485 24259 16543 24265
rect 16485 24225 16497 24259
rect 16531 24256 16543 24259
rect 16758 24256 16764 24268
rect 16531 24228 16764 24256
rect 16531 24225 16543 24228
rect 16485 24219 16543 24225
rect 16758 24216 16764 24228
rect 16816 24216 16822 24268
rect 17589 24259 17647 24265
rect 17589 24225 17601 24259
rect 17635 24256 17647 24259
rect 17678 24256 17684 24268
rect 17635 24228 17684 24256
rect 17635 24225 17647 24228
rect 17589 24219 17647 24225
rect 17678 24216 17684 24228
rect 17736 24216 17742 24268
rect 18785 24259 18843 24265
rect 18785 24225 18797 24259
rect 18831 24256 18843 24259
rect 19058 24256 19064 24268
rect 18831 24228 19064 24256
rect 18831 24225 18843 24228
rect 18785 24219 18843 24225
rect 19058 24216 19064 24228
rect 19116 24216 19122 24268
rect 20806 24216 20812 24268
rect 20864 24256 20870 24268
rect 20901 24259 20959 24265
rect 20901 24256 20913 24259
rect 20864 24228 20913 24256
rect 20864 24216 20870 24228
rect 20901 24225 20913 24228
rect 20947 24225 20959 24259
rect 20901 24219 20959 24225
rect 3053 24191 3111 24197
rect 3053 24157 3065 24191
rect 3099 24157 3111 24191
rect 3053 24151 3111 24157
rect 3068 24120 3096 24151
rect 4246 24148 4252 24200
rect 4304 24188 4310 24200
rect 4617 24191 4675 24197
rect 4617 24188 4629 24191
rect 4304 24160 4629 24188
rect 4304 24148 4310 24160
rect 4617 24157 4629 24160
rect 4663 24157 4675 24191
rect 4617 24151 4675 24157
rect 4801 24191 4859 24197
rect 4801 24157 4813 24191
rect 4847 24188 4859 24191
rect 4890 24188 4896 24200
rect 4847 24160 4896 24188
rect 4847 24157 4859 24160
rect 4801 24151 4859 24157
rect 3326 24120 3332 24132
rect 3068 24092 3332 24120
rect 3326 24080 3332 24092
rect 3384 24120 3390 24132
rect 3881 24123 3939 24129
rect 3881 24120 3893 24123
rect 3384 24092 3893 24120
rect 3384 24080 3390 24092
rect 3881 24089 3893 24092
rect 3927 24120 3939 24123
rect 4816 24120 4844 24151
rect 4890 24148 4896 24160
rect 4948 24148 4954 24200
rect 6549 24191 6607 24197
rect 6549 24157 6561 24191
rect 6595 24188 6607 24191
rect 7190 24188 7196 24200
rect 6595 24160 7196 24188
rect 6595 24157 6607 24160
rect 6549 24151 6607 24157
rect 7190 24148 7196 24160
rect 7248 24148 7254 24200
rect 7929 24191 7987 24197
rect 7929 24157 7941 24191
rect 7975 24157 7987 24191
rect 8110 24188 8116 24200
rect 8071 24160 8116 24188
rect 7929 24151 7987 24157
rect 3927 24092 4844 24120
rect 5905 24123 5963 24129
rect 3927 24089 3939 24092
rect 3881 24083 3939 24089
rect 5905 24089 5917 24123
rect 5951 24120 5963 24123
rect 7374 24120 7380 24132
rect 5951 24092 7380 24120
rect 5951 24089 5963 24092
rect 5905 24083 5963 24089
rect 7374 24080 7380 24092
rect 7432 24120 7438 24132
rect 7944 24120 7972 24151
rect 8110 24148 8116 24160
rect 8168 24148 8174 24200
rect 12250 24120 12256 24132
rect 7432 24092 7972 24120
rect 12211 24092 12256 24120
rect 7432 24080 7438 24092
rect 12250 24080 12256 24092
rect 12308 24080 12314 24132
rect 17770 24120 17776 24132
rect 17731 24092 17776 24120
rect 17770 24080 17776 24092
rect 17828 24080 17834 24132
rect 2317 24055 2375 24061
rect 2317 24021 2329 24055
rect 2363 24052 2375 24055
rect 2498 24052 2504 24064
rect 2363 24024 2504 24052
rect 2363 24021 2375 24024
rect 2317 24015 2375 24021
rect 2498 24012 2504 24024
rect 2556 24012 2562 24064
rect 4157 24055 4215 24061
rect 4157 24021 4169 24055
rect 4203 24052 4215 24055
rect 4982 24052 4988 24064
rect 4203 24024 4988 24052
rect 4203 24021 4215 24024
rect 4157 24015 4215 24021
rect 4982 24012 4988 24024
rect 5040 24012 5046 24064
rect 5261 24055 5319 24061
rect 5261 24021 5273 24055
rect 5307 24052 5319 24055
rect 5442 24052 5448 24064
rect 5307 24024 5448 24052
rect 5307 24021 5319 24024
rect 5261 24015 5319 24021
rect 5442 24012 5448 24024
rect 5500 24012 5506 24064
rect 7098 24052 7104 24064
rect 7059 24024 7104 24052
rect 7098 24012 7104 24024
rect 7156 24012 7162 24064
rect 7466 24052 7472 24064
rect 7427 24024 7472 24052
rect 7466 24012 7472 24024
rect 7524 24012 7530 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2038 23848 2044 23860
rect 1999 23820 2044 23848
rect 2038 23808 2044 23820
rect 2096 23808 2102 23860
rect 3050 23808 3056 23860
rect 3108 23848 3114 23860
rect 3145 23851 3203 23857
rect 3145 23848 3157 23851
rect 3108 23820 3157 23848
rect 3108 23808 3114 23820
rect 3145 23817 3157 23820
rect 3191 23817 3203 23851
rect 3694 23848 3700 23860
rect 3655 23820 3700 23848
rect 3145 23811 3203 23817
rect 1670 23740 1676 23792
rect 1728 23780 1734 23792
rect 2498 23780 2504 23792
rect 1728 23752 2504 23780
rect 1728 23740 1734 23752
rect 2498 23740 2504 23752
rect 2556 23780 2562 23792
rect 3160 23780 3188 23811
rect 3694 23808 3700 23820
rect 3752 23808 3758 23860
rect 4890 23808 4896 23860
rect 4948 23848 4954 23860
rect 5629 23851 5687 23857
rect 5629 23848 5641 23851
rect 4948 23820 5641 23848
rect 4948 23808 4954 23820
rect 5629 23817 5641 23820
rect 5675 23817 5687 23851
rect 6178 23848 6184 23860
rect 6139 23820 6184 23848
rect 5629 23811 5687 23817
rect 6178 23808 6184 23820
rect 6236 23808 6242 23860
rect 13081 23851 13139 23857
rect 13081 23817 13093 23851
rect 13127 23848 13139 23851
rect 13354 23848 13360 23860
rect 13127 23820 13360 23848
rect 13127 23817 13139 23820
rect 13081 23811 13139 23817
rect 3786 23780 3792 23792
rect 2556 23752 2728 23780
rect 3160 23752 3792 23780
rect 2556 23740 2562 23752
rect 2590 23712 2596 23724
rect 2551 23684 2596 23712
rect 2590 23672 2596 23684
rect 2648 23672 2654 23724
rect 2700 23721 2728 23752
rect 3786 23740 3792 23752
rect 3844 23740 3850 23792
rect 4157 23783 4215 23789
rect 4157 23749 4169 23783
rect 4203 23780 4215 23783
rect 4246 23780 4252 23792
rect 4203 23752 4252 23780
rect 4203 23749 4215 23752
rect 4157 23743 4215 23749
rect 4246 23740 4252 23752
rect 4304 23740 4310 23792
rect 5994 23740 6000 23792
rect 6052 23780 6058 23792
rect 6549 23783 6607 23789
rect 6549 23780 6561 23783
rect 6052 23752 6561 23780
rect 6052 23740 6058 23752
rect 6549 23749 6561 23752
rect 6595 23780 6607 23783
rect 6730 23780 6736 23792
rect 6595 23752 6736 23780
rect 6595 23749 6607 23752
rect 6549 23743 6607 23749
rect 6730 23740 6736 23752
rect 6788 23740 6794 23792
rect 2685 23715 2743 23721
rect 2685 23681 2697 23715
rect 2731 23681 2743 23715
rect 2685 23675 2743 23681
rect 2222 23604 2228 23656
rect 2280 23644 2286 23656
rect 2501 23647 2559 23653
rect 2501 23644 2513 23647
rect 2280 23616 2513 23644
rect 2280 23604 2286 23616
rect 2501 23613 2513 23616
rect 2547 23613 2559 23647
rect 4246 23644 4252 23656
rect 4207 23616 4252 23644
rect 2501 23607 2559 23613
rect 4246 23604 4252 23616
rect 4304 23604 4310 23656
rect 6270 23604 6276 23656
rect 6328 23644 6334 23656
rect 7098 23644 7104 23656
rect 6328 23616 7104 23644
rect 6328 23604 6334 23616
rect 7098 23604 7104 23616
rect 7156 23604 7162 23656
rect 9858 23604 9864 23656
rect 9916 23644 9922 23656
rect 10594 23644 10600 23656
rect 9916 23616 10600 23644
rect 9916 23604 9922 23616
rect 10594 23604 10600 23616
rect 10652 23604 10658 23656
rect 11241 23647 11299 23653
rect 11241 23613 11253 23647
rect 11287 23644 11299 23647
rect 11330 23644 11336 23656
rect 11287 23616 11336 23644
rect 11287 23613 11299 23616
rect 11241 23607 11299 23613
rect 11330 23604 11336 23616
rect 11388 23644 11394 23656
rect 11793 23647 11851 23653
rect 11793 23644 11805 23647
rect 11388 23616 11805 23644
rect 11388 23604 11394 23616
rect 11793 23613 11805 23616
rect 11839 23613 11851 23647
rect 11793 23607 11851 23613
rect 12437 23647 12495 23653
rect 12437 23613 12449 23647
rect 12483 23644 12495 23647
rect 13096 23644 13124 23811
rect 13354 23808 13360 23820
rect 13412 23808 13418 23860
rect 13725 23851 13783 23857
rect 13725 23817 13737 23851
rect 13771 23848 13783 23851
rect 14090 23848 14096 23860
rect 13771 23820 14096 23848
rect 13771 23817 13783 23820
rect 13725 23811 13783 23817
rect 14090 23808 14096 23820
rect 14148 23808 14154 23860
rect 14461 23851 14519 23857
rect 14461 23817 14473 23851
rect 14507 23848 14519 23851
rect 15654 23848 15660 23860
rect 14507 23820 15660 23848
rect 14507 23817 14519 23820
rect 14461 23811 14519 23817
rect 12483 23616 13124 23644
rect 13817 23647 13875 23653
rect 12483 23613 12495 23616
rect 12437 23607 12495 23613
rect 13817 23613 13829 23647
rect 13863 23644 13875 23647
rect 14476 23644 14504 23811
rect 15654 23808 15660 23820
rect 15712 23808 15718 23860
rect 18322 23848 18328 23860
rect 18283 23820 18328 23848
rect 18322 23808 18328 23820
rect 18380 23808 18386 23860
rect 19518 23848 19524 23860
rect 19479 23820 19524 23848
rect 19518 23808 19524 23820
rect 19576 23808 19582 23860
rect 21266 23848 21272 23860
rect 21227 23820 21272 23848
rect 21266 23808 21272 23820
rect 21324 23808 21330 23860
rect 23845 23851 23903 23857
rect 23845 23817 23857 23851
rect 23891 23848 23903 23851
rect 25314 23848 25320 23860
rect 23891 23820 25320 23848
rect 23891 23817 23903 23820
rect 23845 23811 23903 23817
rect 25314 23808 25320 23820
rect 25372 23808 25378 23860
rect 15194 23780 15200 23792
rect 15155 23752 15200 23780
rect 15194 23740 15200 23752
rect 15252 23740 15258 23792
rect 16945 23783 17003 23789
rect 16945 23749 16957 23783
rect 16991 23780 17003 23783
rect 19702 23780 19708 23792
rect 16991 23752 19708 23780
rect 16991 23749 17003 23752
rect 16945 23743 17003 23749
rect 19702 23740 19708 23752
rect 19760 23740 19766 23792
rect 15013 23647 15071 23653
rect 15013 23644 15025 23647
rect 13863 23616 14504 23644
rect 14844 23616 15025 23644
rect 13863 23613 13875 23616
rect 13817 23607 13875 23613
rect 1673 23579 1731 23585
rect 1673 23545 1685 23579
rect 1719 23576 1731 23579
rect 3326 23576 3332 23588
rect 1719 23548 3332 23576
rect 1719 23545 1731 23548
rect 1673 23539 1731 23545
rect 3326 23536 3332 23548
rect 3384 23536 3390 23588
rect 4516 23579 4574 23585
rect 4516 23545 4528 23579
rect 4562 23576 4574 23579
rect 4798 23576 4804 23588
rect 4562 23548 4804 23576
rect 4562 23545 4574 23548
rect 4516 23539 4574 23545
rect 4798 23536 4804 23548
rect 4856 23536 4862 23588
rect 7190 23536 7196 23588
rect 7248 23576 7254 23588
rect 7368 23579 7426 23585
rect 7368 23576 7380 23579
rect 7248 23548 7380 23576
rect 7248 23536 7254 23548
rect 7368 23545 7380 23548
rect 7414 23576 7426 23579
rect 7742 23576 7748 23588
rect 7414 23548 7748 23576
rect 7414 23545 7426 23548
rect 7368 23539 7426 23545
rect 7742 23536 7748 23548
rect 7800 23536 7806 23588
rect 1394 23468 1400 23520
rect 1452 23508 1458 23520
rect 1578 23508 1584 23520
rect 1452 23480 1584 23508
rect 1452 23468 1458 23480
rect 1578 23468 1584 23480
rect 1636 23468 1642 23520
rect 2130 23508 2136 23520
rect 2091 23480 2136 23508
rect 2130 23468 2136 23480
rect 2188 23468 2194 23520
rect 6638 23468 6644 23520
rect 6696 23508 6702 23520
rect 8110 23508 8116 23520
rect 6696 23480 8116 23508
rect 6696 23468 6702 23480
rect 8110 23468 8116 23480
rect 8168 23508 8174 23520
rect 8481 23511 8539 23517
rect 8481 23508 8493 23511
rect 8168 23480 8493 23508
rect 8168 23468 8174 23480
rect 8481 23477 8493 23480
rect 8527 23508 8539 23511
rect 9033 23511 9091 23517
rect 9033 23508 9045 23511
rect 8527 23480 9045 23508
rect 8527 23477 8539 23480
rect 8481 23471 8539 23477
rect 9033 23477 9045 23480
rect 9079 23477 9091 23511
rect 11422 23508 11428 23520
rect 11383 23480 11428 23508
rect 9033 23471 9091 23477
rect 11422 23468 11428 23480
rect 11480 23468 11486 23520
rect 11974 23468 11980 23520
rect 12032 23508 12038 23520
rect 12161 23511 12219 23517
rect 12161 23508 12173 23511
rect 12032 23480 12173 23508
rect 12032 23468 12038 23480
rect 12161 23477 12173 23480
rect 12207 23477 12219 23511
rect 12618 23508 12624 23520
rect 12579 23480 12624 23508
rect 12161 23471 12219 23477
rect 12618 23468 12624 23480
rect 12676 23468 12682 23520
rect 13814 23468 13820 23520
rect 13872 23508 13878 23520
rect 14001 23511 14059 23517
rect 14001 23508 14013 23511
rect 13872 23480 14013 23508
rect 13872 23468 13878 23480
rect 14001 23477 14013 23480
rect 14047 23477 14059 23511
rect 14001 23471 14059 23477
rect 14642 23468 14648 23520
rect 14700 23508 14706 23520
rect 14844 23517 14872 23616
rect 15013 23613 15025 23616
rect 15059 23613 15071 23647
rect 15013 23607 15071 23613
rect 16574 23604 16580 23656
rect 16632 23644 16638 23656
rect 16761 23647 16819 23653
rect 16761 23644 16773 23647
rect 16632 23616 16773 23644
rect 16632 23604 16638 23616
rect 16761 23613 16773 23616
rect 16807 23644 16819 23647
rect 17313 23647 17371 23653
rect 17313 23644 17325 23647
rect 16807 23616 17325 23644
rect 16807 23613 16819 23616
rect 16761 23607 16819 23613
rect 17313 23613 17325 23616
rect 17359 23613 17371 23647
rect 17313 23607 17371 23613
rect 18141 23647 18199 23653
rect 18141 23613 18153 23647
rect 18187 23644 18199 23647
rect 19334 23644 19340 23656
rect 18187 23616 18736 23644
rect 19295 23616 19340 23644
rect 18187 23613 18199 23616
rect 18141 23607 18199 23613
rect 18708 23520 18736 23616
rect 19334 23604 19340 23616
rect 19392 23644 19398 23656
rect 19889 23647 19947 23653
rect 19889 23644 19901 23647
rect 19392 23616 19901 23644
rect 19392 23604 19398 23616
rect 19889 23613 19901 23616
rect 19935 23613 19947 23647
rect 21082 23644 21088 23656
rect 20995 23616 21088 23644
rect 19889 23607 19947 23613
rect 21082 23604 21088 23616
rect 21140 23644 21146 23656
rect 21637 23647 21695 23653
rect 21637 23644 21649 23647
rect 21140 23616 21649 23644
rect 21140 23604 21146 23616
rect 21637 23613 21649 23616
rect 21683 23613 21695 23647
rect 21637 23607 21695 23613
rect 23474 23604 23480 23656
rect 23532 23644 23538 23656
rect 23661 23647 23719 23653
rect 23661 23644 23673 23647
rect 23532 23616 23673 23644
rect 23532 23604 23538 23616
rect 23661 23613 23673 23616
rect 23707 23644 23719 23647
rect 24213 23647 24271 23653
rect 24213 23644 24225 23647
rect 23707 23616 24225 23644
rect 23707 23613 23719 23616
rect 23661 23607 23719 23613
rect 24213 23613 24225 23616
rect 24259 23613 24271 23647
rect 24213 23607 24271 23613
rect 14829 23511 14887 23517
rect 14829 23508 14841 23511
rect 14700 23480 14841 23508
rect 14700 23468 14706 23480
rect 14829 23477 14841 23480
rect 14875 23477 14887 23511
rect 14829 23471 14887 23477
rect 15470 23468 15476 23520
rect 15528 23508 15534 23520
rect 15565 23511 15623 23517
rect 15565 23508 15577 23511
rect 15528 23480 15577 23508
rect 15528 23468 15534 23480
rect 15565 23477 15577 23480
rect 15611 23477 15623 23511
rect 15565 23471 15623 23477
rect 16577 23511 16635 23517
rect 16577 23477 16589 23511
rect 16623 23508 16635 23511
rect 16758 23508 16764 23520
rect 16623 23480 16764 23508
rect 16623 23477 16635 23480
rect 16577 23471 16635 23477
rect 16758 23468 16764 23480
rect 16816 23468 16822 23520
rect 17678 23508 17684 23520
rect 17639 23480 17684 23508
rect 17678 23468 17684 23480
rect 17736 23468 17742 23520
rect 18690 23508 18696 23520
rect 18651 23480 18696 23508
rect 18690 23468 18696 23480
rect 18748 23468 18754 23520
rect 19058 23508 19064 23520
rect 19019 23480 19064 23508
rect 19058 23468 19064 23480
rect 19116 23468 19122 23520
rect 20806 23468 20812 23520
rect 20864 23508 20870 23520
rect 20901 23511 20959 23517
rect 20901 23508 20913 23511
rect 20864 23480 20913 23508
rect 20864 23468 20870 23480
rect 20901 23477 20913 23480
rect 20947 23477 20959 23511
rect 20901 23471 20959 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 2774 23264 2780 23316
rect 2832 23304 2838 23316
rect 3145 23307 3203 23313
rect 3145 23304 3157 23307
rect 2832 23276 3157 23304
rect 2832 23264 2838 23276
rect 3145 23273 3157 23276
rect 3191 23273 3203 23307
rect 3145 23267 3203 23273
rect 5997 23307 6055 23313
rect 5997 23273 6009 23307
rect 6043 23304 6055 23307
rect 7190 23304 7196 23316
rect 6043 23276 7196 23304
rect 6043 23273 6055 23276
rect 5997 23267 6055 23273
rect 7190 23264 7196 23276
rect 7248 23264 7254 23316
rect 9858 23304 9864 23316
rect 9819 23276 9864 23304
rect 9858 23264 9864 23276
rect 9916 23264 9922 23316
rect 14001 23307 14059 23313
rect 14001 23273 14013 23307
rect 14047 23304 14059 23307
rect 14090 23304 14096 23316
rect 14047 23276 14096 23304
rect 14047 23273 14059 23276
rect 14001 23267 14059 23273
rect 14090 23264 14096 23276
rect 14148 23264 14154 23316
rect 17218 23304 17224 23316
rect 17179 23276 17224 23304
rect 17218 23264 17224 23276
rect 17276 23264 17282 23316
rect 18325 23307 18383 23313
rect 18325 23273 18337 23307
rect 18371 23304 18383 23307
rect 19058 23304 19064 23316
rect 18371 23276 19064 23304
rect 18371 23273 18383 23276
rect 18325 23267 18383 23273
rect 19058 23264 19064 23276
rect 19116 23264 19122 23316
rect 21082 23304 21088 23316
rect 21043 23276 21088 23304
rect 21082 23264 21088 23276
rect 21140 23264 21146 23316
rect 22557 23307 22615 23313
rect 22557 23273 22569 23307
rect 22603 23304 22615 23307
rect 23474 23304 23480 23316
rect 22603 23276 23480 23304
rect 22603 23273 22615 23276
rect 22557 23267 22615 23273
rect 23474 23264 23480 23276
rect 23532 23264 23538 23316
rect 2869 23239 2927 23245
rect 2869 23205 2881 23239
rect 2915 23236 2927 23239
rect 3326 23236 3332 23248
rect 2915 23208 3332 23236
rect 2915 23205 2927 23208
rect 2869 23199 2927 23205
rect 3326 23196 3332 23208
rect 3384 23196 3390 23248
rect 5077 23239 5135 23245
rect 5077 23205 5089 23239
rect 5123 23236 5135 23239
rect 5166 23236 5172 23248
rect 5123 23208 5172 23236
rect 5123 23205 5135 23208
rect 5077 23199 5135 23205
rect 5166 23196 5172 23208
rect 5224 23196 5230 23248
rect 6540 23239 6598 23245
rect 6540 23205 6552 23239
rect 6586 23236 6598 23239
rect 6638 23236 6644 23248
rect 6586 23208 6644 23236
rect 6586 23205 6598 23208
rect 6540 23199 6598 23205
rect 6638 23196 6644 23208
rect 6696 23196 6702 23248
rect 2130 23168 2136 23180
rect 2091 23140 2136 23168
rect 2130 23128 2136 23140
rect 2188 23128 2194 23180
rect 4246 23128 4252 23180
rect 4304 23168 4310 23180
rect 4341 23171 4399 23177
rect 4341 23168 4353 23171
rect 4304 23140 4353 23168
rect 4304 23128 4310 23140
rect 4341 23137 4353 23140
rect 4387 23168 4399 23171
rect 9674 23168 9680 23180
rect 4387 23140 6316 23168
rect 9635 23140 9680 23168
rect 4387 23137 4399 23140
rect 4341 23131 4399 23137
rect 6288 23112 6316 23140
rect 9674 23128 9680 23140
rect 9732 23128 9738 23180
rect 12713 23171 12771 23177
rect 12713 23137 12725 23171
rect 12759 23168 12771 23171
rect 13078 23168 13084 23180
rect 12759 23140 13084 23168
rect 12759 23137 12771 23140
rect 12713 23131 12771 23137
rect 13078 23128 13084 23140
rect 13136 23128 13142 23180
rect 13817 23171 13875 23177
rect 13817 23137 13829 23171
rect 13863 23168 13875 23171
rect 14274 23168 14280 23180
rect 13863 23140 14280 23168
rect 13863 23137 13875 23140
rect 13817 23131 13875 23137
rect 14274 23128 14280 23140
rect 14332 23128 14338 23180
rect 15286 23168 15292 23180
rect 15247 23140 15292 23168
rect 15286 23128 15292 23140
rect 15344 23128 15350 23180
rect 17034 23168 17040 23180
rect 16995 23140 17040 23168
rect 17034 23128 17040 23140
rect 17092 23128 17098 23180
rect 18138 23168 18144 23180
rect 18099 23140 18144 23168
rect 18138 23128 18144 23140
rect 18196 23128 18202 23180
rect 20898 23168 20904 23180
rect 20859 23140 20904 23168
rect 20898 23128 20904 23140
rect 20956 23128 20962 23180
rect 22370 23168 22376 23180
rect 22331 23140 22376 23168
rect 22370 23128 22376 23140
rect 22428 23128 22434 23180
rect 2222 23100 2228 23112
rect 2183 23072 2228 23100
rect 2222 23060 2228 23072
rect 2280 23060 2286 23112
rect 2409 23103 2467 23109
rect 2409 23069 2421 23103
rect 2455 23100 2467 23103
rect 2682 23100 2688 23112
rect 2455 23072 2688 23100
rect 2455 23069 2467 23072
rect 2409 23063 2467 23069
rect 1673 23035 1731 23041
rect 1673 23001 1685 23035
rect 1719 23032 1731 23035
rect 2424 23032 2452 23063
rect 2682 23060 2688 23072
rect 2740 23060 2746 23112
rect 3970 23060 3976 23112
rect 4028 23100 4034 23112
rect 5169 23103 5227 23109
rect 5169 23100 5181 23103
rect 4028 23072 5181 23100
rect 4028 23060 4034 23072
rect 5169 23069 5181 23072
rect 5215 23100 5227 23103
rect 5258 23100 5264 23112
rect 5215 23072 5264 23100
rect 5215 23069 5227 23072
rect 5169 23063 5227 23069
rect 5258 23060 5264 23072
rect 5316 23060 5322 23112
rect 5353 23103 5411 23109
rect 5353 23069 5365 23103
rect 5399 23069 5411 23103
rect 6270 23100 6276 23112
rect 6231 23072 6276 23100
rect 5353 23063 5411 23069
rect 1719 23004 2452 23032
rect 3881 23035 3939 23041
rect 1719 23001 1731 23004
rect 1673 22995 1731 23001
rect 3881 23001 3893 23035
rect 3927 23032 3939 23035
rect 4798 23032 4804 23044
rect 3927 23004 4804 23032
rect 3927 23001 3939 23004
rect 3881 22995 3939 23001
rect 4798 22992 4804 23004
rect 4856 23032 4862 23044
rect 5368 23032 5396 23063
rect 6270 23060 6276 23072
rect 6328 23060 6334 23112
rect 12894 23032 12900 23044
rect 4856 23004 6224 23032
rect 12855 23004 12900 23032
rect 4856 22992 4862 23004
rect 1762 22964 1768 22976
rect 1723 22936 1768 22964
rect 1762 22924 1768 22936
rect 1820 22924 1826 22976
rect 4430 22924 4436 22976
rect 4488 22964 4494 22976
rect 4709 22967 4767 22973
rect 4709 22964 4721 22967
rect 4488 22936 4721 22964
rect 4488 22924 4494 22936
rect 4709 22933 4721 22936
rect 4755 22933 4767 22967
rect 6196 22964 6224 23004
rect 12894 22992 12900 23004
rect 12952 22992 12958 23044
rect 7653 22967 7711 22973
rect 7653 22964 7665 22967
rect 6196 22936 7665 22964
rect 4709 22927 4767 22933
rect 7653 22933 7665 22936
rect 7699 22933 7711 22967
rect 8478 22964 8484 22976
rect 8439 22936 8484 22964
rect 7653 22927 7711 22933
rect 8478 22924 8484 22936
rect 8536 22924 8542 22976
rect 13630 22964 13636 22976
rect 13591 22936 13636 22964
rect 13630 22924 13636 22936
rect 13688 22924 13694 22976
rect 14274 22964 14280 22976
rect 14235 22936 14280 22964
rect 14274 22924 14280 22936
rect 14332 22924 14338 22976
rect 15473 22967 15531 22973
rect 15473 22933 15485 22967
rect 15519 22964 15531 22967
rect 15562 22964 15568 22976
rect 15519 22936 15568 22964
rect 15519 22933 15531 22936
rect 15473 22927 15531 22933
rect 15562 22924 15568 22936
rect 15620 22924 15626 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 2038 22760 2044 22772
rect 1999 22732 2044 22760
rect 2038 22720 2044 22732
rect 2096 22720 2102 22772
rect 2593 22763 2651 22769
rect 2593 22729 2605 22763
rect 2639 22760 2651 22763
rect 4246 22760 4252 22772
rect 2639 22732 4252 22760
rect 2639 22729 2651 22732
rect 2593 22723 2651 22729
rect 2590 22584 2596 22636
rect 2648 22624 2654 22636
rect 2700 22633 2728 22732
rect 4246 22720 4252 22732
rect 4304 22720 4310 22772
rect 4798 22760 4804 22772
rect 4759 22732 4804 22760
rect 4798 22720 4804 22732
rect 4856 22720 4862 22772
rect 6086 22720 6092 22772
rect 6144 22760 6150 22772
rect 6181 22763 6239 22769
rect 6181 22760 6193 22763
rect 6144 22732 6193 22760
rect 6144 22720 6150 22732
rect 6181 22729 6193 22732
rect 6227 22729 6239 22763
rect 6181 22723 6239 22729
rect 6362 22720 6368 22772
rect 6420 22760 6426 22772
rect 6549 22763 6607 22769
rect 6549 22760 6561 22763
rect 6420 22732 6561 22760
rect 6420 22720 6426 22732
rect 6549 22729 6561 22732
rect 6595 22760 6607 22763
rect 15654 22760 15660 22772
rect 6595 22732 7328 22760
rect 15615 22732 15660 22760
rect 6595 22729 6607 22732
rect 6549 22723 6607 22729
rect 6825 22695 6883 22701
rect 6825 22692 6837 22695
rect 5644 22664 6837 22692
rect 5644 22636 5672 22664
rect 6825 22661 6837 22664
rect 6871 22661 6883 22695
rect 6825 22655 6883 22661
rect 2685 22627 2743 22633
rect 2685 22624 2697 22627
rect 2648 22596 2697 22624
rect 2648 22584 2654 22596
rect 2685 22593 2697 22596
rect 2731 22593 2743 22627
rect 5626 22624 5632 22636
rect 5539 22596 5632 22624
rect 2685 22587 2743 22593
rect 5626 22584 5632 22596
rect 5684 22584 5690 22636
rect 5813 22627 5871 22633
rect 5813 22593 5825 22627
rect 5859 22624 5871 22627
rect 5994 22624 6000 22636
rect 5859 22596 6000 22624
rect 5859 22593 5871 22596
rect 5813 22587 5871 22593
rect 5994 22584 6000 22596
rect 6052 22624 6058 22636
rect 6638 22624 6644 22636
rect 6052 22596 6644 22624
rect 6052 22584 6058 22596
rect 6638 22584 6644 22596
rect 6696 22584 6702 22636
rect 7300 22633 7328 22732
rect 15654 22720 15660 22732
rect 15712 22720 15718 22772
rect 16758 22760 16764 22772
rect 16719 22732 16764 22760
rect 16758 22720 16764 22732
rect 16816 22720 16822 22772
rect 20898 22760 20904 22772
rect 20859 22732 20904 22760
rect 20898 22720 20904 22732
rect 20956 22720 20962 22772
rect 8386 22692 8392 22704
rect 8347 22664 8392 22692
rect 8386 22652 8392 22664
rect 8444 22652 8450 22704
rect 7285 22627 7343 22633
rect 7285 22593 7297 22627
rect 7331 22593 7343 22627
rect 7285 22587 7343 22593
rect 7469 22627 7527 22633
rect 7469 22593 7481 22627
rect 7515 22624 7527 22627
rect 7742 22624 7748 22636
rect 7515 22596 7748 22624
rect 7515 22593 7527 22596
rect 7469 22587 7527 22593
rect 7742 22584 7748 22596
rect 7800 22624 7806 22636
rect 7929 22627 7987 22633
rect 7929 22624 7941 22627
rect 7800 22596 7941 22624
rect 7800 22584 7806 22596
rect 7929 22593 7941 22596
rect 7975 22624 7987 22627
rect 8941 22627 8999 22633
rect 8941 22624 8953 22627
rect 7975 22596 8953 22624
rect 7975 22593 7987 22596
rect 7929 22587 7987 22593
rect 8941 22593 8953 22596
rect 8987 22593 8999 22627
rect 8941 22587 8999 22593
rect 14185 22627 14243 22633
rect 14185 22593 14197 22627
rect 14231 22624 14243 22627
rect 14231 22596 14688 22624
rect 14231 22593 14243 22596
rect 14185 22587 14243 22593
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22556 1455 22559
rect 2038 22556 2044 22568
rect 1443 22528 2044 22556
rect 1443 22525 1455 22528
rect 1397 22519 1455 22525
rect 2038 22516 2044 22528
rect 2096 22516 2102 22568
rect 2952 22559 3010 22565
rect 2952 22525 2964 22559
rect 2998 22556 3010 22559
rect 3326 22556 3332 22568
rect 2998 22528 3332 22556
rect 2998 22525 3010 22528
rect 2952 22519 3010 22525
rect 3326 22516 3332 22528
rect 3384 22516 3390 22568
rect 5534 22556 5540 22568
rect 5495 22528 5540 22556
rect 5534 22516 5540 22528
rect 5592 22516 5598 22568
rect 6086 22516 6092 22568
rect 6144 22556 6150 22568
rect 7193 22559 7251 22565
rect 7193 22556 7205 22559
rect 6144 22528 7205 22556
rect 6144 22516 6150 22528
rect 7193 22525 7205 22528
rect 7239 22525 7251 22559
rect 7193 22519 7251 22525
rect 8478 22516 8484 22568
rect 8536 22556 8542 22568
rect 8757 22559 8815 22565
rect 8757 22556 8769 22559
rect 8536 22528 8769 22556
rect 8536 22516 8542 22528
rect 8757 22525 8769 22528
rect 8803 22525 8815 22559
rect 8757 22519 8815 22525
rect 13354 22488 13360 22500
rect 13315 22460 13360 22488
rect 13354 22448 13360 22460
rect 13412 22488 13418 22500
rect 14001 22491 14059 22497
rect 14001 22488 14013 22491
rect 13412 22460 14013 22488
rect 13412 22448 13418 22460
rect 14001 22457 14013 22460
rect 14047 22457 14059 22491
rect 14001 22451 14059 22457
rect 1578 22420 1584 22432
rect 1539 22392 1584 22420
rect 1578 22380 1584 22392
rect 1636 22380 1642 22432
rect 4062 22420 4068 22432
rect 4023 22392 4068 22420
rect 4062 22380 4068 22392
rect 4120 22380 4126 22432
rect 5166 22420 5172 22432
rect 5127 22392 5172 22420
rect 5166 22380 5172 22392
rect 5224 22380 5230 22432
rect 8202 22420 8208 22432
rect 8163 22392 8208 22420
rect 8202 22380 8208 22392
rect 8260 22420 8266 22432
rect 8849 22423 8907 22429
rect 8849 22420 8861 22423
rect 8260 22392 8861 22420
rect 8260 22380 8266 22392
rect 8849 22389 8861 22392
rect 8895 22389 8907 22423
rect 8849 22383 8907 22389
rect 9306 22380 9312 22432
rect 9364 22420 9370 22432
rect 9674 22420 9680 22432
rect 9364 22392 9680 22420
rect 9364 22380 9370 22392
rect 9674 22380 9680 22392
rect 9732 22380 9738 22432
rect 10873 22423 10931 22429
rect 10873 22389 10885 22423
rect 10919 22420 10931 22423
rect 10962 22420 10968 22432
rect 10919 22392 10968 22420
rect 10919 22389 10931 22392
rect 10873 22383 10931 22389
rect 10962 22380 10968 22392
rect 11020 22380 11026 22432
rect 12805 22423 12863 22429
rect 12805 22389 12817 22423
rect 12851 22420 12863 22423
rect 13078 22420 13084 22432
rect 12851 22392 13084 22420
rect 12851 22389 12863 22392
rect 12805 22383 12863 22389
rect 13078 22380 13084 22392
rect 13136 22380 13142 22432
rect 13538 22420 13544 22432
rect 13499 22392 13544 22420
rect 13538 22380 13544 22392
rect 13596 22380 13602 22432
rect 13630 22380 13636 22432
rect 13688 22420 13694 22432
rect 14660 22429 14688 22596
rect 15194 22516 15200 22568
rect 15252 22556 15258 22568
rect 15473 22559 15531 22565
rect 15473 22556 15485 22559
rect 15252 22528 15485 22556
rect 15252 22516 15258 22528
rect 15473 22525 15485 22528
rect 15519 22556 15531 22559
rect 16025 22559 16083 22565
rect 16025 22556 16037 22559
rect 15519 22528 16037 22556
rect 15519 22525 15531 22528
rect 15473 22519 15531 22525
rect 16025 22525 16037 22528
rect 16071 22525 16083 22559
rect 16025 22519 16083 22525
rect 16577 22559 16635 22565
rect 16577 22525 16589 22559
rect 16623 22556 16635 22559
rect 16623 22528 17540 22556
rect 16623 22525 16635 22528
rect 16577 22519 16635 22525
rect 15286 22448 15292 22500
rect 15344 22488 15350 22500
rect 15381 22491 15439 22497
rect 15381 22488 15393 22491
rect 15344 22460 15393 22488
rect 15344 22448 15350 22460
rect 15381 22457 15393 22460
rect 15427 22488 15439 22491
rect 15746 22488 15752 22500
rect 15427 22460 15752 22488
rect 15427 22457 15439 22460
rect 15381 22451 15439 22457
rect 15746 22448 15752 22460
rect 15804 22448 15810 22500
rect 17512 22432 17540 22528
rect 13909 22423 13967 22429
rect 13909 22420 13921 22423
rect 13688 22392 13921 22420
rect 13688 22380 13694 22392
rect 13909 22389 13921 22392
rect 13955 22389 13967 22423
rect 13909 22383 13967 22389
rect 14645 22423 14703 22429
rect 14645 22389 14657 22423
rect 14691 22420 14703 22423
rect 15102 22420 15108 22432
rect 14691 22392 15108 22420
rect 14691 22389 14703 22392
rect 14645 22383 14703 22389
rect 15102 22380 15108 22392
rect 15160 22380 15166 22432
rect 17034 22420 17040 22432
rect 16995 22392 17040 22420
rect 17034 22380 17040 22392
rect 17092 22380 17098 22432
rect 17494 22420 17500 22432
rect 17455 22392 17500 22420
rect 17494 22380 17500 22392
rect 17552 22380 17558 22432
rect 18138 22380 18144 22432
rect 18196 22420 18202 22432
rect 18233 22423 18291 22429
rect 18233 22420 18245 22423
rect 18196 22392 18245 22420
rect 18196 22380 18202 22392
rect 18233 22389 18245 22392
rect 18279 22389 18291 22423
rect 22370 22420 22376 22432
rect 22331 22392 22376 22420
rect 18233 22383 18291 22389
rect 22370 22380 22376 22392
rect 22428 22380 22434 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 5166 22216 5172 22228
rect 4356 22188 5172 22216
rect 4356 22148 4384 22188
rect 5166 22176 5172 22188
rect 5224 22176 5230 22228
rect 5626 22216 5632 22228
rect 5587 22188 5632 22216
rect 5626 22176 5632 22188
rect 5684 22176 5690 22228
rect 5994 22216 6000 22228
rect 5955 22188 6000 22216
rect 5994 22176 6000 22188
rect 6052 22176 6058 22228
rect 8021 22219 8079 22225
rect 8021 22185 8033 22219
rect 8067 22216 8079 22219
rect 8478 22216 8484 22228
rect 8067 22188 8484 22216
rect 8067 22185 8079 22188
rect 8021 22179 8079 22185
rect 8478 22176 8484 22188
rect 8536 22176 8542 22228
rect 10870 22216 10876 22228
rect 10783 22188 10876 22216
rect 10870 22176 10876 22188
rect 10928 22216 10934 22228
rect 13078 22216 13084 22228
rect 10928 22188 13084 22216
rect 10928 22176 10934 22188
rect 13078 22176 13084 22188
rect 13136 22176 13142 22228
rect 13265 22219 13323 22225
rect 13265 22185 13277 22219
rect 13311 22216 13323 22219
rect 13538 22216 13544 22228
rect 13311 22188 13544 22216
rect 13311 22185 13323 22188
rect 13265 22179 13323 22185
rect 13538 22176 13544 22188
rect 13596 22216 13602 22228
rect 13725 22219 13783 22225
rect 13725 22216 13737 22219
rect 13596 22188 13737 22216
rect 13596 22176 13602 22188
rect 13725 22185 13737 22188
rect 13771 22185 13783 22219
rect 13725 22179 13783 22185
rect 4080 22120 4384 22148
rect 4433 22151 4491 22157
rect 1670 22089 1676 22092
rect 1664 22080 1676 22089
rect 1631 22052 1676 22080
rect 1664 22043 1676 22052
rect 1670 22040 1676 22043
rect 1728 22040 1734 22092
rect 2222 22040 2228 22092
rect 2280 22080 2286 22092
rect 2498 22080 2504 22092
rect 2280 22052 2504 22080
rect 2280 22040 2286 22052
rect 2498 22040 2504 22052
rect 2556 22080 2562 22092
rect 3881 22083 3939 22089
rect 2556 22052 2912 22080
rect 2556 22040 2562 22052
rect 1302 21972 1308 22024
rect 1360 22012 1366 22024
rect 1397 22015 1455 22021
rect 1397 22012 1409 22015
rect 1360 21984 1409 22012
rect 1360 21972 1366 21984
rect 1397 21981 1409 21984
rect 1443 21981 1455 22015
rect 1397 21975 1455 21981
rect 2406 21972 2412 22024
rect 2464 22012 2470 22024
rect 2682 22012 2688 22024
rect 2464 21984 2688 22012
rect 2464 21972 2470 21984
rect 2682 21972 2688 21984
rect 2740 22012 2746 22024
rect 2740 21984 2820 22012
rect 2740 21972 2746 21984
rect 2792 21953 2820 21984
rect 2777 21947 2835 21953
rect 2777 21913 2789 21947
rect 2823 21913 2835 21947
rect 2884 21944 2912 22052
rect 3881 22049 3893 22083
rect 3927 22080 3939 22083
rect 3970 22080 3976 22092
rect 3927 22052 3976 22080
rect 3927 22049 3939 22052
rect 3881 22043 3939 22049
rect 3970 22040 3976 22052
rect 4028 22040 4034 22092
rect 3513 22015 3571 22021
rect 3513 21981 3525 22015
rect 3559 22012 3571 22015
rect 4080 22012 4108 22120
rect 4433 22117 4445 22151
rect 4479 22148 4491 22151
rect 4982 22148 4988 22160
rect 4479 22120 4988 22148
rect 4479 22117 4491 22120
rect 4433 22111 4491 22117
rect 4982 22108 4988 22120
rect 5040 22148 5046 22160
rect 5534 22148 5540 22160
rect 5040 22120 5540 22148
rect 5040 22108 5046 22120
rect 5534 22108 5540 22120
rect 5592 22108 5598 22160
rect 5261 22083 5319 22089
rect 5261 22049 5273 22083
rect 5307 22080 5319 22083
rect 6012 22080 6040 22176
rect 12345 22151 12403 22157
rect 12345 22117 12357 22151
rect 12391 22148 12403 22151
rect 13630 22148 13636 22160
rect 12391 22120 13636 22148
rect 12391 22117 12403 22120
rect 12345 22111 12403 22117
rect 13630 22108 13636 22120
rect 13688 22108 13694 22160
rect 5307 22052 6040 22080
rect 5307 22049 5319 22052
rect 5261 22043 5319 22049
rect 6638 22040 6644 22092
rect 6696 22080 6702 22092
rect 6825 22083 6883 22089
rect 6825 22080 6837 22083
rect 6696 22052 6837 22080
rect 6696 22040 6702 22052
rect 6825 22049 6837 22052
rect 6871 22049 6883 22083
rect 6825 22043 6883 22049
rect 15102 22040 15108 22092
rect 15160 22080 15166 22092
rect 15562 22089 15568 22092
rect 15545 22083 15568 22089
rect 15545 22080 15557 22083
rect 15160 22052 15557 22080
rect 15160 22040 15166 22052
rect 15545 22049 15557 22052
rect 15620 22080 15626 22092
rect 15620 22052 15693 22080
rect 15545 22043 15568 22049
rect 15562 22040 15568 22043
rect 15620 22040 15626 22052
rect 3559 21984 4108 22012
rect 3559 21981 3571 21984
rect 3513 21975 3571 21981
rect 4154 21972 4160 22024
rect 4212 22012 4218 22024
rect 4522 22012 4528 22024
rect 4212 21984 4528 22012
rect 4212 21972 4218 21984
rect 4522 21972 4528 21984
rect 4580 21972 4586 22024
rect 4617 22015 4675 22021
rect 4617 21981 4629 22015
rect 4663 21981 4675 22015
rect 4617 21975 4675 21981
rect 4065 21947 4123 21953
rect 4065 21944 4077 21947
rect 2884 21916 4077 21944
rect 2777 21907 2835 21913
rect 4065 21913 4077 21916
rect 4111 21913 4123 21947
rect 4632 21944 4660 21975
rect 6546 21972 6552 22024
rect 6604 22012 6610 22024
rect 6917 22015 6975 22021
rect 6917 22012 6929 22015
rect 6604 21984 6929 22012
rect 6604 21972 6610 21984
rect 6917 21981 6929 21984
rect 6963 21981 6975 22015
rect 6917 21975 6975 21981
rect 7101 22015 7159 22021
rect 7101 21981 7113 22015
rect 7147 21981 7159 22015
rect 10962 22012 10968 22024
rect 10923 21984 10968 22012
rect 7101 21975 7159 21981
rect 4065 21907 4123 21913
rect 4172 21916 4660 21944
rect 6457 21947 6515 21953
rect 4172 21888 4200 21916
rect 6457 21913 6469 21947
rect 6503 21944 6515 21947
rect 6822 21944 6828 21956
rect 6503 21916 6828 21944
rect 6503 21913 6515 21916
rect 6457 21907 6515 21913
rect 6822 21904 6828 21916
rect 6880 21904 6886 21956
rect 7116 21944 7144 21975
rect 10962 21972 10968 21984
rect 11020 21972 11026 22024
rect 11057 22015 11115 22021
rect 11057 21981 11069 22015
rect 11103 21981 11115 22015
rect 11057 21975 11115 21981
rect 7561 21947 7619 21953
rect 7561 21944 7573 21947
rect 7116 21916 7573 21944
rect 7561 21913 7573 21916
rect 7607 21944 7619 21947
rect 7742 21944 7748 21956
rect 7607 21916 7748 21944
rect 7607 21913 7619 21916
rect 7561 21907 7619 21913
rect 7742 21904 7748 21916
rect 7800 21904 7806 21956
rect 9582 21904 9588 21956
rect 9640 21944 9646 21956
rect 10505 21947 10563 21953
rect 10505 21944 10517 21947
rect 9640 21916 10517 21944
rect 9640 21904 9646 21916
rect 10505 21913 10517 21916
rect 10551 21913 10563 21947
rect 11072 21944 11100 21975
rect 13630 21972 13636 22024
rect 13688 22012 13694 22024
rect 13817 22015 13875 22021
rect 13817 22012 13829 22015
rect 13688 21984 13829 22012
rect 13688 21972 13694 21984
rect 13817 21981 13829 21984
rect 13863 21981 13875 22015
rect 13817 21975 13875 21981
rect 13909 22015 13967 22021
rect 13909 21981 13921 22015
rect 13955 21981 13967 22015
rect 15286 22012 15292 22024
rect 15247 21984 15292 22012
rect 13909 21975 13967 21981
rect 10505 21907 10563 21913
rect 10980 21916 11100 21944
rect 4154 21836 4160 21888
rect 4212 21836 4218 21888
rect 4338 21836 4344 21888
rect 4396 21876 4402 21888
rect 4614 21876 4620 21888
rect 4396 21848 4620 21876
rect 4396 21836 4402 21848
rect 4614 21836 4620 21848
rect 4672 21836 4678 21888
rect 6270 21836 6276 21888
rect 6328 21876 6334 21888
rect 6365 21879 6423 21885
rect 6365 21876 6377 21879
rect 6328 21848 6377 21876
rect 6328 21836 6334 21848
rect 6365 21845 6377 21848
rect 6411 21876 6423 21879
rect 7098 21876 7104 21888
rect 6411 21848 7104 21876
rect 6411 21845 6423 21848
rect 6365 21839 6423 21845
rect 7098 21836 7104 21848
rect 7156 21836 7162 21888
rect 7650 21836 7656 21888
rect 7708 21876 7714 21888
rect 7837 21879 7895 21885
rect 7837 21876 7849 21879
rect 7708 21848 7849 21876
rect 7708 21836 7714 21848
rect 7837 21845 7849 21848
rect 7883 21845 7895 21879
rect 9030 21876 9036 21888
rect 8991 21848 9036 21876
rect 7837 21839 7895 21845
rect 9030 21836 9036 21848
rect 9088 21876 9094 21888
rect 9950 21876 9956 21888
rect 9088 21848 9956 21876
rect 9088 21836 9094 21848
rect 9950 21836 9956 21848
rect 10008 21876 10014 21888
rect 10321 21879 10379 21885
rect 10321 21876 10333 21879
rect 10008 21848 10333 21876
rect 10008 21836 10014 21848
rect 10321 21845 10333 21848
rect 10367 21876 10379 21879
rect 10980 21876 11008 21916
rect 13722 21904 13728 21956
rect 13780 21944 13786 21956
rect 13924 21944 13952 21975
rect 15286 21972 15292 21984
rect 15344 21972 15350 22024
rect 16666 21944 16672 21956
rect 13780 21916 13952 21944
rect 16627 21916 16672 21944
rect 13780 21904 13786 21916
rect 16666 21904 16672 21916
rect 16724 21904 16730 21956
rect 11514 21876 11520 21888
rect 10367 21848 11008 21876
rect 11475 21848 11520 21876
rect 10367 21845 10379 21848
rect 10321 21839 10379 21845
rect 11514 21836 11520 21848
rect 11572 21836 11578 21888
rect 13354 21876 13360 21888
rect 13315 21848 13360 21876
rect 13354 21836 13360 21848
rect 13412 21836 13418 21888
rect 14458 21876 14464 21888
rect 14419 21848 14464 21876
rect 14458 21836 14464 21848
rect 14516 21836 14522 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1302 21632 1308 21684
rect 1360 21672 1366 21684
rect 1673 21675 1731 21681
rect 1673 21672 1685 21675
rect 1360 21644 1685 21672
rect 1360 21632 1366 21644
rect 1673 21641 1685 21644
rect 1719 21672 1731 21675
rect 2133 21675 2191 21681
rect 2133 21672 2145 21675
rect 1719 21644 2145 21672
rect 1719 21641 1731 21644
rect 1673 21635 1731 21641
rect 2133 21641 2145 21644
rect 2179 21672 2191 21675
rect 2590 21672 2596 21684
rect 2179 21644 2596 21672
rect 2179 21641 2191 21644
rect 2133 21635 2191 21641
rect 2240 21545 2268 21644
rect 2590 21632 2596 21644
rect 2648 21632 2654 21684
rect 3602 21632 3608 21684
rect 3660 21672 3666 21684
rect 4709 21675 4767 21681
rect 4709 21672 4721 21675
rect 3660 21644 4721 21672
rect 3660 21632 3666 21644
rect 4709 21641 4721 21644
rect 4755 21672 4767 21675
rect 8202 21672 8208 21684
rect 4755 21644 8208 21672
rect 4755 21641 4767 21644
rect 4709 21635 4767 21641
rect 5368 21545 5396 21644
rect 8202 21632 8208 21644
rect 8260 21632 8266 21684
rect 10597 21675 10655 21681
rect 10597 21641 10609 21675
rect 10643 21672 10655 21675
rect 10870 21672 10876 21684
rect 10643 21644 10876 21672
rect 10643 21641 10655 21644
rect 10597 21635 10655 21641
rect 10870 21632 10876 21644
rect 10928 21632 10934 21684
rect 13541 21675 13599 21681
rect 13541 21641 13553 21675
rect 13587 21672 13599 21675
rect 13722 21672 13728 21684
rect 13587 21644 13728 21672
rect 13587 21641 13599 21644
rect 13541 21635 13599 21641
rect 13722 21632 13728 21644
rect 13780 21632 13786 21684
rect 15562 21672 15568 21684
rect 15523 21644 15568 21672
rect 15562 21632 15568 21644
rect 15620 21632 15626 21684
rect 2225 21539 2283 21545
rect 2225 21505 2237 21539
rect 2271 21505 2283 21539
rect 2225 21499 2283 21505
rect 5353 21539 5411 21545
rect 5353 21505 5365 21539
rect 5399 21505 5411 21539
rect 5353 21499 5411 21505
rect 5442 21496 5448 21548
rect 5500 21536 5506 21548
rect 7653 21539 7711 21545
rect 5500 21508 5545 21536
rect 5500 21496 5506 21508
rect 7653 21505 7665 21539
rect 7699 21536 7711 21539
rect 8021 21539 8079 21545
rect 8021 21536 8033 21539
rect 7699 21508 8033 21536
rect 7699 21505 7711 21508
rect 7653 21499 7711 21505
rect 8021 21505 8033 21508
rect 8067 21536 8079 21539
rect 8202 21536 8208 21548
rect 8067 21508 8208 21536
rect 8067 21505 8079 21508
rect 8021 21499 8079 21505
rect 8202 21496 8208 21508
rect 8260 21496 8266 21548
rect 9030 21496 9036 21548
rect 9088 21536 9094 21548
rect 9493 21539 9551 21545
rect 9493 21536 9505 21539
rect 9088 21508 9505 21536
rect 9088 21496 9094 21508
rect 9493 21505 9505 21508
rect 9539 21505 9551 21539
rect 9493 21499 9551 21505
rect 11054 21496 11060 21548
rect 11112 21536 11118 21548
rect 11333 21539 11391 21545
rect 11333 21536 11345 21539
rect 11112 21508 11345 21536
rect 11112 21496 11118 21508
rect 11333 21505 11345 21508
rect 11379 21536 11391 21539
rect 12066 21536 12072 21548
rect 11379 21508 12072 21536
rect 11379 21505 11391 21508
rect 11333 21499 11391 21505
rect 12066 21496 12072 21508
rect 12124 21536 12130 21548
rect 12989 21539 13047 21545
rect 12989 21536 13001 21539
rect 12124 21508 13001 21536
rect 12124 21496 12130 21508
rect 12989 21505 13001 21508
rect 13035 21505 13047 21539
rect 12989 21499 13047 21505
rect 13722 21496 13728 21548
rect 13780 21536 13786 21548
rect 13906 21536 13912 21548
rect 13780 21508 13912 21536
rect 13780 21496 13786 21508
rect 13906 21496 13912 21508
rect 13964 21496 13970 21548
rect 1854 21428 1860 21480
rect 1912 21468 1918 21480
rect 6089 21471 6147 21477
rect 6089 21468 6101 21471
rect 1912 21440 6101 21468
rect 1912 21428 1918 21440
rect 6089 21437 6101 21440
rect 6135 21468 6147 21471
rect 6638 21468 6644 21480
rect 6135 21440 6644 21468
rect 6135 21437 6147 21440
rect 6089 21431 6147 21437
rect 6638 21428 6644 21440
rect 6696 21428 6702 21480
rect 11149 21471 11207 21477
rect 11149 21437 11161 21471
rect 11195 21468 11207 21471
rect 11238 21468 11244 21480
rect 11195 21440 11244 21468
rect 11195 21437 11207 21440
rect 11149 21431 11207 21437
rect 11238 21428 11244 21440
rect 11296 21428 11302 21480
rect 12253 21471 12311 21477
rect 12253 21437 12265 21471
rect 12299 21468 12311 21471
rect 12805 21471 12863 21477
rect 12805 21468 12817 21471
rect 12299 21440 12817 21468
rect 12299 21437 12311 21440
rect 12253 21431 12311 21437
rect 12805 21437 12817 21440
rect 12851 21468 12863 21471
rect 13998 21468 14004 21480
rect 12851 21440 14004 21468
rect 12851 21437 12863 21440
rect 12805 21431 12863 21437
rect 13998 21428 14004 21440
rect 14056 21428 14062 21480
rect 14182 21468 14188 21480
rect 14143 21440 14188 21468
rect 14182 21428 14188 21440
rect 14240 21428 14246 21480
rect 2314 21360 2320 21412
rect 2372 21400 2378 21412
rect 2470 21403 2528 21409
rect 2470 21400 2482 21403
rect 2372 21372 2482 21400
rect 2372 21360 2378 21372
rect 2470 21369 2482 21372
rect 2516 21369 2528 21403
rect 2470 21363 2528 21369
rect 4433 21403 4491 21409
rect 4433 21369 4445 21403
rect 4479 21400 4491 21403
rect 7377 21403 7435 21409
rect 4479 21372 5304 21400
rect 4479 21369 4491 21372
rect 4433 21363 4491 21369
rect 5276 21344 5304 21372
rect 7377 21369 7389 21403
rect 7423 21400 7435 21403
rect 7558 21400 7564 21412
rect 7423 21372 7564 21400
rect 7423 21369 7435 21372
rect 7377 21363 7435 21369
rect 7558 21360 7564 21372
rect 7616 21400 7622 21412
rect 8389 21403 8447 21409
rect 8389 21400 8401 21403
rect 7616 21372 8401 21400
rect 7616 21360 7622 21372
rect 8389 21369 8401 21372
rect 8435 21369 8447 21403
rect 8389 21363 8447 21369
rect 8478 21360 8484 21412
rect 8536 21400 8542 21412
rect 8849 21403 8907 21409
rect 8849 21400 8861 21403
rect 8536 21372 8861 21400
rect 8536 21360 8542 21372
rect 8849 21369 8861 21372
rect 8895 21400 8907 21403
rect 9401 21403 9459 21409
rect 9401 21400 9413 21403
rect 8895 21372 9413 21400
rect 8895 21369 8907 21372
rect 8849 21363 8907 21369
rect 9401 21369 9413 21372
rect 9447 21369 9459 21403
rect 9401 21363 9459 21369
rect 10229 21403 10287 21409
rect 10229 21369 10241 21403
rect 10275 21400 10287 21403
rect 10870 21400 10876 21412
rect 10275 21372 10876 21400
rect 10275 21369 10287 21372
rect 10229 21363 10287 21369
rect 10870 21360 10876 21372
rect 10928 21360 10934 21412
rect 11885 21403 11943 21409
rect 11885 21369 11897 21403
rect 11931 21400 11943 21403
rect 11931 21372 12940 21400
rect 11931 21369 11943 21372
rect 11885 21363 11943 21369
rect 3602 21332 3608 21344
rect 3563 21304 3608 21332
rect 3602 21292 3608 21304
rect 3660 21292 3666 21344
rect 4893 21335 4951 21341
rect 4893 21301 4905 21335
rect 4939 21332 4951 21335
rect 5166 21332 5172 21344
rect 4939 21304 5172 21332
rect 4939 21301 4951 21304
rect 4893 21295 4951 21301
rect 5166 21292 5172 21304
rect 5224 21292 5230 21344
rect 5258 21292 5264 21344
rect 5316 21332 5322 21344
rect 6546 21332 6552 21344
rect 5316 21304 5361 21332
rect 6507 21304 6552 21332
rect 5316 21292 5322 21304
rect 6546 21292 6552 21304
rect 6604 21292 6610 21344
rect 7006 21332 7012 21344
rect 6967 21304 7012 21332
rect 7006 21292 7012 21304
rect 7064 21292 7070 21344
rect 7469 21335 7527 21341
rect 7469 21301 7481 21335
rect 7515 21332 7527 21335
rect 7650 21332 7656 21344
rect 7515 21304 7656 21332
rect 7515 21301 7527 21304
rect 7469 21295 7527 21301
rect 7650 21292 7656 21304
rect 7708 21292 7714 21344
rect 8938 21332 8944 21344
rect 8899 21304 8944 21332
rect 8938 21292 8944 21304
rect 8996 21292 9002 21344
rect 9030 21292 9036 21344
rect 9088 21332 9094 21344
rect 9309 21335 9367 21341
rect 9309 21332 9321 21335
rect 9088 21304 9321 21332
rect 9088 21292 9094 21304
rect 9309 21301 9321 21304
rect 9355 21301 9367 21335
rect 9309 21295 9367 21301
rect 10781 21335 10839 21341
rect 10781 21301 10793 21335
rect 10827 21332 10839 21335
rect 10962 21332 10968 21344
rect 10827 21304 10968 21332
rect 10827 21301 10839 21304
rect 10781 21295 10839 21301
rect 10962 21292 10968 21304
rect 11020 21292 11026 21344
rect 11241 21335 11299 21341
rect 11241 21301 11253 21335
rect 11287 21332 11299 21335
rect 11514 21332 11520 21344
rect 11287 21304 11520 21332
rect 11287 21301 11299 21304
rect 11241 21295 11299 21301
rect 11514 21292 11520 21304
rect 11572 21292 11578 21344
rect 12342 21292 12348 21344
rect 12400 21332 12406 21344
rect 12912 21341 12940 21372
rect 13906 21360 13912 21412
rect 13964 21400 13970 21412
rect 14458 21409 14464 21412
rect 14430 21403 14464 21409
rect 14430 21400 14442 21403
rect 13964 21372 14442 21400
rect 13964 21360 13970 21372
rect 14430 21369 14442 21372
rect 14516 21400 14522 21412
rect 14516 21372 14578 21400
rect 14430 21363 14464 21369
rect 14458 21360 14464 21363
rect 14516 21360 14522 21372
rect 26234 21360 26240 21412
rect 26292 21400 26298 21412
rect 27614 21400 27620 21412
rect 26292 21372 27620 21400
rect 26292 21360 26298 21372
rect 27614 21360 27620 21372
rect 27672 21360 27678 21412
rect 12437 21335 12495 21341
rect 12437 21332 12449 21335
rect 12400 21304 12449 21332
rect 12400 21292 12406 21304
rect 12437 21301 12449 21304
rect 12483 21301 12495 21335
rect 12437 21295 12495 21301
rect 12897 21335 12955 21341
rect 12897 21301 12909 21335
rect 12943 21332 12955 21335
rect 13722 21332 13728 21344
rect 12943 21304 13728 21332
rect 12943 21301 12955 21304
rect 12897 21295 12955 21301
rect 13722 21292 13728 21304
rect 13780 21292 13786 21344
rect 14093 21335 14151 21341
rect 14093 21301 14105 21335
rect 14139 21332 14151 21335
rect 14182 21332 14188 21344
rect 14139 21304 14188 21332
rect 14139 21301 14151 21304
rect 14093 21295 14151 21301
rect 14182 21292 14188 21304
rect 14240 21332 14246 21344
rect 15286 21332 15292 21344
rect 14240 21304 15292 21332
rect 14240 21292 14246 21304
rect 15286 21292 15292 21304
rect 15344 21332 15350 21344
rect 16117 21335 16175 21341
rect 16117 21332 16129 21335
rect 15344 21304 16129 21332
rect 15344 21292 15350 21304
rect 16117 21301 16129 21304
rect 16163 21301 16175 21335
rect 16117 21295 16175 21301
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1670 21128 1676 21140
rect 1631 21100 1676 21128
rect 1670 21088 1676 21100
rect 1728 21088 1734 21140
rect 2314 21128 2320 21140
rect 2275 21100 2320 21128
rect 2314 21088 2320 21100
rect 2372 21088 2378 21140
rect 2498 21088 2504 21140
rect 2556 21128 2562 21140
rect 2593 21131 2651 21137
rect 2593 21128 2605 21131
rect 2556 21100 2605 21128
rect 2556 21088 2562 21100
rect 2593 21097 2605 21100
rect 2639 21097 2651 21131
rect 2593 21091 2651 21097
rect 3513 21131 3571 21137
rect 3513 21097 3525 21131
rect 3559 21128 3571 21131
rect 4522 21128 4528 21140
rect 3559 21100 4528 21128
rect 3559 21097 3571 21100
rect 3513 21091 3571 21097
rect 4522 21088 4528 21100
rect 4580 21088 4586 21140
rect 5534 21088 5540 21140
rect 5592 21128 5598 21140
rect 5721 21131 5779 21137
rect 5721 21128 5733 21131
rect 5592 21100 5733 21128
rect 5592 21088 5598 21100
rect 5721 21097 5733 21100
rect 5767 21097 5779 21131
rect 5721 21091 5779 21097
rect 6086 21088 6092 21140
rect 6144 21128 6150 21140
rect 6273 21131 6331 21137
rect 6273 21128 6285 21131
rect 6144 21100 6285 21128
rect 6144 21088 6150 21100
rect 6273 21097 6285 21100
rect 6319 21097 6331 21131
rect 6273 21091 6331 21097
rect 7469 21131 7527 21137
rect 7469 21097 7481 21131
rect 7515 21128 7527 21131
rect 7558 21128 7564 21140
rect 7515 21100 7564 21128
rect 7515 21097 7527 21100
rect 7469 21091 7527 21097
rect 7558 21088 7564 21100
rect 7616 21088 7622 21140
rect 9030 21128 9036 21140
rect 8991 21100 9036 21128
rect 9030 21088 9036 21100
rect 9088 21088 9094 21140
rect 13449 21131 13507 21137
rect 13449 21097 13461 21131
rect 13495 21128 13507 21131
rect 13630 21128 13636 21140
rect 13495 21100 13636 21128
rect 13495 21097 13507 21100
rect 13449 21091 13507 21097
rect 13630 21088 13636 21100
rect 13688 21088 13694 21140
rect 15562 21128 15568 21140
rect 15523 21100 15568 21128
rect 15562 21088 15568 21100
rect 15620 21088 15626 21140
rect 9950 21069 9956 21072
rect 9944 21060 9956 21069
rect 9911 21032 9956 21060
rect 9944 21023 9956 21032
rect 9950 21020 9956 21023
rect 10008 21020 10014 21072
rect 13081 21063 13139 21069
rect 13081 21060 13093 21063
rect 12084 21032 13093 21060
rect 4062 20992 4068 21004
rect 3804 20964 4068 20992
rect 1670 20884 1676 20936
rect 1728 20924 1734 20936
rect 3804 20933 3832 20964
rect 4062 20952 4068 20964
rect 4120 20952 4126 21004
rect 4709 20995 4767 21001
rect 4709 20961 4721 20995
rect 4755 20992 4767 20995
rect 5166 20992 5172 21004
rect 4755 20964 5172 20992
rect 4755 20961 4767 20964
rect 4709 20955 4767 20961
rect 5166 20952 5172 20964
rect 5224 20952 5230 21004
rect 7282 20952 7288 21004
rect 7340 20992 7346 21004
rect 7837 20995 7895 21001
rect 7837 20992 7849 20995
rect 7340 20964 7849 20992
rect 7340 20952 7346 20964
rect 7837 20961 7849 20964
rect 7883 20961 7895 20995
rect 7837 20955 7895 20961
rect 9677 20995 9735 21001
rect 9677 20961 9689 20995
rect 9723 20992 9735 20995
rect 9766 20992 9772 21004
rect 9723 20964 9772 20992
rect 9723 20961 9735 20964
rect 9677 20955 9735 20961
rect 9766 20952 9772 20964
rect 9824 20952 9830 21004
rect 12084 20992 12112 21032
rect 13081 21029 13093 21032
rect 13127 21060 13139 21063
rect 13354 21060 13360 21072
rect 13127 21032 13360 21060
rect 13127 21029 13139 21032
rect 13081 21023 13139 21029
rect 13354 21020 13360 21032
rect 13412 21020 13418 21072
rect 12153 20995 12211 21001
rect 12153 20992 12165 20995
rect 12084 20964 12165 20992
rect 12153 20961 12165 20964
rect 12199 20961 12211 20995
rect 13998 20992 14004 21004
rect 13959 20964 14004 20992
rect 12153 20955 12211 20961
rect 13998 20952 14004 20964
rect 14056 20952 14062 21004
rect 14093 20995 14151 21001
rect 14093 20961 14105 20995
rect 14139 20992 14151 20995
rect 14734 20992 14740 21004
rect 14139 20964 14740 20992
rect 14139 20961 14151 20964
rect 14093 20955 14151 20961
rect 14734 20952 14740 20964
rect 14792 20952 14798 21004
rect 3789 20927 3847 20933
rect 3789 20924 3801 20927
rect 1728 20896 3801 20924
rect 1728 20884 1734 20896
rect 3789 20893 3801 20896
rect 3835 20893 3847 20927
rect 3789 20887 3847 20893
rect 4154 20884 4160 20936
rect 4212 20924 4218 20936
rect 4801 20927 4859 20933
rect 4801 20924 4813 20927
rect 4212 20896 4813 20924
rect 4212 20884 4218 20896
rect 4801 20893 4813 20896
rect 4847 20893 4859 20927
rect 4801 20887 4859 20893
rect 3602 20816 3608 20868
rect 3660 20856 3666 20868
rect 4816 20856 4844 20887
rect 4890 20884 4896 20936
rect 4948 20924 4954 20936
rect 4948 20896 4993 20924
rect 4948 20884 4954 20896
rect 5994 20884 6000 20936
rect 6052 20924 6058 20936
rect 6362 20924 6368 20936
rect 6052 20896 6368 20924
rect 6052 20884 6058 20896
rect 6362 20884 6368 20896
rect 6420 20884 6426 20936
rect 6457 20927 6515 20933
rect 6457 20893 6469 20927
rect 6503 20893 6515 20927
rect 6457 20887 6515 20893
rect 5905 20859 5963 20865
rect 5905 20856 5917 20859
rect 3660 20828 4752 20856
rect 4816 20828 5917 20856
rect 3660 20816 3666 20828
rect 1486 20748 1492 20800
rect 1544 20788 1550 20800
rect 2314 20788 2320 20800
rect 1544 20760 2320 20788
rect 1544 20748 1550 20760
rect 2314 20748 2320 20760
rect 2372 20748 2378 20800
rect 4154 20748 4160 20800
rect 4212 20788 4218 20800
rect 4341 20791 4399 20797
rect 4341 20788 4353 20791
rect 4212 20760 4353 20788
rect 4212 20748 4218 20760
rect 4341 20757 4353 20760
rect 4387 20757 4399 20791
rect 4724 20788 4752 20828
rect 5905 20825 5917 20828
rect 5951 20825 5963 20859
rect 5905 20819 5963 20825
rect 5353 20791 5411 20797
rect 5353 20788 5365 20791
rect 4724 20760 5365 20788
rect 4341 20751 4399 20757
rect 5353 20757 5365 20760
rect 5399 20788 5411 20791
rect 5442 20788 5448 20800
rect 5399 20760 5448 20788
rect 5399 20757 5411 20760
rect 5353 20751 5411 20757
rect 5442 20748 5448 20760
rect 5500 20788 5506 20800
rect 6178 20788 6184 20800
rect 5500 20760 6184 20788
rect 5500 20748 5506 20760
rect 6178 20748 6184 20760
rect 6236 20788 6242 20800
rect 6472 20788 6500 20887
rect 7190 20884 7196 20936
rect 7248 20924 7254 20936
rect 7929 20927 7987 20933
rect 7929 20924 7941 20927
rect 7248 20896 7941 20924
rect 7248 20884 7254 20896
rect 7929 20893 7941 20896
rect 7975 20893 7987 20927
rect 7929 20887 7987 20893
rect 8113 20927 8171 20933
rect 8113 20893 8125 20927
rect 8159 20924 8171 20927
rect 8159 20896 8524 20924
rect 8159 20893 8171 20896
rect 8113 20887 8171 20893
rect 7282 20856 7288 20868
rect 7243 20828 7288 20856
rect 7282 20816 7288 20828
rect 7340 20816 7346 20868
rect 8496 20800 8524 20896
rect 12066 20884 12072 20936
rect 12124 20924 12130 20936
rect 12621 20927 12679 20933
rect 12621 20924 12633 20927
rect 12124 20896 12633 20924
rect 12124 20884 12130 20896
rect 12621 20893 12633 20896
rect 12667 20893 12679 20927
rect 12621 20887 12679 20893
rect 14277 20927 14335 20933
rect 14277 20893 14289 20927
rect 14323 20924 14335 20927
rect 15562 20924 15568 20936
rect 14323 20896 15568 20924
rect 14323 20893 14335 20896
rect 14277 20887 14335 20893
rect 15562 20884 15568 20896
rect 15620 20884 15626 20936
rect 6236 20760 6500 20788
rect 7009 20791 7067 20797
rect 6236 20748 6242 20760
rect 7009 20757 7021 20791
rect 7055 20788 7067 20791
rect 7742 20788 7748 20800
rect 7055 20760 7748 20788
rect 7055 20757 7067 20760
rect 7009 20751 7067 20757
rect 7742 20748 7748 20760
rect 7800 20748 7806 20800
rect 8478 20788 8484 20800
rect 8439 20760 8484 20788
rect 8478 20748 8484 20760
rect 8536 20748 8542 20800
rect 11054 20788 11060 20800
rect 11015 20760 11060 20788
rect 11054 20748 11060 20760
rect 11112 20748 11118 20800
rect 11238 20748 11244 20800
rect 11296 20788 11302 20800
rect 11609 20791 11667 20797
rect 11609 20788 11621 20791
rect 11296 20760 11621 20788
rect 11296 20748 11302 20760
rect 11609 20757 11621 20760
rect 11655 20757 11667 20791
rect 11609 20751 11667 20757
rect 11698 20748 11704 20800
rect 11756 20788 11762 20800
rect 12345 20791 12403 20797
rect 12345 20788 12357 20791
rect 11756 20760 12357 20788
rect 11756 20748 11762 20760
rect 12345 20757 12357 20760
rect 12391 20757 12403 20791
rect 12345 20751 12403 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1486 20544 1492 20596
rect 1544 20584 1550 20596
rect 1946 20584 1952 20596
rect 1544 20556 1952 20584
rect 1544 20544 1550 20556
rect 1946 20544 1952 20556
rect 2004 20544 2010 20596
rect 2130 20544 2136 20596
rect 2188 20584 2194 20596
rect 2317 20587 2375 20593
rect 2317 20584 2329 20587
rect 2188 20556 2329 20584
rect 2188 20544 2194 20556
rect 2317 20553 2329 20556
rect 2363 20553 2375 20587
rect 2317 20547 2375 20553
rect 4801 20587 4859 20593
rect 4801 20553 4813 20587
rect 4847 20584 4859 20587
rect 4890 20584 4896 20596
rect 4847 20556 4896 20584
rect 4847 20553 4859 20556
rect 4801 20547 4859 20553
rect 4890 20544 4896 20556
rect 4948 20544 4954 20596
rect 5534 20584 5540 20596
rect 5495 20556 5540 20584
rect 5534 20544 5540 20556
rect 5592 20544 5598 20596
rect 6086 20544 6092 20596
rect 6144 20584 6150 20596
rect 6273 20587 6331 20593
rect 6273 20584 6285 20587
rect 6144 20556 6285 20584
rect 6144 20544 6150 20556
rect 6273 20553 6285 20556
rect 6319 20584 6331 20587
rect 7190 20584 7196 20596
rect 6319 20556 7196 20584
rect 6319 20553 6331 20556
rect 6273 20547 6331 20553
rect 7190 20544 7196 20556
rect 7248 20544 7254 20596
rect 8294 20544 8300 20596
rect 8352 20584 8358 20596
rect 8757 20587 8815 20593
rect 8757 20584 8769 20587
rect 8352 20556 8769 20584
rect 8352 20544 8358 20556
rect 8757 20553 8769 20556
rect 8803 20584 8815 20587
rect 9309 20587 9367 20593
rect 9309 20584 9321 20587
rect 8803 20556 9321 20584
rect 8803 20553 8815 20556
rect 8757 20547 8815 20553
rect 9309 20553 9321 20556
rect 9355 20553 9367 20587
rect 9309 20547 9367 20553
rect 3329 20451 3387 20457
rect 3329 20417 3341 20451
rect 3375 20448 3387 20451
rect 3418 20448 3424 20460
rect 3375 20420 3424 20448
rect 3375 20417 3387 20420
rect 3329 20411 3387 20417
rect 3418 20408 3424 20420
rect 3476 20408 3482 20460
rect 9324 20448 9352 20547
rect 10042 20544 10048 20596
rect 10100 20584 10106 20596
rect 11241 20587 11299 20593
rect 11241 20584 11253 20587
rect 10100 20556 11253 20584
rect 10100 20544 10106 20556
rect 11241 20553 11253 20556
rect 11287 20553 11299 20587
rect 11241 20547 11299 20553
rect 11885 20587 11943 20593
rect 11885 20553 11897 20587
rect 11931 20584 11943 20587
rect 12066 20584 12072 20596
rect 11931 20556 12072 20584
rect 11931 20553 11943 20556
rect 11885 20547 11943 20553
rect 12066 20544 12072 20556
rect 12124 20544 12130 20596
rect 15197 20587 15255 20593
rect 15197 20553 15209 20587
rect 15243 20584 15255 20587
rect 15562 20584 15568 20596
rect 15243 20556 15568 20584
rect 15243 20553 15255 20556
rect 15197 20547 15255 20553
rect 15562 20544 15568 20556
rect 15620 20544 15626 20596
rect 9324 20420 9996 20448
rect 1489 20383 1547 20389
rect 1489 20349 1501 20383
rect 1535 20380 1547 20383
rect 2961 20383 3019 20389
rect 1535 20352 2084 20380
rect 1535 20349 1547 20352
rect 1489 20343 1547 20349
rect 2056 20256 2084 20352
rect 2961 20349 2973 20383
rect 3007 20380 3019 20383
rect 4062 20380 4068 20392
rect 3007 20352 4068 20380
rect 3007 20349 3019 20352
rect 2961 20343 3019 20349
rect 4062 20340 4068 20352
rect 4120 20340 4126 20392
rect 7098 20340 7104 20392
rect 7156 20380 7162 20392
rect 7377 20383 7435 20389
rect 7377 20380 7389 20383
rect 7156 20352 7389 20380
rect 7156 20340 7162 20352
rect 7377 20349 7389 20352
rect 7423 20380 7435 20383
rect 8018 20380 8024 20392
rect 7423 20352 8024 20380
rect 7423 20349 7435 20352
rect 7377 20343 7435 20349
rect 8018 20340 8024 20352
rect 8076 20340 8082 20392
rect 9861 20383 9919 20389
rect 9861 20380 9873 20383
rect 9784 20352 9873 20380
rect 3602 20272 3608 20324
rect 3660 20321 3666 20324
rect 3660 20315 3724 20321
rect 3660 20281 3678 20315
rect 3712 20281 3724 20315
rect 3660 20275 3724 20281
rect 7644 20315 7702 20321
rect 7644 20281 7656 20315
rect 7690 20312 7702 20315
rect 8478 20312 8484 20324
rect 7690 20284 8484 20312
rect 7690 20281 7702 20284
rect 7644 20275 7702 20281
rect 3660 20272 3666 20275
rect 8478 20272 8484 20284
rect 8536 20272 8542 20324
rect 9784 20256 9812 20352
rect 9861 20349 9873 20352
rect 9907 20349 9919 20383
rect 9968 20380 9996 20420
rect 10117 20383 10175 20389
rect 10117 20380 10129 20383
rect 9968 20352 10129 20380
rect 9861 20343 9919 20349
rect 10117 20349 10129 20352
rect 10163 20349 10175 20383
rect 10117 20343 10175 20349
rect 12253 20383 12311 20389
rect 12253 20349 12265 20383
rect 12299 20380 12311 20383
rect 12434 20380 12440 20392
rect 12299 20352 12440 20380
rect 12299 20349 12311 20352
rect 12253 20343 12311 20349
rect 12434 20340 12440 20352
rect 12492 20380 12498 20392
rect 12492 20352 12585 20380
rect 12492 20340 12498 20352
rect 12066 20272 12072 20324
rect 12124 20312 12130 20324
rect 12682 20315 12740 20321
rect 12682 20312 12694 20315
rect 12124 20284 12694 20312
rect 12124 20272 12130 20284
rect 12682 20281 12694 20284
rect 12728 20281 12740 20315
rect 12682 20275 12740 20281
rect 13998 20272 14004 20324
rect 14056 20312 14062 20324
rect 14461 20315 14519 20321
rect 14461 20312 14473 20315
rect 14056 20284 14473 20312
rect 14056 20272 14062 20284
rect 14461 20281 14473 20284
rect 14507 20312 14519 20315
rect 14642 20312 14648 20324
rect 14507 20284 14648 20312
rect 14507 20281 14519 20284
rect 14461 20275 14519 20281
rect 14642 20272 14648 20284
rect 14700 20312 14706 20324
rect 14826 20312 14832 20324
rect 14700 20284 14832 20312
rect 14700 20272 14706 20284
rect 14826 20272 14832 20284
rect 14884 20272 14890 20324
rect 1670 20244 1676 20256
rect 1631 20216 1676 20244
rect 1670 20204 1676 20216
rect 1728 20204 1734 20256
rect 2038 20244 2044 20256
rect 1999 20216 2044 20244
rect 2038 20204 2044 20216
rect 2096 20204 2102 20256
rect 5994 20244 6000 20256
rect 5955 20216 6000 20244
rect 5994 20204 6000 20216
rect 6052 20204 6058 20256
rect 9766 20244 9772 20256
rect 9727 20216 9772 20244
rect 9766 20204 9772 20216
rect 9824 20204 9830 20256
rect 13630 20204 13636 20256
rect 13688 20244 13694 20256
rect 13817 20247 13875 20253
rect 13817 20244 13829 20247
rect 13688 20216 13829 20244
rect 13688 20204 13694 20216
rect 13817 20213 13829 20216
rect 13863 20213 13875 20247
rect 14734 20244 14740 20256
rect 14695 20216 14740 20244
rect 13817 20207 13875 20213
rect 14734 20204 14740 20216
rect 14792 20204 14798 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 2958 20040 2964 20052
rect 2919 20012 2964 20040
rect 2958 20000 2964 20012
rect 3016 20000 3022 20052
rect 3513 20043 3571 20049
rect 3513 20009 3525 20043
rect 3559 20040 3571 20043
rect 3602 20040 3608 20052
rect 3559 20012 3608 20040
rect 3559 20009 3571 20012
rect 3513 20003 3571 20009
rect 3602 20000 3608 20012
rect 3660 20000 3666 20052
rect 6638 20000 6644 20052
rect 6696 20040 6702 20052
rect 6914 20040 6920 20052
rect 6696 20012 6920 20040
rect 6696 20000 6702 20012
rect 6914 20000 6920 20012
rect 6972 20000 6978 20052
rect 7745 20043 7803 20049
rect 7745 20009 7757 20043
rect 7791 20040 7803 20043
rect 7834 20040 7840 20052
rect 7791 20012 7840 20040
rect 7791 20009 7803 20012
rect 7745 20003 7803 20009
rect 7834 20000 7840 20012
rect 7892 20000 7898 20052
rect 8018 20040 8024 20052
rect 7979 20012 8024 20040
rect 8018 20000 8024 20012
rect 8076 20000 8082 20052
rect 8573 20043 8631 20049
rect 8573 20009 8585 20043
rect 8619 20040 8631 20043
rect 9030 20040 9036 20052
rect 8619 20012 9036 20040
rect 8619 20009 8631 20012
rect 8573 20003 8631 20009
rect 9030 20000 9036 20012
rect 9088 20000 9094 20052
rect 10042 20000 10048 20052
rect 10100 20040 10106 20052
rect 10229 20043 10287 20049
rect 10229 20040 10241 20043
rect 10100 20012 10241 20040
rect 10100 20000 10106 20012
rect 10229 20009 10241 20012
rect 10275 20009 10287 20043
rect 10229 20003 10287 20009
rect 11885 20043 11943 20049
rect 11885 20009 11897 20043
rect 11931 20040 11943 20043
rect 12066 20040 12072 20052
rect 11931 20012 12072 20040
rect 11931 20009 11943 20012
rect 11885 20003 11943 20009
rect 12066 20000 12072 20012
rect 12124 20000 12130 20052
rect 3326 19932 3332 19984
rect 3384 19972 3390 19984
rect 3881 19975 3939 19981
rect 3881 19972 3893 19975
rect 3384 19944 3893 19972
rect 3384 19932 3390 19944
rect 3881 19941 3893 19944
rect 3927 19972 3939 19975
rect 4332 19975 4390 19981
rect 4332 19972 4344 19975
rect 3927 19944 4344 19972
rect 3927 19941 3939 19944
rect 3881 19935 3939 19941
rect 4332 19941 4344 19944
rect 4378 19972 4390 19975
rect 4890 19972 4896 19984
rect 4378 19944 4896 19972
rect 4378 19941 4390 19944
rect 4332 19935 4390 19941
rect 4890 19932 4896 19944
rect 4948 19932 4954 19984
rect 7098 19972 7104 19984
rect 5000 19944 7104 19972
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 1443 19876 2084 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 2056 19780 2084 19876
rect 2130 19864 2136 19916
rect 2188 19904 2194 19916
rect 3050 19904 3056 19916
rect 2188 19876 3056 19904
rect 2188 19864 2194 19876
rect 3050 19864 3056 19876
rect 3108 19864 3114 19916
rect 3418 19864 3424 19916
rect 3476 19904 3482 19916
rect 4065 19907 4123 19913
rect 4065 19904 4077 19907
rect 3476 19876 4077 19904
rect 3476 19864 3482 19876
rect 4065 19873 4077 19876
rect 4111 19904 4123 19907
rect 5000 19904 5028 19944
rect 7098 19932 7104 19944
rect 7156 19932 7162 19984
rect 8938 19932 8944 19984
rect 8996 19972 9002 19984
rect 9217 19975 9275 19981
rect 9217 19972 9229 19975
rect 8996 19944 9229 19972
rect 8996 19932 9002 19944
rect 9217 19941 9229 19944
rect 9263 19941 9275 19975
rect 9217 19935 9275 19941
rect 10772 19975 10830 19981
rect 10772 19941 10784 19975
rect 10818 19972 10830 19975
rect 11054 19972 11060 19984
rect 10818 19944 11060 19972
rect 10818 19941 10830 19944
rect 10772 19935 10830 19941
rect 11054 19932 11060 19944
rect 11112 19932 11118 19984
rect 4111 19876 5028 19904
rect 7009 19907 7067 19913
rect 4111 19873 4123 19876
rect 4065 19867 4123 19873
rect 7009 19873 7021 19907
rect 7055 19904 7067 19907
rect 7282 19904 7288 19916
rect 7055 19876 7288 19904
rect 7055 19873 7067 19876
rect 7009 19867 7067 19873
rect 7282 19864 7288 19876
rect 7340 19864 7346 19916
rect 13725 19907 13783 19913
rect 13725 19873 13737 19907
rect 13771 19904 13783 19907
rect 13998 19904 14004 19916
rect 13771 19876 14004 19904
rect 13771 19873 13783 19876
rect 13725 19867 13783 19873
rect 13998 19864 14004 19876
rect 14056 19904 14062 19916
rect 14737 19907 14795 19913
rect 14737 19904 14749 19907
rect 14056 19876 14749 19904
rect 14056 19864 14062 19876
rect 14737 19873 14749 19876
rect 14783 19873 14795 19907
rect 14737 19867 14795 19873
rect 7101 19839 7159 19845
rect 7101 19805 7113 19839
rect 7147 19805 7159 19839
rect 7101 19799 7159 19805
rect 2038 19768 2044 19780
rect 1999 19740 2044 19768
rect 2038 19728 2044 19740
rect 2096 19728 2102 19780
rect 6178 19728 6184 19780
rect 6236 19768 6242 19780
rect 7116 19768 7144 19799
rect 9766 19796 9772 19848
rect 9824 19836 9830 19848
rect 9953 19839 10011 19845
rect 9953 19836 9965 19839
rect 9824 19808 9965 19836
rect 9824 19796 9830 19808
rect 9953 19805 9965 19808
rect 9999 19836 10011 19839
rect 10502 19836 10508 19848
rect 9999 19808 10508 19836
rect 9999 19805 10011 19808
rect 9953 19799 10011 19805
rect 10502 19796 10508 19808
rect 10560 19796 10566 19848
rect 12713 19839 12771 19845
rect 12713 19805 12725 19839
rect 12759 19836 12771 19839
rect 13262 19836 13268 19848
rect 12759 19808 13268 19836
rect 12759 19805 12771 19808
rect 12713 19799 12771 19805
rect 13262 19796 13268 19808
rect 13320 19796 13326 19848
rect 13817 19839 13875 19845
rect 13817 19836 13829 19839
rect 13740 19808 13829 19836
rect 13740 19780 13768 19808
rect 13817 19805 13829 19808
rect 13863 19805 13875 19839
rect 13817 19799 13875 19805
rect 13906 19796 13912 19848
rect 13964 19836 13970 19848
rect 13964 19808 14009 19836
rect 13964 19796 13970 19808
rect 6236 19740 7144 19768
rect 13188 19740 13676 19768
rect 6236 19728 6242 19740
rect 13188 19712 13216 19740
rect 1394 19660 1400 19712
rect 1452 19700 1458 19712
rect 1581 19703 1639 19709
rect 1581 19700 1593 19703
rect 1452 19672 1593 19700
rect 1452 19660 1458 19672
rect 1581 19669 1593 19672
rect 1627 19669 1639 19703
rect 5442 19700 5448 19712
rect 5403 19672 5448 19700
rect 1581 19663 1639 19669
rect 5442 19660 5448 19672
rect 5500 19660 5506 19712
rect 5534 19660 5540 19712
rect 5592 19700 5598 19712
rect 6549 19703 6607 19709
rect 6549 19700 6561 19703
rect 5592 19672 6561 19700
rect 5592 19660 5598 19672
rect 6549 19669 6561 19672
rect 6595 19669 6607 19703
rect 8478 19700 8484 19712
rect 8439 19672 8484 19700
rect 6549 19663 6607 19669
rect 8478 19660 8484 19672
rect 8536 19660 8542 19712
rect 13081 19703 13139 19709
rect 13081 19669 13093 19703
rect 13127 19700 13139 19703
rect 13170 19700 13176 19712
rect 13127 19672 13176 19700
rect 13127 19669 13139 19672
rect 13081 19663 13139 19669
rect 13170 19660 13176 19672
rect 13228 19660 13234 19712
rect 13354 19700 13360 19712
rect 13315 19672 13360 19700
rect 13354 19660 13360 19672
rect 13412 19660 13418 19712
rect 13648 19700 13676 19740
rect 13722 19728 13728 19780
rect 13780 19728 13786 19780
rect 14369 19703 14427 19709
rect 14369 19700 14381 19703
rect 13648 19672 14381 19700
rect 14369 19669 14381 19672
rect 14415 19700 14427 19703
rect 14458 19700 14464 19712
rect 14415 19672 14464 19700
rect 14415 19669 14427 19672
rect 14369 19663 14427 19669
rect 14458 19660 14464 19672
rect 14516 19660 14522 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 3326 19496 3332 19508
rect 3287 19468 3332 19496
rect 3326 19456 3332 19468
rect 3384 19456 3390 19508
rect 6178 19496 6184 19508
rect 6139 19468 6184 19496
rect 6178 19456 6184 19468
rect 6236 19456 6242 19508
rect 7650 19496 7656 19508
rect 7611 19468 7656 19496
rect 7650 19456 7656 19468
rect 7708 19456 7714 19508
rect 10502 19456 10508 19508
rect 10560 19496 10566 19508
rect 10597 19499 10655 19505
rect 10597 19496 10609 19499
rect 10560 19468 10609 19496
rect 10560 19456 10566 19468
rect 10597 19465 10609 19468
rect 10643 19496 10655 19499
rect 12434 19496 12440 19508
rect 10643 19468 12440 19496
rect 10643 19465 10655 19468
rect 10597 19459 10655 19465
rect 12434 19456 12440 19468
rect 12492 19496 12498 19508
rect 12710 19496 12716 19508
rect 12492 19468 12716 19496
rect 12492 19456 12498 19468
rect 12710 19456 12716 19468
rect 12768 19456 12774 19508
rect 9125 19431 9183 19437
rect 9125 19397 9137 19431
rect 9171 19428 9183 19431
rect 11054 19428 11060 19440
rect 9171 19400 11060 19428
rect 9171 19397 9183 19400
rect 9125 19391 9183 19397
rect 4338 19360 4344 19372
rect 3988 19332 4344 19360
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 2409 19295 2467 19301
rect 1443 19264 2084 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 1578 19156 1584 19168
rect 1539 19128 1584 19156
rect 1578 19116 1584 19128
rect 1636 19116 1642 19168
rect 2056 19165 2084 19264
rect 2409 19261 2421 19295
rect 2455 19292 2467 19295
rect 2498 19292 2504 19304
rect 2455 19264 2504 19292
rect 2455 19261 2467 19264
rect 2409 19255 2467 19261
rect 2498 19252 2504 19264
rect 2556 19252 2562 19304
rect 3697 19295 3755 19301
rect 3697 19261 3709 19295
rect 3743 19292 3755 19295
rect 3988 19292 4016 19332
rect 4338 19320 4344 19332
rect 4396 19360 4402 19372
rect 4433 19363 4491 19369
rect 4433 19360 4445 19363
rect 4396 19332 4445 19360
rect 4396 19320 4402 19332
rect 4433 19329 4445 19332
rect 4479 19360 4491 19363
rect 5442 19360 5448 19372
rect 4479 19332 5448 19360
rect 4479 19329 4491 19332
rect 4433 19323 4491 19329
rect 5442 19320 5448 19332
rect 5500 19320 5506 19372
rect 7098 19360 7104 19372
rect 6840 19332 7104 19360
rect 4154 19292 4160 19304
rect 3743 19264 4016 19292
rect 4115 19264 4160 19292
rect 3743 19261 3755 19264
rect 3697 19255 3755 19261
rect 4154 19252 4160 19264
rect 4212 19252 4218 19304
rect 5166 19292 5172 19304
rect 5127 19264 5172 19292
rect 5166 19252 5172 19264
rect 5224 19252 5230 19304
rect 5258 19252 5264 19304
rect 5316 19292 5322 19304
rect 5353 19295 5411 19301
rect 5353 19292 5365 19295
rect 5316 19264 5365 19292
rect 5316 19252 5322 19264
rect 5353 19261 5365 19264
rect 5399 19261 5411 19295
rect 5353 19255 5411 19261
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19292 6699 19295
rect 6840 19292 6868 19332
rect 7098 19320 7104 19332
rect 7156 19360 7162 19372
rect 7282 19360 7288 19372
rect 7156 19332 7288 19360
rect 7156 19320 7162 19332
rect 7282 19320 7288 19332
rect 7340 19320 7346 19372
rect 7834 19320 7840 19372
rect 7892 19360 7898 19372
rect 8113 19363 8171 19369
rect 8113 19360 8125 19363
rect 7892 19332 8125 19360
rect 7892 19320 7898 19332
rect 8113 19329 8125 19332
rect 8159 19329 8171 19363
rect 8113 19323 8171 19329
rect 8297 19363 8355 19369
rect 8297 19329 8309 19363
rect 8343 19360 8355 19363
rect 8478 19360 8484 19372
rect 8343 19332 8484 19360
rect 8343 19329 8355 19332
rect 8297 19323 8355 19329
rect 8478 19320 8484 19332
rect 8536 19320 8542 19372
rect 9876 19369 9904 19400
rect 11054 19388 11060 19400
rect 11112 19388 11118 19440
rect 12621 19431 12679 19437
rect 12621 19397 12633 19431
rect 12667 19428 12679 19431
rect 13722 19428 13728 19440
rect 12667 19400 13728 19428
rect 12667 19397 12679 19400
rect 12621 19391 12679 19397
rect 13722 19388 13728 19400
rect 13780 19388 13786 19440
rect 9861 19363 9919 19369
rect 9861 19329 9873 19363
rect 9907 19329 9919 19363
rect 9861 19323 9919 19329
rect 11425 19363 11483 19369
rect 11425 19329 11437 19363
rect 11471 19360 11483 19363
rect 13170 19360 13176 19372
rect 11471 19332 11928 19360
rect 13131 19332 13176 19360
rect 11471 19329 11483 19332
rect 11425 19323 11483 19329
rect 6687 19264 6868 19292
rect 6687 19261 6699 19264
rect 6641 19255 6699 19261
rect 8938 19252 8944 19304
rect 8996 19292 9002 19304
rect 9585 19295 9643 19301
rect 9585 19292 9597 19295
rect 8996 19264 9597 19292
rect 8996 19252 9002 19264
rect 9585 19261 9597 19264
rect 9631 19261 9643 19295
rect 9585 19255 9643 19261
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 11149 19295 11207 19301
rect 11149 19292 11161 19295
rect 11112 19264 11161 19292
rect 11112 19252 11118 19264
rect 11149 19261 11161 19264
rect 11195 19261 11207 19295
rect 11149 19255 11207 19261
rect 11900 19233 11928 19332
rect 13170 19320 13176 19332
rect 13228 19320 13234 19372
rect 13906 19320 13912 19372
rect 13964 19320 13970 19372
rect 13081 19295 13139 19301
rect 13081 19261 13093 19295
rect 13127 19292 13139 19295
rect 13262 19292 13268 19304
rect 13127 19264 13268 19292
rect 13127 19261 13139 19264
rect 13081 19255 13139 19261
rect 13262 19252 13268 19264
rect 13320 19252 13326 19304
rect 11885 19227 11943 19233
rect 11885 19193 11897 19227
rect 11931 19224 11943 19227
rect 13630 19224 13636 19236
rect 11931 19196 13636 19224
rect 11931 19193 11943 19196
rect 11885 19187 11943 19193
rect 13630 19184 13636 19196
rect 13688 19184 13694 19236
rect 13725 19227 13783 19233
rect 13725 19193 13737 19227
rect 13771 19224 13783 19227
rect 13924 19224 13952 19320
rect 14182 19292 14188 19304
rect 14143 19264 14188 19292
rect 14182 19252 14188 19264
rect 14240 19252 14246 19304
rect 14458 19301 14464 19304
rect 14452 19292 14464 19301
rect 14419 19264 14464 19292
rect 14452 19255 14464 19264
rect 14458 19252 14464 19255
rect 14516 19252 14522 19304
rect 13771 19196 15608 19224
rect 13771 19193 13783 19196
rect 13725 19187 13783 19193
rect 2041 19159 2099 19165
rect 2041 19125 2053 19159
rect 2087 19156 2099 19159
rect 2685 19159 2743 19165
rect 2685 19156 2697 19159
rect 2087 19128 2697 19156
rect 2087 19125 2099 19128
rect 2041 19119 2099 19125
rect 2685 19125 2697 19128
rect 2731 19125 2743 19159
rect 2685 19119 2743 19125
rect 3694 19116 3700 19168
rect 3752 19156 3758 19168
rect 3789 19159 3847 19165
rect 3789 19156 3801 19159
rect 3752 19128 3801 19156
rect 3752 19116 3758 19128
rect 3789 19125 3801 19128
rect 3835 19125 3847 19159
rect 4246 19156 4252 19168
rect 4207 19128 4252 19156
rect 3789 19119 3847 19125
rect 4246 19116 4252 19128
rect 4304 19116 4310 19168
rect 4706 19116 4712 19168
rect 4764 19156 4770 19168
rect 4801 19159 4859 19165
rect 4801 19156 4813 19159
rect 4764 19128 4813 19156
rect 4764 19116 4770 19128
rect 4801 19125 4813 19128
rect 4847 19125 4859 19159
rect 4801 19119 4859 19125
rect 6638 19116 6644 19168
rect 6696 19156 6702 19168
rect 6914 19156 6920 19168
rect 6696 19128 6920 19156
rect 6696 19116 6702 19128
rect 6914 19116 6920 19128
rect 6972 19156 6978 19168
rect 7009 19159 7067 19165
rect 7009 19156 7021 19159
rect 6972 19128 7021 19156
rect 6972 19116 6978 19128
rect 7009 19125 7021 19128
rect 7055 19125 7067 19159
rect 7009 19119 7067 19125
rect 7561 19159 7619 19165
rect 7561 19125 7573 19159
rect 7607 19156 7619 19159
rect 7926 19156 7932 19168
rect 7607 19128 7932 19156
rect 7607 19125 7619 19128
rect 7561 19119 7619 19125
rect 7926 19116 7932 19128
rect 7984 19156 7990 19168
rect 8021 19159 8079 19165
rect 8021 19156 8033 19159
rect 7984 19128 8033 19156
rect 7984 19116 7990 19128
rect 8021 19125 8033 19128
rect 8067 19125 8079 19159
rect 8021 19119 8079 19125
rect 8478 19116 8484 19168
rect 8536 19156 8542 19168
rect 8665 19159 8723 19165
rect 8665 19156 8677 19159
rect 8536 19128 8677 19156
rect 8536 19116 8542 19128
rect 8665 19125 8677 19128
rect 8711 19125 8723 19159
rect 9214 19156 9220 19168
rect 9175 19128 9220 19156
rect 8665 19119 8723 19125
rect 9214 19116 9220 19128
rect 9272 19116 9278 19168
rect 9582 19116 9588 19168
rect 9640 19156 9646 19168
rect 9677 19159 9735 19165
rect 9677 19156 9689 19159
rect 9640 19128 9689 19156
rect 9640 19116 9646 19128
rect 9677 19125 9689 19128
rect 9723 19125 9735 19159
rect 10778 19156 10784 19168
rect 10739 19128 10784 19156
rect 9677 19119 9735 19125
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 11241 19159 11299 19165
rect 11241 19125 11253 19159
rect 11287 19156 11299 19159
rect 11790 19156 11796 19168
rect 11287 19128 11796 19156
rect 11287 19125 11299 19128
rect 11241 19119 11299 19125
rect 11790 19116 11796 19128
rect 11848 19116 11854 19168
rect 12253 19159 12311 19165
rect 12253 19125 12265 19159
rect 12299 19156 12311 19159
rect 12894 19156 12900 19168
rect 12299 19128 12900 19156
rect 12299 19125 12311 19128
rect 12253 19119 12311 19125
rect 12894 19116 12900 19128
rect 12952 19156 12958 19168
rect 12989 19159 13047 19165
rect 12989 19156 13001 19159
rect 12952 19128 13001 19156
rect 12952 19116 12958 19128
rect 12989 19125 13001 19128
rect 13035 19125 13047 19159
rect 12989 19119 13047 19125
rect 13262 19116 13268 19168
rect 13320 19156 13326 19168
rect 14001 19159 14059 19165
rect 14001 19156 14013 19159
rect 13320 19128 14013 19156
rect 13320 19116 13326 19128
rect 14001 19125 14013 19128
rect 14047 19156 14059 19159
rect 14182 19156 14188 19168
rect 14047 19128 14188 19156
rect 14047 19125 14059 19128
rect 14001 19119 14059 19125
rect 14182 19116 14188 19128
rect 14240 19116 14246 19168
rect 15580 19165 15608 19196
rect 15565 19159 15623 19165
rect 15565 19125 15577 19159
rect 15611 19125 15623 19159
rect 15565 19119 15623 19125
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1670 18912 1676 18964
rect 1728 18952 1734 18964
rect 1949 18955 2007 18961
rect 1949 18952 1961 18955
rect 1728 18924 1961 18952
rect 1728 18912 1734 18924
rect 1949 18921 1961 18924
rect 1995 18921 2007 18955
rect 2682 18952 2688 18964
rect 2643 18924 2688 18952
rect 1949 18915 2007 18921
rect 2682 18912 2688 18924
rect 2740 18912 2746 18964
rect 3145 18955 3203 18961
rect 3145 18921 3157 18955
rect 3191 18952 3203 18955
rect 3418 18952 3424 18964
rect 3191 18924 3424 18952
rect 3191 18921 3203 18924
rect 3145 18915 3203 18921
rect 3418 18912 3424 18924
rect 3476 18912 3482 18964
rect 3881 18955 3939 18961
rect 3881 18921 3893 18955
rect 3927 18952 3939 18955
rect 4246 18952 4252 18964
rect 3927 18924 4252 18952
rect 3927 18921 3939 18924
rect 3881 18915 3939 18921
rect 4246 18912 4252 18924
rect 4304 18952 4310 18964
rect 4525 18955 4583 18961
rect 4525 18952 4537 18955
rect 4304 18924 4537 18952
rect 4304 18912 4310 18924
rect 4525 18921 4537 18924
rect 4571 18921 4583 18955
rect 4525 18915 4583 18921
rect 4985 18955 5043 18961
rect 4985 18921 4997 18955
rect 5031 18952 5043 18955
rect 5166 18952 5172 18964
rect 5031 18924 5172 18952
rect 5031 18921 5043 18924
rect 4985 18915 5043 18921
rect 5166 18912 5172 18924
rect 5224 18952 5230 18964
rect 6089 18955 6147 18961
rect 6089 18952 6101 18955
rect 5224 18924 6101 18952
rect 5224 18912 5230 18924
rect 6089 18921 6101 18924
rect 6135 18921 6147 18955
rect 7466 18952 7472 18964
rect 7427 18924 7472 18952
rect 6089 18915 6147 18921
rect 7466 18912 7472 18924
rect 7524 18952 7530 18964
rect 8113 18955 8171 18961
rect 8113 18952 8125 18955
rect 7524 18924 8125 18952
rect 7524 18912 7530 18924
rect 8113 18921 8125 18924
rect 8159 18921 8171 18955
rect 8113 18915 8171 18921
rect 9309 18955 9367 18961
rect 9309 18921 9321 18955
rect 9355 18952 9367 18955
rect 9582 18952 9588 18964
rect 9355 18924 9588 18952
rect 9355 18921 9367 18924
rect 9309 18915 9367 18921
rect 9582 18912 9588 18924
rect 9640 18912 9646 18964
rect 11238 18952 11244 18964
rect 11199 18924 11244 18952
rect 11238 18912 11244 18924
rect 11296 18912 11302 18964
rect 11790 18952 11796 18964
rect 11703 18924 11796 18952
rect 11790 18912 11796 18924
rect 11848 18952 11854 18964
rect 12342 18952 12348 18964
rect 11848 18924 12348 18952
rect 11848 18912 11854 18924
rect 12342 18912 12348 18924
rect 12400 18912 12406 18964
rect 13722 18912 13728 18964
rect 13780 18952 13786 18964
rect 14645 18955 14703 18961
rect 14645 18952 14657 18955
rect 13780 18924 14657 18952
rect 13780 18912 13786 18924
rect 14645 18921 14657 18924
rect 14691 18921 14703 18955
rect 14645 18915 14703 18921
rect 3513 18887 3571 18893
rect 3513 18853 3525 18887
rect 3559 18884 3571 18887
rect 4154 18884 4160 18896
rect 3559 18856 4160 18884
rect 3559 18853 3571 18856
rect 3513 18847 3571 18853
rect 4154 18844 4160 18856
rect 4212 18844 4218 18896
rect 4338 18884 4344 18896
rect 4299 18856 4344 18884
rect 4338 18844 4344 18856
rect 4396 18844 4402 18896
rect 4893 18887 4951 18893
rect 4893 18853 4905 18887
rect 4939 18884 4951 18887
rect 5534 18884 5540 18896
rect 4939 18856 5540 18884
rect 4939 18853 4951 18856
rect 4893 18847 4951 18853
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18816 1455 18819
rect 2222 18816 2228 18828
rect 1443 18788 2228 18816
rect 1443 18785 1455 18788
rect 1397 18779 1455 18785
rect 2222 18776 2228 18788
rect 2280 18776 2286 18828
rect 2498 18816 2504 18828
rect 2459 18788 2504 18816
rect 2498 18776 2504 18788
rect 2556 18776 2562 18828
rect 4246 18776 4252 18828
rect 4304 18816 4310 18828
rect 4908 18816 4936 18847
rect 5534 18844 5540 18856
rect 5592 18844 5598 18896
rect 6457 18887 6515 18893
rect 6457 18853 6469 18887
rect 6503 18884 6515 18887
rect 6638 18884 6644 18896
rect 6503 18856 6644 18884
rect 6503 18853 6515 18856
rect 6457 18847 6515 18853
rect 6638 18844 6644 18856
rect 6696 18844 6702 18896
rect 10045 18887 10103 18893
rect 10045 18853 10057 18887
rect 10091 18884 10103 18887
rect 10134 18884 10140 18896
rect 10091 18856 10140 18884
rect 10091 18853 10103 18856
rect 10045 18847 10103 18853
rect 10134 18844 10140 18856
rect 10192 18844 10198 18896
rect 11054 18844 11060 18896
rect 11112 18884 11118 18896
rect 12986 18893 12992 18896
rect 12069 18887 12127 18893
rect 12069 18884 12081 18887
rect 11112 18856 12081 18884
rect 11112 18844 11118 18856
rect 12069 18853 12081 18856
rect 12115 18853 12127 18887
rect 12980 18884 12992 18893
rect 12899 18856 12992 18884
rect 12069 18847 12127 18853
rect 12980 18847 12992 18856
rect 13044 18884 13050 18896
rect 13630 18884 13636 18896
rect 13044 18856 13636 18884
rect 12986 18844 12992 18847
rect 13044 18844 13050 18856
rect 13630 18844 13636 18856
rect 13688 18844 13694 18896
rect 14090 18844 14096 18896
rect 14148 18884 14154 18896
rect 14550 18884 14556 18896
rect 14148 18856 14556 18884
rect 14148 18844 14154 18856
rect 14550 18844 14556 18856
rect 14608 18844 14614 18896
rect 4304 18788 4936 18816
rect 4304 18776 4310 18788
rect 6178 18776 6184 18828
rect 6236 18816 6242 18828
rect 8018 18816 8024 18828
rect 6236 18788 6684 18816
rect 7979 18788 8024 18816
rect 6236 18776 6242 18788
rect 4890 18708 4896 18760
rect 4948 18748 4954 18760
rect 6656 18757 6684 18788
rect 8018 18776 8024 18788
rect 8076 18776 8082 18828
rect 11146 18816 11152 18828
rect 11107 18788 11152 18816
rect 11146 18776 11152 18788
rect 11204 18776 11210 18828
rect 12710 18816 12716 18828
rect 12623 18788 12716 18816
rect 12710 18776 12716 18788
rect 12768 18816 12774 18828
rect 13262 18816 13268 18828
rect 12768 18788 13268 18816
rect 12768 18776 12774 18788
rect 13262 18776 13268 18788
rect 13320 18776 13326 18828
rect 5077 18751 5135 18757
rect 5077 18748 5089 18751
rect 4948 18720 5089 18748
rect 4948 18708 4954 18720
rect 5077 18717 5089 18720
rect 5123 18717 5135 18751
rect 5077 18711 5135 18717
rect 6549 18751 6607 18757
rect 6549 18717 6561 18751
rect 6595 18717 6607 18751
rect 6549 18711 6607 18717
rect 6641 18751 6699 18757
rect 6641 18717 6653 18751
rect 6687 18717 6699 18751
rect 6641 18711 6699 18717
rect 6564 18680 6592 18711
rect 8202 18708 8208 18760
rect 8260 18748 8266 18760
rect 10137 18751 10195 18757
rect 8260 18720 8305 18748
rect 8260 18708 8266 18720
rect 10137 18717 10149 18751
rect 10183 18717 10195 18751
rect 10318 18748 10324 18760
rect 10279 18720 10324 18748
rect 10137 18711 10195 18717
rect 6822 18680 6828 18692
rect 6564 18652 6828 18680
rect 6822 18640 6828 18652
rect 6880 18640 6886 18692
rect 10152 18680 10180 18711
rect 10318 18708 10324 18720
rect 10376 18708 10382 18760
rect 15286 18748 15292 18760
rect 15247 18720 15292 18748
rect 15286 18708 15292 18720
rect 15344 18708 15350 18760
rect 11330 18680 11336 18692
rect 10152 18652 11336 18680
rect 11330 18640 11336 18652
rect 11388 18640 11394 18692
rect 14093 18683 14151 18689
rect 14093 18649 14105 18683
rect 14139 18680 14151 18683
rect 14458 18680 14464 18692
rect 14139 18652 14464 18680
rect 14139 18649 14151 18652
rect 14093 18643 14151 18649
rect 14458 18640 14464 18652
rect 14516 18640 14522 18692
rect 1394 18572 1400 18624
rect 1452 18612 1458 18624
rect 1581 18615 1639 18621
rect 1581 18612 1593 18615
rect 1452 18584 1593 18612
rect 1452 18572 1458 18584
rect 1581 18581 1593 18584
rect 1627 18581 1639 18615
rect 1581 18575 1639 18581
rect 2409 18615 2467 18621
rect 2409 18581 2421 18615
rect 2455 18612 2467 18615
rect 2590 18612 2596 18624
rect 2455 18584 2596 18612
rect 2455 18581 2467 18584
rect 2409 18575 2467 18581
rect 2590 18572 2596 18584
rect 2648 18572 2654 18624
rect 7006 18572 7012 18624
rect 7064 18612 7070 18624
rect 7101 18615 7159 18621
rect 7101 18612 7113 18615
rect 7064 18584 7113 18612
rect 7064 18572 7070 18584
rect 7101 18581 7113 18584
rect 7147 18581 7159 18615
rect 7650 18612 7656 18624
rect 7611 18584 7656 18612
rect 7101 18575 7159 18581
rect 7650 18572 7656 18584
rect 7708 18572 7714 18624
rect 9677 18615 9735 18621
rect 9677 18581 9689 18615
rect 9723 18612 9735 18615
rect 9858 18612 9864 18624
rect 9723 18584 9864 18612
rect 9723 18581 9735 18584
rect 9677 18575 9735 18581
rect 9858 18572 9864 18584
rect 9916 18572 9922 18624
rect 10686 18612 10692 18624
rect 10647 18584 10692 18612
rect 10686 18572 10692 18584
rect 10744 18572 10750 18624
rect 12529 18615 12587 18621
rect 12529 18581 12541 18615
rect 12575 18612 12587 18615
rect 12710 18612 12716 18624
rect 12575 18584 12716 18612
rect 12575 18581 12587 18584
rect 12529 18575 12587 18581
rect 12710 18572 12716 18584
rect 12768 18572 12774 18624
rect 13814 18572 13820 18624
rect 13872 18612 13878 18624
rect 17586 18612 17592 18624
rect 13872 18584 17592 18612
rect 13872 18572 13878 18584
rect 17586 18572 17592 18584
rect 17644 18572 17650 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 2498 18408 2504 18420
rect 2459 18380 2504 18408
rect 2498 18368 2504 18380
rect 2556 18368 2562 18420
rect 3789 18411 3847 18417
rect 3789 18377 3801 18411
rect 3835 18408 3847 18411
rect 4890 18408 4896 18420
rect 3835 18380 4896 18408
rect 3835 18377 3847 18380
rect 3789 18371 3847 18377
rect 4890 18368 4896 18380
rect 4948 18368 4954 18420
rect 8478 18408 8484 18420
rect 8439 18380 8484 18408
rect 8478 18368 8484 18380
rect 8536 18368 8542 18420
rect 10042 18368 10048 18420
rect 10100 18408 10106 18420
rect 10318 18408 10324 18420
rect 10100 18380 10324 18408
rect 10100 18368 10106 18380
rect 10318 18368 10324 18380
rect 10376 18408 10382 18420
rect 10965 18411 11023 18417
rect 10965 18408 10977 18411
rect 10376 18380 10977 18408
rect 10376 18368 10382 18380
rect 10965 18377 10977 18380
rect 11011 18377 11023 18411
rect 13998 18408 14004 18420
rect 13959 18380 14004 18408
rect 10965 18371 11023 18377
rect 13998 18368 14004 18380
rect 14056 18368 14062 18420
rect 9401 18343 9459 18349
rect 9401 18309 9413 18343
rect 9447 18340 9459 18343
rect 9766 18340 9772 18352
rect 9447 18312 9772 18340
rect 9447 18309 9459 18312
rect 9401 18303 9459 18309
rect 9766 18300 9772 18312
rect 9824 18340 9830 18352
rect 9861 18343 9919 18349
rect 9861 18340 9873 18343
rect 9824 18312 9873 18340
rect 9824 18300 9830 18312
rect 9861 18309 9873 18312
rect 9907 18309 9919 18343
rect 9861 18303 9919 18309
rect 10594 18300 10600 18352
rect 10652 18340 10658 18352
rect 13817 18343 13875 18349
rect 13817 18340 13829 18343
rect 10652 18312 13829 18340
rect 10652 18300 10658 18312
rect 13817 18309 13829 18312
rect 13863 18309 13875 18343
rect 13817 18303 13875 18309
rect 2225 18275 2283 18281
rect 2225 18241 2237 18275
rect 2271 18272 2283 18275
rect 3145 18275 3203 18281
rect 3145 18272 3157 18275
rect 2271 18244 3157 18272
rect 2271 18241 2283 18244
rect 2225 18235 2283 18241
rect 3145 18241 3157 18244
rect 3191 18272 3203 18275
rect 3234 18272 3240 18284
rect 3191 18244 3240 18272
rect 3191 18241 3203 18244
rect 3145 18235 3203 18241
rect 3234 18232 3240 18244
rect 3292 18232 3298 18284
rect 3329 18275 3387 18281
rect 3329 18241 3341 18275
rect 3375 18272 3387 18275
rect 3510 18272 3516 18284
rect 3375 18244 3516 18272
rect 3375 18241 3387 18244
rect 3329 18235 3387 18241
rect 3510 18232 3516 18244
rect 3568 18232 3574 18284
rect 9674 18232 9680 18284
rect 9732 18272 9738 18284
rect 10505 18275 10563 18281
rect 10505 18272 10517 18275
rect 9732 18244 10517 18272
rect 9732 18232 9738 18244
rect 10505 18241 10517 18244
rect 10551 18272 10563 18275
rect 10686 18272 10692 18284
rect 10551 18244 10692 18272
rect 10551 18241 10563 18244
rect 10505 18235 10563 18241
rect 10686 18232 10692 18244
rect 10744 18232 10750 18284
rect 12250 18272 12256 18284
rect 12163 18244 12256 18272
rect 12250 18232 12256 18244
rect 12308 18272 12314 18284
rect 12897 18275 12955 18281
rect 12897 18272 12909 18275
rect 12308 18244 12909 18272
rect 12308 18232 12314 18244
rect 12897 18241 12909 18244
rect 12943 18241 12955 18275
rect 12897 18235 12955 18241
rect 12989 18275 13047 18281
rect 12989 18241 13001 18275
rect 13035 18241 13047 18275
rect 12989 18235 13047 18241
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18204 1455 18207
rect 1670 18204 1676 18216
rect 1443 18176 1676 18204
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 1670 18164 1676 18176
rect 1728 18164 1734 18216
rect 3053 18207 3111 18213
rect 3053 18173 3065 18207
rect 3099 18204 3111 18207
rect 3418 18204 3424 18216
rect 3099 18176 3424 18204
rect 3099 18173 3111 18176
rect 3053 18167 3111 18173
rect 3418 18164 3424 18176
rect 3476 18164 3482 18216
rect 4249 18207 4307 18213
rect 4249 18204 4261 18207
rect 4172 18176 4261 18204
rect 4172 18136 4200 18176
rect 4249 18173 4261 18176
rect 4295 18173 4307 18207
rect 4249 18167 4307 18173
rect 4338 18164 4344 18216
rect 4396 18204 4402 18216
rect 4505 18207 4563 18213
rect 4505 18204 4517 18207
rect 4396 18176 4517 18204
rect 4396 18164 4402 18176
rect 4505 18173 4517 18176
rect 4551 18173 4563 18207
rect 4505 18167 4563 18173
rect 7006 18164 7012 18216
rect 7064 18204 7070 18216
rect 7101 18207 7159 18213
rect 7101 18204 7113 18207
rect 7064 18176 7113 18204
rect 7064 18164 7070 18176
rect 7101 18173 7113 18176
rect 7147 18173 7159 18207
rect 7101 18167 7159 18173
rect 9861 18207 9919 18213
rect 9861 18173 9873 18207
rect 9907 18204 9919 18207
rect 10321 18207 10379 18213
rect 10321 18204 10333 18207
rect 9907 18176 10333 18204
rect 9907 18173 9919 18176
rect 9861 18167 9919 18173
rect 10321 18173 10333 18176
rect 10367 18204 10379 18207
rect 11238 18204 11244 18216
rect 10367 18176 11244 18204
rect 10367 18173 10379 18176
rect 10321 18167 10379 18173
rect 11238 18164 11244 18176
rect 11296 18164 11302 18216
rect 11885 18207 11943 18213
rect 11885 18173 11897 18207
rect 11931 18204 11943 18207
rect 13004 18204 13032 18235
rect 13722 18204 13728 18216
rect 11931 18176 13728 18204
rect 11931 18173 11943 18176
rect 11885 18167 11943 18173
rect 13722 18164 13728 18176
rect 13780 18164 13786 18216
rect 4706 18136 4712 18148
rect 4172 18108 4712 18136
rect 4172 18080 4200 18108
rect 4706 18096 4712 18108
rect 4764 18096 4770 18148
rect 6273 18139 6331 18145
rect 6273 18105 6285 18139
rect 6319 18136 6331 18139
rect 6638 18136 6644 18148
rect 6319 18108 6644 18136
rect 6319 18105 6331 18108
rect 6273 18099 6331 18105
rect 6638 18096 6644 18108
rect 6696 18096 6702 18148
rect 7374 18145 7380 18148
rect 7368 18136 7380 18145
rect 7335 18108 7380 18136
rect 7368 18099 7380 18108
rect 7374 18096 7380 18099
rect 7432 18096 7438 18148
rect 9769 18139 9827 18145
rect 9769 18105 9781 18139
rect 9815 18136 9827 18139
rect 10134 18136 10140 18148
rect 9815 18108 10140 18136
rect 9815 18105 9827 18108
rect 9769 18099 9827 18105
rect 10134 18096 10140 18108
rect 10192 18136 10198 18148
rect 10962 18136 10968 18148
rect 10192 18108 10968 18136
rect 10192 18096 10198 18108
rect 10962 18096 10968 18108
rect 11020 18096 11026 18148
rect 1486 18028 1492 18080
rect 1544 18068 1550 18080
rect 1581 18071 1639 18077
rect 1581 18068 1593 18071
rect 1544 18040 1593 18068
rect 1544 18028 1550 18040
rect 1581 18037 1593 18040
rect 1627 18037 1639 18071
rect 1581 18031 1639 18037
rect 2498 18028 2504 18080
rect 2556 18068 2562 18080
rect 2685 18071 2743 18077
rect 2685 18068 2697 18071
rect 2556 18040 2697 18068
rect 2556 18028 2562 18040
rect 2685 18037 2697 18040
rect 2731 18037 2743 18071
rect 4154 18068 4160 18080
rect 4115 18040 4160 18068
rect 2685 18031 2743 18037
rect 4154 18028 4160 18040
rect 4212 18028 4218 18080
rect 4982 18028 4988 18080
rect 5040 18068 5046 18080
rect 5629 18071 5687 18077
rect 5629 18068 5641 18071
rect 5040 18040 5641 18068
rect 5040 18028 5046 18040
rect 5629 18037 5641 18040
rect 5675 18037 5687 18071
rect 5629 18031 5687 18037
rect 6549 18071 6607 18077
rect 6549 18037 6561 18071
rect 6595 18068 6607 18071
rect 6822 18068 6828 18080
rect 6595 18040 6828 18068
rect 6595 18037 6607 18040
rect 6549 18031 6607 18037
rect 6822 18028 6828 18040
rect 6880 18028 6886 18080
rect 9950 18068 9956 18080
rect 9911 18040 9956 18068
rect 9950 18028 9956 18040
rect 10008 18028 10014 18080
rect 10413 18071 10471 18077
rect 10413 18037 10425 18071
rect 10459 18068 10471 18071
rect 10870 18068 10876 18080
rect 10459 18040 10876 18068
rect 10459 18037 10471 18040
rect 10413 18031 10471 18037
rect 10870 18028 10876 18040
rect 10928 18028 10934 18080
rect 11330 18068 11336 18080
rect 11291 18040 11336 18068
rect 11330 18028 11336 18040
rect 11388 18028 11394 18080
rect 11606 18028 11612 18080
rect 11664 18068 11670 18080
rect 12437 18071 12495 18077
rect 12437 18068 12449 18071
rect 11664 18040 12449 18068
rect 11664 18028 11670 18040
rect 12437 18037 12449 18040
rect 12483 18037 12495 18071
rect 12802 18068 12808 18080
rect 12763 18040 12808 18068
rect 12437 18031 12495 18037
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 13262 18028 13268 18080
rect 13320 18068 13326 18080
rect 13449 18071 13507 18077
rect 13449 18068 13461 18071
rect 13320 18040 13461 18068
rect 13320 18028 13326 18040
rect 13449 18037 13461 18040
rect 13495 18037 13507 18071
rect 13832 18068 13860 18303
rect 14458 18300 14464 18352
rect 14516 18340 14522 18352
rect 15013 18343 15071 18349
rect 15013 18340 15025 18343
rect 14516 18312 15025 18340
rect 14516 18300 14522 18312
rect 14568 18281 14596 18312
rect 15013 18309 15025 18312
rect 15059 18309 15071 18343
rect 15013 18303 15071 18309
rect 14553 18275 14611 18281
rect 14553 18241 14565 18275
rect 14599 18241 14611 18275
rect 14553 18235 14611 18241
rect 14369 18207 14427 18213
rect 14369 18173 14381 18207
rect 14415 18204 14427 18207
rect 14458 18204 14464 18216
rect 14415 18176 14464 18204
rect 14415 18173 14427 18176
rect 14369 18167 14427 18173
rect 14458 18164 14464 18176
rect 14516 18204 14522 18216
rect 15286 18204 15292 18216
rect 14516 18176 15292 18204
rect 14516 18164 14522 18176
rect 15286 18164 15292 18176
rect 15344 18164 15350 18216
rect 14461 18071 14519 18077
rect 14461 18068 14473 18071
rect 13832 18040 14473 18068
rect 13449 18031 13507 18037
rect 14461 18037 14473 18040
rect 14507 18037 14519 18071
rect 14461 18031 14519 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2038 17824 2044 17876
rect 2096 17864 2102 17876
rect 2777 17867 2835 17873
rect 2777 17864 2789 17867
rect 2096 17836 2789 17864
rect 2096 17824 2102 17836
rect 2777 17833 2789 17836
rect 2823 17864 2835 17867
rect 4065 17867 4123 17873
rect 4065 17864 4077 17867
rect 2823 17836 4077 17864
rect 2823 17833 2835 17836
rect 2777 17827 2835 17833
rect 4065 17833 4077 17836
rect 4111 17833 4123 17867
rect 4522 17864 4528 17876
rect 4483 17836 4528 17864
rect 4065 17827 4123 17833
rect 4522 17824 4528 17836
rect 4580 17824 4586 17876
rect 5166 17864 5172 17876
rect 5127 17836 5172 17864
rect 5166 17824 5172 17836
rect 5224 17824 5230 17876
rect 6178 17864 6184 17876
rect 6139 17836 6184 17864
rect 6178 17824 6184 17836
rect 6236 17824 6242 17876
rect 10686 17824 10692 17876
rect 10744 17864 10750 17876
rect 12345 17867 12403 17873
rect 12345 17864 12357 17867
rect 10744 17836 12357 17864
rect 10744 17824 10750 17836
rect 12345 17833 12357 17836
rect 12391 17833 12403 17867
rect 12986 17864 12992 17876
rect 12947 17836 12992 17864
rect 12345 17827 12403 17833
rect 12986 17824 12992 17836
rect 13044 17824 13050 17876
rect 13446 17824 13452 17876
rect 13504 17864 13510 17876
rect 13630 17864 13636 17876
rect 13504 17836 13636 17864
rect 13504 17824 13510 17836
rect 13630 17824 13636 17836
rect 13688 17864 13694 17876
rect 13909 17867 13967 17873
rect 13909 17864 13921 17867
rect 13688 17836 13921 17864
rect 13688 17824 13694 17836
rect 13909 17833 13921 17836
rect 13955 17833 13967 17867
rect 14458 17864 14464 17876
rect 14419 17836 14464 17864
rect 13909 17827 13967 17833
rect 14458 17824 14464 17836
rect 14516 17824 14522 17876
rect 2222 17796 2228 17808
rect 2183 17768 2228 17796
rect 2222 17756 2228 17768
rect 2280 17756 2286 17808
rect 3881 17799 3939 17805
rect 3881 17765 3893 17799
rect 3927 17796 3939 17799
rect 4246 17796 4252 17808
rect 3927 17768 4252 17796
rect 3927 17765 3939 17768
rect 3881 17759 3939 17765
rect 4246 17756 4252 17768
rect 4304 17756 4310 17808
rect 5629 17799 5687 17805
rect 5629 17765 5641 17799
rect 5675 17796 5687 17799
rect 8018 17796 8024 17808
rect 5675 17768 8024 17796
rect 5675 17765 5687 17768
rect 5629 17759 5687 17765
rect 8018 17756 8024 17768
rect 8076 17756 8082 17808
rect 11232 17799 11290 17805
rect 11232 17765 11244 17799
rect 11278 17796 11290 17799
rect 11422 17796 11428 17808
rect 11278 17768 11428 17796
rect 11278 17765 11290 17768
rect 11232 17759 11290 17765
rect 11422 17756 11428 17768
rect 11480 17756 11486 17808
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 4433 17731 4491 17737
rect 4433 17728 4445 17731
rect 1443 17700 4445 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 4433 17697 4445 17700
rect 4479 17728 4491 17731
rect 5258 17728 5264 17740
rect 4479 17700 5264 17728
rect 4479 17697 4491 17700
rect 4433 17691 4491 17697
rect 5258 17688 5264 17700
rect 5316 17688 5322 17740
rect 6908 17731 6966 17737
rect 6908 17697 6920 17731
rect 6954 17728 6966 17731
rect 8202 17728 8208 17740
rect 6954 17700 8208 17728
rect 6954 17697 6966 17700
rect 6908 17691 6966 17697
rect 8202 17688 8208 17700
rect 8260 17688 8266 17740
rect 9953 17731 10011 17737
rect 9953 17697 9965 17731
rect 9999 17728 10011 17731
rect 10778 17728 10784 17740
rect 9999 17700 10784 17728
rect 9999 17697 10011 17700
rect 9953 17691 10011 17697
rect 10778 17688 10784 17700
rect 10836 17688 10842 17740
rect 13354 17688 13360 17740
rect 13412 17728 13418 17740
rect 13814 17728 13820 17740
rect 13412 17700 13820 17728
rect 13412 17688 13418 17700
rect 13814 17688 13820 17700
rect 13872 17688 13878 17740
rect 2498 17620 2504 17672
rect 2556 17660 2562 17672
rect 2869 17663 2927 17669
rect 2869 17660 2881 17663
rect 2556 17632 2881 17660
rect 2556 17620 2562 17632
rect 2869 17629 2881 17632
rect 2915 17629 2927 17663
rect 3050 17660 3056 17672
rect 3011 17632 3056 17660
rect 2869 17623 2927 17629
rect 3050 17620 3056 17632
rect 3108 17620 3114 17672
rect 3510 17660 3516 17672
rect 3423 17632 3516 17660
rect 3510 17620 3516 17632
rect 3568 17660 3574 17672
rect 4709 17663 4767 17669
rect 4709 17660 4721 17663
rect 3568 17632 4721 17660
rect 3568 17620 3574 17632
rect 4709 17629 4721 17632
rect 4755 17660 4767 17663
rect 4982 17660 4988 17672
rect 4755 17632 4988 17660
rect 4755 17629 4767 17632
rect 4709 17623 4767 17629
rect 4982 17620 4988 17632
rect 5040 17620 5046 17672
rect 6362 17620 6368 17672
rect 6420 17660 6426 17672
rect 6641 17663 6699 17669
rect 6641 17660 6653 17663
rect 6420 17632 6653 17660
rect 6420 17620 6426 17632
rect 6641 17629 6653 17632
rect 6687 17629 6699 17663
rect 6641 17623 6699 17629
rect 2774 17552 2780 17604
rect 2832 17592 2838 17604
rect 3528 17592 3556 17620
rect 2832 17564 3556 17592
rect 2832 17552 2838 17564
rect 1946 17524 1952 17536
rect 1907 17496 1952 17524
rect 1946 17484 1952 17496
rect 2004 17484 2010 17536
rect 2409 17527 2467 17533
rect 2409 17493 2421 17527
rect 2455 17524 2467 17527
rect 2682 17524 2688 17536
rect 2455 17496 2688 17524
rect 2455 17493 2467 17496
rect 2409 17487 2467 17493
rect 2682 17484 2688 17496
rect 2740 17484 2746 17536
rect 5534 17524 5540 17536
rect 5495 17496 5540 17524
rect 5534 17484 5540 17496
rect 5592 17484 5598 17536
rect 6454 17524 6460 17536
rect 6415 17496 6460 17524
rect 6454 17484 6460 17496
rect 6512 17484 6518 17536
rect 6656 17524 6684 17623
rect 9398 17620 9404 17672
rect 9456 17660 9462 17672
rect 10965 17663 11023 17669
rect 10965 17660 10977 17663
rect 9456 17632 10977 17660
rect 9456 17620 9462 17632
rect 10965 17629 10977 17632
rect 11011 17629 11023 17663
rect 10965 17623 11023 17629
rect 10134 17592 10140 17604
rect 10095 17564 10140 17592
rect 10134 17552 10140 17564
rect 10192 17552 10198 17604
rect 7006 17524 7012 17536
rect 6656 17496 7012 17524
rect 7006 17484 7012 17496
rect 7064 17484 7070 17536
rect 7374 17484 7380 17536
rect 7432 17524 7438 17536
rect 8021 17527 8079 17533
rect 8021 17524 8033 17527
rect 7432 17496 8033 17524
rect 7432 17484 7438 17496
rect 8021 17493 8033 17496
rect 8067 17493 8079 17527
rect 8021 17487 8079 17493
rect 8202 17484 8208 17536
rect 8260 17524 8266 17536
rect 8665 17527 8723 17533
rect 8665 17524 8677 17527
rect 8260 17496 8677 17524
rect 8260 17484 8266 17496
rect 8665 17493 8677 17496
rect 8711 17524 8723 17527
rect 8754 17524 8760 17536
rect 8711 17496 8760 17524
rect 8711 17493 8723 17496
rect 8665 17487 8723 17493
rect 8754 17484 8760 17496
rect 8812 17484 8818 17536
rect 10505 17527 10563 17533
rect 10505 17493 10517 17527
rect 10551 17524 10563 17527
rect 10686 17524 10692 17536
rect 10551 17496 10692 17524
rect 10551 17493 10563 17496
rect 10505 17487 10563 17493
rect 10686 17484 10692 17496
rect 10744 17524 10750 17536
rect 10870 17524 10876 17536
rect 10744 17496 10876 17524
rect 10744 17484 10750 17496
rect 10870 17484 10876 17496
rect 10928 17484 10934 17536
rect 10980 17524 11008 17623
rect 13998 17620 14004 17672
rect 14056 17660 14062 17672
rect 14056 17632 14101 17660
rect 14056 17620 14062 17632
rect 11238 17524 11244 17536
rect 10980 17496 11244 17524
rect 11238 17484 11244 17496
rect 11296 17484 11302 17536
rect 13262 17524 13268 17536
rect 13223 17496 13268 17524
rect 13262 17484 13268 17496
rect 13320 17484 13326 17536
rect 13446 17524 13452 17536
rect 13407 17496 13452 17524
rect 13446 17484 13452 17496
rect 13504 17484 13510 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 2682 17280 2688 17332
rect 2740 17280 2746 17332
rect 4522 17280 4528 17332
rect 4580 17320 4586 17332
rect 4893 17323 4951 17329
rect 4893 17320 4905 17323
rect 4580 17292 4905 17320
rect 4580 17280 4586 17292
rect 4893 17289 4905 17292
rect 4939 17289 4951 17323
rect 5258 17320 5264 17332
rect 5219 17292 5264 17320
rect 4893 17283 4951 17289
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 6273 17323 6331 17329
rect 6273 17289 6285 17323
rect 6319 17320 6331 17323
rect 6454 17320 6460 17332
rect 6319 17292 6460 17320
rect 6319 17289 6331 17292
rect 6273 17283 6331 17289
rect 6454 17280 6460 17292
rect 6512 17280 6518 17332
rect 7929 17323 7987 17329
rect 7929 17289 7941 17323
rect 7975 17320 7987 17323
rect 8018 17320 8024 17332
rect 7975 17292 8024 17320
rect 7975 17289 7987 17292
rect 7929 17283 7987 17289
rect 8018 17280 8024 17292
rect 8076 17280 8082 17332
rect 11238 17280 11244 17332
rect 11296 17320 11302 17332
rect 11333 17323 11391 17329
rect 11333 17320 11345 17323
rect 11296 17292 11345 17320
rect 11296 17280 11302 17292
rect 11333 17289 11345 17292
rect 11379 17289 11391 17323
rect 11333 17283 11391 17289
rect 13906 17280 13912 17332
rect 13964 17320 13970 17332
rect 14645 17323 14703 17329
rect 14645 17320 14657 17323
rect 13964 17292 14657 17320
rect 13964 17280 13970 17292
rect 14645 17289 14657 17292
rect 14691 17289 14703 17323
rect 14645 17283 14703 17289
rect 2314 17212 2320 17264
rect 2372 17252 2378 17264
rect 2700 17252 2728 17280
rect 2372 17224 2728 17252
rect 2372 17212 2378 17224
rect 6472 17184 6500 17280
rect 7374 17184 7380 17196
rect 6472 17156 7380 17184
rect 7374 17144 7380 17156
rect 7432 17144 7438 17196
rect 8849 17187 8907 17193
rect 8849 17184 8861 17187
rect 7668 17156 8861 17184
rect 7668 17128 7696 17156
rect 8849 17153 8861 17156
rect 8895 17153 8907 17187
rect 8849 17147 8907 17153
rect 9125 17187 9183 17193
rect 9125 17153 9137 17187
rect 9171 17184 9183 17187
rect 9398 17184 9404 17196
rect 9171 17156 9404 17184
rect 9171 17153 9183 17156
rect 9125 17147 9183 17153
rect 9398 17144 9404 17156
rect 9456 17144 9462 17196
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 1946 17116 1952 17128
rect 1443 17088 1952 17116
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 1946 17076 1952 17088
rect 2004 17076 2010 17128
rect 2869 17119 2927 17125
rect 2869 17085 2881 17119
rect 2915 17116 2927 17119
rect 2958 17116 2964 17128
rect 2915 17088 2964 17116
rect 2915 17085 2927 17088
rect 2869 17079 2927 17085
rect 2958 17076 2964 17088
rect 3016 17076 3022 17128
rect 3228 17119 3286 17125
rect 3228 17085 3240 17119
rect 3274 17116 3286 17119
rect 3510 17116 3516 17128
rect 3274 17088 3516 17116
rect 3274 17085 3286 17088
rect 3228 17079 3286 17085
rect 3510 17076 3516 17088
rect 3568 17076 3574 17128
rect 5445 17119 5503 17125
rect 5445 17085 5457 17119
rect 5491 17116 5503 17119
rect 5718 17116 5724 17128
rect 5491 17088 5724 17116
rect 5491 17085 5503 17088
rect 5445 17079 5503 17085
rect 5718 17076 5724 17088
rect 5776 17076 5782 17128
rect 7193 17119 7251 17125
rect 7193 17085 7205 17119
rect 7239 17116 7251 17119
rect 7650 17116 7656 17128
rect 7239 17088 7656 17116
rect 7239 17085 7251 17088
rect 7193 17079 7251 17085
rect 7650 17076 7656 17088
rect 7708 17076 7714 17128
rect 8389 17119 8447 17125
rect 8389 17085 8401 17119
rect 8435 17116 8447 17119
rect 8662 17116 8668 17128
rect 8435 17088 8668 17116
rect 8435 17085 8447 17088
rect 8389 17079 8447 17085
rect 8662 17076 8668 17088
rect 8720 17116 8726 17128
rect 9214 17116 9220 17128
rect 8720 17088 9220 17116
rect 8720 17076 8726 17088
rect 9214 17076 9220 17088
rect 9272 17076 9278 17128
rect 13262 17116 13268 17128
rect 13223 17088 13268 17116
rect 13262 17076 13268 17088
rect 13320 17076 13326 17128
rect 2501 17051 2559 17057
rect 2501 17017 2513 17051
rect 2547 17048 2559 17051
rect 2774 17048 2780 17060
rect 2547 17020 2780 17048
rect 2547 17017 2559 17020
rect 2501 17011 2559 17017
rect 2774 17008 2780 17020
rect 2832 17008 2838 17060
rect 2976 17048 3004 17076
rect 4062 17048 4068 17060
rect 2976 17020 4068 17048
rect 4062 17008 4068 17020
rect 4120 17008 4126 17060
rect 5534 17008 5540 17060
rect 5592 17048 5598 17060
rect 8297 17051 8355 17057
rect 5592 17020 6868 17048
rect 5592 17008 5598 17020
rect 1578 16980 1584 16992
rect 1539 16952 1584 16980
rect 1578 16940 1584 16952
rect 1636 16940 1642 16992
rect 2133 16983 2191 16989
rect 2133 16949 2145 16983
rect 2179 16980 2191 16983
rect 2406 16980 2412 16992
rect 2179 16952 2412 16980
rect 2179 16949 2191 16952
rect 2133 16943 2191 16949
rect 2406 16940 2412 16952
rect 2464 16980 2470 16992
rect 3050 16980 3056 16992
rect 2464 16952 3056 16980
rect 2464 16940 2470 16952
rect 3050 16940 3056 16952
rect 3108 16980 3114 16992
rect 4341 16983 4399 16989
rect 4341 16980 4353 16983
rect 3108 16952 4353 16980
rect 3108 16940 3114 16952
rect 4341 16949 4353 16952
rect 4387 16980 4399 16983
rect 4798 16980 4804 16992
rect 4387 16952 4804 16980
rect 4387 16949 4399 16952
rect 4341 16943 4399 16949
rect 4798 16940 4804 16952
rect 4856 16940 4862 16992
rect 5626 16980 5632 16992
rect 5587 16952 5632 16980
rect 5626 16940 5632 16952
rect 5684 16940 5690 16992
rect 6362 16940 6368 16992
rect 6420 16980 6426 16992
rect 6840 16989 6868 17020
rect 8297 17017 8309 17051
rect 8343 17048 8355 17051
rect 8754 17048 8760 17060
rect 8343 17020 8760 17048
rect 8343 17017 8355 17020
rect 8297 17011 8355 17017
rect 8754 17008 8760 17020
rect 8812 17048 8818 17060
rect 8812 17020 9352 17048
rect 8812 17008 8818 17020
rect 6549 16983 6607 16989
rect 6549 16980 6561 16983
rect 6420 16952 6561 16980
rect 6420 16940 6426 16952
rect 6549 16949 6561 16952
rect 6595 16949 6607 16983
rect 6549 16943 6607 16949
rect 6825 16983 6883 16989
rect 6825 16949 6837 16983
rect 6871 16949 6883 16983
rect 6825 16943 6883 16949
rect 7282 16940 7288 16992
rect 7340 16980 7346 16992
rect 8570 16980 8576 16992
rect 7340 16952 7385 16980
rect 8531 16952 8576 16980
rect 7340 16940 7346 16952
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 9125 16983 9183 16989
rect 9125 16949 9137 16983
rect 9171 16980 9183 16983
rect 9214 16980 9220 16992
rect 9171 16952 9220 16980
rect 9171 16949 9183 16952
rect 9125 16943 9183 16949
rect 9214 16940 9220 16952
rect 9272 16940 9278 16992
rect 9324 16980 9352 17020
rect 9582 17008 9588 17060
rect 9640 17057 9646 17060
rect 9640 17051 9704 17057
rect 9640 17017 9658 17051
rect 9692 17017 9704 17051
rect 9640 17011 9704 17017
rect 12805 17051 12863 17057
rect 12805 17017 12817 17051
rect 12851 17048 12863 17051
rect 13532 17051 13590 17057
rect 13532 17048 13544 17051
rect 12851 17020 13544 17048
rect 12851 17017 12863 17020
rect 12805 17011 12863 17017
rect 13532 17017 13544 17020
rect 13578 17048 13590 17051
rect 13998 17048 14004 17060
rect 13578 17020 14004 17048
rect 13578 17017 13590 17020
rect 13532 17011 13590 17017
rect 9640 17008 9646 17011
rect 13998 17008 14004 17020
rect 14056 17008 14062 17060
rect 10134 16980 10140 16992
rect 9324 16952 10140 16980
rect 10134 16940 10140 16952
rect 10192 16980 10198 16992
rect 10781 16983 10839 16989
rect 10781 16980 10793 16983
rect 10192 16952 10793 16980
rect 10192 16940 10198 16952
rect 10781 16949 10793 16952
rect 10827 16949 10839 16983
rect 10781 16943 10839 16949
rect 11422 16940 11428 16992
rect 11480 16980 11486 16992
rect 11701 16983 11759 16989
rect 11701 16980 11713 16983
rect 11480 16952 11713 16980
rect 11480 16940 11486 16952
rect 11701 16949 11713 16952
rect 11747 16949 11759 16983
rect 11701 16943 11759 16949
rect 12066 16940 12072 16992
rect 12124 16980 12130 16992
rect 13081 16983 13139 16989
rect 13081 16980 13093 16983
rect 12124 16952 13093 16980
rect 12124 16940 12130 16952
rect 13081 16949 13093 16952
rect 13127 16980 13139 16983
rect 13354 16980 13360 16992
rect 13127 16952 13360 16980
rect 13127 16949 13139 16952
rect 13081 16943 13139 16949
rect 13354 16940 13360 16952
rect 13412 16940 13418 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1394 16736 1400 16788
rect 1452 16776 1458 16788
rect 1581 16779 1639 16785
rect 1581 16776 1593 16779
rect 1452 16748 1593 16776
rect 1452 16736 1458 16748
rect 1581 16745 1593 16748
rect 1627 16745 1639 16779
rect 2038 16776 2044 16788
rect 1999 16748 2044 16776
rect 1581 16739 1639 16745
rect 2038 16736 2044 16748
rect 2096 16736 2102 16788
rect 2409 16779 2467 16785
rect 2409 16745 2421 16779
rect 2455 16776 2467 16779
rect 2498 16776 2504 16788
rect 2455 16748 2504 16776
rect 2455 16745 2467 16748
rect 2409 16739 2467 16745
rect 2498 16736 2504 16748
rect 2556 16736 2562 16788
rect 2682 16776 2688 16788
rect 2643 16748 2688 16776
rect 2682 16736 2688 16748
rect 2740 16736 2746 16788
rect 3142 16776 3148 16788
rect 3103 16748 3148 16776
rect 3142 16736 3148 16748
rect 3200 16736 3206 16788
rect 3970 16736 3976 16788
rect 4028 16776 4034 16788
rect 4433 16779 4491 16785
rect 4433 16776 4445 16779
rect 4028 16748 4445 16776
rect 4028 16736 4034 16748
rect 4433 16745 4445 16748
rect 4479 16776 4491 16779
rect 5629 16779 5687 16785
rect 5629 16776 5641 16779
rect 4479 16748 5641 16776
rect 4479 16745 4491 16748
rect 4433 16739 4491 16745
rect 5629 16745 5641 16748
rect 5675 16745 5687 16779
rect 5994 16776 6000 16788
rect 5955 16748 6000 16776
rect 5629 16739 5687 16745
rect 5994 16736 6000 16748
rect 6052 16736 6058 16788
rect 7193 16779 7251 16785
rect 7193 16745 7205 16779
rect 7239 16745 7251 16779
rect 7193 16739 7251 16745
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 1486 16640 1492 16652
rect 1443 16612 1492 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 1486 16600 1492 16612
rect 1544 16600 1550 16652
rect 2501 16643 2559 16649
rect 2501 16609 2513 16643
rect 2547 16640 2559 16643
rect 3160 16640 3188 16736
rect 4522 16708 4528 16720
rect 4435 16680 4528 16708
rect 4522 16668 4528 16680
rect 4580 16708 4586 16720
rect 7208 16708 7236 16739
rect 7282 16736 7288 16788
rect 7340 16776 7346 16788
rect 8205 16779 8263 16785
rect 8205 16776 8217 16779
rect 7340 16748 8217 16776
rect 7340 16736 7346 16748
rect 8205 16745 8217 16748
rect 8251 16745 8263 16779
rect 8662 16776 8668 16788
rect 8623 16748 8668 16776
rect 8205 16739 8263 16745
rect 4580 16680 7236 16708
rect 7653 16711 7711 16717
rect 4580 16668 4586 16680
rect 7653 16677 7665 16711
rect 7699 16708 7711 16711
rect 7834 16708 7840 16720
rect 7699 16680 7840 16708
rect 7699 16677 7711 16680
rect 7653 16671 7711 16677
rect 7834 16668 7840 16680
rect 7892 16708 7898 16720
rect 8110 16708 8116 16720
rect 7892 16680 8116 16708
rect 7892 16668 7898 16680
rect 8110 16668 8116 16680
rect 8168 16668 8174 16720
rect 8220 16708 8248 16739
rect 8662 16736 8668 16748
rect 8720 16736 8726 16788
rect 9493 16779 9551 16785
rect 9493 16745 9505 16779
rect 9539 16776 9551 16779
rect 9582 16776 9588 16788
rect 9539 16748 9588 16776
rect 9539 16745 9551 16748
rect 9493 16739 9551 16745
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 9677 16779 9735 16785
rect 9677 16745 9689 16779
rect 9723 16745 9735 16779
rect 9677 16739 9735 16745
rect 9692 16708 9720 16739
rect 9950 16736 9956 16788
rect 10008 16776 10014 16788
rect 10137 16779 10195 16785
rect 10137 16776 10149 16779
rect 10008 16748 10149 16776
rect 10008 16736 10014 16748
rect 10137 16745 10149 16748
rect 10183 16745 10195 16779
rect 10778 16776 10784 16788
rect 10739 16748 10784 16776
rect 10137 16739 10195 16745
rect 10778 16736 10784 16748
rect 10836 16736 10842 16788
rect 13081 16779 13139 16785
rect 13081 16745 13093 16779
rect 13127 16776 13139 16779
rect 13998 16776 14004 16788
rect 13127 16748 14004 16776
rect 13127 16745 13139 16748
rect 13081 16739 13139 16745
rect 13998 16736 14004 16748
rect 14056 16736 14062 16788
rect 13630 16708 13636 16720
rect 8220 16680 9720 16708
rect 13591 16680 13636 16708
rect 13630 16668 13636 16680
rect 13688 16668 13694 16720
rect 3418 16640 3424 16652
rect 2547 16612 3188 16640
rect 3379 16612 3424 16640
rect 2547 16609 2559 16612
rect 2501 16603 2559 16609
rect 3418 16600 3424 16612
rect 3476 16600 3482 16652
rect 4890 16600 4896 16652
rect 4948 16640 4954 16652
rect 5077 16643 5135 16649
rect 5077 16640 5089 16643
rect 4948 16612 5089 16640
rect 4948 16600 4954 16612
rect 5077 16609 5089 16612
rect 5123 16609 5135 16643
rect 5077 16603 5135 16609
rect 5537 16643 5595 16649
rect 5537 16609 5549 16643
rect 5583 16640 5595 16643
rect 5718 16640 5724 16652
rect 5583 16612 5724 16640
rect 5583 16609 5595 16612
rect 5537 16603 5595 16609
rect 5718 16600 5724 16612
rect 5776 16600 5782 16652
rect 6733 16643 6791 16649
rect 6733 16609 6745 16643
rect 6779 16640 6791 16643
rect 6779 16612 6868 16640
rect 6779 16609 6791 16612
rect 6733 16603 6791 16609
rect 4709 16575 4767 16581
rect 4709 16541 4721 16575
rect 4755 16572 4767 16575
rect 4798 16572 4804 16584
rect 4755 16544 4804 16572
rect 4755 16541 4767 16544
rect 4709 16535 4767 16541
rect 4798 16532 4804 16544
rect 4856 16532 4862 16584
rect 6089 16575 6147 16581
rect 6089 16541 6101 16575
rect 6135 16572 6147 16575
rect 6178 16572 6184 16584
rect 6135 16544 6184 16572
rect 6135 16541 6147 16544
rect 6089 16535 6147 16541
rect 6178 16532 6184 16544
rect 6236 16532 6242 16584
rect 6273 16575 6331 16581
rect 6273 16541 6285 16575
rect 6319 16541 6331 16575
rect 6840 16572 6868 16612
rect 7006 16600 7012 16652
rect 7064 16640 7070 16652
rect 11974 16649 11980 16652
rect 7561 16643 7619 16649
rect 7561 16640 7573 16643
rect 7064 16612 7573 16640
rect 7064 16600 7070 16612
rect 7561 16609 7573 16612
rect 7607 16609 7619 16643
rect 7561 16603 7619 16609
rect 10045 16643 10103 16649
rect 10045 16609 10057 16643
rect 10091 16609 10103 16643
rect 10045 16603 10103 16609
rect 11968 16603 11980 16649
rect 12032 16640 12038 16652
rect 12032 16612 12068 16640
rect 7190 16572 7196 16584
rect 6840 16544 7196 16572
rect 6273 16535 6331 16541
rect 3881 16507 3939 16513
rect 3881 16473 3893 16507
rect 3927 16504 3939 16507
rect 4982 16504 4988 16516
rect 3927 16476 4988 16504
rect 3927 16473 3939 16476
rect 3881 16467 3939 16473
rect 4982 16464 4988 16476
rect 5040 16504 5046 16516
rect 5258 16504 5264 16516
rect 5040 16476 5264 16504
rect 5040 16464 5046 16476
rect 5258 16464 5264 16476
rect 5316 16504 5322 16516
rect 6288 16504 6316 16535
rect 7190 16532 7196 16544
rect 7248 16532 7254 16584
rect 7837 16575 7895 16581
rect 7837 16541 7849 16575
rect 7883 16572 7895 16575
rect 8018 16572 8024 16584
rect 7883 16544 8024 16572
rect 7883 16541 7895 16544
rect 7837 16535 7895 16541
rect 7852 16504 7880 16535
rect 8018 16532 8024 16544
rect 8076 16532 8082 16584
rect 9674 16532 9680 16584
rect 9732 16572 9738 16584
rect 10060 16572 10088 16603
rect 11974 16600 11980 16603
rect 12032 16600 12038 16612
rect 9732 16544 10088 16572
rect 9732 16532 9738 16544
rect 10134 16532 10140 16584
rect 10192 16572 10198 16584
rect 10229 16575 10287 16581
rect 10229 16572 10241 16575
rect 10192 16544 10241 16572
rect 10192 16532 10198 16544
rect 10229 16541 10241 16544
rect 10275 16541 10287 16575
rect 10229 16535 10287 16541
rect 11238 16532 11244 16584
rect 11296 16572 11302 16584
rect 11698 16572 11704 16584
rect 11296 16544 11704 16572
rect 11296 16532 11302 16544
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 5316 16476 7880 16504
rect 5316 16464 5322 16476
rect 4062 16436 4068 16448
rect 4023 16408 4068 16436
rect 4062 16396 4068 16408
rect 4120 16396 4126 16448
rect 6362 16396 6368 16448
rect 6420 16436 6426 16448
rect 7009 16439 7067 16445
rect 7009 16436 7021 16439
rect 6420 16408 7021 16436
rect 6420 16396 6426 16408
rect 7009 16405 7021 16408
rect 7055 16405 7067 16439
rect 7009 16399 7067 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2038 16232 2044 16244
rect 1999 16204 2044 16232
rect 2038 16192 2044 16204
rect 2096 16192 2102 16244
rect 4798 16232 4804 16244
rect 4759 16204 4804 16232
rect 4798 16192 4804 16204
rect 4856 16192 4862 16244
rect 5258 16232 5264 16244
rect 5219 16204 5264 16232
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 5629 16235 5687 16241
rect 5629 16201 5641 16235
rect 5675 16232 5687 16235
rect 5994 16232 6000 16244
rect 5675 16204 6000 16232
rect 5675 16201 5687 16204
rect 5629 16195 5687 16201
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 11054 16192 11060 16244
rect 11112 16232 11118 16244
rect 11149 16235 11207 16241
rect 11149 16232 11161 16235
rect 11112 16204 11161 16232
rect 11112 16192 11118 16204
rect 11149 16201 11161 16204
rect 11195 16232 11207 16235
rect 11974 16232 11980 16244
rect 11195 16204 11980 16232
rect 11195 16201 11207 16204
rect 11149 16195 11207 16201
rect 11974 16192 11980 16204
rect 12032 16232 12038 16244
rect 12069 16235 12127 16241
rect 12069 16232 12081 16235
rect 12032 16204 12081 16232
rect 12032 16192 12038 16204
rect 12069 16201 12081 16204
rect 12115 16201 12127 16235
rect 12069 16195 12127 16201
rect 11698 16164 11704 16176
rect 11659 16136 11704 16164
rect 11698 16124 11704 16136
rect 11756 16124 11762 16176
rect 2406 16096 2412 16108
rect 2367 16068 2412 16096
rect 2406 16056 2412 16068
rect 2464 16096 2470 16108
rect 2464 16068 2995 16096
rect 2464 16056 2470 16068
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 2038 16028 2044 16040
rect 1443 16000 2044 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 2038 15988 2044 16000
rect 2096 15988 2102 16040
rect 2869 16031 2927 16037
rect 2869 15997 2881 16031
rect 2915 15997 2927 16031
rect 2967 16028 2995 16068
rect 6362 16056 6368 16108
rect 6420 16096 6426 16108
rect 7101 16099 7159 16105
rect 7101 16096 7113 16099
rect 6420 16068 7113 16096
rect 6420 16056 6426 16068
rect 7101 16065 7113 16068
rect 7147 16065 7159 16099
rect 7101 16059 7159 16065
rect 9214 16056 9220 16108
rect 9272 16096 9278 16108
rect 9769 16099 9827 16105
rect 9769 16096 9781 16099
rect 9272 16068 9781 16096
rect 9272 16056 9278 16068
rect 9769 16065 9781 16068
rect 9815 16065 9827 16099
rect 9769 16059 9827 16065
rect 3125 16031 3183 16037
rect 3125 16028 3137 16031
rect 2967 16000 3137 16028
rect 2869 15991 2927 15997
rect 3125 15997 3137 16000
rect 3171 15997 3183 16031
rect 3125 15991 3183 15997
rect 1578 15892 1584 15904
rect 1539 15864 1584 15892
rect 1578 15852 1584 15864
rect 1636 15852 1642 15904
rect 2777 15895 2835 15901
rect 2777 15861 2789 15895
rect 2823 15892 2835 15895
rect 2884 15892 2912 15991
rect 7190 15988 7196 16040
rect 7248 16028 7254 16040
rect 7357 16031 7415 16037
rect 7357 16028 7369 16031
rect 7248 16000 7369 16028
rect 7248 15988 7254 16000
rect 7357 15997 7369 16000
rect 7403 15997 7415 16031
rect 9674 16028 9680 16040
rect 9635 16000 9680 16028
rect 7357 15991 7415 15997
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 10042 16037 10048 16040
rect 10036 16028 10048 16037
rect 10003 16000 10048 16028
rect 10036 15991 10048 16000
rect 10042 15988 10048 15991
rect 10100 15988 10106 16040
rect 11716 16028 11744 16124
rect 12437 16099 12495 16105
rect 12437 16065 12449 16099
rect 12483 16096 12495 16099
rect 12802 16096 12808 16108
rect 12483 16068 12808 16096
rect 12483 16065 12495 16068
rect 12437 16059 12495 16065
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 13262 16028 13268 16040
rect 11716 16000 13268 16028
rect 13262 15988 13268 16000
rect 13320 16028 13326 16040
rect 13725 16031 13783 16037
rect 13725 16028 13737 16031
rect 13320 16000 13737 16028
rect 13320 15988 13326 16000
rect 13725 15997 13737 16000
rect 13771 15997 13783 16031
rect 13725 15991 13783 15997
rect 13740 15904 13768 15991
rect 13906 15920 13912 15972
rect 13964 15969 13970 15972
rect 13964 15963 14028 15969
rect 13964 15929 13982 15963
rect 14016 15929 14028 15963
rect 13964 15923 14028 15929
rect 13964 15920 13970 15923
rect 2958 15892 2964 15904
rect 2823 15864 2964 15892
rect 2823 15861 2835 15864
rect 2777 15855 2835 15861
rect 2958 15852 2964 15864
rect 3016 15852 3022 15904
rect 4249 15895 4307 15901
rect 4249 15861 4261 15895
rect 4295 15892 4307 15895
rect 4338 15892 4344 15904
rect 4295 15864 4344 15892
rect 4295 15861 4307 15864
rect 4249 15855 4307 15861
rect 4338 15852 4344 15864
rect 4396 15852 4402 15904
rect 5718 15892 5724 15904
rect 5679 15864 5724 15892
rect 5718 15852 5724 15864
rect 5776 15852 5782 15904
rect 6270 15892 6276 15904
rect 6231 15864 6276 15892
rect 6270 15852 6276 15864
rect 6328 15852 6334 15904
rect 6641 15895 6699 15901
rect 6641 15861 6653 15895
rect 6687 15892 6699 15895
rect 6914 15892 6920 15904
rect 6687 15864 6920 15892
rect 6687 15861 6699 15864
rect 6641 15855 6699 15861
rect 6914 15852 6920 15864
rect 6972 15852 6978 15904
rect 8481 15895 8539 15901
rect 8481 15861 8493 15895
rect 8527 15892 8539 15895
rect 8754 15892 8760 15904
rect 8527 15864 8760 15892
rect 8527 15861 8539 15864
rect 8481 15855 8539 15861
rect 8754 15852 8760 15864
rect 8812 15852 8818 15904
rect 9214 15892 9220 15904
rect 9175 15864 9220 15892
rect 9214 15852 9220 15864
rect 9272 15852 9278 15904
rect 13633 15895 13691 15901
rect 13633 15861 13645 15895
rect 13679 15892 13691 15895
rect 13722 15892 13728 15904
rect 13679 15864 13728 15892
rect 13679 15861 13691 15864
rect 13633 15855 13691 15861
rect 13722 15852 13728 15864
rect 13780 15852 13786 15904
rect 15102 15892 15108 15904
rect 15063 15864 15108 15892
rect 15102 15852 15108 15864
rect 15160 15852 15166 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1486 15648 1492 15700
rect 1544 15688 1550 15700
rect 1581 15691 1639 15697
rect 1581 15688 1593 15691
rect 1544 15660 1593 15688
rect 1544 15648 1550 15660
rect 1581 15657 1593 15660
rect 1627 15688 1639 15691
rect 1857 15691 1915 15697
rect 1857 15688 1869 15691
rect 1627 15660 1869 15688
rect 1627 15657 1639 15660
rect 1581 15651 1639 15657
rect 1857 15657 1869 15660
rect 1903 15657 1915 15691
rect 2314 15688 2320 15700
rect 2275 15660 2320 15688
rect 1857 15651 1915 15657
rect 2314 15648 2320 15660
rect 2372 15688 2378 15700
rect 2777 15691 2835 15697
rect 2777 15688 2789 15691
rect 2372 15660 2789 15688
rect 2372 15648 2378 15660
rect 2777 15657 2789 15660
rect 2823 15657 2835 15691
rect 2777 15651 2835 15657
rect 2869 15691 2927 15697
rect 2869 15657 2881 15691
rect 2915 15688 2927 15691
rect 4062 15688 4068 15700
rect 2915 15660 4068 15688
rect 2915 15657 2927 15660
rect 2869 15651 2927 15657
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 4246 15688 4252 15700
rect 4207 15660 4252 15688
rect 4246 15648 4252 15660
rect 4304 15648 4310 15700
rect 4522 15688 4528 15700
rect 4483 15660 4528 15688
rect 4522 15648 4528 15660
rect 4580 15648 4586 15700
rect 5261 15691 5319 15697
rect 5261 15657 5273 15691
rect 5307 15688 5319 15691
rect 5534 15688 5540 15700
rect 5307 15660 5540 15688
rect 5307 15657 5319 15660
rect 5261 15651 5319 15657
rect 5534 15648 5540 15660
rect 5592 15688 5598 15700
rect 5718 15688 5724 15700
rect 5592 15660 5724 15688
rect 5592 15648 5598 15660
rect 5718 15648 5724 15660
rect 5776 15648 5782 15700
rect 7101 15691 7159 15697
rect 7101 15657 7113 15691
rect 7147 15688 7159 15691
rect 7190 15688 7196 15700
rect 7147 15660 7196 15688
rect 7147 15657 7159 15660
rect 7101 15651 7159 15657
rect 7190 15648 7196 15660
rect 7248 15648 7254 15700
rect 7745 15691 7803 15697
rect 7745 15657 7757 15691
rect 7791 15688 7803 15691
rect 7834 15688 7840 15700
rect 7791 15660 7840 15688
rect 7791 15657 7803 15660
rect 7745 15651 7803 15657
rect 7834 15648 7840 15660
rect 7892 15648 7898 15700
rect 8018 15688 8024 15700
rect 7979 15660 8024 15688
rect 8018 15648 8024 15660
rect 8076 15648 8082 15700
rect 9493 15691 9551 15697
rect 9493 15657 9505 15691
rect 9539 15688 9551 15691
rect 9950 15688 9956 15700
rect 9539 15660 9956 15688
rect 9539 15657 9551 15660
rect 9493 15651 9551 15657
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 10134 15648 10140 15700
rect 10192 15688 10198 15700
rect 10229 15691 10287 15697
rect 10229 15688 10241 15691
rect 10192 15660 10241 15688
rect 10192 15648 10198 15660
rect 10229 15657 10241 15660
rect 10275 15657 10287 15691
rect 10778 15688 10784 15700
rect 10739 15660 10784 15688
rect 10229 15651 10287 15657
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 11238 15688 11244 15700
rect 11151 15660 11244 15688
rect 11238 15648 11244 15660
rect 11296 15688 11302 15700
rect 12345 15691 12403 15697
rect 12345 15688 12357 15691
rect 11296 15660 12357 15688
rect 11296 15648 11302 15660
rect 12345 15657 12357 15660
rect 12391 15657 12403 15691
rect 12345 15651 12403 15657
rect 13817 15691 13875 15697
rect 13817 15657 13829 15691
rect 13863 15688 13875 15691
rect 13906 15688 13912 15700
rect 13863 15660 13912 15688
rect 13863 15657 13875 15660
rect 13817 15651 13875 15657
rect 3881 15623 3939 15629
rect 3881 15589 3893 15623
rect 3927 15620 3939 15623
rect 3970 15620 3976 15632
rect 3927 15592 3976 15620
rect 3927 15589 3939 15592
rect 3881 15583 3939 15589
rect 3970 15580 3976 15592
rect 4028 15580 4034 15632
rect 6178 15620 6184 15632
rect 5736 15592 6184 15620
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15552 1455 15555
rect 2038 15552 2044 15564
rect 1443 15524 2044 15552
rect 1443 15521 1455 15524
rect 1397 15515 1455 15521
rect 2038 15512 2044 15524
rect 2096 15512 2102 15564
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15552 4123 15555
rect 4154 15552 4160 15564
rect 4111 15524 4160 15552
rect 4111 15521 4123 15524
rect 4065 15515 4123 15521
rect 4154 15512 4160 15524
rect 4212 15512 4218 15564
rect 5736 15561 5764 15592
rect 6178 15580 6184 15592
rect 6236 15620 6242 15632
rect 6362 15620 6368 15632
rect 6236 15592 6368 15620
rect 6236 15580 6242 15592
rect 6362 15580 6368 15592
rect 6420 15620 6426 15632
rect 8478 15620 8484 15632
rect 6420 15592 8484 15620
rect 6420 15580 6426 15592
rect 8478 15580 8484 15592
rect 8536 15580 8542 15632
rect 11149 15623 11207 15629
rect 11149 15589 11161 15623
rect 11195 15620 11207 15623
rect 11606 15620 11612 15632
rect 11195 15592 11612 15620
rect 11195 15589 11207 15592
rect 11149 15583 11207 15589
rect 11606 15580 11612 15592
rect 11664 15580 11670 15632
rect 12713 15623 12771 15629
rect 12713 15589 12725 15623
rect 12759 15620 12771 15623
rect 12802 15620 12808 15632
rect 12759 15592 12808 15620
rect 12759 15589 12771 15592
rect 12713 15583 12771 15589
rect 12802 15580 12808 15592
rect 12860 15580 12866 15632
rect 5994 15561 6000 15564
rect 5721 15555 5779 15561
rect 5721 15521 5733 15555
rect 5767 15521 5779 15555
rect 5988 15552 6000 15561
rect 5955 15524 6000 15552
rect 5721 15515 5779 15521
rect 5988 15515 6000 15524
rect 5994 15512 6000 15515
rect 6052 15512 6058 15564
rect 9953 15555 10011 15561
rect 9953 15521 9965 15555
rect 9999 15552 10011 15555
rect 10042 15552 10048 15564
rect 9999 15524 10048 15552
rect 9999 15521 10011 15524
rect 9953 15515 10011 15521
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 13446 15552 13452 15564
rect 12820 15524 13452 15552
rect 3050 15484 3056 15496
rect 3011 15456 3056 15484
rect 3050 15444 3056 15456
rect 3108 15444 3114 15496
rect 8570 15484 8576 15496
rect 8531 15456 8576 15484
rect 8570 15444 8576 15456
rect 8628 15444 8634 15496
rect 10962 15444 10968 15496
rect 11020 15484 11026 15496
rect 11422 15484 11428 15496
rect 11020 15456 11428 15484
rect 11020 15444 11026 15456
rect 11422 15444 11428 15456
rect 11480 15444 11486 15496
rect 12434 15444 12440 15496
rect 12492 15484 12498 15496
rect 12820 15493 12848 15524
rect 13446 15512 13452 15524
rect 13504 15512 13510 15564
rect 12805 15487 12863 15493
rect 12805 15484 12817 15487
rect 12492 15456 12817 15484
rect 12492 15444 12498 15456
rect 12805 15453 12817 15456
rect 12851 15453 12863 15487
rect 12805 15447 12863 15453
rect 12989 15487 13047 15493
rect 12989 15453 13001 15487
rect 13035 15484 13047 15487
rect 13170 15484 13176 15496
rect 13035 15456 13176 15484
rect 13035 15453 13047 15456
rect 12989 15447 13047 15453
rect 13170 15444 13176 15456
rect 13228 15484 13234 15496
rect 13832 15484 13860 15651
rect 13906 15648 13912 15660
rect 13964 15648 13970 15700
rect 14366 15688 14372 15700
rect 14327 15660 14372 15688
rect 14366 15648 14372 15660
rect 14424 15648 14430 15700
rect 15105 15623 15163 15629
rect 15105 15589 15117 15623
rect 15151 15620 15163 15623
rect 15749 15623 15807 15629
rect 15749 15620 15761 15623
rect 15151 15592 15761 15620
rect 15151 15589 15163 15592
rect 15105 15583 15163 15589
rect 15749 15589 15761 15592
rect 15795 15620 15807 15623
rect 16298 15620 16304 15632
rect 15795 15592 16304 15620
rect 15795 15589 15807 15592
rect 15749 15583 15807 15589
rect 16298 15580 16304 15592
rect 16356 15580 16362 15632
rect 14182 15552 14188 15564
rect 14143 15524 14188 15552
rect 14182 15512 14188 15524
rect 14240 15512 14246 15564
rect 15657 15555 15715 15561
rect 15657 15552 15669 15555
rect 14660 15524 15669 15552
rect 13228 15456 13860 15484
rect 13228 15444 13234 15456
rect 14660 15428 14688 15524
rect 15657 15521 15669 15524
rect 15703 15521 15715 15555
rect 15657 15515 15715 15521
rect 15933 15487 15991 15493
rect 15933 15453 15945 15487
rect 15979 15453 15991 15487
rect 15933 15447 15991 15453
rect 2498 15376 2504 15428
rect 2556 15416 2562 15428
rect 3421 15419 3479 15425
rect 3421 15416 3433 15419
rect 2556 15388 3433 15416
rect 2556 15376 2562 15388
rect 3421 15385 3433 15388
rect 3467 15385 3479 15419
rect 14642 15416 14648 15428
rect 14603 15388 14648 15416
rect 3421 15379 3479 15385
rect 14642 15376 14648 15388
rect 14700 15376 14706 15428
rect 15838 15376 15844 15428
rect 15896 15416 15902 15428
rect 15948 15416 15976 15447
rect 15896 15388 15976 15416
rect 15896 15376 15902 15388
rect 2409 15351 2467 15357
rect 2409 15317 2421 15351
rect 2455 15348 2467 15351
rect 2774 15348 2780 15360
rect 2455 15320 2780 15348
rect 2455 15317 2467 15320
rect 2409 15311 2467 15317
rect 2774 15308 2780 15320
rect 2832 15308 2838 15360
rect 5442 15308 5448 15360
rect 5500 15348 5506 15360
rect 5629 15351 5687 15357
rect 5629 15348 5641 15351
rect 5500 15320 5641 15348
rect 5500 15308 5506 15320
rect 5629 15317 5641 15320
rect 5675 15348 5687 15351
rect 6822 15348 6828 15360
rect 5675 15320 6828 15348
rect 5675 15317 5687 15320
rect 5629 15311 5687 15317
rect 6822 15308 6828 15320
rect 6880 15308 6886 15360
rect 8294 15308 8300 15360
rect 8352 15348 8358 15360
rect 8389 15351 8447 15357
rect 8389 15348 8401 15351
rect 8352 15320 8401 15348
rect 8352 15308 8358 15320
rect 8389 15317 8401 15320
rect 8435 15317 8447 15351
rect 9030 15348 9036 15360
rect 8991 15320 9036 15348
rect 8389 15311 8447 15317
rect 9030 15308 9036 15320
rect 9088 15308 9094 15360
rect 15289 15351 15347 15357
rect 15289 15317 15301 15351
rect 15335 15348 15347 15351
rect 15470 15348 15476 15360
rect 15335 15320 15476 15348
rect 15335 15317 15347 15320
rect 15289 15311 15347 15317
rect 15470 15308 15476 15320
rect 15528 15308 15534 15360
rect 16482 15348 16488 15360
rect 16443 15320 16488 15348
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2038 15144 2044 15156
rect 1999 15116 2044 15144
rect 2038 15104 2044 15116
rect 2096 15104 2102 15156
rect 3513 15147 3571 15153
rect 3513 15113 3525 15147
rect 3559 15144 3571 15147
rect 4062 15144 4068 15156
rect 3559 15116 4068 15144
rect 3559 15113 3571 15116
rect 3513 15107 3571 15113
rect 4062 15104 4068 15116
rect 4120 15104 4126 15156
rect 5169 15147 5227 15153
rect 5169 15113 5181 15147
rect 5215 15144 5227 15147
rect 5442 15144 5448 15156
rect 5215 15116 5448 15144
rect 5215 15113 5227 15116
rect 5169 15107 5227 15113
rect 5442 15104 5448 15116
rect 5500 15104 5506 15156
rect 6641 15147 6699 15153
rect 6641 15113 6653 15147
rect 6687 15144 6699 15147
rect 7190 15144 7196 15156
rect 6687 15116 7196 15144
rect 6687 15113 6699 15116
rect 6641 15107 6699 15113
rect 7190 15104 7196 15116
rect 7248 15104 7254 15156
rect 8478 15144 8484 15156
rect 8439 15116 8484 15144
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 10042 15144 10048 15156
rect 10003 15116 10048 15144
rect 10042 15104 10048 15116
rect 10100 15104 10106 15156
rect 10873 15147 10931 15153
rect 10873 15113 10885 15147
rect 10919 15144 10931 15147
rect 10962 15144 10968 15156
rect 10919 15116 10968 15144
rect 10919 15113 10931 15116
rect 10873 15107 10931 15113
rect 10962 15104 10968 15116
rect 11020 15104 11026 15156
rect 11238 15144 11244 15156
rect 11199 15116 11244 15144
rect 11238 15104 11244 15116
rect 11296 15104 11302 15156
rect 11606 15144 11612 15156
rect 11567 15116 11612 15144
rect 11606 15104 11612 15116
rect 11664 15104 11670 15156
rect 12253 15147 12311 15153
rect 12253 15113 12265 15147
rect 12299 15144 12311 15147
rect 12342 15144 12348 15156
rect 12299 15116 12348 15144
rect 12299 15113 12311 15116
rect 12253 15107 12311 15113
rect 12342 15104 12348 15116
rect 12400 15104 12406 15156
rect 13081 15147 13139 15153
rect 13081 15113 13093 15147
rect 13127 15144 13139 15147
rect 13170 15144 13176 15156
rect 13127 15116 13176 15144
rect 13127 15113 13139 15116
rect 13081 15107 13139 15113
rect 13170 15104 13176 15116
rect 13228 15104 13234 15156
rect 16298 15104 16304 15156
rect 16356 15144 16362 15156
rect 16393 15147 16451 15153
rect 16393 15144 16405 15147
rect 16356 15116 16405 15144
rect 16356 15104 16362 15116
rect 16393 15113 16405 15116
rect 16439 15113 16451 15147
rect 16393 15107 16451 15113
rect 2409 15079 2467 15085
rect 2409 15045 2421 15079
rect 2455 15076 2467 15079
rect 3789 15079 3847 15085
rect 3789 15076 3801 15079
rect 2455 15048 3801 15076
rect 2455 15045 2467 15048
rect 2409 15039 2467 15045
rect 3789 15045 3801 15048
rect 3835 15045 3847 15079
rect 4154 15076 4160 15088
rect 4067 15048 4160 15076
rect 3789 15039 3847 15045
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14940 1455 14943
rect 2424 14940 2452 15039
rect 4154 15036 4160 15048
rect 4212 15076 4218 15088
rect 5350 15076 5356 15088
rect 4212 15048 5356 15076
rect 4212 15036 4218 15048
rect 5350 15036 5356 15048
rect 5408 15036 5414 15088
rect 2590 14968 2596 15020
rect 2648 15008 2654 15020
rect 2866 15008 2872 15020
rect 2648 14980 2872 15008
rect 2648 14968 2654 14980
rect 2866 14968 2872 14980
rect 2924 14968 2930 15020
rect 4709 15011 4767 15017
rect 4709 14977 4721 15011
rect 4755 15008 4767 15011
rect 5721 15011 5779 15017
rect 5721 15008 5733 15011
rect 4755 14980 5733 15008
rect 4755 14977 4767 14980
rect 4709 14971 4767 14977
rect 5721 14977 5733 14980
rect 5767 15008 5779 15011
rect 5994 15008 6000 15020
rect 5767 14980 6000 15008
rect 5767 14977 5779 14980
rect 5721 14971 5779 14977
rect 5994 14968 6000 14980
rect 6052 14968 6058 15020
rect 7208 15008 7236 15104
rect 7377 15011 7435 15017
rect 7377 15008 7389 15011
rect 7208 14980 7389 15008
rect 7377 14977 7389 14980
rect 7423 14977 7435 15011
rect 8496 15008 8524 15104
rect 8665 15011 8723 15017
rect 8665 15008 8677 15011
rect 8496 14980 8677 15008
rect 7377 14971 7435 14977
rect 8665 14977 8677 14980
rect 8711 14977 8723 15011
rect 8665 14971 8723 14977
rect 1443 14912 2452 14940
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 2498 14900 2504 14952
rect 2556 14940 2562 14952
rect 2556 14912 2601 14940
rect 2556 14900 2562 14912
rect 2774 14900 2780 14952
rect 2832 14940 2838 14952
rect 3602 14940 3608 14952
rect 2832 14912 3608 14940
rect 2832 14900 2838 14912
rect 3602 14900 3608 14912
rect 3660 14900 3666 14952
rect 5534 14940 5540 14952
rect 5495 14912 5540 14940
rect 5534 14900 5540 14912
rect 5592 14900 5598 14952
rect 6822 14900 6828 14952
rect 6880 14940 6886 14952
rect 7193 14943 7251 14949
rect 7193 14940 7205 14943
rect 6880 14912 7205 14940
rect 6880 14900 6886 14912
rect 7193 14909 7205 14912
rect 7239 14909 7251 14943
rect 7193 14903 7251 14909
rect 7282 14900 7288 14952
rect 7340 14940 7346 14952
rect 8202 14940 8208 14952
rect 7340 14912 8208 14940
rect 7340 14900 7346 14912
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 8680 14940 8708 14971
rect 16482 14968 16488 15020
rect 16540 15008 16546 15020
rect 17037 15011 17095 15017
rect 17037 15008 17049 15011
rect 16540 14980 17049 15008
rect 16540 14968 16546 14980
rect 17037 14977 17049 14980
rect 17083 15008 17095 15011
rect 17862 15008 17868 15020
rect 17083 14980 17868 15008
rect 17083 14977 17095 14980
rect 17037 14971 17095 14977
rect 17862 14968 17868 14980
rect 17920 14968 17926 15020
rect 9214 14940 9220 14952
rect 8680 14912 9220 14940
rect 9214 14900 9220 14912
rect 9272 14900 9278 14952
rect 13722 14900 13728 14952
rect 13780 14940 13786 14952
rect 13909 14943 13967 14949
rect 13909 14940 13921 14943
rect 13780 14912 13921 14940
rect 13780 14900 13786 14912
rect 13909 14909 13921 14912
rect 13955 14940 13967 14943
rect 13955 14912 14320 14940
rect 13955 14909 13967 14912
rect 13909 14903 13967 14909
rect 3050 14832 3056 14884
rect 3108 14872 3114 14884
rect 3145 14875 3203 14881
rect 3145 14872 3157 14875
rect 3108 14844 3157 14872
rect 3108 14832 3114 14844
rect 3145 14841 3157 14844
rect 3191 14872 3203 14875
rect 4338 14872 4344 14884
rect 3191 14844 4344 14872
rect 3191 14841 3203 14844
rect 3145 14835 3203 14841
rect 4338 14832 4344 14844
rect 4396 14832 4402 14884
rect 5077 14875 5135 14881
rect 5077 14841 5089 14875
rect 5123 14872 5135 14875
rect 5629 14875 5687 14881
rect 5629 14872 5641 14875
rect 5123 14844 5641 14872
rect 5123 14841 5135 14844
rect 5077 14835 5135 14841
rect 5629 14841 5641 14844
rect 5675 14872 5687 14875
rect 6546 14872 6552 14884
rect 5675 14844 6552 14872
rect 5675 14841 5687 14844
rect 5629 14835 5687 14841
rect 6546 14832 6552 14844
rect 6604 14832 6610 14884
rect 8754 14832 8760 14884
rect 8812 14872 8818 14884
rect 8910 14875 8968 14881
rect 8910 14872 8922 14875
rect 8812 14844 8922 14872
rect 8812 14832 8818 14844
rect 8910 14841 8922 14844
rect 8956 14841 8968 14875
rect 8910 14835 8968 14841
rect 13170 14832 13176 14884
rect 13228 14872 13234 14884
rect 13449 14875 13507 14881
rect 13449 14872 13461 14875
rect 13228 14844 13461 14872
rect 13228 14832 13234 14844
rect 13449 14841 13461 14844
rect 13495 14872 13507 14875
rect 14090 14872 14096 14884
rect 13495 14844 14096 14872
rect 13495 14841 13507 14844
rect 13449 14835 13507 14841
rect 14090 14832 14096 14844
rect 14148 14881 14154 14884
rect 14148 14875 14212 14881
rect 14148 14841 14166 14875
rect 14200 14841 14212 14875
rect 14148 14835 14212 14841
rect 14148 14832 14154 14835
rect 1394 14764 1400 14816
rect 1452 14804 1458 14816
rect 1581 14807 1639 14813
rect 1581 14804 1593 14807
rect 1452 14776 1593 14804
rect 1452 14764 1458 14776
rect 1581 14773 1593 14776
rect 1627 14773 1639 14807
rect 2682 14804 2688 14816
rect 2643 14776 2688 14804
rect 1581 14767 1639 14773
rect 2682 14764 2688 14776
rect 2740 14764 2746 14816
rect 4154 14764 4160 14816
rect 4212 14804 4218 14816
rect 6178 14804 6184 14816
rect 4212 14776 6184 14804
rect 4212 14764 4218 14776
rect 6178 14764 6184 14776
rect 6236 14764 6242 14816
rect 6822 14804 6828 14816
rect 6783 14776 6828 14804
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7834 14804 7840 14816
rect 7795 14776 7840 14804
rect 7834 14764 7840 14776
rect 7892 14764 7898 14816
rect 12713 14807 12771 14813
rect 12713 14773 12725 14807
rect 12759 14804 12771 14807
rect 12802 14804 12808 14816
rect 12759 14776 12808 14804
rect 12759 14773 12771 14776
rect 12713 14767 12771 14773
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 13817 14807 13875 14813
rect 13817 14773 13829 14807
rect 13863 14804 13875 14807
rect 14292 14804 14320 14912
rect 16853 14875 16911 14881
rect 16853 14872 16865 14875
rect 16224 14844 16865 14872
rect 16224 14816 16252 14844
rect 16853 14841 16865 14844
rect 16899 14841 16911 14875
rect 16853 14835 16911 14841
rect 14366 14804 14372 14816
rect 13863 14776 14372 14804
rect 13863 14773 13875 14776
rect 13817 14767 13875 14773
rect 14366 14764 14372 14776
rect 14424 14764 14430 14816
rect 15289 14807 15347 14813
rect 15289 14773 15301 14807
rect 15335 14804 15347 14807
rect 15378 14804 15384 14816
rect 15335 14776 15384 14804
rect 15335 14773 15347 14776
rect 15289 14767 15347 14773
rect 15378 14764 15384 14776
rect 15436 14764 15442 14816
rect 15838 14804 15844 14816
rect 15799 14776 15844 14804
rect 15838 14764 15844 14776
rect 15896 14764 15902 14816
rect 16206 14804 16212 14816
rect 16167 14776 16212 14804
rect 16206 14764 16212 14776
rect 16264 14764 16270 14816
rect 16390 14764 16396 14816
rect 16448 14804 16454 14816
rect 16761 14807 16819 14813
rect 16761 14804 16773 14807
rect 16448 14776 16773 14804
rect 16448 14764 16454 14776
rect 16761 14773 16773 14776
rect 16807 14773 16819 14807
rect 16761 14767 16819 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1581 14603 1639 14609
rect 1581 14569 1593 14603
rect 1627 14600 1639 14603
rect 2498 14600 2504 14612
rect 1627 14572 2504 14600
rect 1627 14569 1639 14572
rect 1581 14563 1639 14569
rect 2498 14560 2504 14572
rect 2556 14560 2562 14612
rect 3602 14600 3608 14612
rect 3563 14572 3608 14600
rect 3602 14560 3608 14572
rect 3660 14560 3666 14612
rect 5445 14603 5503 14609
rect 5445 14569 5457 14603
rect 5491 14569 5503 14603
rect 5994 14600 6000 14612
rect 5955 14572 6000 14600
rect 5445 14563 5503 14569
rect 5460 14532 5488 14563
rect 5994 14560 6000 14572
rect 6052 14600 6058 14612
rect 7374 14600 7380 14612
rect 6052 14572 7380 14600
rect 6052 14560 6058 14572
rect 7374 14560 7380 14572
rect 7432 14600 7438 14612
rect 7929 14603 7987 14609
rect 7929 14600 7941 14603
rect 7432 14572 7941 14600
rect 7432 14560 7438 14572
rect 7929 14569 7941 14572
rect 7975 14569 7987 14603
rect 7929 14563 7987 14569
rect 9677 14603 9735 14609
rect 9677 14569 9689 14603
rect 9723 14600 9735 14603
rect 9766 14600 9772 14612
rect 9723 14572 9772 14600
rect 9723 14569 9735 14572
rect 9677 14563 9735 14569
rect 9766 14560 9772 14572
rect 9824 14560 9830 14612
rect 9858 14560 9864 14612
rect 9916 14600 9922 14612
rect 10137 14603 10195 14609
rect 10137 14600 10149 14603
rect 9916 14572 10149 14600
rect 9916 14560 9922 14572
rect 10137 14569 10149 14572
rect 10183 14569 10195 14603
rect 14090 14600 14096 14612
rect 14051 14572 14096 14600
rect 10137 14563 10195 14569
rect 14090 14560 14096 14572
rect 14148 14560 14154 14612
rect 15749 14603 15807 14609
rect 15749 14569 15761 14603
rect 15795 14600 15807 14603
rect 16298 14600 16304 14612
rect 15795 14572 16304 14600
rect 15795 14569 15807 14572
rect 15749 14563 15807 14569
rect 16298 14560 16304 14572
rect 16356 14600 16362 14612
rect 16853 14603 16911 14609
rect 16853 14600 16865 14603
rect 16356 14572 16865 14600
rect 16356 14560 16362 14572
rect 16853 14569 16865 14572
rect 16899 14569 16911 14603
rect 16853 14563 16911 14569
rect 6546 14532 6552 14544
rect 5460 14504 6552 14532
rect 6546 14492 6552 14504
rect 6604 14532 6610 14544
rect 6794 14535 6852 14541
rect 6794 14532 6806 14535
rect 6604 14504 6806 14532
rect 6604 14492 6610 14504
rect 6794 14501 6806 14504
rect 6840 14501 6852 14535
rect 6794 14495 6852 14501
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 2038 14464 2044 14476
rect 1443 14436 2044 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 2038 14424 2044 14436
rect 2096 14424 2102 14476
rect 2222 14424 2228 14476
rect 2280 14464 2286 14476
rect 2777 14467 2835 14473
rect 2777 14464 2789 14467
rect 2280 14436 2789 14464
rect 2280 14424 2286 14436
rect 2777 14433 2789 14436
rect 2823 14433 2835 14467
rect 2777 14427 2835 14433
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 4154 14464 4160 14476
rect 4111 14436 4160 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 4154 14424 4160 14436
rect 4212 14424 4218 14476
rect 4338 14473 4344 14476
rect 4332 14464 4344 14473
rect 4299 14436 4344 14464
rect 4332 14427 4344 14436
rect 4338 14424 4344 14427
rect 4396 14424 4402 14476
rect 9493 14467 9551 14473
rect 9493 14433 9505 14467
rect 9539 14464 9551 14467
rect 9950 14464 9956 14476
rect 9539 14436 9956 14464
rect 9539 14433 9551 14436
rect 9493 14427 9551 14433
rect 9950 14424 9956 14436
rect 10008 14464 10014 14476
rect 10045 14467 10103 14473
rect 10045 14464 10057 14467
rect 10008 14436 10057 14464
rect 10008 14424 10014 14436
rect 10045 14433 10057 14436
rect 10091 14433 10103 14467
rect 10045 14427 10103 14433
rect 12980 14467 13038 14473
rect 12980 14433 12992 14467
rect 13026 14464 13038 14467
rect 13354 14464 13360 14476
rect 13026 14436 13360 14464
rect 13026 14433 13038 14436
rect 12980 14427 13038 14433
rect 13354 14424 13360 14436
rect 13412 14464 13418 14476
rect 15013 14467 15071 14473
rect 15013 14464 15025 14467
rect 13412 14436 15025 14464
rect 13412 14424 13418 14436
rect 15013 14433 15025 14436
rect 15059 14433 15071 14467
rect 15654 14464 15660 14476
rect 15615 14436 15660 14464
rect 15013 14427 15071 14433
rect 2866 14396 2872 14408
rect 2827 14368 2872 14396
rect 2866 14356 2872 14368
rect 2924 14356 2930 14408
rect 3053 14399 3111 14405
rect 3053 14365 3065 14399
rect 3099 14396 3111 14399
rect 3510 14396 3516 14408
rect 3099 14368 3516 14396
rect 3099 14365 3111 14368
rect 3053 14359 3111 14365
rect 2317 14331 2375 14337
rect 2317 14297 2329 14331
rect 2363 14328 2375 14331
rect 3068 14328 3096 14359
rect 3510 14356 3516 14368
rect 3568 14356 3574 14408
rect 6178 14356 6184 14408
rect 6236 14396 6242 14408
rect 6549 14399 6607 14405
rect 6549 14396 6561 14399
rect 6236 14368 6561 14396
rect 6236 14356 6242 14368
rect 6549 14365 6561 14368
rect 6595 14365 6607 14399
rect 6549 14359 6607 14365
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14396 10379 14399
rect 11054 14396 11060 14408
rect 10367 14368 11060 14396
rect 10367 14365 10379 14368
rect 10321 14359 10379 14365
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 12710 14396 12716 14408
rect 12671 14368 12716 14396
rect 12710 14356 12716 14368
rect 12768 14356 12774 14408
rect 15028 14396 15056 14427
rect 15654 14424 15660 14436
rect 15712 14424 15718 14476
rect 17218 14464 17224 14476
rect 17179 14436 17224 14464
rect 17218 14424 17224 14436
rect 17276 14424 17282 14476
rect 15838 14396 15844 14408
rect 15028 14368 15844 14396
rect 15838 14356 15844 14368
rect 15896 14356 15902 14408
rect 16390 14396 16396 14408
rect 16351 14368 16396 14396
rect 16390 14356 16396 14368
rect 16448 14356 16454 14408
rect 16850 14356 16856 14408
rect 16908 14396 16914 14408
rect 17313 14399 17371 14405
rect 17313 14396 17325 14399
rect 16908 14368 17325 14396
rect 16908 14356 16914 14368
rect 17313 14365 17325 14368
rect 17359 14365 17371 14399
rect 17313 14359 17371 14365
rect 17497 14399 17555 14405
rect 17497 14365 17509 14399
rect 17543 14396 17555 14399
rect 17862 14396 17868 14408
rect 17543 14368 17868 14396
rect 17543 14365 17555 14368
rect 17497 14359 17555 14365
rect 17862 14356 17868 14368
rect 17920 14356 17926 14408
rect 2363 14300 3096 14328
rect 2363 14297 2375 14300
rect 2317 14291 2375 14297
rect 14090 14288 14096 14340
rect 14148 14328 14154 14340
rect 16206 14328 16212 14340
rect 14148 14300 16212 14328
rect 14148 14288 14154 14300
rect 16206 14288 16212 14300
rect 16264 14288 16270 14340
rect 1854 14260 1860 14272
rect 1815 14232 1860 14260
rect 1854 14220 1860 14232
rect 1912 14220 1918 14272
rect 2406 14260 2412 14272
rect 2367 14232 2412 14260
rect 2406 14220 2412 14232
rect 2464 14220 2470 14272
rect 6362 14260 6368 14272
rect 6323 14232 6368 14260
rect 6362 14220 6368 14232
rect 6420 14220 6426 14272
rect 8754 14260 8760 14272
rect 8715 14232 8760 14260
rect 8754 14220 8760 14232
rect 8812 14220 8818 14272
rect 9125 14263 9183 14269
rect 9125 14229 9137 14263
rect 9171 14260 9183 14263
rect 9582 14260 9588 14272
rect 9171 14232 9588 14260
rect 9171 14229 9183 14232
rect 9125 14223 9183 14229
rect 9582 14220 9588 14232
rect 9640 14220 9646 14272
rect 12526 14260 12532 14272
rect 12487 14232 12532 14260
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 14642 14260 14648 14272
rect 14603 14232 14648 14260
rect 14642 14220 14648 14232
rect 14700 14220 14706 14272
rect 15286 14260 15292 14272
rect 15247 14232 15292 14260
rect 15286 14220 15292 14232
rect 15344 14220 15350 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 4338 14016 4344 14068
rect 4396 14056 4402 14068
rect 4433 14059 4491 14065
rect 4433 14056 4445 14059
rect 4396 14028 4445 14056
rect 4396 14016 4402 14028
rect 4433 14025 4445 14028
rect 4479 14025 4491 14059
rect 4433 14019 4491 14025
rect 4798 14016 4804 14068
rect 4856 14056 4862 14068
rect 4985 14059 5043 14065
rect 4985 14056 4997 14059
rect 4856 14028 4997 14056
rect 4856 14016 4862 14028
rect 4985 14025 4997 14028
rect 5031 14025 5043 14059
rect 5166 14056 5172 14068
rect 5127 14028 5172 14056
rect 4985 14019 5043 14025
rect 1578 13988 1584 14000
rect 1539 13960 1584 13988
rect 1578 13948 1584 13960
rect 1636 13948 1642 14000
rect 2869 13991 2927 13997
rect 2869 13957 2881 13991
rect 2915 13988 2927 13991
rect 3786 13988 3792 14000
rect 2915 13960 3792 13988
rect 2915 13957 2927 13960
rect 2869 13951 2927 13957
rect 3786 13948 3792 13960
rect 3844 13948 3850 14000
rect 3326 13920 3332 13932
rect 3287 13892 3332 13920
rect 3326 13880 3332 13892
rect 3384 13880 3390 13932
rect 3510 13920 3516 13932
rect 3471 13892 3516 13920
rect 3510 13880 3516 13892
rect 3568 13880 3574 13932
rect 5000 13920 5028 14019
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 6178 14056 6184 14068
rect 6139 14028 6184 14056
rect 6178 14016 6184 14028
rect 6236 14016 6242 14068
rect 6825 14059 6883 14065
rect 6825 14025 6837 14059
rect 6871 14056 6883 14059
rect 7282 14056 7288 14068
rect 6871 14028 7288 14056
rect 6871 14025 6883 14028
rect 6825 14019 6883 14025
rect 7282 14016 7288 14028
rect 7340 14016 7346 14068
rect 8570 14016 8576 14068
rect 8628 14056 8634 14068
rect 9401 14059 9459 14065
rect 9401 14056 9413 14059
rect 8628 14028 9413 14056
rect 8628 14016 8634 14028
rect 9401 14025 9413 14028
rect 9447 14025 9459 14059
rect 9766 14056 9772 14068
rect 9727 14028 9772 14056
rect 9401 14019 9459 14025
rect 6086 13948 6092 14000
rect 6144 13988 6150 14000
rect 6730 13988 6736 14000
rect 6144 13960 6736 13988
rect 6144 13948 6150 13960
rect 6730 13948 6736 13960
rect 6788 13948 6794 14000
rect 8202 13948 8208 14000
rect 8260 13988 8266 14000
rect 8389 13991 8447 13997
rect 8389 13988 8401 13991
rect 8260 13960 8401 13988
rect 8260 13948 8266 13960
rect 8389 13957 8401 13960
rect 8435 13957 8447 13991
rect 8389 13951 8447 13957
rect 5442 13920 5448 13932
rect 5000 13892 5448 13920
rect 5442 13880 5448 13892
rect 5500 13920 5506 13932
rect 5629 13923 5687 13929
rect 5629 13920 5641 13923
rect 5500 13892 5641 13920
rect 5500 13880 5506 13892
rect 5629 13889 5641 13892
rect 5675 13889 5687 13923
rect 5629 13883 5687 13889
rect 5813 13923 5871 13929
rect 5813 13889 5825 13923
rect 5859 13920 5871 13923
rect 6362 13920 6368 13932
rect 5859 13892 6368 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 6362 13880 6368 13892
rect 6420 13880 6426 13932
rect 7374 13920 7380 13932
rect 7335 13892 7380 13920
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 7929 13923 7987 13929
rect 7929 13889 7941 13923
rect 7975 13920 7987 13923
rect 9030 13920 9036 13932
rect 7975 13892 9036 13920
rect 7975 13889 7987 13892
rect 7929 13883 7987 13889
rect 9030 13880 9036 13892
rect 9088 13880 9094 13932
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 1854 13852 1860 13864
rect 1443 13824 1860 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 1854 13812 1860 13824
rect 1912 13812 1918 13864
rect 2222 13812 2228 13864
rect 2280 13852 2286 13864
rect 2409 13855 2467 13861
rect 2409 13852 2421 13855
rect 2280 13824 2421 13852
rect 2280 13812 2286 13824
rect 2409 13821 2421 13824
rect 2455 13821 2467 13855
rect 2958 13852 2964 13864
rect 2409 13815 2467 13821
rect 2700 13824 2964 13852
rect 2130 13716 2136 13728
rect 2091 13688 2136 13716
rect 2130 13676 2136 13688
rect 2188 13676 2194 13728
rect 2314 13676 2320 13728
rect 2372 13716 2378 13728
rect 2700 13716 2728 13824
rect 2958 13812 2964 13824
rect 3016 13852 3022 13864
rect 4157 13855 4215 13861
rect 4157 13852 4169 13855
rect 3016 13824 4169 13852
rect 3016 13812 3022 13824
rect 4157 13821 4169 13824
rect 4203 13852 4215 13855
rect 4246 13852 4252 13864
rect 4203 13824 4252 13852
rect 4203 13821 4215 13824
rect 4157 13815 4215 13821
rect 4246 13812 4252 13824
rect 4304 13812 4310 13864
rect 6641 13855 6699 13861
rect 6641 13821 6653 13855
rect 6687 13852 6699 13855
rect 6687 13824 6868 13852
rect 6687 13821 6699 13824
rect 6641 13815 6699 13821
rect 3234 13784 3240 13796
rect 3195 13756 3240 13784
rect 3234 13744 3240 13756
rect 3292 13744 3298 13796
rect 4522 13744 4528 13796
rect 4580 13784 4586 13796
rect 4706 13784 4712 13796
rect 4580 13756 4712 13784
rect 4580 13744 4586 13756
rect 4706 13744 4712 13756
rect 4764 13744 4770 13796
rect 6840 13784 6868 13824
rect 7190 13812 7196 13864
rect 7248 13852 7254 13864
rect 7285 13855 7343 13861
rect 7285 13852 7297 13855
rect 7248 13824 7297 13852
rect 7248 13812 7254 13824
rect 7285 13821 7297 13824
rect 7331 13852 7343 13855
rect 7834 13852 7840 13864
rect 7331 13824 7840 13852
rect 7331 13821 7343 13824
rect 7285 13815 7343 13821
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 8297 13855 8355 13861
rect 8297 13821 8309 13855
rect 8343 13852 8355 13855
rect 8386 13852 8392 13864
rect 8343 13824 8392 13852
rect 8343 13821 8355 13824
rect 8297 13815 8355 13821
rect 8386 13812 8392 13824
rect 8444 13852 8450 13864
rect 8846 13852 8852 13864
rect 8444 13824 8852 13852
rect 8444 13812 8450 13824
rect 8846 13812 8852 13824
rect 8904 13812 8910 13864
rect 9416 13852 9444 14019
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 9950 14056 9956 14068
rect 9911 14028 9956 14056
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 11054 14056 11060 14068
rect 11015 14028 11060 14056
rect 11054 14016 11060 14028
rect 11112 14016 11118 14068
rect 13265 14059 13323 14065
rect 13265 14025 13277 14059
rect 13311 14056 13323 14059
rect 14182 14056 14188 14068
rect 13311 14028 14188 14056
rect 13311 14025 13323 14028
rect 13265 14019 13323 14025
rect 14182 14016 14188 14028
rect 14240 14056 14246 14068
rect 14642 14056 14648 14068
rect 14240 14028 14648 14056
rect 14240 14016 14246 14028
rect 14642 14016 14648 14028
rect 14700 14016 14706 14068
rect 9784 13852 9812 14016
rect 9858 13948 9864 14000
rect 9916 13988 9922 14000
rect 11333 13991 11391 13997
rect 11333 13988 11345 13991
rect 9916 13960 11345 13988
rect 9916 13948 9922 13960
rect 11333 13957 11345 13960
rect 11379 13957 11391 13991
rect 11333 13951 11391 13957
rect 12710 13948 12716 14000
rect 12768 13988 12774 14000
rect 12805 13991 12863 13997
rect 12805 13988 12817 13991
rect 12768 13960 12817 13988
rect 12768 13948 12774 13960
rect 12805 13957 12817 13960
rect 12851 13988 12863 13991
rect 14366 13988 14372 14000
rect 12851 13960 14372 13988
rect 12851 13957 12863 13960
rect 12805 13951 12863 13957
rect 14366 13948 14372 13960
rect 14424 13948 14430 14000
rect 10042 13880 10048 13932
rect 10100 13920 10106 13932
rect 10505 13923 10563 13929
rect 10505 13920 10517 13923
rect 10100 13892 10517 13920
rect 10100 13880 10106 13892
rect 10505 13889 10517 13892
rect 10551 13920 10563 13923
rect 10686 13920 10692 13932
rect 10551 13892 10692 13920
rect 10551 13889 10563 13892
rect 10505 13883 10563 13889
rect 10686 13880 10692 13892
rect 10744 13880 10750 13932
rect 12250 13920 12256 13932
rect 12211 13892 12256 13920
rect 12250 13880 12256 13892
rect 12308 13880 12314 13932
rect 13173 13923 13231 13929
rect 13173 13889 13185 13923
rect 13219 13920 13231 13923
rect 13909 13923 13967 13929
rect 13909 13920 13921 13923
rect 13219 13892 13921 13920
rect 13219 13889 13231 13892
rect 13173 13883 13231 13889
rect 13909 13889 13921 13892
rect 13955 13920 13967 13923
rect 13955 13892 14964 13920
rect 13955 13889 13967 13892
rect 13909 13883 13967 13889
rect 14936 13864 14964 13892
rect 10413 13855 10471 13861
rect 10413 13852 10425 13855
rect 9416 13824 9628 13852
rect 9784 13824 10425 13852
rect 8662 13784 8668 13796
rect 6840 13756 8668 13784
rect 5534 13716 5540 13728
rect 2372 13688 2728 13716
rect 5495 13688 5540 13716
rect 2372 13676 2378 13688
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 7208 13725 7236 13756
rect 8662 13744 8668 13756
rect 8720 13744 8726 13796
rect 9600 13784 9628 13824
rect 10413 13821 10425 13824
rect 10459 13821 10471 13855
rect 14277 13855 14335 13861
rect 14277 13852 14289 13855
rect 10413 13815 10471 13821
rect 13740 13824 14289 13852
rect 10321 13787 10379 13793
rect 10321 13784 10333 13787
rect 9600 13756 10333 13784
rect 10321 13753 10333 13756
rect 10367 13753 10379 13787
rect 13740 13784 13768 13824
rect 14277 13821 14289 13824
rect 14323 13821 14335 13855
rect 14277 13815 14335 13821
rect 14366 13812 14372 13864
rect 14424 13852 14430 13864
rect 14737 13855 14795 13861
rect 14737 13852 14749 13855
rect 14424 13824 14749 13852
rect 14424 13812 14430 13824
rect 14737 13821 14749 13824
rect 14783 13852 14795 13855
rect 14829 13855 14887 13861
rect 14829 13852 14841 13855
rect 14783 13824 14841 13852
rect 14783 13821 14795 13824
rect 14737 13815 14795 13821
rect 14829 13821 14841 13824
rect 14875 13821 14887 13855
rect 14829 13815 14887 13821
rect 10321 13747 10379 13753
rect 13648 13756 13768 13784
rect 14844 13784 14872 13815
rect 14918 13812 14924 13864
rect 14976 13852 14982 13864
rect 15096 13855 15154 13861
rect 15096 13852 15108 13855
rect 14976 13824 15108 13852
rect 14976 13812 14982 13824
rect 15096 13821 15108 13824
rect 15142 13852 15154 13855
rect 15378 13852 15384 13864
rect 15142 13824 15384 13852
rect 15142 13821 15154 13824
rect 15096 13815 15154 13821
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 16850 13852 16856 13864
rect 16811 13824 16856 13852
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 17218 13852 17224 13864
rect 17179 13824 17224 13852
rect 17218 13812 17224 13824
rect 17276 13812 17282 13864
rect 15286 13784 15292 13796
rect 14844 13756 15292 13784
rect 13648 13728 13676 13756
rect 15286 13744 15292 13756
rect 15344 13744 15350 13796
rect 7193 13719 7251 13725
rect 7193 13685 7205 13719
rect 7239 13685 7251 13719
rect 7193 13679 7251 13685
rect 8386 13676 8392 13728
rect 8444 13716 8450 13728
rect 8757 13719 8815 13725
rect 8757 13716 8769 13719
rect 8444 13688 8769 13716
rect 8444 13676 8450 13688
rect 8757 13685 8769 13688
rect 8803 13685 8815 13719
rect 13630 13716 13636 13728
rect 13591 13688 13636 13716
rect 8757 13679 8815 13685
rect 13630 13676 13636 13688
rect 13688 13676 13694 13728
rect 13722 13676 13728 13728
rect 13780 13716 13786 13728
rect 13780 13688 13825 13716
rect 13780 13676 13786 13688
rect 15378 13676 15384 13728
rect 15436 13716 15442 13728
rect 15562 13716 15568 13728
rect 15436 13688 15568 13716
rect 15436 13676 15442 13688
rect 15562 13676 15568 13688
rect 15620 13676 15626 13728
rect 16206 13716 16212 13728
rect 16167 13688 16212 13716
rect 16206 13676 16212 13688
rect 16264 13676 16270 13728
rect 17681 13719 17739 13725
rect 17681 13685 17693 13719
rect 17727 13716 17739 13719
rect 17862 13716 17868 13728
rect 17727 13688 17868 13716
rect 17727 13685 17739 13688
rect 17681 13679 17739 13685
rect 17862 13676 17868 13688
rect 17920 13676 17926 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1581 13515 1639 13521
rect 1581 13481 1593 13515
rect 1627 13512 1639 13515
rect 1854 13512 1860 13524
rect 1627 13484 1860 13512
rect 1627 13481 1639 13484
rect 1581 13475 1639 13481
rect 1854 13472 1860 13484
rect 1912 13472 1918 13524
rect 2130 13472 2136 13524
rect 2188 13512 2194 13524
rect 2225 13515 2283 13521
rect 2225 13512 2237 13515
rect 2188 13484 2237 13512
rect 2188 13472 2194 13484
rect 2225 13481 2237 13484
rect 2271 13481 2283 13515
rect 2225 13475 2283 13481
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 4065 13515 4123 13521
rect 4065 13512 4077 13515
rect 2832 13484 2877 13512
rect 3436 13484 4077 13512
rect 2832 13472 2838 13484
rect 3436 13456 3464 13484
rect 4065 13481 4077 13484
rect 4111 13481 4123 13515
rect 4065 13475 4123 13481
rect 4154 13472 4160 13524
rect 4212 13512 4218 13524
rect 4433 13515 4491 13521
rect 4433 13512 4445 13515
rect 4212 13484 4445 13512
rect 4212 13472 4218 13484
rect 4433 13481 4445 13484
rect 4479 13481 4491 13515
rect 4433 13475 4491 13481
rect 2869 13447 2927 13453
rect 2869 13413 2881 13447
rect 2915 13444 2927 13447
rect 3418 13444 3424 13456
rect 2915 13416 3424 13444
rect 2915 13413 2927 13416
rect 2869 13407 2927 13413
rect 3418 13404 3424 13416
rect 3476 13404 3482 13456
rect 3878 13444 3884 13456
rect 3839 13416 3884 13444
rect 3878 13404 3884 13416
rect 3936 13404 3942 13456
rect 4448 13444 4476 13475
rect 4522 13472 4528 13524
rect 4580 13512 4586 13524
rect 5997 13515 6055 13521
rect 5997 13512 6009 13515
rect 4580 13484 6009 13512
rect 4580 13472 4586 13484
rect 5997 13481 6009 13484
rect 6043 13481 6055 13515
rect 5997 13475 6055 13481
rect 6546 13472 6552 13524
rect 6604 13512 6610 13524
rect 6641 13515 6699 13521
rect 6641 13512 6653 13515
rect 6604 13484 6653 13512
rect 6604 13472 6610 13484
rect 6641 13481 6653 13484
rect 6687 13481 6699 13515
rect 7190 13512 7196 13524
rect 7151 13484 7196 13512
rect 6641 13475 6699 13481
rect 6089 13447 6147 13453
rect 6089 13444 6101 13447
rect 4448 13416 6101 13444
rect 6089 13413 6101 13416
rect 6135 13444 6147 13447
rect 6178 13444 6184 13456
rect 6135 13416 6184 13444
rect 6135 13413 6147 13416
rect 6089 13407 6147 13413
rect 6178 13404 6184 13416
rect 6236 13404 6242 13456
rect 6656 13444 6684 13475
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 7466 13472 7472 13524
rect 7524 13512 7530 13524
rect 7653 13515 7711 13521
rect 7653 13512 7665 13515
rect 7524 13484 7665 13512
rect 7524 13472 7530 13484
rect 7653 13481 7665 13484
rect 7699 13512 7711 13515
rect 8570 13512 8576 13524
rect 7699 13484 8576 13512
rect 7699 13481 7711 13484
rect 7653 13475 7711 13481
rect 8570 13472 8576 13484
rect 8628 13472 8634 13524
rect 9398 13512 9404 13524
rect 9359 13484 9404 13512
rect 9398 13472 9404 13484
rect 9456 13512 9462 13524
rect 10045 13515 10103 13521
rect 10045 13512 10057 13515
rect 9456 13484 10057 13512
rect 9456 13472 9462 13484
rect 10045 13481 10057 13484
rect 10091 13481 10103 13515
rect 10686 13512 10692 13524
rect 10647 13484 10692 13512
rect 10045 13475 10103 13481
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 11241 13515 11299 13521
rect 11241 13481 11253 13515
rect 11287 13512 11299 13515
rect 11330 13512 11336 13524
rect 11287 13484 11336 13512
rect 11287 13481 11299 13484
rect 11241 13475 11299 13481
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 11514 13472 11520 13524
rect 11572 13512 11578 13524
rect 11701 13515 11759 13521
rect 11701 13512 11713 13515
rect 11572 13484 11713 13512
rect 11572 13472 11578 13484
rect 11701 13481 11713 13484
rect 11747 13481 11759 13515
rect 11701 13475 11759 13481
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 12710 13512 12716 13524
rect 12492 13484 12716 13512
rect 12492 13472 12498 13484
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 13170 13512 13176 13524
rect 13131 13484 13176 13512
rect 13170 13472 13176 13484
rect 13228 13472 13234 13524
rect 13446 13472 13452 13524
rect 13504 13512 13510 13524
rect 13541 13515 13599 13521
rect 13541 13512 13553 13515
rect 13504 13484 13553 13512
rect 13504 13472 13510 13484
rect 13541 13481 13553 13484
rect 13587 13512 13599 13515
rect 13722 13512 13728 13524
rect 13587 13484 13728 13512
rect 13587 13481 13599 13484
rect 13541 13475 13599 13481
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 13998 13512 14004 13524
rect 13959 13484 14004 13512
rect 13998 13472 14004 13484
rect 14056 13472 14062 13524
rect 14918 13512 14924 13524
rect 14879 13484 14924 13512
rect 14918 13472 14924 13484
rect 14976 13472 14982 13524
rect 16298 13512 16304 13524
rect 16259 13484 16304 13512
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 6656 13416 7696 13444
rect 1394 13376 1400 13388
rect 1355 13348 1400 13376
rect 1394 13336 1400 13348
rect 1452 13336 1458 13388
rect 1946 13376 1952 13388
rect 1859 13348 1952 13376
rect 1946 13336 1952 13348
rect 2004 13376 2010 13388
rect 4525 13379 4583 13385
rect 2004 13348 3740 13376
rect 2004 13336 2010 13348
rect 2961 13311 3019 13317
rect 2961 13277 2973 13311
rect 3007 13277 3019 13311
rect 3712 13308 3740 13348
rect 4525 13345 4537 13379
rect 4571 13376 4583 13379
rect 4798 13376 4804 13388
rect 4571 13348 4804 13376
rect 4571 13345 4583 13348
rect 4525 13339 4583 13345
rect 4798 13336 4804 13348
rect 4856 13336 4862 13388
rect 7101 13379 7159 13385
rect 7101 13345 7113 13379
rect 7147 13376 7159 13379
rect 7374 13376 7380 13388
rect 7147 13348 7380 13376
rect 7147 13345 7159 13348
rect 7101 13339 7159 13345
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 7558 13376 7564 13388
rect 7519 13348 7564 13376
rect 7558 13336 7564 13348
rect 7616 13336 7622 13388
rect 7668 13376 7696 13416
rect 15562 13404 15568 13456
rect 15620 13444 15626 13456
rect 16206 13444 16212 13456
rect 15620 13416 16212 13444
rect 15620 13404 15626 13416
rect 16206 13404 16212 13416
rect 16264 13404 16270 13456
rect 18230 13453 18236 13456
rect 18224 13444 18236 13453
rect 18191 13416 18236 13444
rect 18224 13407 18236 13416
rect 18230 13404 18236 13407
rect 18288 13404 18294 13456
rect 11606 13376 11612 13388
rect 7668 13348 7788 13376
rect 11567 13348 11612 13376
rect 4706 13308 4712 13320
rect 3712 13280 4712 13308
rect 2961 13271 3019 13277
rect 2130 13200 2136 13252
rect 2188 13240 2194 13252
rect 2976 13240 3004 13271
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 6273 13311 6331 13317
rect 6273 13277 6285 13311
rect 6319 13308 6331 13311
rect 6362 13308 6368 13320
rect 6319 13280 6368 13308
rect 6319 13277 6331 13280
rect 6273 13271 6331 13277
rect 6362 13268 6368 13280
rect 6420 13268 6426 13320
rect 7760 13317 7788 13348
rect 11606 13336 11612 13348
rect 11664 13336 11670 13388
rect 15657 13379 15715 13385
rect 15657 13345 15669 13379
rect 15703 13376 15715 13379
rect 15838 13376 15844 13388
rect 15703 13348 15844 13376
rect 15703 13345 15715 13348
rect 15657 13339 15715 13345
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 17957 13379 18015 13385
rect 17957 13345 17969 13379
rect 18003 13376 18015 13379
rect 18506 13376 18512 13388
rect 18003 13348 18512 13376
rect 18003 13345 18015 13348
rect 17957 13339 18015 13345
rect 18506 13336 18512 13348
rect 18564 13336 18570 13388
rect 7745 13311 7803 13317
rect 7745 13277 7757 13311
rect 7791 13277 7803 13311
rect 7745 13271 7803 13277
rect 10042 13268 10048 13320
rect 10100 13308 10106 13320
rect 10137 13311 10195 13317
rect 10137 13308 10149 13311
rect 10100 13280 10149 13308
rect 10100 13268 10106 13280
rect 10137 13277 10149 13280
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 11790 13308 11796 13320
rect 10367 13280 11796 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 3510 13240 3516 13252
rect 2188 13212 3004 13240
rect 3423 13212 3516 13240
rect 2188 13200 2194 13212
rect 3510 13200 3516 13212
rect 3568 13240 3574 13252
rect 4062 13240 4068 13252
rect 3568 13212 4068 13240
rect 3568 13200 3574 13212
rect 4062 13200 4068 13212
rect 4120 13200 4126 13252
rect 5626 13240 5632 13252
rect 5587 13212 5632 13240
rect 5626 13200 5632 13212
rect 5684 13200 5690 13252
rect 9030 13200 9036 13252
rect 9088 13240 9094 13252
rect 9125 13243 9183 13249
rect 9125 13240 9137 13243
rect 9088 13212 9137 13240
rect 9088 13200 9094 13212
rect 9125 13209 9137 13212
rect 9171 13240 9183 13243
rect 10336 13240 10364 13271
rect 11790 13268 11796 13280
rect 11848 13268 11854 13320
rect 11885 13311 11943 13317
rect 11885 13277 11897 13311
rect 11931 13308 11943 13311
rect 11974 13308 11980 13320
rect 11931 13280 11980 13308
rect 11931 13277 11943 13280
rect 11885 13271 11943 13277
rect 11974 13268 11980 13280
rect 12032 13268 12038 13320
rect 14090 13308 14096 13320
rect 14051 13280 14096 13308
rect 14090 13268 14096 13280
rect 14148 13268 14154 13320
rect 14274 13308 14280 13320
rect 14235 13280 14280 13308
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 15749 13311 15807 13317
rect 15749 13277 15761 13311
rect 15795 13277 15807 13311
rect 15930 13308 15936 13320
rect 15891 13280 15936 13308
rect 15749 13271 15807 13277
rect 9171 13212 10364 13240
rect 13633 13243 13691 13249
rect 9171 13209 9183 13212
rect 9125 13203 9183 13209
rect 13633 13209 13645 13243
rect 13679 13240 13691 13243
rect 15764 13240 15792 13271
rect 15930 13268 15936 13280
rect 15988 13268 15994 13320
rect 16666 13308 16672 13320
rect 16627 13280 16672 13308
rect 16666 13268 16672 13280
rect 16724 13268 16730 13320
rect 17402 13240 17408 13252
rect 13679 13212 17408 13240
rect 13679 13209 13691 13212
rect 13633 13203 13691 13209
rect 17402 13200 17408 13212
rect 17460 13200 17466 13252
rect 2409 13175 2467 13181
rect 2409 13141 2421 13175
rect 2455 13172 2467 13175
rect 2590 13172 2596 13184
rect 2455 13144 2596 13172
rect 2455 13141 2467 13144
rect 2409 13135 2467 13141
rect 2590 13132 2596 13144
rect 2648 13132 2654 13184
rect 3142 13132 3148 13184
rect 3200 13172 3206 13184
rect 5261 13175 5319 13181
rect 5261 13172 5273 13175
rect 3200 13144 5273 13172
rect 3200 13132 3206 13144
rect 5261 13141 5273 13144
rect 5307 13172 5319 13175
rect 5534 13172 5540 13184
rect 5307 13144 5540 13172
rect 5307 13141 5319 13144
rect 5261 13135 5319 13141
rect 5534 13132 5540 13144
rect 5592 13172 5598 13184
rect 6822 13172 6828 13184
rect 5592 13144 6828 13172
rect 5592 13132 5598 13144
rect 6822 13132 6828 13144
rect 6880 13132 6886 13184
rect 8386 13172 8392 13184
rect 8347 13144 8392 13172
rect 8386 13132 8392 13144
rect 8444 13132 8450 13184
rect 8478 13132 8484 13184
rect 8536 13172 8542 13184
rect 9677 13175 9735 13181
rect 9677 13172 9689 13175
rect 8536 13144 9689 13172
rect 8536 13132 8542 13144
rect 9677 13141 9689 13144
rect 9723 13141 9735 13175
rect 9677 13135 9735 13141
rect 9858 13132 9864 13184
rect 9916 13172 9922 13184
rect 10870 13172 10876 13184
rect 9916 13144 10876 13172
rect 9916 13132 9922 13144
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 10962 13132 10968 13184
rect 11020 13172 11026 13184
rect 11057 13175 11115 13181
rect 11057 13172 11069 13175
rect 11020 13144 11069 13172
rect 11020 13132 11026 13144
rect 11057 13141 11069 13144
rect 11103 13141 11115 13175
rect 11057 13135 11115 13141
rect 12434 13132 12440 13184
rect 12492 13172 12498 13184
rect 12805 13175 12863 13181
rect 12492 13144 12537 13172
rect 12492 13132 12498 13144
rect 12805 13141 12817 13175
rect 12851 13172 12863 13175
rect 13354 13172 13360 13184
rect 12851 13144 13360 13172
rect 12851 13141 12863 13144
rect 12805 13135 12863 13141
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 15289 13175 15347 13181
rect 15289 13141 15301 13175
rect 15335 13172 15347 13175
rect 16022 13172 16028 13184
rect 15335 13144 16028 13172
rect 15335 13141 15347 13144
rect 15289 13135 15347 13141
rect 16022 13132 16028 13144
rect 16080 13132 16086 13184
rect 19334 13172 19340 13184
rect 19295 13144 19340 13172
rect 19334 13132 19340 13144
rect 19392 13132 19398 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1949 12971 2007 12977
rect 1949 12937 1961 12971
rect 1995 12968 2007 12971
rect 2314 12968 2320 12980
rect 1995 12940 2320 12968
rect 1995 12937 2007 12940
rect 1949 12931 2007 12937
rect 2056 12841 2084 12940
rect 2314 12928 2320 12940
rect 2372 12928 2378 12980
rect 4522 12928 4528 12980
rect 4580 12968 4586 12980
rect 4985 12971 5043 12977
rect 4985 12968 4997 12971
rect 4580 12940 4997 12968
rect 4580 12928 4586 12940
rect 4985 12937 4997 12940
rect 5031 12937 5043 12971
rect 5166 12968 5172 12980
rect 5127 12940 5172 12968
rect 4985 12931 5043 12937
rect 4157 12903 4215 12909
rect 4157 12869 4169 12903
rect 4203 12900 4215 12903
rect 4798 12900 4804 12912
rect 4203 12872 4804 12900
rect 4203 12869 4215 12872
rect 4157 12863 4215 12869
rect 4798 12860 4804 12872
rect 4856 12860 4862 12912
rect 5000 12900 5028 12931
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 6178 12968 6184 12980
rect 6139 12940 6184 12968
rect 6178 12928 6184 12940
rect 6236 12928 6242 12980
rect 6546 12968 6552 12980
rect 6507 12940 6552 12968
rect 6546 12928 6552 12940
rect 6604 12928 6610 12980
rect 7558 12928 7564 12980
rect 7616 12968 7622 12980
rect 7837 12971 7895 12977
rect 7837 12968 7849 12971
rect 7616 12940 7849 12968
rect 7616 12928 7622 12940
rect 7837 12937 7849 12940
rect 7883 12968 7895 12971
rect 7926 12968 7932 12980
rect 7883 12940 7932 12968
rect 7883 12937 7895 12940
rect 7837 12931 7895 12937
rect 7926 12928 7932 12940
rect 7984 12928 7990 12980
rect 8297 12971 8355 12977
rect 8297 12937 8309 12971
rect 8343 12968 8355 12971
rect 8386 12968 8392 12980
rect 8343 12940 8392 12968
rect 8343 12937 8355 12940
rect 8297 12931 8355 12937
rect 8386 12928 8392 12940
rect 8444 12928 8450 12980
rect 8941 12971 8999 12977
rect 8941 12937 8953 12971
rect 8987 12968 8999 12971
rect 9214 12968 9220 12980
rect 8987 12940 9220 12968
rect 8987 12937 8999 12940
rect 8941 12931 8999 12937
rect 6362 12900 6368 12912
rect 5000 12872 6368 12900
rect 6362 12860 6368 12872
rect 6420 12860 6426 12912
rect 2041 12835 2099 12841
rect 2041 12801 2053 12835
rect 2087 12801 2099 12835
rect 5718 12832 5724 12844
rect 5679 12804 5724 12832
rect 2041 12795 2099 12801
rect 2056 12628 2084 12795
rect 5718 12792 5724 12804
rect 5776 12792 5782 12844
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 6914 12832 6920 12844
rect 6604 12804 6920 12832
rect 6604 12792 6610 12804
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 7466 12832 7472 12844
rect 7427 12804 7472 12832
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 9048 12841 9076 12940
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 11238 12928 11244 12980
rect 11296 12968 11302 12980
rect 11333 12971 11391 12977
rect 11333 12968 11345 12971
rect 11296 12940 11345 12968
rect 11296 12928 11302 12940
rect 11333 12937 11345 12940
rect 11379 12968 11391 12971
rect 11606 12968 11612 12980
rect 11379 12940 11612 12968
rect 11379 12937 11391 12940
rect 11333 12931 11391 12937
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 11974 12968 11980 12980
rect 11935 12940 11980 12968
rect 11974 12928 11980 12940
rect 12032 12928 12038 12980
rect 12437 12971 12495 12977
rect 12437 12937 12449 12971
rect 12483 12968 12495 12971
rect 13630 12968 13636 12980
rect 12483 12940 13636 12968
rect 12483 12937 12495 12940
rect 12437 12931 12495 12937
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 13998 12968 14004 12980
rect 13959 12940 14004 12968
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 14642 12928 14648 12980
rect 14700 12968 14706 12980
rect 15013 12971 15071 12977
rect 15013 12968 15025 12971
rect 14700 12940 15025 12968
rect 14700 12928 14706 12940
rect 15013 12937 15025 12940
rect 15059 12968 15071 12971
rect 15838 12968 15844 12980
rect 15059 12940 15844 12968
rect 15059 12937 15071 12940
rect 15013 12931 15071 12937
rect 15838 12928 15844 12940
rect 15896 12928 15902 12980
rect 17402 12968 17408 12980
rect 17363 12940 17408 12968
rect 17402 12928 17408 12940
rect 17460 12928 17466 12980
rect 18230 12968 18236 12980
rect 18191 12940 18236 12968
rect 18230 12928 18236 12940
rect 18288 12928 18294 12980
rect 18506 12928 18512 12980
rect 18564 12968 18570 12980
rect 18601 12971 18659 12977
rect 18601 12968 18613 12971
rect 18564 12940 18613 12968
rect 18564 12928 18570 12940
rect 18601 12937 18613 12940
rect 18647 12937 18659 12971
rect 18601 12931 18659 12937
rect 12894 12860 12900 12912
rect 12952 12900 12958 12912
rect 12952 12872 13400 12900
rect 12952 12860 12958 12872
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12801 9091 12835
rect 9033 12795 9091 12801
rect 11514 12792 11520 12844
rect 11572 12832 11578 12844
rect 11609 12835 11667 12841
rect 11609 12832 11621 12835
rect 11572 12804 11621 12832
rect 11572 12792 11578 12804
rect 11609 12801 11621 12804
rect 11655 12801 11667 12835
rect 11609 12795 11667 12801
rect 13081 12835 13139 12841
rect 13081 12801 13093 12835
rect 13127 12832 13139 12835
rect 13170 12832 13176 12844
rect 13127 12804 13176 12832
rect 13127 12801 13139 12804
rect 13081 12795 13139 12801
rect 13170 12792 13176 12804
rect 13228 12792 13234 12844
rect 2130 12724 2136 12776
rect 2188 12764 2194 12776
rect 2297 12767 2355 12773
rect 2297 12764 2309 12767
rect 2188 12736 2309 12764
rect 2188 12724 2194 12736
rect 2297 12733 2309 12736
rect 2343 12764 2355 12767
rect 2343 12736 2452 12764
rect 2343 12733 2355 12736
rect 2297 12727 2355 12733
rect 2424 12696 2452 12736
rect 4154 12724 4160 12776
rect 4212 12764 4218 12776
rect 4433 12767 4491 12773
rect 4433 12764 4445 12767
rect 4212 12736 4445 12764
rect 4212 12724 4218 12736
rect 4433 12733 4445 12736
rect 4479 12733 4491 12767
rect 7190 12764 7196 12776
rect 7151 12736 7196 12764
rect 4433 12727 4491 12733
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 12492 12736 12817 12764
rect 12492 12724 12498 12736
rect 12805 12733 12817 12736
rect 12851 12764 12863 12767
rect 12894 12764 12900 12776
rect 12851 12736 12900 12764
rect 12851 12733 12863 12736
rect 12805 12727 12863 12733
rect 12894 12724 12900 12736
rect 12952 12724 12958 12776
rect 2774 12696 2780 12708
rect 2424 12668 2780 12696
rect 2774 12656 2780 12668
rect 2832 12656 2838 12708
rect 5644 12668 6868 12696
rect 5644 12640 5672 12668
rect 2130 12628 2136 12640
rect 2056 12600 2136 12628
rect 2130 12588 2136 12600
rect 2188 12588 2194 12640
rect 3418 12628 3424 12640
rect 3379 12600 3424 12628
rect 3418 12588 3424 12600
rect 3476 12588 3482 12640
rect 5534 12628 5540 12640
rect 5495 12600 5540 12628
rect 5534 12588 5540 12600
rect 5592 12588 5598 12640
rect 5626 12588 5632 12640
rect 5684 12628 5690 12640
rect 6840 12637 6868 12668
rect 9030 12656 9036 12708
rect 9088 12696 9094 12708
rect 9278 12699 9336 12705
rect 9278 12696 9290 12699
rect 9088 12668 9290 12696
rect 9088 12656 9094 12668
rect 9278 12665 9290 12668
rect 9324 12665 9336 12699
rect 9278 12659 9336 12665
rect 12710 12656 12716 12708
rect 12768 12696 12774 12708
rect 13170 12696 13176 12708
rect 12768 12668 13176 12696
rect 12768 12656 12774 12668
rect 13170 12656 13176 12668
rect 13228 12656 13234 12708
rect 13372 12696 13400 12872
rect 14274 12792 14280 12844
rect 14332 12832 14338 12844
rect 14461 12835 14519 12841
rect 14461 12832 14473 12835
rect 14332 12804 14473 12832
rect 14332 12792 14338 12804
rect 14461 12801 14473 12804
rect 14507 12832 14519 12835
rect 14507 12804 15608 12832
rect 14507 12801 14519 12804
rect 14461 12795 14519 12801
rect 15580 12776 15608 12804
rect 17954 12792 17960 12844
rect 18012 12832 18018 12844
rect 18230 12832 18236 12844
rect 18012 12804 18236 12832
rect 18012 12792 18018 12804
rect 18230 12792 18236 12804
rect 18288 12792 18294 12844
rect 13630 12764 13636 12776
rect 13591 12736 13636 12764
rect 13630 12724 13636 12736
rect 13688 12764 13694 12776
rect 14090 12764 14096 12776
rect 13688 12736 14096 12764
rect 13688 12724 13694 12736
rect 14090 12724 14096 12736
rect 14148 12724 14154 12776
rect 15286 12724 15292 12776
rect 15344 12764 15350 12776
rect 15381 12767 15439 12773
rect 15381 12764 15393 12767
rect 15344 12736 15393 12764
rect 15344 12724 15350 12736
rect 15381 12733 15393 12736
rect 15427 12764 15439 12767
rect 15473 12767 15531 12773
rect 15473 12764 15485 12767
rect 15427 12736 15485 12764
rect 15427 12733 15439 12736
rect 15381 12727 15439 12733
rect 15473 12733 15485 12736
rect 15519 12733 15531 12767
rect 15473 12727 15531 12733
rect 15488 12696 15516 12727
rect 15562 12724 15568 12776
rect 15620 12764 15626 12776
rect 15740 12767 15798 12773
rect 15740 12764 15752 12767
rect 15620 12736 15752 12764
rect 15620 12724 15626 12736
rect 15740 12733 15752 12736
rect 15786 12733 15798 12767
rect 15740 12727 15798 12733
rect 15654 12696 15660 12708
rect 13372 12668 13676 12696
rect 15488 12668 15660 12696
rect 13648 12640 13676 12668
rect 15654 12656 15660 12668
rect 15712 12656 15718 12708
rect 6825 12631 6883 12637
rect 5684 12600 5729 12628
rect 5684 12588 5690 12600
rect 6825 12597 6837 12631
rect 6871 12597 6883 12631
rect 6825 12591 6883 12597
rect 7282 12588 7288 12640
rect 7340 12628 7346 12640
rect 7340 12600 7385 12628
rect 7340 12588 7346 12600
rect 9950 12588 9956 12640
rect 10008 12628 10014 12640
rect 10413 12631 10471 12637
rect 10413 12628 10425 12631
rect 10008 12600 10425 12628
rect 10008 12588 10014 12600
rect 10413 12597 10425 12600
rect 10459 12597 10471 12631
rect 10413 12591 10471 12597
rect 12526 12588 12532 12640
rect 12584 12628 12590 12640
rect 12897 12631 12955 12637
rect 12897 12628 12909 12631
rect 12584 12600 12909 12628
rect 12584 12588 12590 12600
rect 12897 12597 12909 12600
rect 12943 12628 12955 12631
rect 13538 12628 13544 12640
rect 12943 12600 13544 12628
rect 12943 12597 12955 12600
rect 12897 12591 12955 12597
rect 13538 12588 13544 12600
rect 13596 12588 13602 12640
rect 13630 12588 13636 12640
rect 13688 12588 13694 12640
rect 16850 12628 16856 12640
rect 16811 12600 16856 12628
rect 16850 12588 16856 12600
rect 16908 12588 16914 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 3694 12424 3700 12436
rect 3655 12396 3700 12424
rect 3694 12384 3700 12396
rect 3752 12384 3758 12436
rect 5261 12427 5319 12433
rect 5261 12393 5273 12427
rect 5307 12424 5319 12427
rect 5718 12424 5724 12436
rect 5307 12396 5724 12424
rect 5307 12393 5319 12396
rect 5261 12387 5319 12393
rect 5718 12384 5724 12396
rect 5776 12424 5782 12436
rect 6178 12424 6184 12436
rect 5776 12396 6184 12424
rect 5776 12384 5782 12396
rect 6178 12384 6184 12396
rect 6236 12384 6242 12436
rect 6454 12384 6460 12436
rect 6512 12424 6518 12436
rect 6546 12424 6552 12436
rect 6512 12396 6552 12424
rect 6512 12384 6518 12396
rect 6546 12384 6552 12396
rect 6604 12384 6610 12436
rect 7374 12424 7380 12436
rect 7335 12396 7380 12424
rect 7374 12384 7380 12396
rect 7432 12384 7438 12436
rect 7466 12384 7472 12436
rect 7524 12424 7530 12436
rect 7653 12427 7711 12433
rect 7653 12424 7665 12427
rect 7524 12396 7665 12424
rect 7524 12384 7530 12396
rect 7653 12393 7665 12396
rect 7699 12393 7711 12427
rect 7653 12387 7711 12393
rect 8297 12427 8355 12433
rect 8297 12393 8309 12427
rect 8343 12424 8355 12427
rect 8478 12424 8484 12436
rect 8343 12396 8484 12424
rect 8343 12393 8355 12396
rect 8297 12387 8355 12393
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 9030 12424 9036 12436
rect 8991 12396 9036 12424
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 9398 12424 9404 12436
rect 9359 12396 9404 12424
rect 9398 12384 9404 12396
rect 9456 12384 9462 12436
rect 9677 12427 9735 12433
rect 9677 12393 9689 12427
rect 9723 12424 9735 12427
rect 9858 12424 9864 12436
rect 9723 12396 9864 12424
rect 9723 12393 9735 12396
rect 9677 12387 9735 12393
rect 9858 12384 9864 12396
rect 9916 12384 9922 12436
rect 12342 12384 12348 12436
rect 12400 12424 12406 12436
rect 12526 12424 12532 12436
rect 12400 12396 12532 12424
rect 12400 12384 12406 12396
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 13170 12424 13176 12436
rect 13131 12396 13176 12424
rect 13170 12384 13176 12396
rect 13228 12384 13234 12436
rect 13354 12384 13360 12436
rect 13412 12424 13418 12436
rect 13906 12424 13912 12436
rect 13412 12396 13912 12424
rect 13412 12384 13418 12396
rect 13906 12384 13912 12396
rect 13964 12384 13970 12436
rect 15562 12424 15568 12436
rect 15523 12396 15568 12424
rect 15562 12384 15568 12396
rect 15620 12384 15626 12436
rect 16301 12427 16359 12433
rect 16301 12393 16313 12427
rect 16347 12424 16359 12427
rect 16482 12424 16488 12436
rect 16347 12396 16488 12424
rect 16347 12393 16359 12396
rect 16301 12387 16359 12393
rect 16482 12384 16488 12396
rect 16540 12384 16546 12436
rect 1664 12359 1722 12365
rect 1664 12325 1676 12359
rect 1710 12356 1722 12359
rect 1946 12356 1952 12368
rect 1710 12328 1952 12356
rect 1710 12325 1722 12328
rect 1664 12319 1722 12325
rect 1946 12316 1952 12328
rect 2004 12316 2010 12368
rect 10045 12359 10103 12365
rect 10045 12325 10057 12359
rect 10091 12356 10103 12359
rect 10870 12356 10876 12368
rect 10091 12328 10876 12356
rect 10091 12325 10103 12328
rect 10045 12319 10103 12325
rect 10870 12316 10876 12328
rect 10928 12316 10934 12368
rect 13265 12359 13323 12365
rect 13265 12325 13277 12359
rect 13311 12356 13323 12359
rect 14277 12359 14335 12365
rect 14277 12356 14289 12359
rect 13311 12328 14289 12356
rect 13311 12325 13323 12328
rect 13265 12319 13323 12325
rect 14277 12325 14289 12328
rect 14323 12356 14335 12359
rect 15470 12356 15476 12368
rect 14323 12328 15476 12356
rect 14323 12325 14335 12328
rect 14277 12319 14335 12325
rect 15470 12316 15476 12328
rect 15528 12316 15534 12368
rect 4065 12291 4123 12297
rect 4065 12257 4077 12291
rect 4111 12288 4123 12291
rect 4798 12288 4804 12300
rect 4111 12260 4804 12288
rect 4111 12257 4123 12260
rect 4065 12251 4123 12257
rect 4798 12248 4804 12260
rect 4856 12248 4862 12300
rect 5442 12248 5448 12300
rect 5500 12288 5506 12300
rect 5609 12291 5667 12297
rect 5609 12288 5621 12291
rect 5500 12260 5621 12288
rect 5500 12248 5506 12260
rect 5609 12257 5621 12260
rect 5655 12288 5667 12291
rect 8202 12288 8208 12300
rect 5655 12260 7604 12288
rect 8163 12260 8208 12288
rect 5655 12257 5667 12260
rect 5609 12251 5667 12257
rect 1397 12223 1455 12229
rect 1397 12189 1409 12223
rect 1443 12189 1455 12223
rect 1397 12183 1455 12189
rect 1412 12084 1440 12183
rect 4246 12180 4252 12232
rect 4304 12220 4310 12232
rect 5350 12220 5356 12232
rect 4304 12192 5356 12220
rect 4304 12180 4310 12192
rect 5350 12180 5356 12192
rect 5408 12180 5414 12232
rect 7576 12220 7604 12260
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 9950 12248 9956 12300
rect 10008 12248 10014 12300
rect 10137 12291 10195 12297
rect 10137 12257 10149 12291
rect 10183 12288 10195 12291
rect 10689 12291 10747 12297
rect 10689 12288 10701 12291
rect 10183 12260 10701 12288
rect 10183 12257 10195 12260
rect 10137 12251 10195 12257
rect 10689 12257 10701 12260
rect 10735 12257 10747 12291
rect 11606 12288 11612 12300
rect 11567 12260 11612 12288
rect 10689 12251 10747 12257
rect 8389 12223 8447 12229
rect 8389 12220 8401 12223
rect 7576 12192 8401 12220
rect 8389 12189 8401 12192
rect 8435 12220 8447 12223
rect 8754 12220 8760 12232
rect 8435 12192 8760 12220
rect 8435 12189 8447 12192
rect 8389 12183 8447 12189
rect 8754 12180 8760 12192
rect 8812 12220 8818 12232
rect 9968 12220 9996 12248
rect 10229 12223 10287 12229
rect 10229 12220 10241 12223
rect 8812 12192 10241 12220
rect 8812 12180 8818 12192
rect 10229 12189 10241 12192
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 6914 12112 6920 12164
rect 6972 12152 6978 12164
rect 7282 12152 7288 12164
rect 6972 12124 7288 12152
rect 6972 12112 6978 12124
rect 7282 12112 7288 12124
rect 7340 12152 7346 12164
rect 7837 12155 7895 12161
rect 7837 12152 7849 12155
rect 7340 12124 7849 12152
rect 7340 12112 7346 12124
rect 7837 12121 7849 12124
rect 7883 12121 7895 12155
rect 10704 12152 10732 12251
rect 11606 12248 11612 12260
rect 11664 12248 11670 12300
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 11756 12260 11801 12288
rect 11756 12248 11762 12260
rect 12342 12248 12348 12300
rect 12400 12288 12406 12300
rect 15013 12291 15071 12297
rect 15013 12288 15025 12291
rect 12400 12260 15025 12288
rect 12400 12248 12406 12260
rect 15013 12257 15025 12260
rect 15059 12288 15071 12291
rect 15562 12288 15568 12300
rect 15059 12260 15568 12288
rect 15059 12257 15071 12260
rect 15013 12251 15071 12257
rect 15562 12248 15568 12260
rect 15620 12248 15626 12300
rect 16206 12288 16212 12300
rect 16167 12260 16212 12288
rect 16206 12248 16212 12260
rect 16264 12248 16270 12300
rect 17494 12248 17500 12300
rect 17552 12288 17558 12300
rect 17773 12291 17831 12297
rect 17773 12288 17785 12291
rect 17552 12260 17785 12288
rect 17552 12248 17558 12260
rect 17773 12257 17785 12260
rect 17819 12257 17831 12291
rect 17773 12251 17831 12257
rect 11882 12220 11888 12232
rect 11843 12192 11888 12220
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 13354 12180 13360 12232
rect 13412 12220 13418 12232
rect 14458 12220 14464 12232
rect 13412 12192 14464 12220
rect 13412 12180 13418 12192
rect 14458 12180 14464 12192
rect 14516 12180 14522 12232
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12220 16451 12223
rect 17865 12223 17923 12229
rect 16439 12192 16473 12220
rect 16439 12189 16451 12192
rect 16393 12183 16451 12189
rect 17865 12189 17877 12223
rect 17911 12189 17923 12223
rect 17865 12183 17923 12189
rect 11241 12155 11299 12161
rect 11241 12152 11253 12155
rect 10704 12124 11253 12152
rect 7837 12115 7895 12121
rect 11241 12121 11253 12124
rect 11287 12121 11299 12155
rect 11241 12115 11299 12121
rect 12805 12155 12863 12161
rect 12805 12121 12817 12155
rect 12851 12152 12863 12155
rect 13446 12152 13452 12164
rect 12851 12124 13452 12152
rect 12851 12121 12863 12124
rect 12805 12115 12863 12121
rect 13446 12112 13452 12124
rect 13504 12112 13510 12164
rect 15654 12112 15660 12164
rect 15712 12152 15718 12164
rect 15930 12152 15936 12164
rect 15712 12124 15936 12152
rect 15712 12112 15718 12124
rect 15930 12112 15936 12124
rect 15988 12152 15994 12164
rect 16408 12152 16436 12183
rect 16850 12152 16856 12164
rect 15988 12124 16856 12152
rect 15988 12112 15994 12124
rect 16850 12112 16856 12124
rect 16908 12112 16914 12164
rect 17770 12112 17776 12164
rect 17828 12152 17834 12164
rect 17880 12152 17908 12183
rect 17954 12180 17960 12232
rect 18012 12220 18018 12232
rect 18785 12223 18843 12229
rect 18785 12220 18797 12223
rect 18012 12192 18797 12220
rect 18012 12180 18018 12192
rect 18785 12189 18797 12192
rect 18831 12189 18843 12223
rect 18785 12183 18843 12189
rect 17828 12124 17908 12152
rect 17828 12112 17834 12124
rect 2130 12084 2136 12096
rect 1412 12056 2136 12084
rect 2130 12044 2136 12056
rect 2188 12044 2194 12096
rect 2774 12044 2780 12096
rect 2832 12084 2838 12096
rect 3421 12087 3479 12093
rect 2832 12056 2877 12084
rect 2832 12044 2838 12056
rect 3421 12053 3433 12087
rect 3467 12084 3479 12087
rect 3970 12084 3976 12096
rect 3467 12056 3976 12084
rect 3467 12053 3479 12056
rect 3421 12047 3479 12053
rect 3970 12044 3976 12056
rect 4028 12044 4034 12096
rect 4246 12084 4252 12096
rect 4207 12056 4252 12084
rect 4246 12044 4252 12056
rect 4304 12044 4310 12096
rect 4706 12084 4712 12096
rect 4619 12056 4712 12084
rect 4706 12044 4712 12056
rect 4764 12084 4770 12096
rect 5994 12084 6000 12096
rect 4764 12056 6000 12084
rect 4764 12044 4770 12056
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6730 12084 6736 12096
rect 6643 12056 6736 12084
rect 6730 12044 6736 12056
rect 6788 12084 6794 12096
rect 7466 12084 7472 12096
rect 6788 12056 7472 12084
rect 6788 12044 6794 12056
rect 7466 12044 7472 12056
rect 7524 12044 7530 12096
rect 9214 12044 9220 12096
rect 9272 12084 9278 12096
rect 9582 12084 9588 12096
rect 9272 12056 9588 12084
rect 9272 12044 9278 12056
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 11057 12087 11115 12093
rect 11057 12084 11069 12087
rect 9732 12056 11069 12084
rect 9732 12044 9738 12056
rect 11057 12053 11069 12056
rect 11103 12053 11115 12087
rect 11057 12047 11115 12053
rect 13354 12044 13360 12096
rect 13412 12084 13418 12096
rect 13817 12087 13875 12093
rect 13817 12084 13829 12087
rect 13412 12056 13829 12084
rect 13412 12044 13418 12056
rect 13817 12053 13829 12056
rect 13863 12053 13875 12087
rect 13817 12047 13875 12053
rect 14737 12087 14795 12093
rect 14737 12053 14749 12087
rect 14783 12084 14795 12087
rect 15672 12084 15700 12112
rect 15838 12084 15844 12096
rect 14783 12056 15700 12084
rect 15799 12056 15844 12084
rect 14783 12053 14795 12056
rect 14737 12047 14795 12053
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 17402 12084 17408 12096
rect 17363 12056 17408 12084
rect 17402 12044 17408 12056
rect 17460 12044 17466 12096
rect 18414 12084 18420 12096
rect 18375 12056 18420 12084
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1578 11880 1584 11892
rect 1539 11852 1584 11880
rect 1578 11840 1584 11852
rect 1636 11840 1642 11892
rect 3970 11880 3976 11892
rect 2332 11852 3976 11880
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 2332 11676 2360 11852
rect 3970 11840 3976 11852
rect 4028 11840 4034 11892
rect 4798 11880 4804 11892
rect 4759 11852 4804 11880
rect 4798 11840 4804 11852
rect 4856 11880 4862 11892
rect 5537 11883 5595 11889
rect 5537 11880 5549 11883
rect 4856 11852 5549 11880
rect 4856 11840 4862 11852
rect 5537 11849 5549 11852
rect 5583 11849 5595 11883
rect 6178 11880 6184 11892
rect 6139 11852 6184 11880
rect 5537 11843 5595 11849
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 8754 11880 8760 11892
rect 8715 11852 8760 11880
rect 8754 11840 8760 11852
rect 8812 11880 8818 11892
rect 9125 11883 9183 11889
rect 9125 11880 9137 11883
rect 8812 11852 9137 11880
rect 8812 11840 8818 11852
rect 9125 11849 9137 11852
rect 9171 11849 9183 11883
rect 9306 11880 9312 11892
rect 9267 11852 9312 11880
rect 9125 11843 9183 11849
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 11241 11883 11299 11889
rect 11241 11849 11253 11883
rect 11287 11880 11299 11883
rect 11698 11880 11704 11892
rect 11287 11852 11704 11880
rect 11287 11849 11299 11852
rect 11241 11843 11299 11849
rect 11698 11840 11704 11852
rect 11756 11840 11762 11892
rect 13906 11880 13912 11892
rect 13867 11852 13912 11880
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 14458 11880 14464 11892
rect 14419 11852 14464 11880
rect 14458 11840 14464 11852
rect 14516 11840 14522 11892
rect 16482 11880 16488 11892
rect 16443 11852 16488 11880
rect 16482 11840 16488 11852
rect 16540 11840 16546 11892
rect 17770 11880 17776 11892
rect 17731 11852 17776 11880
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 19150 11880 19156 11892
rect 18524 11852 19156 11880
rect 5350 11772 5356 11824
rect 5408 11812 5414 11824
rect 5813 11815 5871 11821
rect 5813 11812 5825 11815
rect 5408 11784 5825 11812
rect 5408 11772 5414 11784
rect 5813 11781 5825 11784
rect 5859 11781 5871 11815
rect 5813 11775 5871 11781
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11744 2467 11747
rect 2455 11716 2995 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 1443 11648 2360 11676
rect 2869 11679 2927 11685
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 2869 11645 2881 11679
rect 2915 11645 2927 11679
rect 2967 11676 2995 11716
rect 3136 11679 3194 11685
rect 3136 11676 3148 11679
rect 2967 11648 3148 11676
rect 2869 11639 2927 11645
rect 3136 11645 3148 11648
rect 3182 11676 3194 11679
rect 3418 11676 3424 11688
rect 3182 11648 3424 11676
rect 3182 11645 3194 11648
rect 3136 11639 3194 11645
rect 2884 11608 2912 11639
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 4430 11636 4436 11688
rect 4488 11676 4494 11688
rect 5258 11676 5264 11688
rect 4488 11648 5264 11676
rect 4488 11636 4494 11648
rect 5258 11636 5264 11648
rect 5316 11676 5322 11688
rect 5353 11679 5411 11685
rect 5353 11676 5365 11679
rect 5316 11648 5365 11676
rect 5316 11636 5322 11648
rect 5353 11645 5365 11648
rect 5399 11645 5411 11679
rect 5828 11676 5856 11775
rect 6196 11744 6224 11840
rect 10873 11815 10931 11821
rect 10873 11781 10885 11815
rect 10919 11812 10931 11815
rect 11882 11812 11888 11824
rect 10919 11784 11888 11812
rect 10919 11781 10931 11784
rect 10873 11775 10931 11781
rect 11882 11772 11888 11784
rect 11940 11772 11946 11824
rect 14550 11772 14556 11824
rect 14608 11812 14614 11824
rect 16025 11815 16083 11821
rect 16025 11812 16037 11815
rect 14608 11784 16037 11812
rect 14608 11772 14614 11784
rect 16025 11781 16037 11784
rect 16071 11812 16083 11815
rect 16206 11812 16212 11824
rect 16071 11784 16212 11812
rect 16071 11781 16083 11784
rect 16025 11775 16083 11781
rect 16206 11772 16212 11784
rect 16264 11772 16270 11824
rect 9858 11744 9864 11756
rect 6196 11716 6951 11744
rect 9819 11716 9864 11744
rect 6923 11688 6951 11716
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 15562 11744 15568 11756
rect 13924 11716 15424 11744
rect 15523 11716 15568 11744
rect 6178 11676 6184 11688
rect 5828 11648 6184 11676
rect 5353 11639 5411 11645
rect 6178 11636 6184 11648
rect 6236 11676 6242 11688
rect 6549 11679 6607 11685
rect 6549 11676 6561 11679
rect 6236 11648 6561 11676
rect 6236 11636 6242 11648
rect 6549 11645 6561 11648
rect 6595 11676 6607 11679
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 6595 11648 6837 11676
rect 6595 11645 6607 11648
rect 6549 11639 6607 11645
rect 6825 11645 6837 11648
rect 6871 11645 6883 11679
rect 6825 11639 6883 11645
rect 6914 11636 6920 11688
rect 6972 11676 6978 11688
rect 7081 11679 7139 11685
rect 7081 11676 7093 11679
rect 6972 11648 7093 11676
rect 6972 11636 6978 11648
rect 7081 11645 7093 11648
rect 7127 11645 7139 11679
rect 7081 11639 7139 11645
rect 9674 11636 9680 11688
rect 9732 11676 9738 11688
rect 9769 11679 9827 11685
rect 9769 11676 9781 11679
rect 9732 11648 9781 11676
rect 9732 11636 9738 11648
rect 9769 11645 9781 11648
rect 9815 11645 9827 11679
rect 9769 11639 9827 11645
rect 11606 11636 11612 11688
rect 11664 11676 11670 11688
rect 11793 11679 11851 11685
rect 11793 11676 11805 11679
rect 11664 11648 11805 11676
rect 11664 11636 11670 11648
rect 11793 11645 11805 11648
rect 11839 11645 11851 11679
rect 11793 11639 11851 11645
rect 11882 11636 11888 11688
rect 11940 11676 11946 11688
rect 12161 11679 12219 11685
rect 12161 11676 12173 11679
rect 11940 11648 12173 11676
rect 11940 11636 11946 11648
rect 12161 11645 12173 11648
rect 12207 11676 12219 11679
rect 12529 11679 12587 11685
rect 12529 11676 12541 11679
rect 12207 11648 12541 11676
rect 12207 11645 12219 11648
rect 12161 11639 12219 11645
rect 12529 11645 12541 11648
rect 12575 11645 12587 11679
rect 13924 11676 13952 11716
rect 12529 11639 12587 11645
rect 12820 11648 13952 11676
rect 10042 11608 10048 11620
rect 2700 11580 2912 11608
rect 9692 11580 10048 11608
rect 2041 11543 2099 11549
rect 2041 11509 2053 11543
rect 2087 11540 2099 11543
rect 2130 11540 2136 11552
rect 2087 11512 2136 11540
rect 2087 11509 2099 11512
rect 2041 11503 2099 11509
rect 2130 11500 2136 11512
rect 2188 11540 2194 11552
rect 2700 11549 2728 11580
rect 2685 11543 2743 11549
rect 2685 11540 2697 11543
rect 2188 11512 2697 11540
rect 2188 11500 2194 11512
rect 2685 11509 2697 11512
rect 2731 11509 2743 11543
rect 4246 11540 4252 11552
rect 4207 11512 4252 11540
rect 2685 11503 2743 11509
rect 4246 11500 4252 11512
rect 4304 11500 4310 11552
rect 5261 11543 5319 11549
rect 5261 11509 5273 11543
rect 5307 11540 5319 11543
rect 5442 11540 5448 11552
rect 5307 11512 5448 11540
rect 5307 11509 5319 11512
rect 5261 11503 5319 11509
rect 5442 11500 5448 11512
rect 5500 11500 5506 11552
rect 8202 11540 8208 11552
rect 8163 11512 8208 11540
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 9692 11549 9720 11580
rect 10042 11568 10048 11580
rect 10100 11608 10106 11620
rect 10962 11608 10968 11620
rect 10100 11580 10968 11608
rect 10100 11568 10106 11580
rect 10962 11568 10968 11580
rect 11020 11568 11026 11620
rect 12820 11617 12848 11648
rect 13998 11636 14004 11688
rect 14056 11676 14062 11688
rect 14734 11676 14740 11688
rect 14056 11648 14740 11676
rect 14056 11636 14062 11648
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 15396 11676 15424 11716
rect 15562 11704 15568 11716
rect 15620 11704 15626 11756
rect 18524 11753 18552 11852
rect 19150 11840 19156 11852
rect 19208 11840 19214 11892
rect 18509 11747 18567 11753
rect 18509 11713 18521 11747
rect 18555 11713 18567 11747
rect 18509 11707 18567 11713
rect 18601 11747 18659 11753
rect 18601 11713 18613 11747
rect 18647 11713 18659 11747
rect 18601 11707 18659 11713
rect 17037 11679 17095 11685
rect 17037 11676 17049 11679
rect 15396 11648 17049 11676
rect 17037 11645 17049 11648
rect 17083 11676 17095 11679
rect 17954 11676 17960 11688
rect 17083 11648 17960 11676
rect 17083 11645 17095 11648
rect 17037 11639 17095 11645
rect 17954 11636 17960 11648
rect 18012 11636 18018 11688
rect 18414 11676 18420 11688
rect 18375 11648 18420 11676
rect 18414 11636 18420 11648
rect 18472 11636 18478 11688
rect 12796 11611 12854 11617
rect 12796 11577 12808 11611
rect 12842 11577 12854 11611
rect 15381 11611 15439 11617
rect 15381 11608 15393 11611
rect 12796 11571 12854 11577
rect 14844 11580 15393 11608
rect 9677 11543 9735 11549
rect 9677 11509 9689 11543
rect 9723 11509 9735 11543
rect 9677 11503 9735 11509
rect 10413 11543 10471 11549
rect 10413 11509 10425 11543
rect 10459 11540 10471 11543
rect 10870 11540 10876 11552
rect 10459 11512 10876 11540
rect 10459 11509 10471 11512
rect 10413 11503 10471 11509
rect 10870 11500 10876 11512
rect 10928 11500 10934 11552
rect 11330 11540 11336 11552
rect 11291 11512 11336 11540
rect 11330 11500 11336 11512
rect 11388 11500 11394 11552
rect 12526 11500 12532 11552
rect 12584 11540 12590 11552
rect 12820 11540 12848 11571
rect 12584 11512 12848 11540
rect 12584 11500 12590 11512
rect 14734 11500 14740 11552
rect 14792 11540 14798 11552
rect 14844 11549 14872 11580
rect 15381 11577 15393 11580
rect 15427 11577 15439 11611
rect 17972 11608 18000 11636
rect 18616 11608 18644 11707
rect 18690 11608 18696 11620
rect 17972 11580 18696 11608
rect 15381 11571 15439 11577
rect 18690 11568 18696 11580
rect 18748 11568 18754 11620
rect 14829 11543 14887 11549
rect 14829 11540 14841 11543
rect 14792 11512 14841 11540
rect 14792 11500 14798 11512
rect 14829 11509 14841 11512
rect 14875 11509 14887 11543
rect 15010 11540 15016 11552
rect 14971 11512 15016 11540
rect 14829 11503 14887 11509
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 15102 11500 15108 11552
rect 15160 11540 15166 11552
rect 15473 11543 15531 11549
rect 15473 11540 15485 11543
rect 15160 11512 15485 11540
rect 15160 11500 15166 11512
rect 15473 11509 15485 11512
rect 15519 11540 15531 11543
rect 15746 11540 15752 11552
rect 15519 11512 15752 11540
rect 15519 11509 15531 11512
rect 15473 11503 15531 11509
rect 15746 11500 15752 11512
rect 15804 11500 15810 11552
rect 17494 11540 17500 11552
rect 17455 11512 17500 11540
rect 17494 11500 17500 11512
rect 17552 11500 17558 11552
rect 18046 11540 18052 11552
rect 18007 11512 18052 11540
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 2409 11339 2467 11345
rect 2409 11305 2421 11339
rect 2455 11336 2467 11339
rect 2498 11336 2504 11348
rect 2455 11308 2504 11336
rect 2455 11305 2467 11308
rect 2409 11299 2467 11305
rect 2498 11296 2504 11308
rect 2556 11296 2562 11348
rect 2590 11296 2596 11348
rect 2648 11296 2654 11348
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 2832 11308 3433 11336
rect 2832 11296 2838 11308
rect 3421 11305 3433 11308
rect 3467 11305 3479 11339
rect 3878 11336 3884 11348
rect 3839 11308 3884 11336
rect 3421 11299 3479 11305
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 3970 11296 3976 11348
rect 4028 11336 4034 11348
rect 4249 11339 4307 11345
rect 4249 11336 4261 11339
rect 4028 11308 4261 11336
rect 4028 11296 4034 11308
rect 4249 11305 4261 11308
rect 4295 11305 4307 11339
rect 5258 11336 5264 11348
rect 5219 11308 5264 11336
rect 4249 11299 4307 11305
rect 5258 11296 5264 11308
rect 5316 11296 5322 11348
rect 6825 11339 6883 11345
rect 6825 11305 6837 11339
rect 6871 11336 6883 11339
rect 6914 11336 6920 11348
rect 6871 11308 6920 11336
rect 6871 11305 6883 11308
rect 6825 11299 6883 11305
rect 6914 11296 6920 11308
rect 6972 11296 6978 11348
rect 8294 11336 8300 11348
rect 8255 11308 8300 11336
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 8478 11296 8484 11348
rect 8536 11336 8542 11348
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 8536 11308 8953 11336
rect 8536 11296 8542 11308
rect 8941 11305 8953 11308
rect 8987 11305 8999 11339
rect 8941 11299 8999 11305
rect 9401 11339 9459 11345
rect 9401 11305 9413 11339
rect 9447 11336 9459 11339
rect 9858 11336 9864 11348
rect 9447 11308 9864 11336
rect 9447 11305 9459 11308
rect 9401 11299 9459 11305
rect 9858 11296 9864 11308
rect 9916 11296 9922 11348
rect 9950 11296 9956 11348
rect 10008 11336 10014 11348
rect 11793 11339 11851 11345
rect 10008 11308 10053 11336
rect 10008 11296 10014 11308
rect 11793 11305 11805 11339
rect 11839 11336 11851 11339
rect 12526 11336 12532 11348
rect 11839 11308 12532 11336
rect 11839 11305 11851 11308
rect 11793 11299 11851 11305
rect 12526 11296 12532 11308
rect 12584 11296 12590 11348
rect 12894 11336 12900 11348
rect 12855 11308 12900 11336
rect 12894 11296 12900 11308
rect 12952 11296 12958 11348
rect 13354 11336 13360 11348
rect 13315 11308 13360 11336
rect 13354 11296 13360 11308
rect 13412 11296 13418 11348
rect 15838 11296 15844 11348
rect 15896 11336 15902 11348
rect 17497 11339 17555 11345
rect 17497 11336 17509 11339
rect 15896 11308 17509 11336
rect 15896 11296 15902 11308
rect 17497 11305 17509 11308
rect 17543 11305 17555 11339
rect 18046 11336 18052 11348
rect 18007 11308 18052 11336
rect 17497 11299 17555 11305
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 2608 11268 2636 11296
rect 2866 11268 2872 11280
rect 2608 11240 2872 11268
rect 2866 11228 2872 11240
rect 2924 11228 2930 11280
rect 5712 11271 5770 11277
rect 5712 11237 5724 11271
rect 5758 11268 5770 11271
rect 5994 11268 6000 11280
rect 5758 11240 6000 11268
rect 5758 11237 5770 11240
rect 5712 11231 5770 11237
rect 5994 11228 6000 11240
rect 6052 11268 6058 11280
rect 6730 11268 6736 11280
rect 6052 11240 6736 11268
rect 6052 11228 6058 11240
rect 6730 11228 6736 11240
rect 6788 11228 6794 11280
rect 7469 11271 7527 11277
rect 7469 11237 7481 11271
rect 7515 11268 7527 11271
rect 7837 11271 7895 11277
rect 7837 11268 7849 11271
rect 7515 11240 7849 11268
rect 7515 11237 7527 11240
rect 7469 11231 7527 11237
rect 7837 11237 7849 11240
rect 7883 11268 7895 11271
rect 8202 11268 8208 11280
rect 7883 11240 8208 11268
rect 7883 11237 7895 11240
rect 7837 11231 7895 11237
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 9876 11268 9904 11296
rect 10658 11271 10716 11277
rect 10658 11268 10670 11271
rect 9876 11240 10670 11268
rect 10658 11237 10670 11240
rect 10704 11268 10716 11271
rect 11054 11268 11060 11280
rect 10704 11240 11060 11268
rect 10704 11237 10716 11240
rect 10658 11231 10716 11237
rect 11054 11228 11060 11240
rect 11112 11228 11118 11280
rect 11330 11228 11336 11280
rect 11388 11268 11394 11280
rect 13265 11271 13323 11277
rect 13265 11268 13277 11271
rect 11388 11240 13277 11268
rect 11388 11228 11394 11240
rect 13265 11237 13277 11240
rect 13311 11268 13323 11271
rect 13446 11268 13452 11280
rect 13311 11240 13452 11268
rect 13311 11237 13323 11240
rect 13265 11231 13323 11237
rect 13446 11228 13452 11240
rect 13504 11228 13510 11280
rect 14642 11268 14648 11280
rect 14603 11240 14648 11268
rect 14642 11228 14648 11240
rect 14700 11228 14706 11280
rect 17770 11228 17776 11280
rect 17828 11268 17834 11280
rect 18506 11268 18512 11280
rect 17828 11240 18512 11268
rect 17828 11228 17834 11240
rect 18506 11228 18512 11240
rect 18564 11228 18570 11280
rect 2590 11160 2596 11212
rect 2648 11200 2654 11212
rect 2777 11203 2835 11209
rect 2777 11200 2789 11203
rect 2648 11172 2789 11200
rect 2648 11160 2654 11172
rect 2777 11169 2789 11172
rect 2823 11200 2835 11203
rect 3878 11200 3884 11212
rect 2823 11172 3884 11200
rect 2823 11169 2835 11172
rect 2777 11163 2835 11169
rect 3878 11160 3884 11172
rect 3936 11160 3942 11212
rect 4062 11200 4068 11212
rect 4023 11172 4068 11200
rect 4062 11160 4068 11172
rect 4120 11200 4126 11212
rect 4525 11203 4583 11209
rect 4525 11200 4537 11203
rect 4120 11172 4537 11200
rect 4120 11160 4126 11172
rect 4525 11169 4537 11172
rect 4571 11169 4583 11203
rect 4525 11163 4583 11169
rect 5350 11160 5356 11212
rect 5408 11200 5414 11212
rect 5445 11203 5503 11209
rect 5445 11200 5457 11203
rect 5408 11172 5457 11200
rect 5408 11160 5414 11172
rect 5445 11169 5457 11172
rect 5491 11169 5503 11203
rect 8220 11200 8248 11228
rect 8220 11172 8524 11200
rect 5445 11163 5503 11169
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11132 1455 11135
rect 1762 11132 1768 11144
rect 1443 11104 1768 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 1762 11092 1768 11104
rect 1820 11132 1826 11144
rect 1857 11135 1915 11141
rect 1857 11132 1869 11135
rect 1820 11104 1869 11132
rect 1820 11092 1826 11104
rect 1857 11101 1869 11104
rect 1903 11101 1915 11135
rect 2866 11132 2872 11144
rect 2827 11104 2872 11132
rect 1857 11095 1915 11101
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11132 3111 11135
rect 3418 11132 3424 11144
rect 3099 11104 3424 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 2317 10999 2375 11005
rect 2317 10965 2329 10999
rect 2363 10996 2375 10999
rect 3068 10996 3096 11095
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 7282 11092 7288 11144
rect 7340 11132 7346 11144
rect 8496 11141 8524 11172
rect 9766 11160 9772 11212
rect 9824 11200 9830 11212
rect 10413 11203 10471 11209
rect 10413 11200 10425 11203
rect 9824 11172 10425 11200
rect 9824 11160 9830 11172
rect 10413 11169 10425 11172
rect 10459 11200 10471 11203
rect 11882 11200 11888 11212
rect 10459 11172 11888 11200
rect 10459 11169 10471 11172
rect 10413 11163 10471 11169
rect 11882 11160 11888 11172
rect 11940 11160 11946 11212
rect 13906 11200 13912 11212
rect 13556 11172 13912 11200
rect 13556 11141 13584 11172
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 15654 11160 15660 11212
rect 15712 11200 15718 11212
rect 15821 11203 15879 11209
rect 15821 11200 15833 11203
rect 15712 11172 15833 11200
rect 15712 11160 15718 11172
rect 15821 11169 15833 11172
rect 15867 11169 15879 11203
rect 15821 11163 15879 11169
rect 18322 11160 18328 11212
rect 18380 11200 18386 11212
rect 18417 11203 18475 11209
rect 18417 11200 18429 11203
rect 18380 11172 18429 11200
rect 18380 11160 18386 11172
rect 18417 11169 18429 11172
rect 18463 11169 18475 11203
rect 18417 11163 18475 11169
rect 8389 11135 8447 11141
rect 8389 11132 8401 11135
rect 7340 11104 8401 11132
rect 7340 11092 7346 11104
rect 8389 11101 8401 11104
rect 8435 11101 8447 11135
rect 8389 11095 8447 11101
rect 8481 11135 8539 11141
rect 8481 11101 8493 11135
rect 8527 11101 8539 11135
rect 8481 11095 8539 11101
rect 13541 11135 13599 11141
rect 13541 11101 13553 11135
rect 13587 11101 13599 11135
rect 15010 11132 15016 11144
rect 14971 11104 15016 11132
rect 13541 11095 13599 11101
rect 7929 11067 7987 11073
rect 7929 11033 7941 11067
rect 7975 11064 7987 11067
rect 8294 11064 8300 11076
rect 7975 11036 8300 11064
rect 7975 11033 7987 11036
rect 7929 11027 7987 11033
rect 8294 11024 8300 11036
rect 8352 11024 8358 11076
rect 8404 11064 8432 11095
rect 15010 11092 15016 11104
rect 15068 11092 15074 11144
rect 15470 11092 15476 11144
rect 15528 11132 15534 11144
rect 15565 11135 15623 11141
rect 15565 11132 15577 11135
rect 15528 11104 15577 11132
rect 15528 11092 15534 11104
rect 15565 11101 15577 11104
rect 15611 11101 15623 11135
rect 18690 11132 18696 11144
rect 18651 11104 18696 11132
rect 15565 11095 15623 11101
rect 18690 11092 18696 11104
rect 18748 11092 18754 11144
rect 8570 11064 8576 11076
rect 8404 11036 8576 11064
rect 8570 11024 8576 11036
rect 8628 11024 8634 11076
rect 13906 11064 13912 11076
rect 13867 11036 13912 11064
rect 13906 11024 13912 11036
rect 13964 11024 13970 11076
rect 14274 11064 14280 11076
rect 14235 11036 14280 11064
rect 14274 11024 14280 11036
rect 14332 11024 14338 11076
rect 16945 11067 17003 11073
rect 16945 11064 16957 11067
rect 16500 11036 16957 11064
rect 4982 10996 4988 11008
rect 2363 10968 3096 10996
rect 4943 10968 4988 10996
rect 2363 10965 2375 10968
rect 2317 10959 2375 10965
rect 4982 10956 4988 10968
rect 5040 10956 5046 11008
rect 9950 10956 9956 11008
rect 10008 10996 10014 11008
rect 10134 10996 10140 11008
rect 10008 10968 10140 10996
rect 10008 10956 10014 10968
rect 10134 10956 10140 10968
rect 10192 10956 10198 11008
rect 10321 10999 10379 11005
rect 10321 10965 10333 10999
rect 10367 10996 10379 10999
rect 10778 10996 10784 11008
rect 10367 10968 10784 10996
rect 10367 10965 10379 10968
rect 10321 10959 10379 10965
rect 10778 10956 10784 10968
rect 10836 10956 10842 11008
rect 12529 10999 12587 11005
rect 12529 10965 12541 10999
rect 12575 10996 12587 10999
rect 13170 10996 13176 11008
rect 12575 10968 13176 10996
rect 12575 10965 12587 10968
rect 12529 10959 12587 10965
rect 13170 10956 13176 10968
rect 13228 10956 13234 11008
rect 14642 10956 14648 11008
rect 14700 10996 14706 11008
rect 15746 10996 15752 11008
rect 14700 10968 15752 10996
rect 14700 10956 14706 10968
rect 15746 10956 15752 10968
rect 15804 10956 15810 11008
rect 16206 10956 16212 11008
rect 16264 10996 16270 11008
rect 16500 10996 16528 11036
rect 16945 11033 16957 11036
rect 16991 11033 17003 11067
rect 16945 11027 17003 11033
rect 16264 10968 16528 10996
rect 16264 10956 16270 10968
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1397 10795 1455 10801
rect 1397 10761 1409 10795
rect 1443 10792 1455 10795
rect 2590 10792 2596 10804
rect 1443 10764 2596 10792
rect 1443 10761 1455 10764
rect 1397 10755 1455 10761
rect 2590 10752 2596 10764
rect 2648 10752 2654 10804
rect 3142 10792 3148 10804
rect 3103 10764 3148 10792
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 3237 10795 3295 10801
rect 3237 10761 3249 10795
rect 3283 10792 3295 10795
rect 3326 10792 3332 10804
rect 3283 10764 3332 10792
rect 3283 10761 3295 10764
rect 3237 10755 3295 10761
rect 3326 10752 3332 10764
rect 3384 10752 3390 10804
rect 4890 10752 4896 10804
rect 4948 10792 4954 10804
rect 5169 10795 5227 10801
rect 5169 10792 5181 10795
rect 4948 10764 5181 10792
rect 4948 10752 4954 10764
rect 5169 10761 5181 10764
rect 5215 10792 5227 10795
rect 5442 10792 5448 10804
rect 5215 10764 5448 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 6178 10792 6184 10804
rect 6139 10764 6184 10792
rect 6178 10752 6184 10764
rect 6236 10752 6242 10804
rect 6641 10795 6699 10801
rect 6641 10761 6653 10795
rect 6687 10792 6699 10795
rect 6822 10792 6828 10804
rect 6687 10764 6828 10792
rect 6687 10761 6699 10764
rect 6641 10755 6699 10761
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 9217 10795 9275 10801
rect 9217 10761 9229 10795
rect 9263 10792 9275 10795
rect 9766 10792 9772 10804
rect 9263 10764 9332 10792
rect 9727 10764 9772 10792
rect 9263 10761 9275 10764
rect 9217 10755 9275 10761
rect 1854 10656 1860 10668
rect 1815 10628 1860 10656
rect 1854 10616 1860 10628
rect 1912 10616 1918 10668
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 2682 10656 2688 10668
rect 2087 10628 2688 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 3160 10656 3188 10752
rect 6196 10724 6224 10752
rect 7653 10727 7711 10733
rect 7653 10724 7665 10727
rect 6196 10696 7665 10724
rect 7653 10693 7665 10696
rect 7699 10693 7711 10727
rect 7653 10687 7711 10693
rect 3697 10659 3755 10665
rect 3697 10656 3709 10659
rect 3160 10628 3709 10656
rect 3697 10625 3709 10628
rect 3743 10625 3755 10659
rect 3878 10656 3884 10668
rect 3839 10628 3884 10656
rect 3697 10619 3755 10625
rect 3878 10616 3884 10628
rect 3936 10616 3942 10668
rect 4709 10659 4767 10665
rect 4709 10625 4721 10659
rect 4755 10656 4767 10659
rect 5077 10659 5135 10665
rect 5077 10656 5089 10659
rect 4755 10628 5089 10656
rect 4755 10625 4767 10628
rect 4709 10619 4767 10625
rect 5077 10625 5089 10628
rect 5123 10656 5135 10659
rect 5813 10659 5871 10665
rect 5813 10656 5825 10659
rect 5123 10628 5825 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 5813 10625 5825 10628
rect 5859 10656 5871 10659
rect 5994 10656 6000 10668
rect 5859 10628 6000 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 5994 10616 6000 10628
rect 6052 10616 6058 10668
rect 7668 10656 7696 10687
rect 9304 10668 9332 10764
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 11054 10752 11060 10804
rect 11112 10792 11118 10804
rect 11701 10795 11759 10801
rect 11701 10792 11713 10795
rect 11112 10764 11713 10792
rect 11112 10752 11118 10764
rect 11701 10761 11713 10764
rect 11747 10761 11759 10795
rect 13446 10792 13452 10804
rect 13407 10764 13452 10792
rect 11701 10755 11759 10761
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 13538 10752 13544 10804
rect 13596 10792 13602 10804
rect 14001 10795 14059 10801
rect 14001 10792 14013 10795
rect 13596 10764 14013 10792
rect 13596 10752 13602 10764
rect 14001 10761 14013 10764
rect 14047 10761 14059 10795
rect 14001 10755 14059 10761
rect 15105 10795 15163 10801
rect 15105 10761 15117 10795
rect 15151 10792 15163 10795
rect 16114 10792 16120 10804
rect 15151 10764 16120 10792
rect 15151 10761 15163 10764
rect 15105 10755 15163 10761
rect 16114 10752 16120 10764
rect 16172 10752 16178 10804
rect 16666 10792 16672 10804
rect 16579 10764 16672 10792
rect 16666 10752 16672 10764
rect 16724 10792 16730 10804
rect 17402 10792 17408 10804
rect 16724 10764 17408 10792
rect 16724 10752 16730 10764
rect 17402 10752 17408 10764
rect 17460 10752 17466 10804
rect 18049 10795 18107 10801
rect 18049 10761 18061 10795
rect 18095 10792 18107 10795
rect 18598 10792 18604 10804
rect 18095 10764 18604 10792
rect 18095 10761 18107 10764
rect 18049 10755 18107 10761
rect 18598 10752 18604 10764
rect 18656 10752 18662 10804
rect 9674 10684 9680 10736
rect 9732 10724 9738 10736
rect 10321 10727 10379 10733
rect 10321 10724 10333 10727
rect 9732 10696 10333 10724
rect 9732 10684 9738 10696
rect 10321 10693 10333 10696
rect 10367 10693 10379 10727
rect 13814 10724 13820 10736
rect 13775 10696 13820 10724
rect 10321 10687 10379 10693
rect 13814 10684 13820 10696
rect 13872 10724 13878 10736
rect 15470 10724 15476 10736
rect 13872 10696 14596 10724
rect 15383 10696 15476 10724
rect 13872 10684 13878 10696
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 7668 10628 7849 10656
rect 7837 10625 7849 10628
rect 7883 10625 7895 10659
rect 9304 10628 9312 10668
rect 7837 10619 7895 10625
rect 9306 10616 9312 10628
rect 9364 10656 9370 10668
rect 10778 10656 10784 10668
rect 9364 10628 10784 10656
rect 9364 10616 9370 10628
rect 10778 10616 10784 10628
rect 10836 10656 10842 10668
rect 10873 10659 10931 10665
rect 10873 10656 10885 10659
rect 10836 10628 10885 10656
rect 10836 10616 10842 10628
rect 10873 10625 10885 10628
rect 10919 10625 10931 10659
rect 10873 10619 10931 10625
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10656 13139 10659
rect 13170 10656 13176 10668
rect 13127 10628 13176 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 14458 10656 14464 10668
rect 14419 10628 14464 10656
rect 14458 10616 14464 10628
rect 14516 10616 14522 10668
rect 14568 10665 14596 10696
rect 15470 10684 15476 10696
rect 15528 10724 15534 10736
rect 15930 10724 15936 10736
rect 15528 10696 15936 10724
rect 15528 10684 15534 10696
rect 15930 10684 15936 10696
rect 15988 10684 15994 10736
rect 16945 10727 17003 10733
rect 16945 10724 16957 10727
rect 16040 10696 16957 10724
rect 16040 10668 16068 10696
rect 16945 10693 16957 10696
rect 16991 10693 17003 10727
rect 16945 10687 17003 10693
rect 14553 10659 14611 10665
rect 14553 10625 14565 10659
rect 14599 10625 14611 10659
rect 16022 10656 16028 10668
rect 15983 10628 16028 10656
rect 14553 10619 14611 10625
rect 16022 10616 16028 10628
rect 16080 10616 16086 10668
rect 16114 10616 16120 10668
rect 16172 10656 16178 10668
rect 16172 10628 16217 10656
rect 16172 10616 16178 10628
rect 17402 10616 17408 10668
rect 17460 10656 17466 10668
rect 17497 10659 17555 10665
rect 17497 10656 17509 10659
rect 17460 10628 17509 10656
rect 17460 10616 17466 10628
rect 17497 10625 17509 10628
rect 17543 10656 17555 10659
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 17543 10628 18613 10656
rect 17543 10625 17555 10628
rect 17497 10619 17555 10625
rect 18601 10625 18613 10628
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 1394 10548 1400 10600
rect 1452 10588 1458 10600
rect 1765 10591 1823 10597
rect 1765 10588 1777 10591
rect 1452 10560 1777 10588
rect 1452 10548 1458 10560
rect 1765 10557 1777 10560
rect 1811 10557 1823 10591
rect 1765 10551 1823 10557
rect 2777 10591 2835 10597
rect 2777 10557 2789 10591
rect 2823 10588 2835 10591
rect 3605 10591 3663 10597
rect 3605 10588 3617 10591
rect 2823 10560 3617 10588
rect 2823 10557 2835 10560
rect 2777 10551 2835 10557
rect 3605 10557 3617 10560
rect 3651 10588 3663 10591
rect 4522 10588 4528 10600
rect 3651 10560 4528 10588
rect 3651 10557 3663 10560
rect 3605 10551 3663 10557
rect 4522 10548 4528 10560
rect 4580 10548 4586 10600
rect 4982 10548 4988 10600
rect 5040 10588 5046 10600
rect 5442 10588 5448 10600
rect 5040 10560 5448 10588
rect 5040 10548 5046 10560
rect 5442 10548 5448 10560
rect 5500 10588 5506 10600
rect 5537 10591 5595 10597
rect 5537 10588 5549 10591
rect 5500 10560 5549 10588
rect 5500 10548 5506 10560
rect 5537 10557 5549 10560
rect 5583 10557 5595 10591
rect 12158 10588 12164 10600
rect 12119 10560 12164 10588
rect 5537 10551 5595 10557
rect 12158 10548 12164 10560
rect 12216 10588 12222 10600
rect 12897 10591 12955 10597
rect 12897 10588 12909 10591
rect 12216 10560 12909 10588
rect 12216 10548 12222 10560
rect 12897 10557 12909 10560
rect 12943 10557 12955 10591
rect 14366 10588 14372 10600
rect 14327 10560 14372 10588
rect 12897 10551 12955 10557
rect 14366 10548 14372 10560
rect 14424 10548 14430 10600
rect 15838 10548 15844 10600
rect 15896 10588 15902 10600
rect 15933 10591 15991 10597
rect 15933 10588 15945 10591
rect 15896 10560 15945 10588
rect 15896 10548 15902 10560
rect 15933 10557 15945 10560
rect 15979 10557 15991 10591
rect 15933 10551 15991 10557
rect 842 10480 848 10532
rect 900 10520 906 10532
rect 7282 10520 7288 10532
rect 900 10492 7288 10520
rect 900 10480 906 10492
rect 7282 10480 7288 10492
rect 7340 10480 7346 10532
rect 8104 10523 8162 10529
rect 8104 10489 8116 10523
rect 8150 10520 8162 10523
rect 8202 10520 8208 10532
rect 8150 10492 8208 10520
rect 8150 10489 8162 10492
rect 8104 10483 8162 10489
rect 8202 10480 8208 10492
rect 8260 10480 8266 10532
rect 10594 10480 10600 10532
rect 10652 10520 10658 10532
rect 10781 10523 10839 10529
rect 10781 10520 10793 10523
rect 10652 10492 10793 10520
rect 10652 10480 10658 10492
rect 10781 10489 10793 10492
rect 10827 10520 10839 10523
rect 11333 10523 11391 10529
rect 11333 10520 11345 10523
rect 10827 10492 11345 10520
rect 10827 10489 10839 10492
rect 10781 10483 10839 10489
rect 11333 10489 11345 10492
rect 11379 10489 11391 10523
rect 11333 10483 11391 10489
rect 12805 10523 12863 10529
rect 12805 10489 12817 10523
rect 12851 10520 12863 10523
rect 13078 10520 13084 10532
rect 12851 10492 13084 10520
rect 12851 10489 12863 10492
rect 12805 10483 12863 10489
rect 13078 10480 13084 10492
rect 13136 10480 13142 10532
rect 18509 10523 18567 10529
rect 18509 10520 18521 10523
rect 15580 10492 18521 10520
rect 3878 10412 3884 10464
rect 3936 10452 3942 10464
rect 4246 10452 4252 10464
rect 3936 10424 4252 10452
rect 3936 10412 3942 10424
rect 4246 10412 4252 10424
rect 4304 10412 4310 10464
rect 5258 10412 5264 10464
rect 5316 10452 5322 10464
rect 5629 10455 5687 10461
rect 5629 10452 5641 10455
rect 5316 10424 5641 10452
rect 5316 10412 5322 10424
rect 5629 10421 5641 10424
rect 5675 10421 5687 10455
rect 5629 10415 5687 10421
rect 9490 10412 9496 10464
rect 9548 10452 9554 10464
rect 10137 10455 10195 10461
rect 10137 10452 10149 10455
rect 9548 10424 10149 10452
rect 9548 10412 9554 10424
rect 10137 10421 10149 10424
rect 10183 10452 10195 10455
rect 10689 10455 10747 10461
rect 10689 10452 10701 10455
rect 10183 10424 10701 10452
rect 10183 10421 10195 10424
rect 10137 10415 10195 10421
rect 10689 10421 10701 10424
rect 10735 10421 10747 10455
rect 10689 10415 10747 10421
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 12710 10452 12716 10464
rect 12483 10424 12716 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 15580 10461 15608 10492
rect 18509 10489 18521 10492
rect 18555 10520 18567 10523
rect 19061 10523 19119 10529
rect 19061 10520 19073 10523
rect 18555 10492 19073 10520
rect 18555 10489 18567 10492
rect 18509 10483 18567 10489
rect 19061 10489 19073 10492
rect 19107 10489 19119 10523
rect 19061 10483 19119 10489
rect 15565 10455 15623 10461
rect 15565 10421 15577 10455
rect 15611 10421 15623 10455
rect 15565 10415 15623 10421
rect 15746 10412 15752 10464
rect 15804 10452 15810 10464
rect 17770 10452 17776 10464
rect 15804 10424 17776 10452
rect 15804 10412 15810 10424
rect 17770 10412 17776 10424
rect 17828 10412 17834 10464
rect 18417 10455 18475 10461
rect 18417 10421 18429 10455
rect 18463 10452 18475 10455
rect 18782 10452 18788 10464
rect 18463 10424 18788 10452
rect 18463 10421 18475 10424
rect 18417 10415 18475 10421
rect 18782 10412 18788 10424
rect 18840 10412 18846 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1762 10248 1768 10260
rect 1723 10220 1768 10248
rect 1762 10208 1768 10220
rect 1820 10208 1826 10260
rect 4154 10208 4160 10260
rect 4212 10248 4218 10260
rect 4249 10251 4307 10257
rect 4249 10248 4261 10251
rect 4212 10220 4261 10248
rect 4212 10208 4218 10220
rect 4249 10217 4261 10220
rect 4295 10217 4307 10251
rect 4890 10248 4896 10260
rect 4851 10220 4896 10248
rect 4249 10211 4307 10217
rect 4890 10208 4896 10220
rect 4948 10208 4954 10260
rect 5442 10248 5448 10260
rect 5403 10220 5448 10248
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 7834 10248 7840 10260
rect 7795 10220 7840 10248
rect 7834 10208 7840 10220
rect 7892 10208 7898 10260
rect 8294 10208 8300 10260
rect 8352 10248 8358 10260
rect 8481 10251 8539 10257
rect 8481 10248 8493 10251
rect 8352 10220 8493 10248
rect 8352 10208 8358 10220
rect 8481 10217 8493 10220
rect 8527 10248 8539 10251
rect 9401 10251 9459 10257
rect 9401 10248 9413 10251
rect 8527 10220 9413 10248
rect 8527 10217 8539 10220
rect 8481 10211 8539 10217
rect 9401 10217 9413 10220
rect 9447 10217 9459 10251
rect 9766 10248 9772 10260
rect 9401 10211 9459 10217
rect 9600 10220 9772 10248
rect 3513 10183 3571 10189
rect 3513 10149 3525 10183
rect 3559 10180 3571 10183
rect 4706 10180 4712 10192
rect 3559 10152 4712 10180
rect 3559 10149 3571 10152
rect 3513 10143 3571 10149
rect 3528 10056 3556 10143
rect 4706 10140 4712 10152
rect 4764 10140 4770 10192
rect 5905 10183 5963 10189
rect 5905 10149 5917 10183
rect 5951 10180 5963 10183
rect 5994 10180 6000 10192
rect 5951 10152 6000 10180
rect 5951 10149 5963 10152
rect 5905 10143 5963 10149
rect 5994 10140 6000 10152
rect 6052 10140 6058 10192
rect 5534 10072 5540 10124
rect 5592 10112 5598 10124
rect 5813 10115 5871 10121
rect 5813 10112 5825 10115
rect 5592 10084 5825 10112
rect 5592 10072 5598 10084
rect 5813 10081 5825 10084
rect 5859 10081 5871 10115
rect 5813 10075 5871 10081
rect 8294 10072 8300 10124
rect 8352 10112 8358 10124
rect 8389 10115 8447 10121
rect 8389 10112 8401 10115
rect 8352 10084 8401 10112
rect 8352 10072 8358 10084
rect 8389 10081 8401 10084
rect 8435 10081 8447 10115
rect 9600 10112 9628 10220
rect 9766 10208 9772 10220
rect 9824 10208 9830 10260
rect 11054 10248 11060 10260
rect 11015 10220 11060 10248
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 12805 10251 12863 10257
rect 12805 10217 12817 10251
rect 12851 10248 12863 10251
rect 12894 10248 12900 10260
rect 12851 10220 12900 10248
rect 12851 10217 12863 10220
rect 12805 10211 12863 10217
rect 12894 10208 12900 10220
rect 12952 10208 12958 10260
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 14001 10251 14059 10257
rect 14001 10248 14013 10251
rect 13872 10220 14013 10248
rect 13872 10208 13878 10220
rect 14001 10217 14013 10220
rect 14047 10217 14059 10251
rect 14001 10211 14059 10217
rect 14458 10208 14464 10260
rect 14516 10248 14522 10260
rect 14737 10251 14795 10257
rect 14737 10248 14749 10251
rect 14516 10220 14749 10248
rect 14516 10208 14522 10220
rect 14737 10217 14749 10220
rect 14783 10217 14795 10251
rect 17402 10248 17408 10260
rect 17363 10220 17408 10248
rect 14737 10211 14795 10217
rect 17402 10208 17408 10220
rect 17460 10208 17466 10260
rect 18509 10251 18567 10257
rect 18509 10217 18521 10251
rect 18555 10248 18567 10251
rect 18690 10248 18696 10260
rect 18555 10220 18696 10248
rect 18555 10217 18567 10220
rect 18509 10211 18567 10217
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 9674 10140 9680 10192
rect 9732 10180 9738 10192
rect 11609 10183 11667 10189
rect 11609 10180 11621 10183
rect 9732 10152 11621 10180
rect 9732 10140 9738 10152
rect 11609 10149 11621 10152
rect 11655 10149 11667 10183
rect 12526 10180 12532 10192
rect 12439 10152 12532 10180
rect 11609 10143 11667 10149
rect 12526 10140 12532 10152
rect 12584 10180 12590 10192
rect 13078 10180 13084 10192
rect 12584 10152 13084 10180
rect 12584 10140 12590 10152
rect 13078 10140 13084 10152
rect 13136 10140 13142 10192
rect 14366 10180 14372 10192
rect 14327 10152 14372 10180
rect 14366 10140 14372 10152
rect 14424 10140 14430 10192
rect 16114 10140 16120 10192
rect 16172 10180 16178 10192
rect 16270 10183 16328 10189
rect 16270 10180 16282 10183
rect 16172 10152 16282 10180
rect 16172 10140 16178 10152
rect 16270 10149 16282 10152
rect 16316 10149 16328 10183
rect 16270 10143 16328 10149
rect 9600 10084 9720 10112
rect 8389 10075 8447 10081
rect 1854 10044 1860 10056
rect 1815 10016 1860 10044
rect 1854 10004 1860 10016
rect 1912 10004 1918 10056
rect 2038 10044 2044 10056
rect 1951 10016 2044 10044
rect 2038 10004 2044 10016
rect 2096 10044 2102 10056
rect 3510 10044 3516 10056
rect 2096 10016 3516 10044
rect 2096 10004 2102 10016
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 5350 10004 5356 10056
rect 5408 10044 5414 10056
rect 5997 10047 6055 10053
rect 5997 10044 6009 10047
rect 5408 10016 6009 10044
rect 5408 10004 5414 10016
rect 5997 10013 6009 10016
rect 6043 10044 6055 10047
rect 7193 10047 7251 10053
rect 7193 10044 7205 10047
rect 6043 10016 7205 10044
rect 6043 10013 6055 10016
rect 5997 10007 6055 10013
rect 7193 10013 7205 10016
rect 7239 10044 7251 10047
rect 7374 10044 7380 10056
rect 7239 10016 7380 10044
rect 7239 10013 7251 10016
rect 7193 10007 7251 10013
rect 7374 10004 7380 10016
rect 7432 10004 7438 10056
rect 8478 10004 8484 10056
rect 8536 10044 8542 10056
rect 8665 10047 8723 10053
rect 8665 10044 8677 10047
rect 8536 10016 8677 10044
rect 8536 10004 8542 10016
rect 8665 10013 8677 10016
rect 8711 10044 8723 10047
rect 9306 10044 9312 10056
rect 8711 10016 9312 10044
rect 8711 10013 8723 10016
rect 8665 10007 8723 10013
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 9692 10053 9720 10084
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 9933 10115 9991 10121
rect 9933 10112 9945 10115
rect 9824 10084 9945 10112
rect 9824 10072 9830 10084
rect 9933 10081 9945 10084
rect 9979 10081 9991 10115
rect 9933 10075 9991 10081
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 13173 10115 13231 10121
rect 13173 10112 13185 10115
rect 12492 10084 13185 10112
rect 12492 10072 12498 10084
rect 13173 10081 13185 10084
rect 13219 10081 13231 10115
rect 13173 10075 13231 10081
rect 9677 10047 9735 10053
rect 9677 10013 9689 10047
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 1394 9976 1400 9988
rect 1355 9948 1400 9976
rect 1394 9936 1400 9948
rect 1452 9936 1458 9988
rect 6549 9979 6607 9985
rect 6549 9945 6561 9979
rect 6595 9976 6607 9979
rect 8021 9979 8079 9985
rect 8021 9976 8033 9979
rect 6595 9948 8033 9976
rect 6595 9945 6607 9948
rect 6549 9939 6607 9945
rect 8021 9945 8033 9948
rect 8067 9976 8079 9979
rect 8294 9976 8300 9988
rect 8067 9948 8300 9976
rect 8067 9945 8079 9948
rect 8021 9939 8079 9945
rect 8294 9936 8300 9948
rect 8352 9936 8358 9988
rect 2406 9908 2412 9920
rect 2367 9880 2412 9908
rect 2406 9868 2412 9880
rect 2464 9868 2470 9920
rect 3050 9908 3056 9920
rect 3011 9880 3056 9908
rect 3050 9868 3056 9880
rect 3108 9868 3114 9920
rect 3878 9908 3884 9920
rect 3839 9880 3884 9908
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 5258 9908 5264 9920
rect 5219 9880 5264 9908
rect 5258 9868 5264 9880
rect 5316 9868 5322 9920
rect 6914 9908 6920 9920
rect 6875 9880 6920 9908
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 9033 9911 9091 9917
rect 9033 9908 9045 9911
rect 8444 9880 9045 9908
rect 8444 9868 8450 9880
rect 9033 9877 9045 9880
rect 9079 9877 9091 9911
rect 9692 9908 9720 10007
rect 12894 10004 12900 10056
rect 12952 10044 12958 10056
rect 13262 10044 13268 10056
rect 12952 10016 13268 10044
rect 12952 10004 12958 10016
rect 13262 10004 13268 10016
rect 13320 10004 13326 10056
rect 13446 10044 13452 10056
rect 13407 10016 13452 10044
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 16022 10044 16028 10056
rect 15983 10016 16028 10044
rect 16022 10004 16028 10016
rect 16080 10004 16086 10056
rect 18141 9979 18199 9985
rect 18141 9945 18153 9979
rect 18187 9976 18199 9979
rect 18322 9976 18328 9988
rect 18187 9948 18328 9976
rect 18187 9945 18199 9948
rect 18141 9939 18199 9945
rect 18322 9936 18328 9948
rect 18380 9976 18386 9988
rect 19242 9976 19248 9988
rect 18380 9948 19248 9976
rect 18380 9936 18386 9948
rect 19242 9936 19248 9948
rect 19300 9936 19306 9988
rect 10318 9908 10324 9920
rect 9692 9880 10324 9908
rect 9033 9871 9091 9877
rect 10318 9868 10324 9880
rect 10376 9868 10382 9920
rect 10962 9868 10968 9920
rect 11020 9908 11026 9920
rect 11977 9911 12035 9917
rect 11977 9908 11989 9911
rect 11020 9880 11989 9908
rect 11020 9868 11026 9880
rect 11977 9877 11989 9880
rect 12023 9877 12035 9911
rect 15654 9908 15660 9920
rect 15615 9880 15660 9908
rect 11977 9871 12035 9877
rect 15654 9868 15660 9880
rect 15712 9868 15718 9920
rect 18782 9908 18788 9920
rect 18743 9880 18788 9908
rect 18782 9868 18788 9880
rect 18840 9868 18846 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1397 9707 1455 9713
rect 1397 9673 1409 9707
rect 1443 9704 1455 9707
rect 1762 9704 1768 9716
rect 1443 9676 1768 9704
rect 1443 9673 1455 9676
rect 1397 9667 1455 9673
rect 1762 9664 1768 9676
rect 1820 9664 1826 9716
rect 5258 9664 5264 9716
rect 5316 9704 5322 9716
rect 6825 9707 6883 9713
rect 6825 9704 6837 9707
rect 5316 9676 6837 9704
rect 5316 9664 5322 9676
rect 6825 9673 6837 9676
rect 6871 9673 6883 9707
rect 8478 9704 8484 9716
rect 8439 9676 8484 9704
rect 6825 9667 6883 9673
rect 8478 9664 8484 9676
rect 8536 9664 8542 9716
rect 9769 9707 9827 9713
rect 9769 9673 9781 9707
rect 9815 9704 9827 9707
rect 10318 9704 10324 9716
rect 9815 9676 10324 9704
rect 9815 9673 9827 9676
rect 9769 9667 9827 9673
rect 10318 9664 10324 9676
rect 10376 9664 10382 9716
rect 12894 9704 12900 9716
rect 12360 9676 12900 9704
rect 1854 9596 1860 9648
rect 1912 9636 1918 9648
rect 2409 9639 2467 9645
rect 2409 9636 2421 9639
rect 1912 9608 2421 9636
rect 1912 9596 1918 9608
rect 2409 9605 2421 9608
rect 2455 9605 2467 9639
rect 2409 9599 2467 9605
rect 5077 9639 5135 9645
rect 5077 9605 5089 9639
rect 5123 9636 5135 9639
rect 5350 9636 5356 9648
rect 5123 9608 5356 9636
rect 5123 9605 5135 9608
rect 5077 9599 5135 9605
rect 5350 9596 5356 9608
rect 5408 9596 5414 9648
rect 6638 9596 6644 9648
rect 6696 9596 6702 9648
rect 8110 9636 8116 9648
rect 8071 9608 8116 9636
rect 8110 9596 8116 9608
rect 8168 9596 8174 9648
rect 8665 9639 8723 9645
rect 8665 9605 8677 9639
rect 8711 9636 8723 9639
rect 9582 9636 9588 9648
rect 8711 9608 9588 9636
rect 8711 9605 8723 9608
rect 8665 9599 8723 9605
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 10594 9636 10600 9648
rect 10555 9608 10600 9636
rect 10594 9596 10600 9608
rect 10652 9596 10658 9648
rect 12253 9639 12311 9645
rect 12253 9605 12265 9639
rect 12299 9636 12311 9639
rect 12360 9636 12388 9676
rect 12894 9664 12900 9676
rect 12952 9664 12958 9716
rect 12299 9608 12388 9636
rect 15197 9639 15255 9645
rect 12299 9605 12311 9608
rect 12253 9599 12311 9605
rect 15197 9605 15209 9639
rect 15243 9636 15255 9639
rect 15562 9636 15568 9648
rect 15243 9608 15568 9636
rect 15243 9605 15255 9608
rect 15197 9599 15255 9605
rect 15562 9596 15568 9608
rect 15620 9596 15626 9648
rect 16298 9636 16304 9648
rect 16259 9608 16304 9636
rect 16298 9596 16304 9608
rect 16356 9596 16362 9648
rect 2038 9568 2044 9580
rect 1999 9540 2044 9568
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 2130 9528 2136 9580
rect 2188 9568 2194 9580
rect 3050 9568 3056 9580
rect 2188 9540 3056 9568
rect 2188 9528 2194 9540
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9568 5503 9571
rect 5534 9568 5540 9580
rect 5491 9540 5540 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 1762 9500 1768 9512
rect 1675 9472 1768 9500
rect 1762 9460 1768 9472
rect 1820 9500 1826 9512
rect 2406 9500 2412 9512
rect 1820 9472 2412 9500
rect 1820 9460 1826 9472
rect 2406 9460 2412 9472
rect 2464 9460 2470 9512
rect 2866 9460 2872 9512
rect 2924 9500 2930 9512
rect 3320 9503 3378 9509
rect 3320 9500 3332 9503
rect 2924 9472 3332 9500
rect 2924 9460 2930 9472
rect 3320 9469 3332 9472
rect 3366 9500 3378 9503
rect 4062 9500 4068 9512
rect 3366 9472 4068 9500
rect 3366 9469 3378 9472
rect 3320 9463 3378 9469
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 6546 9460 6552 9512
rect 6604 9500 6610 9512
rect 6656 9500 6684 9596
rect 7374 9568 7380 9580
rect 7335 9540 7380 9568
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 8294 9528 8300 9580
rect 8352 9568 8358 9580
rect 9125 9571 9183 9577
rect 9125 9568 9137 9571
rect 8352 9540 9137 9568
rect 8352 9528 8358 9540
rect 9125 9537 9137 9540
rect 9171 9537 9183 9571
rect 9306 9568 9312 9580
rect 9267 9540 9312 9568
rect 9125 9531 9183 9537
rect 9306 9528 9312 9540
rect 9364 9568 9370 9580
rect 9766 9568 9772 9580
rect 9364 9540 9772 9568
rect 9364 9528 9370 9540
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9568 10379 9571
rect 11333 9571 11391 9577
rect 11333 9568 11345 9571
rect 10367 9540 11345 9568
rect 10367 9537 10379 9540
rect 10321 9531 10379 9537
rect 11333 9537 11345 9540
rect 11379 9568 11391 9571
rect 11882 9568 11888 9580
rect 11379 9540 11888 9568
rect 11379 9537 11391 9540
rect 11333 9531 11391 9537
rect 11882 9528 11888 9540
rect 11940 9528 11946 9580
rect 16114 9528 16120 9580
rect 16172 9568 16178 9580
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16172 9540 16865 9568
rect 16172 9528 16178 9540
rect 16853 9537 16865 9540
rect 16899 9568 16911 9571
rect 17313 9571 17371 9577
rect 17313 9568 17325 9571
rect 16899 9540 17325 9568
rect 16899 9537 16911 9540
rect 16853 9531 16911 9537
rect 17313 9537 17325 9540
rect 17359 9537 17371 9571
rect 17313 9531 17371 9537
rect 6604 9472 6684 9500
rect 9033 9503 9091 9509
rect 6604 9460 6610 9472
rect 9033 9469 9045 9503
rect 9079 9500 9091 9503
rect 9674 9500 9680 9512
rect 9079 9472 9680 9500
rect 9079 9469 9091 9472
rect 9033 9463 9091 9469
rect 9674 9460 9680 9472
rect 9732 9460 9738 9512
rect 10594 9460 10600 9512
rect 10652 9500 10658 9512
rect 11241 9503 11299 9509
rect 11241 9500 11253 9503
rect 10652 9472 11253 9500
rect 10652 9460 10658 9472
rect 11241 9469 11253 9472
rect 11287 9500 11299 9503
rect 11974 9500 11980 9512
rect 11287 9472 11980 9500
rect 11287 9469 11299 9472
rect 11241 9463 11299 9469
rect 11974 9460 11980 9472
rect 12032 9460 12038 9512
rect 13817 9503 13875 9509
rect 13817 9469 13829 9503
rect 13863 9500 13875 9503
rect 13863 9472 14228 9500
rect 13863 9469 13875 9472
rect 13817 9463 13875 9469
rect 6362 9392 6368 9444
rect 6420 9432 6426 9444
rect 6641 9435 6699 9441
rect 6641 9432 6653 9435
rect 6420 9404 6653 9432
rect 6420 9392 6426 9404
rect 6641 9401 6653 9404
rect 6687 9432 6699 9435
rect 7285 9435 7343 9441
rect 7285 9432 7297 9435
rect 6687 9404 7297 9432
rect 6687 9401 6699 9404
rect 6641 9395 6699 9401
rect 7285 9401 7297 9404
rect 7331 9401 7343 9435
rect 7285 9395 7343 9401
rect 12897 9435 12955 9441
rect 12897 9401 12909 9435
rect 12943 9432 12955 9435
rect 13446 9432 13452 9444
rect 12943 9404 13452 9432
rect 12943 9401 12955 9404
rect 12897 9395 12955 9401
rect 13446 9392 13452 9404
rect 13504 9432 13510 9444
rect 13906 9432 13912 9444
rect 13504 9404 13912 9432
rect 13504 9392 13510 9404
rect 13906 9392 13912 9404
rect 13964 9432 13970 9444
rect 14062 9435 14120 9441
rect 14062 9432 14074 9435
rect 13964 9404 14074 9432
rect 13964 9392 13970 9404
rect 14062 9401 14074 9404
rect 14108 9401 14120 9435
rect 14062 9395 14120 9401
rect 1578 9324 1584 9376
rect 1636 9364 1642 9376
rect 1857 9367 1915 9373
rect 1857 9364 1869 9367
rect 1636 9336 1869 9364
rect 1636 9324 1642 9336
rect 1857 9333 1869 9336
rect 1903 9364 1915 9367
rect 2777 9367 2835 9373
rect 2777 9364 2789 9367
rect 1903 9336 2789 9364
rect 1903 9333 1915 9336
rect 1857 9327 1915 9333
rect 2777 9333 2789 9336
rect 2823 9333 2835 9367
rect 2777 9327 2835 9333
rect 4433 9367 4491 9373
rect 4433 9333 4445 9367
rect 4479 9364 4491 9367
rect 4614 9364 4620 9376
rect 4479 9336 4620 9364
rect 4479 9333 4491 9336
rect 4433 9327 4491 9333
rect 4614 9324 4620 9336
rect 4672 9324 4678 9376
rect 5994 9364 6000 9376
rect 5955 9336 6000 9364
rect 5994 9324 6000 9336
rect 6052 9324 6058 9376
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 7193 9367 7251 9373
rect 7193 9364 7205 9367
rect 6972 9336 7205 9364
rect 6972 9324 6978 9336
rect 7193 9333 7205 9336
rect 7239 9333 7251 9367
rect 10778 9364 10784 9376
rect 10739 9336 10784 9364
rect 7193 9327 7251 9333
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 10870 9324 10876 9376
rect 10928 9364 10934 9376
rect 11149 9367 11207 9373
rect 11149 9364 11161 9367
rect 10928 9336 11161 9364
rect 10928 9324 10934 9336
rect 11149 9333 11161 9336
rect 11195 9333 11207 9367
rect 11149 9327 11207 9333
rect 11698 9324 11704 9376
rect 11756 9364 11762 9376
rect 11793 9367 11851 9373
rect 11793 9364 11805 9367
rect 11756 9336 11805 9364
rect 11756 9324 11762 9336
rect 11793 9333 11805 9336
rect 11839 9364 11851 9367
rect 12342 9364 12348 9376
rect 11839 9336 12348 9364
rect 11839 9333 11851 9336
rect 11793 9327 11851 9333
rect 12342 9324 12348 9336
rect 12400 9324 12406 9376
rect 13354 9364 13360 9376
rect 13315 9336 13360 9364
rect 13354 9324 13360 9336
rect 13412 9324 13418 9376
rect 13725 9367 13783 9373
rect 13725 9333 13737 9367
rect 13771 9364 13783 9367
rect 13814 9364 13820 9376
rect 13771 9336 13820 9364
rect 13771 9333 13783 9336
rect 13725 9327 13783 9333
rect 13814 9324 13820 9336
rect 13872 9364 13878 9376
rect 14200 9364 14228 9472
rect 15746 9460 15752 9512
rect 15804 9500 15810 9512
rect 16669 9503 16727 9509
rect 16669 9500 16681 9503
rect 15804 9472 16681 9500
rect 15804 9460 15810 9472
rect 16669 9469 16681 9472
rect 16715 9500 16727 9503
rect 18233 9503 18291 9509
rect 18233 9500 18245 9503
rect 16715 9472 18245 9500
rect 16715 9469 16727 9472
rect 16669 9463 16727 9469
rect 18233 9469 18245 9472
rect 18279 9469 18291 9503
rect 18233 9463 18291 9469
rect 16761 9435 16819 9441
rect 16761 9401 16773 9435
rect 16807 9432 16819 9435
rect 16807 9404 17724 9432
rect 16807 9401 16819 9404
rect 16761 9395 16819 9401
rect 17696 9376 17724 9404
rect 16022 9364 16028 9376
rect 13872 9336 16028 9364
rect 13872 9324 13878 9336
rect 16022 9324 16028 9336
rect 16080 9364 16086 9376
rect 16117 9367 16175 9373
rect 16117 9364 16129 9367
rect 16080 9336 16129 9364
rect 16080 9324 16086 9336
rect 16117 9333 16129 9336
rect 16163 9364 16175 9367
rect 16666 9364 16672 9376
rect 16163 9336 16672 9364
rect 16163 9333 16175 9336
rect 16117 9327 16175 9333
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 17678 9364 17684 9376
rect 17639 9336 17684 9364
rect 17678 9324 17684 9336
rect 17736 9324 17742 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2866 9160 2872 9172
rect 2827 9132 2872 9160
rect 2866 9120 2872 9132
rect 2924 9120 2930 9172
rect 3510 9160 3516 9172
rect 3471 9132 3516 9160
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 4525 9163 4583 9169
rect 4525 9129 4537 9163
rect 4571 9160 4583 9163
rect 4706 9160 4712 9172
rect 4571 9132 4712 9160
rect 4571 9129 4583 9132
rect 4525 9123 4583 9129
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 6454 9120 6460 9172
rect 6512 9160 6518 9172
rect 6638 9160 6644 9172
rect 6512 9132 6644 9160
rect 6512 9120 6518 9132
rect 6638 9120 6644 9132
rect 6696 9120 6702 9172
rect 7742 9160 7748 9172
rect 7703 9132 7748 9160
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 8478 9120 8484 9172
rect 8536 9160 8542 9172
rect 8665 9163 8723 9169
rect 8665 9160 8677 9163
rect 8536 9132 8677 9160
rect 8536 9120 8542 9132
rect 8665 9129 8677 9132
rect 8711 9129 8723 9163
rect 8665 9123 8723 9129
rect 10778 9120 10784 9172
rect 10836 9160 10842 9172
rect 11241 9163 11299 9169
rect 11241 9160 11253 9163
rect 10836 9132 11253 9160
rect 10836 9120 10842 9132
rect 11241 9129 11253 9132
rect 11287 9160 11299 9163
rect 12066 9160 12072 9172
rect 11287 9132 12072 9160
rect 11287 9129 11299 9132
rect 11241 9123 11299 9129
rect 12066 9120 12072 9132
rect 12124 9120 12130 9172
rect 16114 9120 16120 9172
rect 16172 9160 16178 9172
rect 16393 9163 16451 9169
rect 16393 9160 16405 9163
rect 16172 9132 16405 9160
rect 16172 9120 16178 9132
rect 16393 9129 16405 9132
rect 16439 9129 16451 9163
rect 16393 9123 16451 9129
rect 4430 9092 4436 9104
rect 4391 9064 4436 9092
rect 4430 9052 4436 9064
rect 4488 9052 4494 9104
rect 9674 9052 9680 9104
rect 9732 9092 9738 9104
rect 10137 9095 10195 9101
rect 10137 9092 10149 9095
rect 9732 9064 10149 9092
rect 9732 9052 9738 9064
rect 10137 9061 10149 9064
rect 10183 9092 10195 9095
rect 10962 9092 10968 9104
rect 10183 9064 10968 9092
rect 10183 9061 10195 9064
rect 10137 9055 10195 9061
rect 10962 9052 10968 9064
rect 11020 9052 11026 9104
rect 14918 9092 14924 9104
rect 14879 9064 14924 9092
rect 14918 9052 14924 9064
rect 14976 9052 14982 9104
rect 16844 9095 16902 9101
rect 16844 9061 16856 9095
rect 16890 9092 16902 9095
rect 17402 9092 17408 9104
rect 16890 9064 17408 9092
rect 16890 9061 16902 9064
rect 16844 9055 16902 9061
rect 17402 9052 17408 9064
rect 17460 9052 17466 9104
rect 1756 9027 1814 9033
rect 1756 8993 1768 9027
rect 1802 9024 1814 9027
rect 6365 9027 6423 9033
rect 1802 8996 3372 9024
rect 1802 8993 1814 8996
rect 1756 8987 1814 8993
rect 3344 8968 3372 8996
rect 6365 8993 6377 9027
rect 6411 9024 6423 9027
rect 6454 9024 6460 9036
rect 6411 8996 6460 9024
rect 6411 8993 6423 8996
rect 6365 8987 6423 8993
rect 6454 8984 6460 8996
rect 6512 8984 6518 9036
rect 6632 9027 6690 9033
rect 6632 8993 6644 9027
rect 6678 9024 6690 9027
rect 7558 9024 7564 9036
rect 6678 8996 7564 9024
rect 6678 8993 6690 8996
rect 6632 8987 6690 8993
rect 7558 8984 7564 8996
rect 7616 8984 7622 9036
rect 9950 8984 9956 9036
rect 10008 9024 10014 9036
rect 10045 9027 10103 9033
rect 10045 9024 10057 9027
rect 10008 8996 10057 9024
rect 10008 8984 10014 8996
rect 10045 8993 10057 8996
rect 10091 8993 10103 9027
rect 10045 8987 10103 8993
rect 11882 8984 11888 9036
rect 11940 9024 11946 9036
rect 12049 9027 12107 9033
rect 12049 9024 12061 9027
rect 11940 8996 12061 9024
rect 11940 8984 11946 8996
rect 12049 8993 12061 8996
rect 12095 9024 12107 9027
rect 12342 9024 12348 9036
rect 12095 8996 12348 9024
rect 12095 8993 12107 8996
rect 12049 8987 12107 8993
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 16577 9027 16635 9033
rect 16577 8993 16589 9027
rect 16623 9024 16635 9027
rect 16666 9024 16672 9036
rect 16623 8996 16672 9024
rect 16623 8993 16635 8996
rect 16577 8987 16635 8993
rect 16666 8984 16672 8996
rect 16724 8984 16730 9036
rect 1489 8959 1547 8965
rect 1489 8925 1501 8959
rect 1535 8925 1547 8959
rect 1489 8919 1547 8925
rect 1504 8820 1532 8919
rect 3326 8916 3332 8968
rect 3384 8956 3390 8968
rect 3878 8956 3884 8968
rect 3384 8928 3884 8956
rect 3384 8916 3390 8928
rect 3878 8916 3884 8928
rect 3936 8956 3942 8968
rect 4614 8956 4620 8968
rect 3936 8928 4476 8956
rect 4575 8928 4620 8956
rect 3936 8916 3942 8928
rect 4062 8888 4068 8900
rect 4023 8860 4068 8888
rect 4062 8848 4068 8860
rect 4120 8848 4126 8900
rect 4448 8888 4476 8928
rect 4614 8916 4620 8928
rect 4672 8956 4678 8968
rect 5077 8959 5135 8965
rect 5077 8956 5089 8959
rect 4672 8928 5089 8956
rect 4672 8916 4678 8928
rect 5077 8925 5089 8928
rect 5123 8925 5135 8959
rect 5534 8956 5540 8968
rect 5495 8928 5540 8956
rect 5077 8919 5135 8925
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 10226 8916 10232 8968
rect 10284 8956 10290 8968
rect 11790 8956 11796 8968
rect 10284 8928 10329 8956
rect 11751 8928 11796 8956
rect 10284 8916 10290 8928
rect 11790 8916 11796 8928
rect 11848 8916 11854 8968
rect 15286 8916 15292 8968
rect 15344 8956 15350 8968
rect 15565 8959 15623 8965
rect 15565 8956 15577 8959
rect 15344 8928 15577 8956
rect 15344 8916 15350 8928
rect 15565 8925 15577 8928
rect 15611 8925 15623 8959
rect 15565 8919 15623 8925
rect 9125 8891 9183 8897
rect 4448 8860 6316 8888
rect 2130 8820 2136 8832
rect 1504 8792 2136 8820
rect 2130 8780 2136 8792
rect 2188 8780 2194 8832
rect 5534 8780 5540 8832
rect 5592 8820 5598 8832
rect 6288 8829 6316 8860
rect 9125 8857 9137 8891
rect 9171 8888 9183 8891
rect 9306 8888 9312 8900
rect 9171 8860 9312 8888
rect 9171 8857 9183 8860
rect 9125 8851 9183 8857
rect 9306 8848 9312 8860
rect 9364 8888 9370 8900
rect 9493 8891 9551 8897
rect 9493 8888 9505 8891
rect 9364 8860 9505 8888
rect 9364 8848 9370 8860
rect 9493 8857 9505 8860
rect 9539 8888 9551 8891
rect 10244 8888 10272 8916
rect 9539 8860 10272 8888
rect 9539 8857 9551 8860
rect 9493 8851 9551 8857
rect 5813 8823 5871 8829
rect 5813 8820 5825 8823
rect 5592 8792 5825 8820
rect 5592 8780 5598 8792
rect 5813 8789 5825 8792
rect 5859 8789 5871 8823
rect 5813 8783 5871 8789
rect 6273 8823 6331 8829
rect 6273 8789 6285 8823
rect 6319 8820 6331 8823
rect 7374 8820 7380 8832
rect 6319 8792 7380 8820
rect 6319 8789 6331 8792
rect 6273 8783 6331 8789
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 8386 8820 8392 8832
rect 8347 8792 8392 8820
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 9677 8823 9735 8829
rect 9677 8789 9689 8823
rect 9723 8820 9735 8823
rect 10042 8820 10048 8832
rect 9723 8792 10048 8820
rect 9723 8789 9735 8792
rect 9677 8783 9735 8789
rect 10042 8780 10048 8792
rect 10100 8780 10106 8832
rect 10870 8820 10876 8832
rect 10831 8792 10876 8820
rect 10870 8780 10876 8792
rect 10928 8780 10934 8832
rect 11606 8820 11612 8832
rect 11567 8792 11612 8820
rect 11606 8780 11612 8792
rect 11664 8780 11670 8832
rect 13170 8820 13176 8832
rect 13131 8792 13176 8820
rect 13170 8780 13176 8792
rect 13228 8780 13234 8832
rect 13906 8820 13912 8832
rect 13867 8792 13912 8820
rect 13906 8780 13912 8792
rect 13964 8780 13970 8832
rect 14182 8820 14188 8832
rect 14143 8792 14188 8820
rect 14182 8780 14188 8792
rect 14240 8780 14246 8832
rect 14550 8820 14556 8832
rect 14511 8792 14556 8820
rect 14550 8780 14556 8792
rect 14608 8780 14614 8832
rect 15654 8780 15660 8832
rect 15712 8820 15718 8832
rect 16117 8823 16175 8829
rect 16117 8820 16129 8823
rect 15712 8792 16129 8820
rect 15712 8780 15718 8792
rect 16117 8789 16129 8792
rect 16163 8820 16175 8823
rect 16482 8820 16488 8832
rect 16163 8792 16488 8820
rect 16163 8789 16175 8792
rect 16117 8783 16175 8789
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 17954 8820 17960 8832
rect 17915 8792 17960 8820
rect 17954 8780 17960 8792
rect 18012 8780 18018 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 2685 8619 2743 8625
rect 2685 8616 2697 8619
rect 2372 8588 2697 8616
rect 2372 8576 2378 8588
rect 2685 8585 2697 8588
rect 2731 8585 2743 8619
rect 2685 8579 2743 8585
rect 6270 8576 6276 8628
rect 6328 8616 6334 8628
rect 6825 8619 6883 8625
rect 6825 8616 6837 8619
rect 6328 8588 6837 8616
rect 6328 8576 6334 8588
rect 6825 8585 6837 8588
rect 6871 8585 6883 8619
rect 6825 8579 6883 8585
rect 7558 8576 7564 8628
rect 7616 8616 7622 8628
rect 7837 8619 7895 8625
rect 7837 8616 7849 8619
rect 7616 8588 7849 8616
rect 7616 8576 7622 8588
rect 7837 8585 7849 8588
rect 7883 8585 7895 8619
rect 7837 8579 7895 8585
rect 10045 8619 10103 8625
rect 10045 8585 10057 8619
rect 10091 8616 10103 8619
rect 10226 8616 10232 8628
rect 10091 8588 10232 8616
rect 10091 8585 10103 8588
rect 10045 8579 10103 8585
rect 10226 8576 10232 8588
rect 10284 8616 10290 8628
rect 10597 8619 10655 8625
rect 10597 8616 10609 8619
rect 10284 8588 10609 8616
rect 10284 8576 10290 8588
rect 10597 8585 10609 8588
rect 10643 8585 10655 8619
rect 10597 8579 10655 8585
rect 13906 8576 13912 8628
rect 13964 8616 13970 8628
rect 14369 8619 14427 8625
rect 14369 8616 14381 8619
rect 13964 8588 14381 8616
rect 13964 8576 13970 8588
rect 14369 8585 14381 8588
rect 14415 8585 14427 8619
rect 15286 8616 15292 8628
rect 15247 8588 15292 8616
rect 14369 8579 14427 8585
rect 15286 8576 15292 8588
rect 15344 8576 15350 8628
rect 15470 8576 15476 8628
rect 15528 8616 15534 8628
rect 15565 8619 15623 8625
rect 15565 8616 15577 8619
rect 15528 8588 15577 8616
rect 15528 8576 15534 8588
rect 15565 8585 15577 8588
rect 15611 8585 15623 8619
rect 15746 8616 15752 8628
rect 15707 8588 15752 8616
rect 15565 8579 15623 8585
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 2222 8480 2228 8492
rect 1719 8452 2228 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 2222 8440 2228 8452
rect 2280 8440 2286 8492
rect 3326 8480 3332 8492
rect 3287 8452 3332 8480
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 7374 8480 7380 8492
rect 7335 8452 7380 8480
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 10870 8440 10876 8492
rect 10928 8480 10934 8492
rect 11333 8483 11391 8489
rect 11333 8480 11345 8483
rect 10928 8452 11345 8480
rect 10928 8440 10934 8452
rect 11333 8449 11345 8452
rect 11379 8449 11391 8483
rect 11333 8443 11391 8449
rect 4157 8415 4215 8421
rect 4157 8412 4169 8415
rect 2148 8384 4169 8412
rect 2148 8356 2176 8384
rect 4157 8381 4169 8384
rect 4203 8412 4215 8415
rect 4249 8415 4307 8421
rect 4249 8412 4261 8415
rect 4203 8384 4261 8412
rect 4203 8381 4215 8384
rect 4157 8375 4215 8381
rect 4249 8381 4261 8384
rect 4295 8412 4307 8415
rect 6641 8415 6699 8421
rect 4295 8384 6316 8412
rect 4295 8381 4307 8384
rect 4249 8375 4307 8381
rect 2130 8344 2136 8356
rect 2091 8316 2136 8344
rect 2130 8304 2136 8316
rect 2188 8304 2194 8356
rect 3053 8347 3111 8353
rect 3053 8344 3065 8347
rect 2608 8316 3065 8344
rect 2608 8288 2636 8316
rect 3053 8313 3065 8316
rect 3099 8313 3111 8347
rect 3053 8307 3111 8313
rect 3789 8347 3847 8353
rect 3789 8313 3801 8347
rect 3835 8344 3847 8347
rect 4494 8347 4552 8353
rect 4494 8344 4506 8347
rect 3835 8316 4506 8344
rect 3835 8313 3847 8316
rect 3789 8307 3847 8313
rect 4494 8313 4506 8316
rect 4540 8344 4552 8347
rect 4614 8344 4620 8356
rect 4540 8316 4620 8344
rect 4540 8313 4552 8316
rect 4494 8307 4552 8313
rect 4614 8304 4620 8316
rect 4672 8304 4678 8356
rect 2590 8276 2596 8288
rect 2551 8248 2596 8276
rect 2590 8236 2596 8248
rect 2648 8236 2654 8288
rect 3142 8276 3148 8288
rect 3103 8248 3148 8276
rect 3142 8236 3148 8248
rect 3200 8236 3206 8288
rect 5534 8236 5540 8288
rect 5592 8276 5598 8288
rect 6288 8285 6316 8384
rect 6641 8381 6653 8415
rect 6687 8412 6699 8415
rect 7190 8412 7196 8424
rect 6687 8384 7196 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 7190 8372 7196 8384
rect 7248 8372 7254 8424
rect 8573 8415 8631 8421
rect 8573 8381 8585 8415
rect 8619 8412 8631 8415
rect 8665 8415 8723 8421
rect 8665 8412 8677 8415
rect 8619 8384 8677 8412
rect 8619 8381 8631 8384
rect 8573 8375 8631 8381
rect 8665 8381 8677 8384
rect 8711 8412 8723 8415
rect 9398 8412 9404 8424
rect 8711 8384 9404 8412
rect 8711 8381 8723 8384
rect 8665 8375 8723 8381
rect 9398 8372 9404 8384
rect 9456 8412 9462 8424
rect 12989 8415 13047 8421
rect 9456 8384 11836 8412
rect 9456 8372 9462 8384
rect 11808 8356 11836 8384
rect 12989 8381 13001 8415
rect 13035 8412 13047 8415
rect 13814 8412 13820 8424
rect 13035 8384 13820 8412
rect 13035 8381 13047 8384
rect 12989 8375 13047 8381
rect 7098 8304 7104 8356
rect 7156 8344 7162 8356
rect 7466 8344 7472 8356
rect 7156 8316 7472 8344
rect 7156 8304 7162 8316
rect 7466 8304 7472 8316
rect 7524 8304 7530 8356
rect 8478 8304 8484 8356
rect 8536 8344 8542 8356
rect 8910 8347 8968 8353
rect 8910 8344 8922 8347
rect 8536 8316 8922 8344
rect 8536 8304 8542 8316
rect 8910 8313 8922 8316
rect 8956 8313 8968 8347
rect 8910 8307 8968 8313
rect 11057 8347 11115 8353
rect 11057 8313 11069 8347
rect 11103 8344 11115 8347
rect 11422 8344 11428 8356
rect 11103 8316 11428 8344
rect 11103 8313 11115 8316
rect 11057 8307 11115 8313
rect 11422 8304 11428 8316
rect 11480 8304 11486 8356
rect 11790 8304 11796 8356
rect 11848 8344 11854 8356
rect 11885 8347 11943 8353
rect 11885 8344 11897 8347
rect 11848 8316 11897 8344
rect 11848 8304 11854 8316
rect 11885 8313 11897 8316
rect 11931 8344 11943 8347
rect 12897 8347 12955 8353
rect 12897 8344 12909 8347
rect 11931 8316 12909 8344
rect 11931 8313 11943 8316
rect 11885 8307 11943 8313
rect 12897 8313 12909 8316
rect 12943 8344 12955 8347
rect 13004 8344 13032 8375
rect 13814 8372 13820 8384
rect 13872 8372 13878 8424
rect 15304 8412 15332 8576
rect 15580 8480 15608 8579
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 17221 8619 17279 8625
rect 17221 8585 17233 8619
rect 17267 8616 17279 8619
rect 17402 8616 17408 8628
rect 17267 8588 17408 8616
rect 17267 8585 17279 8588
rect 17221 8579 17279 8585
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 16206 8480 16212 8492
rect 15580 8452 16212 8480
rect 16206 8440 16212 8452
rect 16264 8440 16270 8492
rect 16393 8483 16451 8489
rect 16393 8449 16405 8483
rect 16439 8480 16451 8483
rect 16482 8480 16488 8492
rect 16439 8452 16488 8480
rect 16439 8449 16451 8452
rect 16393 8443 16451 8449
rect 16482 8440 16488 8452
rect 16540 8440 16546 8492
rect 16117 8415 16175 8421
rect 16117 8412 16129 8415
rect 15304 8384 16129 8412
rect 16117 8381 16129 8384
rect 16163 8381 16175 8415
rect 16117 8375 16175 8381
rect 12943 8316 13032 8344
rect 12943 8313 12955 8316
rect 12897 8307 12955 8313
rect 13170 8304 13176 8356
rect 13228 8353 13234 8356
rect 13228 8347 13292 8353
rect 13228 8313 13246 8347
rect 13280 8313 13292 8347
rect 17494 8344 17500 8356
rect 17455 8316 17500 8344
rect 13228 8307 13292 8313
rect 13228 8304 13234 8307
rect 17494 8304 17500 8316
rect 17552 8304 17558 8356
rect 5629 8279 5687 8285
rect 5629 8276 5641 8279
rect 5592 8248 5641 8276
rect 5592 8236 5598 8248
rect 5629 8245 5641 8248
rect 5675 8245 5687 8279
rect 5629 8239 5687 8245
rect 6273 8279 6331 8285
rect 6273 8245 6285 8279
rect 6319 8276 6331 8279
rect 6454 8276 6460 8288
rect 6319 8248 6460 8276
rect 6319 8245 6331 8248
rect 6273 8239 6331 8245
rect 6454 8236 6460 8248
rect 6512 8276 6518 8288
rect 6822 8276 6828 8288
rect 6512 8248 6828 8276
rect 6512 8236 6518 8248
rect 6822 8236 6828 8248
rect 6880 8236 6886 8288
rect 6914 8236 6920 8288
rect 6972 8276 6978 8288
rect 7285 8279 7343 8285
rect 7285 8276 7297 8279
rect 6972 8248 7297 8276
rect 6972 8236 6978 8248
rect 7285 8245 7297 8248
rect 7331 8245 7343 8279
rect 7285 8239 7343 8245
rect 12253 8279 12311 8285
rect 12253 8245 12265 8279
rect 12299 8276 12311 8279
rect 12434 8276 12440 8288
rect 12299 8248 12440 8276
rect 12299 8245 12311 8248
rect 12253 8239 12311 8245
rect 12434 8236 12440 8248
rect 12492 8236 12498 8288
rect 16666 8236 16672 8288
rect 16724 8276 16730 8288
rect 16761 8279 16819 8285
rect 16761 8276 16773 8279
rect 16724 8248 16773 8276
rect 16724 8236 16730 8248
rect 16761 8245 16773 8248
rect 16807 8245 16819 8279
rect 16761 8239 16819 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1762 8072 1768 8084
rect 1723 8044 1768 8072
rect 1762 8032 1768 8044
rect 1820 8072 1826 8084
rect 2222 8072 2228 8084
rect 1820 8044 2228 8072
rect 1820 8032 1826 8044
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 2777 8075 2835 8081
rect 2777 8041 2789 8075
rect 2823 8072 2835 8075
rect 3142 8072 3148 8084
rect 2823 8044 3148 8072
rect 2823 8041 2835 8044
rect 2777 8035 2835 8041
rect 3142 8032 3148 8044
rect 3200 8032 3206 8084
rect 5905 8075 5963 8081
rect 5905 8041 5917 8075
rect 5951 8072 5963 8075
rect 7190 8072 7196 8084
rect 5951 8044 7196 8072
rect 5951 8041 5963 8044
rect 5905 8035 5963 8041
rect 7190 8032 7196 8044
rect 7248 8072 7254 8084
rect 9401 8075 9459 8081
rect 9401 8072 9413 8075
rect 7248 8044 9413 8072
rect 7248 8032 7254 8044
rect 9401 8041 9413 8044
rect 9447 8041 9459 8075
rect 9674 8072 9680 8084
rect 9635 8044 9680 8072
rect 9401 8035 9459 8041
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 11698 8072 11704 8084
rect 11659 8044 11704 8072
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 12066 8072 12072 8084
rect 12027 8044 12072 8072
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 13262 8072 13268 8084
rect 13223 8044 13268 8072
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 13354 8032 13360 8084
rect 13412 8072 13418 8084
rect 13633 8075 13691 8081
rect 13633 8072 13645 8075
rect 13412 8044 13645 8072
rect 13412 8032 13418 8044
rect 13633 8041 13645 8044
rect 13679 8041 13691 8075
rect 13633 8035 13691 8041
rect 16206 8032 16212 8084
rect 16264 8072 16270 8084
rect 16577 8075 16635 8081
rect 16577 8072 16589 8075
rect 16264 8044 16589 8072
rect 16264 8032 16270 8044
rect 16577 8041 16589 8044
rect 16623 8072 16635 8075
rect 16758 8072 16764 8084
rect 16623 8044 16764 8072
rect 16623 8041 16635 8044
rect 16577 8035 16635 8041
rect 16758 8032 16764 8044
rect 16816 8032 16822 8084
rect 17678 8072 17684 8084
rect 17639 8044 17684 8072
rect 17678 8032 17684 8044
rect 17736 8032 17742 8084
rect 4706 8004 4712 8016
rect 4619 7976 4712 8004
rect 4706 7964 4712 7976
rect 4764 8004 4770 8016
rect 4764 7976 5120 8004
rect 4764 7964 4770 7976
rect 4801 7939 4859 7945
rect 4801 7905 4813 7939
rect 4847 7936 4859 7939
rect 4982 7936 4988 7948
rect 4847 7908 4988 7936
rect 4847 7905 4859 7908
rect 4801 7899 4859 7905
rect 1578 7828 1584 7880
rect 1636 7868 1642 7880
rect 1857 7871 1915 7877
rect 1857 7868 1869 7871
rect 1636 7840 1869 7868
rect 1636 7828 1642 7840
rect 1857 7837 1869 7840
rect 1903 7837 1915 7871
rect 2038 7868 2044 7880
rect 1999 7840 2044 7868
rect 1857 7831 1915 7837
rect 2038 7828 2044 7840
rect 2096 7828 2102 7880
rect 3881 7871 3939 7877
rect 3881 7837 3893 7871
rect 3927 7868 3939 7871
rect 4522 7868 4528 7880
rect 3927 7840 4528 7868
rect 3927 7837 3939 7840
rect 3881 7831 3939 7837
rect 4522 7828 4528 7840
rect 4580 7868 4586 7880
rect 4816 7868 4844 7899
rect 4982 7896 4988 7908
rect 5040 7896 5046 7948
rect 4580 7840 4844 7868
rect 4893 7871 4951 7877
rect 4580 7828 4586 7840
rect 4893 7837 4905 7871
rect 4939 7837 4951 7871
rect 5092 7868 5120 7976
rect 5166 7964 5172 8016
rect 5224 8004 5230 8016
rect 6365 8007 6423 8013
rect 6365 8004 6377 8007
rect 5224 7976 6377 8004
rect 5224 7964 5230 7976
rect 6365 7973 6377 7976
rect 6411 8004 6423 8007
rect 9033 8007 9091 8013
rect 9033 8004 9045 8007
rect 6411 7976 9045 8004
rect 6411 7973 6423 7976
rect 6365 7967 6423 7973
rect 9033 7973 9045 7976
rect 9079 7973 9091 8007
rect 9033 7967 9091 7973
rect 12710 7964 12716 8016
rect 12768 8004 12774 8016
rect 13725 8007 13783 8013
rect 13725 8004 13737 8007
rect 12768 7976 13737 8004
rect 12768 7964 12774 7976
rect 13725 7973 13737 7976
rect 13771 8004 13783 8007
rect 14277 8007 14335 8013
rect 14277 8004 14289 8007
rect 13771 7976 14289 8004
rect 13771 7973 13783 7976
rect 13725 7967 13783 7973
rect 14277 7973 14289 7976
rect 14323 7973 14335 8007
rect 14277 7967 14335 7973
rect 6270 7936 6276 7948
rect 6231 7908 6276 7936
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 8110 7936 8116 7948
rect 6380 7908 8116 7936
rect 6380 7868 6408 7908
rect 8110 7896 8116 7908
rect 8168 7896 8174 7948
rect 8294 7896 8300 7948
rect 8352 7936 8358 7948
rect 8389 7939 8447 7945
rect 8389 7936 8401 7939
rect 8352 7908 8401 7936
rect 8352 7896 8358 7908
rect 8389 7905 8401 7908
rect 8435 7905 8447 7939
rect 8389 7899 8447 7905
rect 8481 7939 8539 7945
rect 8481 7905 8493 7939
rect 8527 7905 8539 7939
rect 8481 7899 8539 7905
rect 5092 7840 6408 7868
rect 6549 7871 6607 7877
rect 4893 7831 4951 7837
rect 6549 7837 6561 7871
rect 6595 7868 6607 7871
rect 6595 7840 7144 7868
rect 6595 7837 6607 7840
rect 6549 7831 6607 7837
rect 1397 7735 1455 7741
rect 1397 7701 1409 7735
rect 1443 7732 1455 7735
rect 1854 7732 1860 7744
rect 1443 7704 1860 7732
rect 1443 7701 1455 7704
rect 1397 7695 1455 7701
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 3142 7732 3148 7744
rect 3103 7704 3148 7732
rect 3142 7692 3148 7704
rect 3200 7692 3206 7744
rect 3510 7732 3516 7744
rect 3471 7704 3516 7732
rect 3510 7692 3516 7704
rect 3568 7692 3574 7744
rect 4341 7735 4399 7741
rect 4341 7701 4353 7735
rect 4387 7732 4399 7735
rect 4522 7732 4528 7744
rect 4387 7704 4528 7732
rect 4387 7701 4399 7704
rect 4341 7695 4399 7701
rect 4522 7692 4528 7704
rect 4580 7692 4586 7744
rect 4614 7692 4620 7744
rect 4672 7732 4678 7744
rect 4908 7732 4936 7831
rect 7116 7744 7144 7840
rect 8496 7812 8524 7899
rect 9950 7896 9956 7948
rect 10008 7936 10014 7948
rect 10045 7939 10103 7945
rect 10045 7936 10057 7939
rect 10008 7908 10057 7936
rect 10008 7896 10014 7908
rect 10045 7905 10057 7908
rect 10091 7905 10103 7939
rect 16482 7936 16488 7948
rect 16443 7908 16488 7936
rect 10045 7899 10103 7905
rect 16482 7896 16488 7908
rect 16540 7896 16546 7948
rect 18046 7936 18052 7948
rect 18007 7908 18052 7936
rect 18046 7896 18052 7908
rect 18104 7896 18110 7948
rect 8570 7828 8576 7880
rect 8628 7868 8634 7880
rect 10134 7868 10140 7880
rect 8628 7840 8673 7868
rect 10095 7840 10140 7868
rect 8628 7828 8634 7840
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 8018 7800 8024 7812
rect 7979 7772 8024 7800
rect 8018 7760 8024 7772
rect 8076 7760 8082 7812
rect 8478 7760 8484 7812
rect 8536 7760 8542 7812
rect 8588 7800 8616 7828
rect 9858 7800 9864 7812
rect 8588 7772 9864 7800
rect 9858 7760 9864 7772
rect 9916 7800 9922 7812
rect 10244 7800 10272 7831
rect 10778 7828 10784 7880
rect 10836 7868 10842 7880
rect 11606 7868 11612 7880
rect 10836 7840 11612 7868
rect 10836 7828 10842 7840
rect 11606 7828 11612 7840
rect 11664 7868 11670 7880
rect 12161 7871 12219 7877
rect 12161 7868 12173 7871
rect 11664 7840 12173 7868
rect 11664 7828 11670 7840
rect 12161 7837 12173 7840
rect 12207 7837 12219 7871
rect 12161 7831 12219 7837
rect 12250 7828 12256 7880
rect 12308 7868 12314 7880
rect 13081 7871 13139 7877
rect 13081 7868 13093 7871
rect 12308 7840 13093 7868
rect 12308 7828 12314 7840
rect 13081 7837 13093 7840
rect 13127 7868 13139 7871
rect 13170 7868 13176 7880
rect 13127 7840 13176 7868
rect 13127 7837 13139 7840
rect 13081 7831 13139 7837
rect 13170 7828 13176 7840
rect 13228 7868 13234 7880
rect 13906 7868 13912 7880
rect 13228 7840 13912 7868
rect 13228 7828 13234 7840
rect 13906 7828 13912 7840
rect 13964 7828 13970 7880
rect 16390 7828 16396 7880
rect 16448 7868 16454 7880
rect 16669 7871 16727 7877
rect 16669 7868 16681 7871
rect 16448 7840 16681 7868
rect 16448 7828 16454 7840
rect 16669 7837 16681 7840
rect 16715 7837 16727 7871
rect 18138 7868 18144 7880
rect 18099 7840 18144 7868
rect 16669 7831 16727 7837
rect 18138 7828 18144 7840
rect 18196 7828 18202 7880
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7837 18291 7871
rect 18233 7831 18291 7837
rect 9916 7772 10272 7800
rect 14737 7803 14795 7809
rect 9916 7760 9922 7772
rect 14737 7769 14749 7803
rect 14783 7800 14795 7803
rect 15562 7800 15568 7812
rect 14783 7772 15568 7800
rect 14783 7769 14795 7772
rect 14737 7763 14795 7769
rect 15562 7760 15568 7772
rect 15620 7800 15626 7812
rect 16117 7803 16175 7809
rect 16117 7800 16129 7803
rect 15620 7772 16129 7800
rect 15620 7760 15626 7772
rect 16117 7769 16129 7772
rect 16163 7769 16175 7803
rect 16117 7763 16175 7769
rect 16574 7760 16580 7812
rect 16632 7800 16638 7812
rect 17589 7803 17647 7809
rect 17589 7800 17601 7803
rect 16632 7772 17601 7800
rect 16632 7760 16638 7772
rect 17589 7769 17601 7772
rect 17635 7800 17647 7803
rect 18248 7800 18276 7831
rect 17635 7772 18276 7800
rect 19705 7803 19763 7809
rect 17635 7769 17647 7772
rect 17589 7763 17647 7769
rect 19705 7769 19717 7803
rect 19751 7800 19763 7803
rect 20070 7800 20076 7812
rect 19751 7772 20076 7800
rect 19751 7769 19763 7772
rect 19705 7763 19763 7769
rect 20070 7760 20076 7772
rect 20128 7760 20134 7812
rect 5353 7735 5411 7741
rect 5353 7732 5365 7735
rect 4672 7704 5365 7732
rect 4672 7692 4678 7704
rect 5353 7701 5365 7704
rect 5399 7701 5411 7735
rect 5353 7695 5411 7701
rect 5813 7735 5871 7741
rect 5813 7701 5825 7735
rect 5859 7732 5871 7735
rect 6086 7732 6092 7744
rect 5859 7704 6092 7732
rect 5859 7701 5871 7704
rect 5813 7695 5871 7701
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 6914 7732 6920 7744
rect 6875 7704 6920 7732
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 7098 7692 7104 7744
rect 7156 7732 7162 7744
rect 7285 7735 7343 7741
rect 7285 7732 7297 7735
rect 7156 7704 7297 7732
rect 7156 7692 7162 7704
rect 7285 7701 7297 7704
rect 7331 7732 7343 7735
rect 7653 7735 7711 7741
rect 7653 7732 7665 7735
rect 7331 7704 7665 7732
rect 7331 7701 7343 7704
rect 7285 7695 7343 7701
rect 7653 7701 7665 7704
rect 7699 7701 7711 7735
rect 10870 7732 10876 7744
rect 10831 7704 10876 7732
rect 7653 7695 7711 7701
rect 10870 7692 10876 7704
rect 10928 7692 10934 7744
rect 11238 7732 11244 7744
rect 11199 7704 11244 7732
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 11330 7692 11336 7744
rect 11388 7732 11394 7744
rect 11517 7735 11575 7741
rect 11517 7732 11529 7735
rect 11388 7704 11529 7732
rect 11388 7692 11394 7704
rect 11517 7701 11529 7704
rect 11563 7701 11575 7735
rect 11517 7695 11575 7701
rect 15105 7735 15163 7741
rect 15105 7701 15117 7735
rect 15151 7732 15163 7735
rect 15654 7732 15660 7744
rect 15151 7704 15660 7732
rect 15151 7701 15163 7704
rect 15105 7695 15163 7701
rect 15654 7692 15660 7704
rect 15712 7692 15718 7744
rect 15746 7692 15752 7744
rect 15804 7732 15810 7744
rect 15804 7704 15849 7732
rect 15804 7692 15810 7704
rect 16850 7692 16856 7744
rect 16908 7732 16914 7744
rect 17129 7735 17187 7741
rect 17129 7732 17141 7735
rect 16908 7704 17141 7732
rect 16908 7692 16914 7704
rect 17129 7701 17141 7704
rect 17175 7701 17187 7735
rect 19978 7732 19984 7744
rect 19939 7704 19984 7732
rect 17129 7695 17187 7701
rect 19978 7692 19984 7704
rect 20036 7692 20042 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1394 7528 1400 7540
rect 1355 7500 1400 7528
rect 1394 7488 1400 7500
rect 1452 7488 1458 7540
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 4985 7531 5043 7537
rect 4985 7528 4997 7531
rect 4212 7500 4997 7528
rect 4212 7488 4218 7500
rect 4985 7497 4997 7500
rect 5031 7497 5043 7531
rect 5166 7528 5172 7540
rect 5127 7500 5172 7528
rect 4985 7491 5043 7497
rect 3605 7463 3663 7469
rect 3605 7429 3617 7463
rect 3651 7460 3663 7463
rect 4430 7460 4436 7472
rect 3651 7432 4436 7460
rect 3651 7429 3663 7432
rect 3605 7423 3663 7429
rect 4430 7420 4436 7432
rect 4488 7420 4494 7472
rect 4706 7460 4712 7472
rect 4667 7432 4712 7460
rect 4706 7420 4712 7432
rect 4764 7420 4770 7472
rect 2038 7392 2044 7404
rect 1999 7364 2044 7392
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 3510 7352 3516 7404
rect 3568 7392 3574 7404
rect 4249 7395 4307 7401
rect 4249 7392 4261 7395
rect 3568 7364 4261 7392
rect 3568 7352 3574 7364
rect 4249 7361 4261 7364
rect 4295 7392 4307 7395
rect 4614 7392 4620 7404
rect 4295 7364 4620 7392
rect 4295 7361 4307 7364
rect 4249 7355 4307 7361
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 1857 7327 1915 7333
rect 1857 7293 1869 7327
rect 1903 7324 1915 7327
rect 1946 7324 1952 7336
rect 1903 7296 1952 7324
rect 1903 7293 1915 7296
rect 1857 7287 1915 7293
rect 1946 7284 1952 7296
rect 2004 7284 2010 7336
rect 5000 7324 5028 7491
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 7558 7488 7564 7540
rect 7616 7528 7622 7540
rect 8205 7531 8263 7537
rect 8205 7528 8217 7531
rect 7616 7500 8217 7528
rect 7616 7488 7622 7500
rect 8205 7497 8217 7500
rect 8251 7497 8263 7531
rect 8205 7491 8263 7497
rect 8478 7488 8484 7540
rect 8536 7528 8542 7540
rect 8757 7531 8815 7537
rect 8757 7528 8769 7531
rect 8536 7500 8769 7528
rect 8536 7488 8542 7500
rect 8757 7497 8769 7500
rect 8803 7497 8815 7531
rect 10778 7528 10784 7540
rect 10739 7500 10784 7528
rect 8757 7491 8815 7497
rect 10778 7488 10784 7500
rect 10836 7488 10842 7540
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 12250 7528 12256 7540
rect 11931 7500 12256 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 13354 7488 13360 7540
rect 13412 7528 13418 7540
rect 13633 7531 13691 7537
rect 13633 7528 13645 7531
rect 13412 7500 13645 7528
rect 13412 7488 13418 7500
rect 13633 7497 13645 7500
rect 13679 7497 13691 7531
rect 13633 7491 13691 7497
rect 15654 7488 15660 7540
rect 15712 7528 15718 7540
rect 15749 7531 15807 7537
rect 15749 7528 15761 7531
rect 15712 7500 15761 7528
rect 15712 7488 15718 7500
rect 15749 7497 15761 7500
rect 15795 7497 15807 7531
rect 16758 7528 16764 7540
rect 16719 7500 16764 7528
rect 15749 7491 15807 7497
rect 16758 7488 16764 7500
rect 16816 7488 16822 7540
rect 8570 7420 8576 7472
rect 8628 7460 8634 7472
rect 9125 7463 9183 7469
rect 9125 7460 9137 7463
rect 8628 7432 9137 7460
rect 8628 7420 8634 7432
rect 9125 7429 9137 7432
rect 9171 7429 9183 7463
rect 9125 7423 9183 7429
rect 13173 7463 13231 7469
rect 13173 7429 13185 7463
rect 13219 7460 13231 7463
rect 17313 7463 17371 7469
rect 17313 7460 17325 7463
rect 13219 7432 14320 7460
rect 13219 7429 13231 7432
rect 13173 7423 13231 7429
rect 5810 7392 5816 7404
rect 5771 7364 5816 7392
rect 5810 7352 5816 7364
rect 5868 7392 5874 7404
rect 6086 7392 6092 7404
rect 5868 7364 6092 7392
rect 5868 7352 5874 7364
rect 6086 7352 6092 7364
rect 6144 7352 6150 7404
rect 10870 7352 10876 7404
rect 10928 7392 10934 7404
rect 11333 7395 11391 7401
rect 11333 7392 11345 7395
rect 10928 7364 11345 7392
rect 10928 7352 10934 7364
rect 11333 7361 11345 7364
rect 11379 7392 11391 7395
rect 12434 7392 12440 7404
rect 11379 7364 12440 7392
rect 11379 7361 11391 7364
rect 11333 7355 11391 7361
rect 12434 7352 12440 7364
rect 12492 7392 12498 7404
rect 13188 7392 13216 7423
rect 14292 7404 14320 7432
rect 16224 7432 17325 7460
rect 12492 7364 13216 7392
rect 13541 7395 13599 7401
rect 12492 7352 12498 7364
rect 13541 7361 13553 7395
rect 13587 7392 13599 7395
rect 13630 7392 13636 7404
rect 13587 7364 13636 7392
rect 13587 7361 13599 7364
rect 13541 7355 13599 7361
rect 13630 7352 13636 7364
rect 13688 7392 13694 7404
rect 13688 7364 14044 7392
rect 13688 7352 13694 7364
rect 5537 7327 5595 7333
rect 5537 7324 5549 7327
rect 5000 7296 5549 7324
rect 5537 7293 5549 7296
rect 5583 7324 5595 7327
rect 5994 7324 6000 7336
rect 5583 7296 6000 7324
rect 5583 7293 5595 7296
rect 5537 7287 5595 7293
rect 5994 7284 6000 7296
rect 6052 7284 6058 7336
rect 6822 7324 6828 7336
rect 6735 7296 6828 7324
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 9674 7284 9680 7336
rect 9732 7324 9738 7336
rect 10597 7327 10655 7333
rect 10597 7324 10609 7327
rect 9732 7296 10609 7324
rect 9732 7284 9738 7296
rect 10597 7293 10609 7296
rect 10643 7324 10655 7327
rect 11149 7327 11207 7333
rect 11149 7324 11161 7327
rect 10643 7296 11161 7324
rect 10643 7293 10655 7296
rect 10597 7287 10655 7293
rect 11149 7293 11161 7296
rect 11195 7324 11207 7327
rect 11790 7324 11796 7336
rect 11195 7296 11796 7324
rect 11195 7293 11207 7296
rect 11149 7287 11207 7293
rect 11790 7284 11796 7296
rect 11848 7284 11854 7336
rect 12802 7284 12808 7336
rect 12860 7324 12866 7336
rect 13354 7324 13360 7336
rect 12860 7296 13360 7324
rect 12860 7284 12866 7296
rect 13354 7284 13360 7296
rect 13412 7284 13418 7336
rect 14016 7333 14044 7364
rect 14090 7352 14096 7404
rect 14148 7392 14154 7404
rect 14274 7392 14280 7404
rect 14148 7364 14193 7392
rect 14235 7364 14280 7392
rect 14148 7352 14154 7364
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 15746 7352 15752 7404
rect 15804 7392 15810 7404
rect 16224 7401 16252 7432
rect 17313 7429 17325 7432
rect 17359 7460 17371 7463
rect 18138 7460 18144 7472
rect 17359 7432 18144 7460
rect 17359 7429 17371 7432
rect 17313 7423 17371 7429
rect 18138 7420 18144 7432
rect 18196 7420 18202 7472
rect 16209 7395 16267 7401
rect 16209 7392 16221 7395
rect 15804 7364 16221 7392
rect 15804 7352 15810 7364
rect 16209 7361 16221 7364
rect 16255 7361 16267 7395
rect 16390 7392 16396 7404
rect 16351 7364 16396 7392
rect 16209 7355 16267 7361
rect 16390 7352 16396 7364
rect 16448 7352 16454 7404
rect 18690 7392 18696 7404
rect 18651 7364 18696 7392
rect 18690 7352 18696 7364
rect 18748 7352 18754 7404
rect 19334 7352 19340 7404
rect 19392 7392 19398 7404
rect 19521 7395 19579 7401
rect 19521 7392 19533 7395
rect 19392 7364 19533 7392
rect 19392 7352 19398 7364
rect 19521 7361 19533 7364
rect 19567 7392 19579 7395
rect 20165 7395 20223 7401
rect 20165 7392 20177 7395
rect 19567 7364 20177 7392
rect 19567 7361 19579 7364
rect 19521 7355 19579 7361
rect 20165 7361 20177 7364
rect 20211 7361 20223 7395
rect 20165 7355 20223 7361
rect 14001 7327 14059 7333
rect 14001 7293 14013 7327
rect 14047 7324 14059 7327
rect 14550 7324 14556 7336
rect 14047 7296 14556 7324
rect 14047 7293 14059 7296
rect 14001 7287 14059 7293
rect 14550 7284 14556 7296
rect 14608 7284 14614 7336
rect 15470 7284 15476 7336
rect 15528 7324 15534 7336
rect 15565 7327 15623 7333
rect 15565 7324 15577 7327
rect 15528 7296 15577 7324
rect 15528 7284 15534 7296
rect 15565 7293 15577 7296
rect 15611 7324 15623 7327
rect 16117 7327 16175 7333
rect 16117 7324 16129 7327
rect 15611 7296 16129 7324
rect 15611 7293 15623 7296
rect 15565 7287 15623 7293
rect 16117 7293 16129 7296
rect 16163 7324 16175 7327
rect 17681 7327 17739 7333
rect 17681 7324 17693 7327
rect 16163 7296 17693 7324
rect 16163 7293 16175 7296
rect 16117 7287 16175 7293
rect 17681 7293 17693 7296
rect 17727 7324 17739 7327
rect 18046 7324 18052 7336
rect 17727 7296 18052 7324
rect 17727 7293 17739 7296
rect 17681 7287 17739 7293
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 18414 7324 18420 7336
rect 18375 7296 18420 7324
rect 18414 7284 18420 7296
rect 18472 7284 18478 7336
rect 18509 7327 18567 7333
rect 18509 7293 18521 7327
rect 18555 7324 18567 7327
rect 18598 7324 18604 7336
rect 18555 7296 18604 7324
rect 18555 7293 18567 7296
rect 18509 7287 18567 7293
rect 18598 7284 18604 7296
rect 18656 7324 18662 7336
rect 19061 7327 19119 7333
rect 19061 7324 19073 7327
rect 18656 7296 19073 7324
rect 18656 7284 18662 7296
rect 19061 7293 19073 7296
rect 19107 7324 19119 7327
rect 19150 7324 19156 7336
rect 19107 7296 19156 7324
rect 19107 7293 19119 7296
rect 19061 7287 19119 7293
rect 19150 7284 19156 7296
rect 19208 7284 19214 7336
rect 1486 7216 1492 7268
rect 1544 7256 1550 7268
rect 1765 7259 1823 7265
rect 1765 7256 1777 7259
rect 1544 7228 1777 7256
rect 1544 7216 1550 7228
rect 1765 7225 1777 7228
rect 1811 7256 1823 7259
rect 2777 7259 2835 7265
rect 2777 7256 2789 7259
rect 1811 7228 2789 7256
rect 1811 7225 1823 7228
rect 1765 7219 1823 7225
rect 2777 7225 2789 7228
rect 2823 7225 2835 7259
rect 2777 7219 2835 7225
rect 3510 7216 3516 7268
rect 3568 7256 3574 7268
rect 3973 7259 4031 7265
rect 3973 7256 3985 7259
rect 3568 7228 3985 7256
rect 3568 7216 3574 7228
rect 3973 7225 3985 7228
rect 4019 7225 4031 7259
rect 6730 7256 6736 7268
rect 3973 7219 4031 7225
rect 5644 7228 6736 7256
rect 1578 7148 1584 7200
rect 1636 7188 1642 7200
rect 2409 7191 2467 7197
rect 2409 7188 2421 7191
rect 1636 7160 2421 7188
rect 1636 7148 1642 7160
rect 2409 7157 2421 7160
rect 2455 7157 2467 7191
rect 3418 7188 3424 7200
rect 3379 7160 3424 7188
rect 2409 7151 2467 7157
rect 3418 7148 3424 7160
rect 3476 7188 3482 7200
rect 4065 7191 4123 7197
rect 4065 7188 4077 7191
rect 3476 7160 4077 7188
rect 3476 7148 3482 7160
rect 4065 7157 4077 7160
rect 4111 7157 4123 7191
rect 4065 7151 4123 7157
rect 5166 7148 5172 7200
rect 5224 7188 5230 7200
rect 5644 7197 5672 7228
rect 6730 7216 6736 7228
rect 6788 7216 6794 7268
rect 5629 7191 5687 7197
rect 5629 7188 5641 7191
rect 5224 7160 5641 7188
rect 5224 7148 5230 7160
rect 5629 7157 5641 7160
rect 5675 7157 5687 7191
rect 6270 7188 6276 7200
rect 6231 7160 6276 7188
rect 5629 7151 5687 7157
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 6454 7148 6460 7200
rect 6512 7188 6518 7200
rect 6549 7191 6607 7197
rect 6549 7188 6561 7191
rect 6512 7160 6561 7188
rect 6512 7148 6518 7160
rect 6549 7157 6561 7160
rect 6595 7188 6607 7191
rect 6840 7188 6868 7284
rect 7098 7265 7104 7268
rect 7092 7256 7104 7265
rect 7059 7228 7104 7256
rect 7092 7219 7104 7228
rect 7098 7216 7104 7219
rect 7156 7216 7162 7268
rect 8294 7216 8300 7268
rect 8352 7256 8358 7268
rect 9309 7259 9367 7265
rect 9309 7256 9321 7259
rect 8352 7228 9321 7256
rect 8352 7216 8358 7228
rect 9309 7225 9321 7228
rect 9355 7225 9367 7259
rect 9309 7219 9367 7225
rect 10134 7216 10140 7268
rect 10192 7256 10198 7268
rect 10229 7259 10287 7265
rect 10229 7256 10241 7259
rect 10192 7228 10241 7256
rect 10192 7216 10198 7228
rect 10229 7225 10241 7228
rect 10275 7256 10287 7259
rect 10778 7256 10784 7268
rect 10275 7228 10784 7256
rect 10275 7225 10287 7228
rect 10229 7219 10287 7225
rect 10778 7216 10784 7228
rect 10836 7216 10842 7268
rect 11054 7216 11060 7268
rect 11112 7256 11118 7268
rect 11241 7259 11299 7265
rect 11241 7256 11253 7259
rect 11112 7228 11253 7256
rect 11112 7216 11118 7228
rect 11241 7225 11253 7228
rect 11287 7225 11299 7259
rect 17034 7256 17040 7268
rect 11241 7219 11299 7225
rect 12176 7228 17040 7256
rect 6595 7160 6868 7188
rect 9861 7191 9919 7197
rect 6595 7157 6607 7160
rect 6549 7151 6607 7157
rect 9861 7157 9873 7191
rect 9907 7188 9919 7191
rect 9950 7188 9956 7200
rect 9907 7160 9956 7188
rect 9907 7157 9919 7160
rect 9861 7151 9919 7157
rect 9950 7148 9956 7160
rect 10008 7188 10014 7200
rect 12176 7188 12204 7228
rect 17034 7216 17040 7228
rect 17092 7216 17098 7268
rect 19978 7256 19984 7268
rect 19891 7228 19984 7256
rect 19978 7216 19984 7228
rect 20036 7256 20042 7268
rect 20622 7256 20628 7268
rect 20036 7228 20628 7256
rect 20036 7216 20042 7228
rect 20622 7216 20628 7228
rect 20680 7216 20686 7268
rect 10008 7160 12204 7188
rect 12253 7191 12311 7197
rect 10008 7148 10014 7160
rect 12253 7157 12265 7191
rect 12299 7188 12311 7191
rect 12342 7188 12348 7200
rect 12299 7160 12348 7188
rect 12299 7157 12311 7160
rect 12253 7151 12311 7157
rect 12342 7148 12348 7160
rect 12400 7148 12406 7200
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 14921 7191 14979 7197
rect 12492 7160 12537 7188
rect 12492 7148 12498 7160
rect 14921 7157 14933 7191
rect 14967 7188 14979 7191
rect 15289 7191 15347 7197
rect 15289 7188 15301 7191
rect 14967 7160 15301 7188
rect 14967 7157 14979 7160
rect 14921 7151 14979 7157
rect 15289 7157 15301 7160
rect 15335 7188 15347 7191
rect 16390 7188 16396 7200
rect 15335 7160 16396 7188
rect 15335 7157 15347 7160
rect 15289 7151 15347 7157
rect 16390 7148 16396 7160
rect 16448 7148 16454 7200
rect 18049 7191 18107 7197
rect 18049 7157 18061 7191
rect 18095 7188 18107 7191
rect 18322 7188 18328 7200
rect 18095 7160 18328 7188
rect 18095 7157 18107 7160
rect 18049 7151 18107 7157
rect 18322 7148 18328 7160
rect 18380 7148 18386 7200
rect 19518 7148 19524 7200
rect 19576 7188 19582 7200
rect 19613 7191 19671 7197
rect 19613 7188 19625 7191
rect 19576 7160 19625 7188
rect 19576 7148 19582 7160
rect 19613 7157 19625 7160
rect 19659 7157 19671 7191
rect 20070 7188 20076 7200
rect 19983 7160 20076 7188
rect 19613 7151 19671 7157
rect 20070 7148 20076 7160
rect 20128 7188 20134 7200
rect 20806 7188 20812 7200
rect 20128 7160 20812 7188
rect 20128 7148 20134 7160
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1397 6987 1455 6993
rect 1397 6953 1409 6987
rect 1443 6984 1455 6987
rect 1486 6984 1492 6996
rect 1443 6956 1492 6984
rect 1443 6953 1455 6956
rect 1397 6947 1455 6953
rect 1486 6944 1492 6956
rect 1544 6944 1550 6996
rect 1946 6984 1952 6996
rect 1907 6956 1952 6984
rect 1946 6944 1952 6956
rect 2004 6944 2010 6996
rect 2038 6944 2044 6996
rect 2096 6984 2102 6996
rect 3142 6984 3148 6996
rect 2096 6956 3148 6984
rect 2096 6944 2102 6956
rect 3142 6944 3148 6956
rect 3200 6984 3206 6996
rect 3602 6984 3608 6996
rect 3200 6956 3608 6984
rect 3200 6944 3206 6956
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 4430 6984 4436 6996
rect 4391 6956 4436 6984
rect 4430 6944 4436 6956
rect 4488 6944 4494 6996
rect 4798 6944 4804 6996
rect 4856 6984 4862 6996
rect 9306 6984 9312 6996
rect 4856 6956 9312 6984
rect 4856 6944 4862 6956
rect 9306 6944 9312 6956
rect 9364 6944 9370 6996
rect 9858 6984 9864 6996
rect 9819 6956 9864 6984
rect 9858 6944 9864 6956
rect 9916 6944 9922 6996
rect 13725 6987 13783 6993
rect 13725 6953 13737 6987
rect 13771 6984 13783 6987
rect 14090 6984 14096 6996
rect 13771 6956 14096 6984
rect 13771 6953 13783 6956
rect 13725 6947 13783 6953
rect 14090 6944 14096 6956
rect 14148 6944 14154 6996
rect 15381 6987 15439 6993
rect 15381 6953 15393 6987
rect 15427 6984 15439 6987
rect 16209 6987 16267 6993
rect 16209 6984 16221 6987
rect 15427 6956 16221 6984
rect 15427 6953 15439 6956
rect 15381 6947 15439 6953
rect 16209 6953 16221 6956
rect 16255 6984 16267 6987
rect 16482 6984 16488 6996
rect 16255 6956 16488 6984
rect 16255 6953 16267 6956
rect 16209 6947 16267 6953
rect 16482 6944 16488 6956
rect 16540 6944 16546 6996
rect 18414 6984 18420 6996
rect 18375 6956 18420 6984
rect 18414 6944 18420 6956
rect 18472 6944 18478 6996
rect 18506 6944 18512 6996
rect 18564 6984 18570 6996
rect 19058 6984 19064 6996
rect 18564 6956 19064 6984
rect 18564 6944 18570 6956
rect 19058 6944 19064 6956
rect 19116 6984 19122 6996
rect 19245 6987 19303 6993
rect 19245 6984 19257 6987
rect 19116 6956 19257 6984
rect 19116 6944 19122 6956
rect 19245 6953 19257 6956
rect 19291 6953 19303 6987
rect 19245 6947 19303 6953
rect 2777 6919 2835 6925
rect 2777 6885 2789 6919
rect 2823 6916 2835 6919
rect 2823 6888 4200 6916
rect 2823 6885 2835 6888
rect 2777 6879 2835 6885
rect 4172 6848 4200 6888
rect 4890 6876 4896 6928
rect 4948 6916 4954 6928
rect 9214 6916 9220 6928
rect 4948 6888 9220 6916
rect 4948 6876 4954 6888
rect 9214 6876 9220 6888
rect 9272 6876 9278 6928
rect 11425 6919 11483 6925
rect 11425 6885 11437 6919
rect 11471 6916 11483 6919
rect 11514 6916 11520 6928
rect 11471 6888 11520 6916
rect 11471 6885 11483 6888
rect 11425 6879 11483 6885
rect 11514 6876 11520 6888
rect 11572 6876 11578 6928
rect 5442 6848 5448 6860
rect 4172 6820 5448 6848
rect 5442 6808 5448 6820
rect 5500 6808 5506 6860
rect 5810 6808 5816 6860
rect 5868 6848 5874 6860
rect 6264 6851 6322 6857
rect 6264 6848 6276 6851
rect 5868 6820 6276 6848
rect 5868 6808 5874 6820
rect 6264 6817 6276 6820
rect 6310 6848 6322 6851
rect 7650 6848 7656 6860
rect 6310 6820 7656 6848
rect 6310 6817 6322 6820
rect 6264 6811 6322 6817
rect 7650 6808 7656 6820
rect 7708 6808 7714 6860
rect 8113 6851 8171 6857
rect 8113 6817 8125 6851
rect 8159 6848 8171 6851
rect 8294 6848 8300 6860
rect 8159 6820 8300 6848
rect 8159 6817 8171 6820
rect 8113 6811 8171 6817
rect 8294 6808 8300 6820
rect 8352 6808 8358 6860
rect 8478 6848 8484 6860
rect 8439 6820 8484 6848
rect 8478 6808 8484 6820
rect 8536 6808 8542 6860
rect 8662 6808 8668 6860
rect 8720 6848 8726 6860
rect 9582 6848 9588 6860
rect 8720 6820 9588 6848
rect 8720 6808 8726 6820
rect 9582 6808 9588 6820
rect 9640 6808 9646 6860
rect 12989 6851 13047 6857
rect 12989 6817 13001 6851
rect 13035 6848 13047 6851
rect 13446 6848 13452 6860
rect 13035 6820 13452 6848
rect 13035 6817 13047 6820
rect 12989 6811 13047 6817
rect 13446 6808 13452 6820
rect 13504 6808 13510 6860
rect 13906 6808 13912 6860
rect 13964 6848 13970 6860
rect 14001 6851 14059 6857
rect 14001 6848 14013 6851
rect 13964 6820 14013 6848
rect 13964 6808 13970 6820
rect 14001 6817 14013 6820
rect 14047 6817 14059 6851
rect 14001 6811 14059 6817
rect 14090 6808 14096 6860
rect 14148 6848 14154 6860
rect 14185 6851 14243 6857
rect 14185 6848 14197 6851
rect 14148 6820 14197 6848
rect 14148 6808 14154 6820
rect 14185 6817 14197 6820
rect 14231 6817 14243 6851
rect 14185 6811 14243 6817
rect 16482 6808 16488 6860
rect 16540 6848 16546 6860
rect 16649 6851 16707 6857
rect 16649 6848 16661 6851
rect 16540 6820 16661 6848
rect 16540 6808 16546 6820
rect 16649 6817 16661 6820
rect 16695 6817 16707 6851
rect 16649 6811 16707 6817
rect 18782 6808 18788 6860
rect 18840 6848 18846 6860
rect 19337 6851 19395 6857
rect 19337 6848 19349 6851
rect 18840 6820 19349 6848
rect 18840 6808 18846 6820
rect 19337 6817 19349 6820
rect 19383 6817 19395 6851
rect 22278 6848 22284 6860
rect 22239 6820 22284 6848
rect 19337 6811 19395 6817
rect 22278 6808 22284 6820
rect 22336 6808 22342 6860
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6749 2927 6783
rect 3050 6780 3056 6792
rect 3011 6752 3056 6780
rect 2869 6743 2927 6749
rect 2884 6712 2912 6743
rect 3050 6740 3056 6752
rect 3108 6740 3114 6792
rect 4522 6780 4528 6792
rect 4483 6752 4528 6780
rect 4522 6740 4528 6752
rect 4580 6740 4586 6792
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6780 4767 6783
rect 5994 6780 6000 6792
rect 4755 6752 5304 6780
rect 5955 6752 6000 6780
rect 4755 6749 4767 6752
rect 4709 6743 4767 6749
rect 2884 6684 4108 6712
rect 4080 6656 4108 6684
rect 4154 6672 4160 6724
rect 4212 6712 4218 6724
rect 5166 6712 5172 6724
rect 4212 6684 5172 6712
rect 4212 6672 4218 6684
rect 5166 6672 5172 6684
rect 5224 6672 5230 6724
rect 5276 6656 5304 6752
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 11054 6740 11060 6792
rect 11112 6780 11118 6792
rect 11517 6783 11575 6789
rect 11517 6780 11529 6783
rect 11112 6752 11529 6780
rect 11112 6740 11118 6752
rect 11517 6749 11529 6752
rect 11563 6749 11575 6783
rect 11517 6743 11575 6749
rect 11606 6740 11612 6792
rect 11664 6780 11670 6792
rect 12529 6783 12587 6789
rect 11664 6752 11709 6780
rect 11664 6740 11670 6752
rect 12529 6749 12541 6783
rect 12575 6780 12587 6783
rect 13078 6780 13084 6792
rect 12575 6752 13084 6780
rect 12575 6749 12587 6752
rect 12529 6743 12587 6749
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 13265 6783 13323 6789
rect 13265 6749 13277 6783
rect 13311 6780 13323 6783
rect 13630 6780 13636 6792
rect 13311 6752 13636 6780
rect 13311 6749 13323 6752
rect 13265 6743 13323 6749
rect 13630 6740 13636 6752
rect 13688 6740 13694 6792
rect 16393 6783 16451 6789
rect 16393 6749 16405 6783
rect 16439 6749 16451 6783
rect 16393 6743 16451 6749
rect 9674 6672 9680 6724
rect 9732 6712 9738 6724
rect 10781 6715 10839 6721
rect 10781 6712 10793 6715
rect 9732 6684 10793 6712
rect 9732 6672 9738 6684
rect 10781 6681 10793 6684
rect 10827 6712 10839 6715
rect 10870 6712 10876 6724
rect 10827 6684 10876 6712
rect 10827 6681 10839 6684
rect 10781 6675 10839 6681
rect 10870 6672 10876 6684
rect 10928 6672 10934 6724
rect 12161 6715 12219 6721
rect 12161 6681 12173 6715
rect 12207 6712 12219 6715
rect 12894 6712 12900 6724
rect 12207 6684 12900 6712
rect 12207 6681 12219 6684
rect 12161 6675 12219 6681
rect 12894 6672 12900 6684
rect 12952 6672 12958 6724
rect 13814 6672 13820 6724
rect 13872 6712 13878 6724
rect 15013 6715 15071 6721
rect 15013 6712 15025 6715
rect 13872 6684 15025 6712
rect 13872 6672 13878 6684
rect 15013 6681 15025 6684
rect 15059 6681 15071 6715
rect 15013 6675 15071 6681
rect 2222 6644 2228 6656
rect 2183 6616 2228 6644
rect 2222 6604 2228 6616
rect 2280 6604 2286 6656
rect 2409 6647 2467 6653
rect 2409 6613 2421 6647
rect 2455 6644 2467 6647
rect 2682 6644 2688 6656
rect 2455 6616 2688 6644
rect 2455 6613 2467 6616
rect 2409 6607 2467 6613
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 3510 6604 3516 6656
rect 3568 6644 3574 6656
rect 3605 6647 3663 6653
rect 3605 6644 3617 6647
rect 3568 6616 3617 6644
rect 3568 6604 3574 6616
rect 3605 6613 3617 6616
rect 3651 6613 3663 6647
rect 4062 6644 4068 6656
rect 4023 6616 4068 6644
rect 3605 6607 3663 6613
rect 4062 6604 4068 6616
rect 4120 6604 4126 6656
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 5537 6647 5595 6653
rect 5537 6644 5549 6647
rect 5316 6616 5549 6644
rect 5316 6604 5322 6616
rect 5537 6613 5549 6616
rect 5583 6613 5595 6647
rect 5537 6607 5595 6613
rect 7098 6604 7104 6656
rect 7156 6644 7162 6656
rect 7377 6647 7435 6653
rect 7377 6644 7389 6647
rect 7156 6616 7389 6644
rect 7156 6604 7162 6616
rect 7377 6613 7389 6616
rect 7423 6613 7435 6647
rect 8938 6644 8944 6656
rect 8899 6616 8944 6644
rect 7377 6607 7435 6613
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 9306 6644 9312 6656
rect 9267 6616 9312 6644
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 10226 6644 10232 6656
rect 10187 6616 10232 6644
rect 10226 6604 10232 6616
rect 10284 6604 10290 6656
rect 11057 6647 11115 6653
rect 11057 6613 11069 6647
rect 11103 6644 11115 6647
rect 12250 6644 12256 6656
rect 11103 6616 12256 6644
rect 11103 6613 11115 6616
rect 11057 6607 11115 6613
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 12618 6644 12624 6656
rect 12579 6616 12624 6644
rect 12618 6604 12624 6616
rect 12676 6604 12682 6656
rect 14366 6644 14372 6656
rect 14327 6616 14372 6644
rect 14366 6604 14372 6616
rect 14424 6604 14430 6656
rect 14642 6644 14648 6656
rect 14603 6616 14648 6644
rect 14642 6604 14648 6616
rect 14700 6604 14706 6656
rect 16408 6644 16436 6743
rect 19426 6740 19432 6792
rect 19484 6780 19490 6792
rect 19889 6783 19947 6789
rect 19889 6780 19901 6783
rect 19484 6752 19901 6780
rect 19484 6740 19490 6752
rect 19889 6749 19901 6752
rect 19935 6749 19947 6783
rect 19889 6743 19947 6749
rect 18877 6715 18935 6721
rect 18877 6681 18889 6715
rect 18923 6712 18935 6715
rect 21177 6715 21235 6721
rect 21177 6712 21189 6715
rect 18923 6684 21189 6712
rect 18923 6681 18935 6684
rect 18877 6675 18935 6681
rect 21177 6681 21189 6684
rect 21223 6712 21235 6715
rect 21634 6712 21640 6724
rect 21223 6684 21640 6712
rect 21223 6681 21235 6684
rect 21177 6675 21235 6681
rect 21634 6672 21640 6684
rect 21692 6672 21698 6724
rect 16574 6644 16580 6656
rect 16408 6616 16580 6644
rect 16574 6604 16580 6616
rect 16632 6604 16638 6656
rect 17770 6644 17776 6656
rect 17731 6616 17776 6644
rect 17770 6604 17776 6616
rect 17828 6604 17834 6656
rect 18690 6644 18696 6656
rect 18651 6616 18696 6644
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 20254 6644 20260 6656
rect 20215 6616 20260 6644
rect 20254 6604 20260 6616
rect 20312 6604 20318 6656
rect 21542 6644 21548 6656
rect 21503 6616 21548 6644
rect 21542 6604 21548 6616
rect 21600 6604 21606 6656
rect 22462 6644 22468 6656
rect 22423 6616 22468 6644
rect 22462 6604 22468 6616
rect 22520 6604 22526 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1673 6443 1731 6449
rect 1673 6409 1685 6443
rect 1719 6440 1731 6443
rect 2038 6440 2044 6452
rect 1719 6412 2044 6440
rect 1719 6409 1731 6412
rect 1673 6403 1731 6409
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 2130 6400 2136 6452
rect 2188 6440 2194 6452
rect 4709 6443 4767 6449
rect 2188 6412 2233 6440
rect 2188 6400 2194 6412
rect 4709 6409 4721 6443
rect 4755 6440 4767 6443
rect 5442 6440 5448 6452
rect 4755 6412 5448 6440
rect 4755 6409 4767 6412
rect 4709 6403 4767 6409
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 5994 6400 6000 6452
rect 6052 6440 6058 6452
rect 6089 6443 6147 6449
rect 6089 6440 6101 6443
rect 6052 6412 6101 6440
rect 6052 6400 6058 6412
rect 6089 6409 6101 6412
rect 6135 6440 6147 6443
rect 6454 6440 6460 6452
rect 6135 6412 6460 6440
rect 6135 6409 6147 6412
rect 6089 6403 6147 6409
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 6822 6440 6828 6452
rect 6783 6412 6828 6440
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 7558 6400 7564 6452
rect 7616 6440 7622 6452
rect 7837 6443 7895 6449
rect 7837 6440 7849 6443
rect 7616 6412 7849 6440
rect 7616 6400 7622 6412
rect 7837 6409 7849 6412
rect 7883 6409 7895 6443
rect 8294 6440 8300 6452
rect 8255 6412 8300 6440
rect 7837 6403 7895 6409
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 8570 6440 8576 6452
rect 8531 6412 8576 6440
rect 8570 6400 8576 6412
rect 8628 6400 8634 6452
rect 9398 6440 9404 6452
rect 9359 6412 9404 6440
rect 9398 6400 9404 6412
rect 9456 6400 9462 6452
rect 11882 6400 11888 6452
rect 11940 6440 11946 6452
rect 15657 6443 15715 6449
rect 15657 6440 15669 6443
rect 11940 6412 15669 6440
rect 11940 6400 11946 6412
rect 15657 6409 15669 6412
rect 15703 6440 15715 6443
rect 16666 6440 16672 6452
rect 15703 6412 16672 6440
rect 15703 6409 15715 6412
rect 15657 6403 15715 6409
rect 16666 6400 16672 6412
rect 16724 6400 16730 6452
rect 17678 6400 17684 6452
rect 17736 6440 17742 6452
rect 17773 6443 17831 6449
rect 17773 6440 17785 6443
rect 17736 6412 17785 6440
rect 17736 6400 17742 6412
rect 17773 6409 17785 6412
rect 17819 6409 17831 6443
rect 18046 6440 18052 6452
rect 18007 6412 18052 6440
rect 17773 6403 17831 6409
rect 18046 6400 18052 6412
rect 18104 6400 18110 6452
rect 19058 6440 19064 6452
rect 19019 6412 19064 6440
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 20714 6400 20720 6452
rect 20772 6440 20778 6452
rect 21177 6443 21235 6449
rect 21177 6440 21189 6443
rect 20772 6412 21189 6440
rect 20772 6400 20778 6412
rect 21177 6409 21189 6412
rect 21223 6409 21235 6443
rect 22278 6440 22284 6452
rect 22239 6412 22284 6440
rect 21177 6403 21235 6409
rect 22278 6400 22284 6412
rect 22336 6400 22342 6452
rect 2148 6304 2176 6400
rect 2225 6307 2283 6313
rect 2225 6304 2237 6307
rect 2148 6276 2237 6304
rect 2225 6273 2237 6276
rect 2271 6273 2283 6307
rect 5258 6304 5264 6316
rect 5219 6276 5264 6304
rect 2225 6267 2283 6273
rect 5258 6264 5264 6276
rect 5316 6304 5322 6316
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 5316 6276 6377 6304
rect 5316 6264 5322 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 7282 6304 7288 6316
rect 7243 6276 7288 6304
rect 6365 6267 6423 6273
rect 7282 6264 7288 6276
rect 7340 6264 7346 6316
rect 7469 6307 7527 6313
rect 7469 6273 7481 6307
rect 7515 6304 7527 6307
rect 7576 6304 7604 6400
rect 7515 6276 7604 6304
rect 9416 6304 9444 6400
rect 13630 6372 13636 6384
rect 11808 6344 13636 6372
rect 9493 6307 9551 6313
rect 9493 6304 9505 6307
rect 9416 6276 9505 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 9493 6273 9505 6276
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 3050 6236 3056 6248
rect 2884 6208 3056 6236
rect 2884 6180 2912 6208
rect 3050 6196 3056 6208
rect 3108 6196 3114 6248
rect 7190 6236 7196 6248
rect 7151 6208 7196 6236
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 10686 6196 10692 6248
rect 10744 6236 10750 6248
rect 11808 6245 11836 6344
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 19426 6332 19432 6384
rect 19484 6372 19490 6384
rect 19484 6344 20208 6372
rect 19484 6332 19490 6344
rect 13081 6307 13139 6313
rect 13081 6273 13093 6307
rect 13127 6273 13139 6307
rect 13081 6267 13139 6273
rect 11793 6239 11851 6245
rect 11793 6236 11805 6239
rect 10744 6208 11805 6236
rect 10744 6196 10750 6208
rect 11793 6205 11805 6208
rect 11839 6205 11851 6239
rect 11793 6199 11851 6205
rect 12253 6239 12311 6245
rect 12253 6205 12265 6239
rect 12299 6236 12311 6239
rect 12299 6208 12471 6236
rect 12299 6205 12311 6208
rect 12253 6199 12311 6205
rect 2492 6171 2550 6177
rect 2492 6137 2504 6171
rect 2538 6168 2550 6171
rect 2866 6168 2872 6180
rect 2538 6140 2872 6168
rect 2538 6137 2550 6140
rect 2492 6131 2550 6137
rect 2866 6128 2872 6140
rect 2924 6128 2930 6180
rect 4249 6171 4307 6177
rect 4249 6137 4261 6171
rect 4295 6168 4307 6171
rect 5077 6171 5135 6177
rect 5077 6168 5089 6171
rect 4295 6140 5089 6168
rect 4295 6137 4307 6140
rect 4249 6131 4307 6137
rect 5077 6137 5089 6140
rect 5123 6168 5135 6171
rect 5442 6168 5448 6180
rect 5123 6140 5448 6168
rect 5123 6137 5135 6140
rect 5077 6131 5135 6137
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 9033 6171 9091 6177
rect 9033 6137 9045 6171
rect 9079 6168 9091 6171
rect 9760 6171 9818 6177
rect 9760 6168 9772 6171
rect 9079 6140 9772 6168
rect 9079 6137 9091 6140
rect 9033 6131 9091 6137
rect 9760 6137 9772 6140
rect 9806 6168 9818 6171
rect 11054 6168 11060 6180
rect 9806 6140 11060 6168
rect 9806 6137 9818 6140
rect 9760 6131 9818 6137
rect 11054 6128 11060 6140
rect 11112 6168 11118 6180
rect 12268 6168 12296 6199
rect 11112 6140 12296 6168
rect 12443 6168 12471 6208
rect 12618 6196 12624 6248
rect 12676 6236 12682 6248
rect 12805 6239 12863 6245
rect 12805 6236 12817 6239
rect 12676 6208 12817 6236
rect 12676 6196 12682 6208
rect 12805 6205 12817 6208
rect 12851 6205 12863 6239
rect 12805 6199 12863 6205
rect 13096 6168 13124 6267
rect 16666 6264 16672 6316
rect 16724 6304 16730 6316
rect 18506 6304 18512 6316
rect 16724 6276 18512 6304
rect 16724 6264 16730 6276
rect 18506 6264 18512 6276
rect 18564 6304 18570 6316
rect 18693 6307 18751 6313
rect 18693 6304 18705 6307
rect 18564 6276 18705 6304
rect 18564 6264 18570 6276
rect 18693 6273 18705 6276
rect 18739 6273 18751 6307
rect 18693 6267 18751 6273
rect 19242 6264 19248 6316
rect 19300 6304 19306 6316
rect 20180 6313 20208 6344
rect 19521 6307 19579 6313
rect 19521 6304 19533 6307
rect 19300 6276 19533 6304
rect 19300 6264 19306 6276
rect 19521 6273 19533 6276
rect 19567 6304 19579 6307
rect 20073 6307 20131 6313
rect 20073 6304 20085 6307
rect 19567 6276 20085 6304
rect 19567 6273 19579 6276
rect 19521 6267 19579 6273
rect 20073 6273 20085 6276
rect 20119 6273 20131 6307
rect 20073 6267 20131 6273
rect 20165 6307 20223 6313
rect 20165 6273 20177 6307
rect 20211 6304 20223 6307
rect 20530 6304 20536 6316
rect 20211 6276 20536 6304
rect 20211 6273 20223 6276
rect 20165 6267 20223 6273
rect 20530 6264 20536 6276
rect 20588 6304 20594 6316
rect 20625 6307 20683 6313
rect 20625 6304 20637 6307
rect 20588 6276 20637 6304
rect 20588 6264 20594 6276
rect 20625 6273 20637 6276
rect 20671 6273 20683 6307
rect 21634 6304 21640 6316
rect 21595 6276 21640 6304
rect 20625 6267 20683 6273
rect 21634 6264 21640 6276
rect 21692 6264 21698 6316
rect 21729 6307 21787 6313
rect 21729 6273 21741 6307
rect 21775 6273 21787 6307
rect 21729 6267 21787 6273
rect 14185 6239 14243 6245
rect 14185 6205 14197 6239
rect 14231 6236 14243 6239
rect 14277 6239 14335 6245
rect 14277 6236 14289 6239
rect 14231 6208 14289 6236
rect 14231 6205 14243 6208
rect 14185 6199 14243 6205
rect 14277 6205 14289 6208
rect 14323 6205 14335 6239
rect 14277 6199 14335 6205
rect 14544 6239 14602 6245
rect 14544 6205 14556 6239
rect 14590 6236 14602 6239
rect 14826 6236 14832 6248
rect 14590 6208 14832 6236
rect 14590 6205 14602 6208
rect 14544 6199 14602 6205
rect 12443 6140 13124 6168
rect 14292 6168 14320 6199
rect 14826 6196 14832 6208
rect 14884 6196 14890 6248
rect 16482 6196 16488 6248
rect 16540 6236 16546 6248
rect 16758 6236 16764 6248
rect 16540 6208 16764 6236
rect 16540 6196 16546 6208
rect 16758 6196 16764 6208
rect 16816 6196 16822 6248
rect 17678 6196 17684 6248
rect 17736 6236 17742 6248
rect 18417 6239 18475 6245
rect 18417 6236 18429 6239
rect 17736 6208 18429 6236
rect 17736 6196 17742 6208
rect 18417 6205 18429 6208
rect 18463 6205 18475 6239
rect 19978 6236 19984 6248
rect 19939 6208 19984 6236
rect 18417 6199 18475 6205
rect 19978 6196 19984 6208
rect 20036 6196 20042 6248
rect 21744 6236 21772 6267
rect 21652 6208 21772 6236
rect 14292 6140 16528 6168
rect 11112 6128 11118 6140
rect 3050 6060 3056 6112
rect 3108 6100 3114 6112
rect 3605 6103 3663 6109
rect 3605 6100 3617 6103
rect 3108 6072 3617 6100
rect 3108 6060 3114 6072
rect 3605 6069 3617 6072
rect 3651 6069 3663 6103
rect 4522 6100 4528 6112
rect 4483 6072 4528 6100
rect 3605 6063 3663 6069
rect 4522 6060 4528 6072
rect 4580 6100 4586 6112
rect 5169 6103 5227 6109
rect 5169 6100 5181 6103
rect 4580 6072 5181 6100
rect 4580 6060 4586 6072
rect 5169 6069 5181 6072
rect 5215 6069 5227 6103
rect 5169 6063 5227 6069
rect 9858 6060 9864 6112
rect 9916 6100 9922 6112
rect 10873 6103 10931 6109
rect 10873 6100 10885 6103
rect 9916 6072 10885 6100
rect 9916 6060 9922 6072
rect 10873 6069 10885 6072
rect 10919 6069 10931 6103
rect 11514 6100 11520 6112
rect 11475 6072 11520 6100
rect 10873 6063 10931 6069
rect 11514 6060 11520 6072
rect 11572 6060 11578 6112
rect 12434 6060 12440 6112
rect 12492 6100 12498 6112
rect 12894 6100 12900 6112
rect 12492 6072 12537 6100
rect 12855 6072 12900 6100
rect 12492 6060 12498 6072
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 13446 6100 13452 6112
rect 13407 6072 13452 6100
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 16500 6109 16528 6140
rect 17034 6128 17040 6180
rect 17092 6168 17098 6180
rect 17497 6171 17555 6177
rect 17497 6168 17509 6171
rect 17092 6140 17509 6168
rect 17092 6128 17098 6140
rect 17497 6137 17509 6140
rect 17543 6168 17555 6171
rect 18509 6171 18567 6177
rect 18509 6168 18521 6171
rect 17543 6140 18521 6168
rect 17543 6137 17555 6140
rect 17497 6131 17555 6137
rect 18509 6137 18521 6140
rect 18555 6137 18567 6171
rect 21542 6168 21548 6180
rect 18509 6131 18567 6137
rect 19628 6140 21548 6168
rect 16485 6103 16543 6109
rect 16485 6069 16497 6103
rect 16531 6100 16543 6103
rect 16574 6100 16580 6112
rect 16531 6072 16580 6100
rect 16531 6069 16543 6072
rect 16485 6063 16543 6069
rect 16574 6060 16580 6072
rect 16632 6060 16638 6112
rect 16942 6100 16948 6112
rect 16903 6072 16948 6100
rect 16942 6060 16948 6072
rect 17000 6060 17006 6112
rect 19628 6109 19656 6140
rect 21542 6128 21548 6140
rect 21600 6128 21606 6180
rect 19613 6103 19671 6109
rect 19613 6069 19625 6103
rect 19659 6069 19671 6103
rect 20990 6100 20996 6112
rect 20951 6072 20996 6100
rect 19613 6063 19671 6069
rect 20990 6060 20996 6072
rect 21048 6100 21054 6112
rect 21652 6100 21680 6208
rect 21048 6072 21680 6100
rect 21048 6060 21054 6072
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 3602 5856 3608 5908
rect 3660 5896 3666 5908
rect 5258 5896 5264 5908
rect 3660 5868 5264 5896
rect 3660 5856 3666 5868
rect 5258 5856 5264 5868
rect 5316 5896 5322 5908
rect 5445 5899 5503 5905
rect 5445 5896 5457 5899
rect 5316 5868 5457 5896
rect 5316 5856 5322 5868
rect 5445 5865 5457 5868
rect 5491 5865 5503 5899
rect 5445 5859 5503 5865
rect 6549 5899 6607 5905
rect 6549 5865 6561 5899
rect 6595 5896 6607 5899
rect 7282 5896 7288 5908
rect 6595 5868 7288 5896
rect 6595 5865 6607 5868
rect 6549 5859 6607 5865
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 7650 5896 7656 5908
rect 7611 5868 7656 5896
rect 7650 5856 7656 5868
rect 7708 5856 7714 5908
rect 8294 5896 8300 5908
rect 8255 5868 8300 5896
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 11054 5896 11060 5908
rect 11015 5868 11060 5896
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 11606 5896 11612 5908
rect 11567 5868 11612 5896
rect 11606 5856 11612 5868
rect 11664 5856 11670 5908
rect 12069 5899 12127 5905
rect 12069 5865 12081 5899
rect 12115 5896 12127 5899
rect 12618 5896 12624 5908
rect 12115 5868 12624 5896
rect 12115 5865 12127 5868
rect 12069 5859 12127 5865
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 14369 5899 14427 5905
rect 14369 5865 14381 5899
rect 14415 5896 14427 5899
rect 14826 5896 14832 5908
rect 14415 5868 14832 5896
rect 14415 5865 14427 5868
rect 14369 5859 14427 5865
rect 14826 5856 14832 5868
rect 14884 5856 14890 5908
rect 15654 5856 15660 5908
rect 15712 5896 15718 5908
rect 15749 5899 15807 5905
rect 15749 5896 15761 5899
rect 15712 5868 15761 5896
rect 15712 5856 15718 5868
rect 15749 5865 15761 5868
rect 15795 5865 15807 5899
rect 16666 5896 16672 5908
rect 16627 5868 16672 5896
rect 15749 5859 15807 5865
rect 16666 5856 16672 5868
rect 16724 5856 16730 5908
rect 19978 5896 19984 5908
rect 19939 5868 19984 5896
rect 19978 5856 19984 5868
rect 20036 5856 20042 5908
rect 20530 5896 20536 5908
rect 20491 5868 20536 5896
rect 20530 5856 20536 5868
rect 20588 5856 20594 5908
rect 20806 5856 20812 5908
rect 20864 5896 20870 5908
rect 20901 5899 20959 5905
rect 20901 5896 20913 5899
rect 20864 5868 20913 5896
rect 20864 5856 20870 5868
rect 20901 5865 20913 5868
rect 20947 5865 20959 5899
rect 21358 5896 21364 5908
rect 21319 5868 21364 5896
rect 20901 5859 20959 5865
rect 21358 5856 21364 5868
rect 21416 5856 21422 5908
rect 1664 5831 1722 5837
rect 1664 5797 1676 5831
rect 1710 5828 1722 5831
rect 2038 5828 2044 5840
rect 1710 5800 2044 5828
rect 1710 5797 1722 5800
rect 1664 5791 1722 5797
rect 2038 5788 2044 5800
rect 2096 5788 2102 5840
rect 6822 5788 6828 5840
rect 6880 5828 6886 5840
rect 6917 5831 6975 5837
rect 6917 5828 6929 5831
rect 6880 5800 6929 5828
rect 6880 5788 6886 5800
rect 6917 5797 6929 5800
rect 6963 5828 6975 5831
rect 9306 5828 9312 5840
rect 6963 5800 9312 5828
rect 6963 5797 6975 5800
rect 6917 5791 6975 5797
rect 9306 5788 9312 5800
rect 9364 5788 9370 5840
rect 17120 5831 17178 5837
rect 17120 5828 17132 5831
rect 9692 5800 12204 5828
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5760 1455 5763
rect 2130 5760 2136 5772
rect 1443 5732 2136 5760
rect 1443 5729 1455 5732
rect 1397 5723 1455 5729
rect 2130 5720 2136 5732
rect 2188 5760 2194 5772
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 2188 5732 4077 5760
rect 2188 5720 2194 5732
rect 4065 5729 4077 5732
rect 4111 5760 4123 5763
rect 4154 5760 4160 5772
rect 4111 5732 4160 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 4154 5720 4160 5732
rect 4212 5720 4218 5772
rect 4332 5763 4390 5769
rect 4332 5729 4344 5763
rect 4378 5760 4390 5763
rect 4614 5760 4620 5772
rect 4378 5732 4620 5760
rect 4378 5729 4390 5732
rect 4332 5723 4390 5729
rect 4614 5720 4620 5732
rect 4672 5720 4678 5772
rect 7009 5763 7067 5769
rect 7009 5729 7021 5763
rect 7055 5760 7067 5763
rect 7558 5760 7564 5772
rect 7055 5732 7564 5760
rect 7055 5729 7067 5732
rect 7009 5723 7067 5729
rect 7558 5720 7564 5732
rect 7616 5720 7622 5772
rect 8570 5760 8576 5772
rect 8531 5732 8576 5760
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 9214 5720 9220 5772
rect 9272 5760 9278 5772
rect 9398 5760 9404 5772
rect 9272 5732 9404 5760
rect 9272 5720 9278 5732
rect 9398 5720 9404 5732
rect 9456 5760 9462 5772
rect 9692 5769 9720 5800
rect 9950 5769 9956 5772
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 9456 5732 9689 5760
rect 9456 5720 9462 5732
rect 9677 5729 9689 5732
rect 9723 5729 9735 5763
rect 9944 5760 9956 5769
rect 9911 5732 9956 5760
rect 9677 5723 9735 5729
rect 9944 5723 9956 5732
rect 9950 5720 9956 5723
rect 10008 5720 10014 5772
rect 12066 5720 12072 5772
rect 12124 5760 12130 5772
rect 12176 5769 12204 5800
rect 15948 5800 17132 5828
rect 12434 5769 12440 5772
rect 12161 5763 12219 5769
rect 12161 5760 12173 5763
rect 12124 5732 12173 5760
rect 12124 5720 12130 5732
rect 12161 5729 12173 5732
rect 12207 5729 12219 5763
rect 12161 5723 12219 5729
rect 12428 5723 12440 5769
rect 12492 5760 12498 5772
rect 12492 5732 12528 5760
rect 12434 5720 12440 5723
rect 12492 5720 12498 5732
rect 15562 5720 15568 5772
rect 15620 5760 15626 5772
rect 15657 5763 15715 5769
rect 15657 5760 15669 5763
rect 15620 5732 15669 5760
rect 15620 5720 15626 5732
rect 15657 5729 15669 5732
rect 15703 5729 15715 5763
rect 15657 5723 15715 5729
rect 15948 5704 15976 5800
rect 17120 5797 17132 5800
rect 17166 5828 17178 5831
rect 17770 5828 17776 5840
rect 17166 5800 17776 5828
rect 17166 5797 17178 5800
rect 17120 5791 17178 5797
rect 17770 5788 17776 5800
rect 17828 5788 17834 5840
rect 16574 5720 16580 5772
rect 16632 5760 16638 5772
rect 16853 5763 16911 5769
rect 16853 5760 16865 5763
rect 16632 5732 16865 5760
rect 16632 5720 16638 5732
rect 16853 5729 16865 5732
rect 16899 5760 16911 5763
rect 17402 5760 17408 5772
rect 16899 5732 17408 5760
rect 16899 5729 16911 5732
rect 16853 5723 16911 5729
rect 17402 5720 17408 5732
rect 17460 5720 17466 5772
rect 19334 5760 19340 5772
rect 19295 5732 19340 5760
rect 19334 5720 19340 5732
rect 19392 5720 19398 5772
rect 21266 5760 21272 5772
rect 21227 5732 21272 5760
rect 21266 5720 21272 5732
rect 21324 5720 21330 5772
rect 22462 5720 22468 5772
rect 22520 5760 22526 5772
rect 23290 5760 23296 5772
rect 22520 5732 23296 5760
rect 22520 5720 22526 5732
rect 23290 5720 23296 5732
rect 23348 5720 23354 5772
rect 7098 5652 7104 5704
rect 7156 5692 7162 5704
rect 15930 5692 15936 5704
rect 7156 5664 7201 5692
rect 15843 5664 15936 5692
rect 7156 5652 7162 5664
rect 15930 5652 15936 5664
rect 15988 5652 15994 5704
rect 20990 5652 20996 5704
rect 21048 5692 21054 5704
rect 21453 5695 21511 5701
rect 21453 5692 21465 5695
rect 21048 5664 21465 5692
rect 21048 5652 21054 5664
rect 21453 5661 21465 5664
rect 21499 5661 21511 5695
rect 21453 5655 21511 5661
rect 2406 5584 2412 5636
rect 2464 5624 2470 5636
rect 2777 5627 2835 5633
rect 2777 5624 2789 5627
rect 2464 5596 2789 5624
rect 2464 5584 2470 5596
rect 2777 5593 2789 5596
rect 2823 5624 2835 5627
rect 2866 5624 2872 5636
rect 2823 5596 2872 5624
rect 2823 5593 2835 5596
rect 2777 5587 2835 5593
rect 2866 5584 2872 5596
rect 2924 5624 2930 5636
rect 9398 5624 9404 5636
rect 2924 5596 3924 5624
rect 2924 5584 2930 5596
rect 3896 5568 3924 5596
rect 5000 5596 6132 5624
rect 9359 5596 9404 5624
rect 3694 5556 3700 5568
rect 3655 5528 3700 5556
rect 3694 5516 3700 5528
rect 3752 5516 3758 5568
rect 3878 5556 3884 5568
rect 3791 5528 3884 5556
rect 3878 5516 3884 5528
rect 3936 5556 3942 5568
rect 5000 5556 5028 5596
rect 6104 5565 6132 5596
rect 9398 5584 9404 5596
rect 9456 5584 9462 5636
rect 13906 5584 13912 5636
rect 13964 5624 13970 5636
rect 14090 5624 14096 5636
rect 13964 5596 14096 5624
rect 13964 5584 13970 5596
rect 14090 5584 14096 5596
rect 14148 5624 14154 5636
rect 14645 5627 14703 5633
rect 14645 5624 14657 5627
rect 14148 5596 14657 5624
rect 14148 5584 14154 5596
rect 14645 5593 14657 5596
rect 14691 5593 14703 5627
rect 14645 5587 14703 5593
rect 15289 5627 15347 5633
rect 15289 5593 15301 5627
rect 15335 5624 15347 5627
rect 16574 5624 16580 5636
rect 15335 5596 16580 5624
rect 15335 5593 15347 5596
rect 15289 5587 15347 5593
rect 16574 5584 16580 5596
rect 16632 5584 16638 5636
rect 19521 5627 19579 5633
rect 19521 5593 19533 5627
rect 19567 5624 19579 5627
rect 20806 5624 20812 5636
rect 19567 5596 20812 5624
rect 19567 5593 19579 5596
rect 19521 5587 19579 5593
rect 20806 5584 20812 5596
rect 20864 5584 20870 5636
rect 3936 5528 5028 5556
rect 6089 5559 6147 5565
rect 3936 5516 3942 5528
rect 6089 5525 6101 5559
rect 6135 5556 6147 5559
rect 6365 5559 6423 5565
rect 6365 5556 6377 5559
rect 6135 5528 6377 5556
rect 6135 5525 6147 5528
rect 6089 5519 6147 5525
rect 6365 5525 6377 5528
rect 6411 5525 6423 5559
rect 6365 5519 6423 5525
rect 7650 5516 7656 5568
rect 7708 5556 7714 5568
rect 7929 5559 7987 5565
rect 7929 5556 7941 5559
rect 7708 5528 7941 5556
rect 7708 5516 7714 5528
rect 7929 5525 7941 5528
rect 7975 5525 7987 5559
rect 7929 5519 7987 5525
rect 13541 5559 13599 5565
rect 13541 5525 13553 5559
rect 13587 5556 13599 5559
rect 13630 5556 13636 5568
rect 13587 5528 13636 5556
rect 13587 5525 13599 5528
rect 13541 5519 13599 5525
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 14734 5516 14740 5568
rect 14792 5556 14798 5568
rect 15013 5559 15071 5565
rect 15013 5556 15025 5559
rect 14792 5528 15025 5556
rect 14792 5516 14798 5528
rect 15013 5525 15025 5528
rect 15059 5525 15071 5559
rect 16390 5556 16396 5568
rect 16351 5528 16396 5556
rect 15013 5519 15071 5525
rect 16390 5516 16396 5528
rect 16448 5516 16454 5568
rect 18138 5516 18144 5568
rect 18196 5556 18202 5568
rect 18233 5559 18291 5565
rect 18233 5556 18245 5559
rect 18196 5528 18245 5556
rect 18196 5516 18202 5528
rect 18233 5525 18245 5528
rect 18279 5525 18291 5559
rect 18233 5519 18291 5525
rect 18782 5516 18788 5568
rect 18840 5556 18846 5568
rect 18877 5559 18935 5565
rect 18877 5556 18889 5559
rect 18840 5528 18889 5556
rect 18840 5516 18846 5528
rect 18877 5525 18889 5528
rect 18923 5525 18935 5559
rect 23474 5556 23480 5568
rect 23435 5528 23480 5556
rect 18877 5519 18935 5525
rect 23474 5516 23480 5528
rect 23532 5516 23538 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 3329 5355 3387 5361
rect 3329 5321 3341 5355
rect 3375 5352 3387 5355
rect 3605 5355 3663 5361
rect 3605 5352 3617 5355
rect 3375 5324 3617 5352
rect 3375 5321 3387 5324
rect 3329 5315 3387 5321
rect 3605 5321 3617 5324
rect 3651 5321 3663 5355
rect 3605 5315 3663 5321
rect 4154 5312 4160 5364
rect 4212 5352 4218 5364
rect 4617 5355 4675 5361
rect 4617 5352 4629 5355
rect 4212 5324 4629 5352
rect 4212 5312 4218 5324
rect 4617 5321 4629 5324
rect 4663 5321 4675 5355
rect 4617 5315 4675 5321
rect 8849 5355 8907 5361
rect 8849 5321 8861 5355
rect 8895 5352 8907 5355
rect 9950 5352 9956 5364
rect 8895 5324 9956 5352
rect 8895 5321 8907 5324
rect 8849 5315 8907 5321
rect 9950 5312 9956 5324
rect 10008 5352 10014 5364
rect 10686 5352 10692 5364
rect 10008 5324 10692 5352
rect 10008 5312 10014 5324
rect 10686 5312 10692 5324
rect 10744 5312 10750 5364
rect 11054 5312 11060 5364
rect 11112 5352 11118 5364
rect 11238 5352 11244 5364
rect 11112 5324 11244 5352
rect 11112 5312 11118 5324
rect 11238 5312 11244 5324
rect 11296 5312 11302 5364
rect 12066 5312 12072 5364
rect 12124 5352 12130 5364
rect 12161 5355 12219 5361
rect 12161 5352 12173 5355
rect 12124 5324 12173 5352
rect 12124 5312 12130 5324
rect 12161 5321 12173 5324
rect 12207 5321 12219 5355
rect 12161 5315 12219 5321
rect 1397 5287 1455 5293
rect 1397 5253 1409 5287
rect 1443 5284 1455 5287
rect 2866 5284 2872 5296
rect 1443 5256 2872 5284
rect 1443 5253 1455 5256
rect 1397 5247 1455 5253
rect 2866 5244 2872 5256
rect 2924 5284 2930 5296
rect 4062 5284 4068 5296
rect 2924 5256 4068 5284
rect 2924 5244 2930 5256
rect 4062 5244 4068 5256
rect 4120 5244 4126 5296
rect 4893 5287 4951 5293
rect 4893 5253 4905 5287
rect 4939 5284 4951 5287
rect 9214 5284 9220 5296
rect 4939 5256 5764 5284
rect 9175 5256 9220 5284
rect 4939 5253 4951 5256
rect 4893 5247 4951 5253
rect 1854 5216 1860 5228
rect 1815 5188 1860 5216
rect 1854 5176 1860 5188
rect 1912 5176 1918 5228
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5216 2099 5219
rect 2406 5216 2412 5228
rect 2087 5188 2412 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 2406 5176 2412 5188
rect 2464 5176 2470 5228
rect 3694 5176 3700 5228
rect 3752 5216 3758 5228
rect 5736 5225 5764 5256
rect 9214 5244 9220 5256
rect 9272 5284 9278 5296
rect 12176 5284 12204 5315
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 12989 5355 13047 5361
rect 12989 5352 13001 5355
rect 12492 5324 13001 5352
rect 12492 5312 12498 5324
rect 12989 5321 13001 5324
rect 13035 5321 13047 5355
rect 12989 5315 13047 5321
rect 14826 5312 14832 5364
rect 14884 5352 14890 5364
rect 14921 5355 14979 5361
rect 14921 5352 14933 5355
rect 14884 5324 14933 5352
rect 14884 5312 14890 5324
rect 14921 5321 14933 5324
rect 14967 5321 14979 5355
rect 14921 5315 14979 5321
rect 15565 5355 15623 5361
rect 15565 5321 15577 5355
rect 15611 5352 15623 5355
rect 15930 5352 15936 5364
rect 15611 5324 15936 5352
rect 15611 5321 15623 5324
rect 15565 5315 15623 5321
rect 15930 5312 15936 5324
rect 15988 5312 15994 5364
rect 16393 5355 16451 5361
rect 16393 5321 16405 5355
rect 16439 5352 16451 5355
rect 16482 5352 16488 5364
rect 16439 5324 16488 5352
rect 16439 5321 16451 5324
rect 16393 5315 16451 5321
rect 16482 5312 16488 5324
rect 16540 5312 16546 5364
rect 19426 5352 19432 5364
rect 19387 5324 19432 5352
rect 19426 5312 19432 5324
rect 19484 5312 19490 5364
rect 21358 5312 21364 5364
rect 21416 5352 21422 5364
rect 21913 5355 21971 5361
rect 21913 5352 21925 5355
rect 21416 5324 21925 5352
rect 21416 5312 21422 5324
rect 21913 5321 21925 5324
rect 21959 5321 21971 5355
rect 23290 5352 23296 5364
rect 23251 5324 23296 5352
rect 21913 5315 21971 5321
rect 23290 5312 23296 5324
rect 23348 5312 23354 5364
rect 13357 5287 13415 5293
rect 13357 5284 13369 5287
rect 9272 5256 9352 5284
rect 12176 5256 13369 5284
rect 9272 5244 9278 5256
rect 9324 5225 9352 5256
rect 13357 5253 13369 5256
rect 13403 5284 13415 5287
rect 13403 5256 13584 5284
rect 13403 5253 13415 5256
rect 13357 5247 13415 5253
rect 4249 5219 4307 5225
rect 4249 5216 4261 5219
rect 3752 5188 4261 5216
rect 3752 5176 3758 5188
rect 4249 5185 4261 5188
rect 4295 5216 4307 5219
rect 5721 5219 5779 5225
rect 4295 5188 5396 5216
rect 4295 5185 4307 5188
rect 4249 5179 4307 5185
rect 5368 5160 5396 5188
rect 5721 5185 5733 5219
rect 5767 5185 5779 5219
rect 5721 5179 5779 5185
rect 9309 5219 9367 5225
rect 9309 5185 9321 5219
rect 9355 5185 9367 5219
rect 11238 5216 11244 5228
rect 11199 5188 11244 5216
rect 9309 5179 9367 5185
rect 1394 5108 1400 5160
rect 1452 5148 1458 5160
rect 1765 5151 1823 5157
rect 1765 5148 1777 5151
rect 1452 5120 1777 5148
rect 1452 5108 1458 5120
rect 1765 5117 1777 5120
rect 1811 5117 1823 5151
rect 1765 5111 1823 5117
rect 2501 5151 2559 5157
rect 2501 5117 2513 5151
rect 2547 5148 2559 5151
rect 3050 5148 3056 5160
rect 2547 5120 3056 5148
rect 2547 5117 2559 5120
rect 2501 5111 2559 5117
rect 3050 5108 3056 5120
rect 3108 5108 3114 5160
rect 3145 5151 3203 5157
rect 3145 5117 3157 5151
rect 3191 5148 3203 5151
rect 4614 5148 4620 5160
rect 3191 5120 4620 5148
rect 3191 5117 3203 5120
rect 3145 5111 3203 5117
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 5350 5108 5356 5160
rect 5408 5148 5414 5160
rect 5534 5148 5540 5160
rect 5408 5120 5540 5148
rect 5408 5108 5414 5120
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 6454 5108 6460 5160
rect 6512 5148 6518 5160
rect 6641 5151 6699 5157
rect 6641 5148 6653 5151
rect 6512 5120 6653 5148
rect 6512 5108 6518 5120
rect 6641 5117 6653 5120
rect 6687 5148 6699 5151
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6687 5120 6837 5148
rect 6687 5117 6699 5120
rect 6641 5111 6699 5117
rect 6825 5117 6837 5120
rect 6871 5148 6883 5151
rect 9324 5148 9352 5179
rect 11238 5176 11244 5188
rect 11296 5176 11302 5228
rect 13556 5225 13584 5256
rect 19334 5244 19340 5296
rect 19392 5284 19398 5296
rect 20073 5287 20131 5293
rect 20073 5284 20085 5287
rect 19392 5256 20085 5284
rect 19392 5244 19398 5256
rect 20073 5253 20085 5256
rect 20119 5284 20131 5287
rect 22281 5287 22339 5293
rect 22281 5284 22293 5287
rect 20119 5256 22293 5284
rect 20119 5253 20131 5256
rect 20073 5247 20131 5253
rect 22281 5253 22293 5256
rect 22327 5253 22339 5287
rect 22281 5247 22339 5253
rect 13541 5219 13599 5225
rect 13541 5185 13553 5219
rect 13587 5185 13599 5219
rect 13541 5179 13599 5185
rect 16301 5219 16359 5225
rect 16301 5185 16313 5219
rect 16347 5216 16359 5219
rect 16945 5219 17003 5225
rect 16945 5216 16957 5219
rect 16347 5188 16957 5216
rect 16347 5185 16359 5188
rect 16301 5179 16359 5185
rect 16945 5185 16957 5188
rect 16991 5216 17003 5219
rect 17862 5216 17868 5228
rect 16991 5188 17868 5216
rect 16991 5185 17003 5188
rect 16945 5179 17003 5185
rect 17862 5176 17868 5188
rect 17920 5216 17926 5228
rect 17920 5188 18184 5216
rect 17920 5176 17926 5188
rect 18156 5160 18184 5188
rect 20530 5176 20536 5228
rect 20588 5216 20594 5228
rect 21085 5219 21143 5225
rect 21085 5216 21097 5219
rect 20588 5188 21097 5216
rect 20588 5176 20594 5188
rect 21085 5185 21097 5188
rect 21131 5185 21143 5219
rect 21085 5179 21143 5185
rect 6871 5120 9352 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 9398 5108 9404 5160
rect 9456 5148 9462 5160
rect 9565 5151 9623 5157
rect 9565 5148 9577 5151
rect 9456 5120 9577 5148
rect 9456 5108 9462 5120
rect 9565 5117 9577 5120
rect 9611 5117 9623 5151
rect 9565 5111 9623 5117
rect 12342 5108 12348 5160
rect 12400 5148 12406 5160
rect 12529 5151 12587 5157
rect 12529 5148 12541 5151
rect 12400 5120 12541 5148
rect 12400 5108 12406 5120
rect 12529 5117 12541 5120
rect 12575 5148 12587 5151
rect 12618 5148 12624 5160
rect 12575 5120 12624 5148
rect 12575 5117 12587 5120
rect 12529 5111 12587 5117
rect 12618 5108 12624 5120
rect 12676 5108 12682 5160
rect 16850 5148 16856 5160
rect 16811 5120 16856 5148
rect 16850 5108 16856 5120
rect 16908 5108 16914 5160
rect 17402 5148 17408 5160
rect 17315 5120 17408 5148
rect 17402 5108 17408 5120
rect 17460 5148 17466 5160
rect 18049 5151 18107 5157
rect 18049 5148 18061 5151
rect 17460 5120 18061 5148
rect 17460 5108 17466 5120
rect 18049 5117 18061 5120
rect 18095 5117 18107 5151
rect 18049 5111 18107 5117
rect 3329 5083 3387 5089
rect 3329 5049 3341 5083
rect 3375 5080 3387 5083
rect 5626 5080 5632 5092
rect 3375 5052 5632 5080
rect 3375 5049 3387 5052
rect 3329 5043 3387 5049
rect 5626 5040 5632 5052
rect 5684 5040 5690 5092
rect 6270 5080 6276 5092
rect 6183 5052 6276 5080
rect 6270 5040 6276 5052
rect 6328 5080 6334 5092
rect 7070 5083 7128 5089
rect 7070 5080 7082 5083
rect 6328 5052 7082 5080
rect 6328 5040 6334 5052
rect 7070 5049 7082 5052
rect 7116 5049 7128 5083
rect 11606 5080 11612 5092
rect 11567 5052 11612 5080
rect 7070 5043 7128 5049
rect 11606 5040 11612 5052
rect 11664 5040 11670 5092
rect 13630 5040 13636 5092
rect 13688 5080 13694 5092
rect 13786 5083 13844 5089
rect 13786 5080 13798 5083
rect 13688 5052 13798 5080
rect 13688 5040 13694 5052
rect 13786 5049 13798 5052
rect 13832 5049 13844 5083
rect 13786 5043 13844 5049
rect 16574 5040 16580 5092
rect 16632 5080 16638 5092
rect 16761 5083 16819 5089
rect 16761 5080 16773 5083
rect 16632 5052 16773 5080
rect 16632 5040 16638 5052
rect 16761 5049 16773 5052
rect 16807 5080 16819 5083
rect 17494 5080 17500 5092
rect 16807 5052 17500 5080
rect 16807 5049 16819 5052
rect 16761 5043 16819 5049
rect 17494 5040 17500 5052
rect 17552 5040 17558 5092
rect 17865 5083 17923 5089
rect 17865 5049 17877 5083
rect 17911 5080 17923 5083
rect 18064 5080 18092 5111
rect 18138 5108 18144 5160
rect 18196 5148 18202 5160
rect 18305 5151 18363 5157
rect 18305 5148 18317 5151
rect 18196 5120 18317 5148
rect 18196 5108 18202 5120
rect 18305 5117 18317 5120
rect 18351 5117 18363 5151
rect 18305 5111 18363 5117
rect 20990 5108 20996 5160
rect 21048 5148 21054 5160
rect 21545 5151 21603 5157
rect 21545 5148 21557 5151
rect 21048 5120 21557 5148
rect 21048 5108 21054 5120
rect 21545 5117 21557 5120
rect 21591 5117 21603 5151
rect 21545 5111 21603 5117
rect 22097 5151 22155 5157
rect 22097 5117 22109 5151
rect 22143 5148 22155 5151
rect 22186 5148 22192 5160
rect 22143 5120 22192 5148
rect 22143 5117 22155 5120
rect 22097 5111 22155 5117
rect 22186 5108 22192 5120
rect 22244 5148 22250 5160
rect 22557 5151 22615 5157
rect 22557 5148 22569 5151
rect 22244 5120 22569 5148
rect 22244 5108 22250 5120
rect 22557 5117 22569 5120
rect 22603 5117 22615 5151
rect 22557 5111 22615 5117
rect 18414 5080 18420 5092
rect 17911 5052 18420 5080
rect 17911 5049 17923 5052
rect 17865 5043 17923 5049
rect 18414 5040 18420 5052
rect 18472 5040 18478 5092
rect 20364 5052 21036 5080
rect 3513 5015 3571 5021
rect 3513 4981 3525 5015
rect 3559 5012 3571 5015
rect 3694 5012 3700 5024
rect 3559 4984 3700 5012
rect 3559 4981 3571 4984
rect 3513 4975 3571 4981
rect 3694 4972 3700 4984
rect 3752 5012 3758 5024
rect 3973 5015 4031 5021
rect 3973 5012 3985 5015
rect 3752 4984 3985 5012
rect 3752 4972 3758 4984
rect 3973 4981 3985 4984
rect 4019 4981 4031 5015
rect 3973 4975 4031 4981
rect 4065 5015 4123 5021
rect 4065 4981 4077 5015
rect 4111 5012 4123 5015
rect 4154 5012 4160 5024
rect 4111 4984 4160 5012
rect 4111 4981 4123 4984
rect 4065 4975 4123 4981
rect 4154 4972 4160 4984
rect 4212 4972 4218 5024
rect 4706 4972 4712 5024
rect 4764 5012 4770 5024
rect 4893 5015 4951 5021
rect 4893 5012 4905 5015
rect 4764 4984 4905 5012
rect 4764 4972 4770 4984
rect 4893 4981 4905 4984
rect 4939 5012 4951 5015
rect 4985 5015 5043 5021
rect 4985 5012 4997 5015
rect 4939 4984 4997 5012
rect 4939 4981 4951 4984
rect 4893 4975 4951 4981
rect 4985 4981 4997 4984
rect 5031 4981 5043 5015
rect 5166 5012 5172 5024
rect 5127 4984 5172 5012
rect 4985 4975 5043 4981
rect 5166 4972 5172 4984
rect 5224 4972 5230 5024
rect 5534 5012 5540 5024
rect 5495 4984 5540 5012
rect 5534 4972 5540 4984
rect 5592 4972 5598 5024
rect 7742 4972 7748 5024
rect 7800 5012 7806 5024
rect 8205 5015 8263 5021
rect 8205 5012 8217 5015
rect 7800 4984 8217 5012
rect 7800 4972 7806 4984
rect 8205 4981 8217 4984
rect 8251 4981 8263 5015
rect 8205 4975 8263 4981
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 12713 5015 12771 5021
rect 12713 5012 12725 5015
rect 12492 4984 12725 5012
rect 12492 4972 12498 4984
rect 12713 4981 12725 4984
rect 12759 4981 12771 5015
rect 12713 4975 12771 4981
rect 19426 4972 19432 5024
rect 19484 5012 19490 5024
rect 20364 5021 20392 5052
rect 20349 5015 20407 5021
rect 20349 5012 20361 5015
rect 19484 4984 20361 5012
rect 19484 4972 19490 4984
rect 20349 4981 20361 4984
rect 20395 4981 20407 5015
rect 20530 5012 20536 5024
rect 20491 4984 20536 5012
rect 20349 4975 20407 4981
rect 20530 4972 20536 4984
rect 20588 4972 20594 5024
rect 20714 4972 20720 5024
rect 20772 5012 20778 5024
rect 21008 5021 21036 5052
rect 20901 5015 20959 5021
rect 20901 5012 20913 5015
rect 20772 4984 20913 5012
rect 20772 4972 20778 4984
rect 20901 4981 20913 4984
rect 20947 4981 20959 5015
rect 20901 4975 20959 4981
rect 20993 5015 21051 5021
rect 20993 4981 21005 5015
rect 21039 4981 21051 5015
rect 20993 4975 21051 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1673 4811 1731 4817
rect 1673 4777 1685 4811
rect 1719 4808 1731 4811
rect 2130 4808 2136 4820
rect 1719 4780 2136 4808
rect 1719 4777 1731 4780
rect 1673 4771 1731 4777
rect 2130 4768 2136 4780
rect 2188 4768 2194 4820
rect 2777 4811 2835 4817
rect 2777 4777 2789 4811
rect 2823 4808 2835 4811
rect 2866 4808 2872 4820
rect 2823 4780 2872 4808
rect 2823 4777 2835 4780
rect 2777 4771 2835 4777
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 4433 4811 4491 4817
rect 4433 4777 4445 4811
rect 4479 4808 4491 4811
rect 5166 4808 5172 4820
rect 4479 4780 5172 4808
rect 4479 4777 4491 4780
rect 4433 4771 4491 4777
rect 5166 4768 5172 4780
rect 5224 4808 5230 4820
rect 5534 4808 5540 4820
rect 5224 4780 5540 4808
rect 5224 4768 5230 4780
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 6362 4808 6368 4820
rect 6323 4780 6368 4808
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 7098 4808 7104 4820
rect 7059 4780 7104 4808
rect 7098 4768 7104 4780
rect 7156 4768 7162 4820
rect 7558 4808 7564 4820
rect 7519 4780 7564 4808
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 8018 4808 8024 4820
rect 7979 4780 8024 4808
rect 8018 4768 8024 4780
rect 8076 4768 8082 4820
rect 8938 4808 8944 4820
rect 8899 4780 8944 4808
rect 8938 4768 8944 4780
rect 8996 4768 9002 4820
rect 9030 4768 9036 4820
rect 9088 4808 9094 4820
rect 9214 4808 9220 4820
rect 9088 4780 9220 4808
rect 9088 4768 9094 4780
rect 9214 4768 9220 4780
rect 9272 4808 9278 4820
rect 9309 4811 9367 4817
rect 9309 4808 9321 4811
rect 9272 4780 9321 4808
rect 9272 4768 9278 4780
rect 9309 4777 9321 4780
rect 9355 4777 9367 4811
rect 10962 4808 10968 4820
rect 10923 4780 10968 4808
rect 9309 4771 9367 4777
rect 10962 4768 10968 4780
rect 11020 4768 11026 4820
rect 11425 4811 11483 4817
rect 11425 4777 11437 4811
rect 11471 4808 11483 4811
rect 11790 4808 11796 4820
rect 11471 4780 11796 4808
rect 11471 4777 11483 4780
rect 11425 4771 11483 4777
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 12802 4768 12808 4820
rect 12860 4808 12866 4820
rect 12989 4811 13047 4817
rect 12989 4808 13001 4811
rect 12860 4780 13001 4808
rect 12860 4768 12866 4780
rect 12989 4777 13001 4780
rect 13035 4808 13047 4811
rect 13722 4808 13728 4820
rect 13035 4780 13728 4808
rect 13035 4777 13047 4780
rect 12989 4771 13047 4777
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 15470 4808 15476 4820
rect 15431 4780 15476 4808
rect 15470 4768 15476 4780
rect 15528 4768 15534 4820
rect 15930 4768 15936 4820
rect 15988 4808 15994 4820
rect 16117 4811 16175 4817
rect 16117 4808 16129 4811
rect 15988 4780 16129 4808
rect 15988 4768 15994 4780
rect 16117 4777 16129 4780
rect 16163 4777 16175 4811
rect 17218 4808 17224 4820
rect 16117 4771 16175 4777
rect 16224 4780 17224 4808
rect 2682 4700 2688 4752
rect 2740 4740 2746 4752
rect 2740 4712 2912 4740
rect 2740 4700 2746 4712
rect 2884 4684 2912 4712
rect 5442 4700 5448 4752
rect 5500 4740 5506 4752
rect 5994 4740 6000 4752
rect 5500 4712 6000 4740
rect 5500 4700 5506 4712
rect 5994 4700 6000 4712
rect 6052 4740 6058 4752
rect 6457 4743 6515 4749
rect 6457 4740 6469 4743
rect 6052 4712 6469 4740
rect 6052 4700 6058 4712
rect 6457 4709 6469 4712
rect 6503 4709 6515 4743
rect 10778 4740 10784 4752
rect 10739 4712 10784 4740
rect 6457 4703 6515 4709
rect 10778 4700 10784 4712
rect 10836 4700 10842 4752
rect 11333 4743 11391 4749
rect 11333 4709 11345 4743
rect 11379 4740 11391 4743
rect 11974 4740 11980 4752
rect 11379 4712 11980 4740
rect 11379 4709 11391 4712
rect 11333 4703 11391 4709
rect 11974 4700 11980 4712
rect 12032 4700 12038 4752
rect 12250 4700 12256 4752
rect 12308 4740 12314 4752
rect 12897 4743 12955 4749
rect 12897 4740 12909 4743
rect 12308 4712 12909 4740
rect 12308 4700 12314 4712
rect 12897 4709 12909 4712
rect 12943 4740 12955 4743
rect 14645 4743 14703 4749
rect 14645 4740 14657 4743
rect 12943 4712 14657 4740
rect 12943 4709 12955 4712
rect 12897 4703 12955 4709
rect 14645 4709 14657 4712
rect 14691 4709 14703 4743
rect 14645 4703 14703 4709
rect 14826 4700 14832 4752
rect 14884 4740 14890 4752
rect 15105 4743 15163 4749
rect 15105 4740 15117 4743
rect 14884 4712 15117 4740
rect 14884 4700 14890 4712
rect 15105 4709 15117 4712
rect 15151 4740 15163 4743
rect 16224 4740 16252 4780
rect 17218 4768 17224 4780
rect 17276 4768 17282 4820
rect 17862 4808 17868 4820
rect 17823 4780 17868 4808
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 19334 4768 19340 4820
rect 19392 4808 19398 4820
rect 19392 4780 19656 4808
rect 19392 4768 19398 4780
rect 15151 4712 16252 4740
rect 15151 4709 15163 4712
rect 15105 4703 15163 4709
rect 16666 4700 16672 4752
rect 16724 4740 16730 4752
rect 16724 4712 17632 4740
rect 16724 4700 16730 4712
rect 2866 4632 2872 4684
rect 2924 4672 2930 4684
rect 2924 4644 2969 4672
rect 2924 4632 2930 4644
rect 4430 4632 4436 4684
rect 4488 4672 4494 4684
rect 4801 4675 4859 4681
rect 4801 4672 4813 4675
rect 4488 4644 4813 4672
rect 4488 4632 4494 4644
rect 4801 4641 4813 4644
rect 4847 4641 4859 4675
rect 4801 4635 4859 4641
rect 4893 4675 4951 4681
rect 4893 4641 4905 4675
rect 4939 4672 4951 4675
rect 5537 4675 5595 4681
rect 4939 4644 5488 4672
rect 4939 4641 4951 4644
rect 4893 4635 4951 4641
rect 3050 4604 3056 4616
rect 3011 4576 3056 4604
rect 3050 4564 3056 4576
rect 3108 4564 3114 4616
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4908 4604 4936 4635
rect 4212 4576 4936 4604
rect 5077 4607 5135 4613
rect 4212 4564 4218 4576
rect 5077 4573 5089 4607
rect 5123 4604 5135 4607
rect 5350 4604 5356 4616
rect 5123 4576 5356 4604
rect 5123 4573 5135 4576
rect 5077 4567 5135 4573
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 5460 4604 5488 4644
rect 5537 4641 5549 4675
rect 5583 4672 5595 4675
rect 5626 4672 5632 4684
rect 5583 4644 5632 4672
rect 5583 4641 5595 4644
rect 5537 4635 5595 4641
rect 5626 4632 5632 4644
rect 5684 4632 5690 4684
rect 7190 4632 7196 4684
rect 7248 4672 7254 4684
rect 7929 4675 7987 4681
rect 7929 4672 7941 4675
rect 7248 4644 7941 4672
rect 7248 4632 7254 4644
rect 7929 4641 7941 4644
rect 7975 4641 7987 4675
rect 7929 4635 7987 4641
rect 9953 4675 10011 4681
rect 9953 4641 9965 4675
rect 9999 4641 10011 4675
rect 12437 4675 12495 4681
rect 12437 4672 12449 4675
rect 9953 4635 10011 4641
rect 11624 4644 12449 4672
rect 5905 4607 5963 4613
rect 5460 4576 5856 4604
rect 3697 4539 3755 4545
rect 3697 4505 3709 4539
rect 3743 4536 3755 4539
rect 4062 4536 4068 4548
rect 3743 4508 4068 4536
rect 3743 4505 3755 4508
rect 3697 4499 3755 4505
rect 4062 4496 4068 4508
rect 4120 4536 4126 4548
rect 5534 4536 5540 4548
rect 4120 4508 5540 4536
rect 4120 4496 4126 4508
rect 5534 4496 5540 4508
rect 5592 4496 5598 4548
rect 2314 4468 2320 4480
rect 2275 4440 2320 4468
rect 2314 4428 2320 4440
rect 2372 4428 2378 4480
rect 2409 4471 2467 4477
rect 2409 4437 2421 4471
rect 2455 4468 2467 4471
rect 2866 4468 2872 4480
rect 2455 4440 2872 4468
rect 2455 4437 2467 4440
rect 2409 4431 2467 4437
rect 2866 4428 2872 4440
rect 2924 4428 2930 4480
rect 4338 4468 4344 4480
rect 4299 4440 4344 4468
rect 4338 4428 4344 4440
rect 4396 4428 4402 4480
rect 5828 4468 5856 4576
rect 5905 4573 5917 4607
rect 5951 4604 5963 4607
rect 6641 4607 6699 4613
rect 6641 4604 6653 4607
rect 5951 4576 6653 4604
rect 5951 4573 5963 4576
rect 5905 4567 5963 4573
rect 6641 4573 6653 4576
rect 6687 4604 6699 4607
rect 8113 4607 8171 4613
rect 6687 4576 7604 4604
rect 6687 4573 6699 4576
rect 6641 4567 6699 4573
rect 7576 4548 7604 4576
rect 8113 4573 8125 4607
rect 8159 4573 8171 4607
rect 9968 4604 9996 4635
rect 10505 4607 10563 4613
rect 10505 4604 10517 4607
rect 9968 4576 10517 4604
rect 8113 4567 8171 4573
rect 10505 4573 10517 4576
rect 10551 4604 10563 4607
rect 10778 4604 10784 4616
rect 10551 4576 10784 4604
rect 10551 4573 10563 4576
rect 10505 4567 10563 4573
rect 5997 4539 6055 4545
rect 5997 4505 6009 4539
rect 6043 4536 6055 4539
rect 6822 4536 6828 4548
rect 6043 4508 6828 4536
rect 6043 4505 6055 4508
rect 5997 4499 6055 4505
rect 6822 4496 6828 4508
rect 6880 4496 6886 4548
rect 7558 4496 7564 4548
rect 7616 4536 7622 4548
rect 7926 4536 7932 4548
rect 7616 4508 7932 4536
rect 7616 4496 7622 4508
rect 7926 4496 7932 4508
rect 7984 4536 7990 4548
rect 8128 4536 8156 4567
rect 10778 4564 10784 4576
rect 10836 4564 10842 4616
rect 11514 4564 11520 4616
rect 11572 4604 11578 4616
rect 11624 4613 11652 4644
rect 12437 4641 12449 4644
rect 12483 4672 12495 4675
rect 13262 4672 13268 4684
rect 12483 4644 13268 4672
rect 12483 4641 12495 4644
rect 12437 4635 12495 4641
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 13630 4672 13636 4684
rect 13591 4644 13636 4672
rect 13630 4632 13636 4644
rect 13688 4632 13694 4684
rect 14090 4672 14096 4684
rect 14051 4644 14096 4672
rect 14090 4632 14096 4644
rect 14148 4632 14154 4684
rect 15289 4675 15347 4681
rect 15289 4641 15301 4675
rect 15335 4672 15347 4675
rect 15378 4672 15384 4684
rect 15335 4644 15384 4672
rect 15335 4641 15347 4644
rect 15289 4635 15347 4641
rect 15378 4632 15384 4644
rect 15436 4672 15442 4684
rect 16298 4672 16304 4684
rect 15436 4644 16304 4672
rect 15436 4632 15442 4644
rect 16298 4632 16304 4644
rect 16356 4632 16362 4684
rect 16853 4675 16911 4681
rect 16853 4641 16865 4675
rect 16899 4672 16911 4675
rect 17034 4672 17040 4684
rect 16899 4644 17040 4672
rect 16899 4641 16911 4644
rect 16853 4635 16911 4641
rect 17034 4632 17040 4644
rect 17092 4632 17098 4684
rect 17604 4681 17632 4712
rect 18046 4700 18052 4752
rect 18104 4740 18110 4752
rect 18417 4743 18475 4749
rect 18417 4740 18429 4743
rect 18104 4712 18429 4740
rect 18104 4700 18110 4712
rect 18417 4709 18429 4712
rect 18463 4740 18475 4743
rect 19429 4743 19487 4749
rect 19429 4740 19441 4743
rect 18463 4712 19441 4740
rect 18463 4709 18475 4712
rect 18417 4703 18475 4709
rect 19429 4709 19441 4712
rect 19475 4709 19487 4743
rect 19429 4703 19487 4709
rect 17589 4675 17647 4681
rect 17589 4641 17601 4675
rect 17635 4672 17647 4675
rect 18509 4675 18567 4681
rect 17635 4644 18276 4672
rect 17635 4641 17647 4644
rect 17589 4635 17647 4641
rect 11609 4607 11667 4613
rect 11609 4604 11621 4607
rect 11572 4576 11621 4604
rect 11572 4564 11578 4576
rect 11609 4573 11621 4576
rect 11655 4573 11667 4607
rect 13170 4604 13176 4616
rect 13131 4576 13176 4604
rect 11609 4567 11667 4573
rect 13170 4564 13176 4576
rect 13228 4564 13234 4616
rect 16942 4604 16948 4616
rect 16903 4576 16948 4604
rect 16942 4564 16948 4576
rect 17000 4564 17006 4616
rect 17129 4607 17187 4613
rect 17129 4573 17141 4607
rect 17175 4604 17187 4607
rect 18138 4604 18144 4616
rect 17175 4576 18144 4604
rect 17175 4573 17187 4576
rect 17129 4567 17187 4573
rect 8662 4536 8668 4548
rect 7984 4508 8156 4536
rect 8575 4508 8668 4536
rect 7984 4496 7990 4508
rect 8662 4496 8668 4508
rect 8720 4536 8726 4548
rect 9766 4536 9772 4548
rect 8720 4508 9772 4536
rect 8720 4496 8726 4508
rect 9766 4496 9772 4508
rect 9824 4496 9830 4548
rect 12069 4539 12127 4545
rect 12069 4505 12081 4539
rect 12115 4536 12127 4539
rect 13188 4536 13216 4564
rect 12115 4508 13216 4536
rect 12115 4505 12127 4508
rect 12069 4499 12127 4505
rect 16390 4496 16396 4548
rect 16448 4536 16454 4548
rect 17144 4536 17172 4567
rect 18138 4564 18144 4576
rect 18196 4564 18202 4616
rect 18248 4604 18276 4644
rect 18509 4641 18521 4675
rect 18555 4672 18567 4675
rect 19061 4675 19119 4681
rect 19061 4672 19073 4675
rect 18555 4644 19073 4672
rect 18555 4641 18567 4644
rect 18509 4635 18567 4641
rect 19061 4641 19073 4644
rect 19107 4672 19119 4675
rect 19334 4672 19340 4684
rect 19107 4644 19340 4672
rect 19107 4641 19119 4644
rect 19061 4635 19119 4641
rect 19334 4632 19340 4644
rect 19392 4632 19398 4684
rect 19628 4681 19656 4780
rect 20530 4768 20536 4820
rect 20588 4808 20594 4820
rect 21266 4808 21272 4820
rect 20588 4780 21272 4808
rect 20588 4768 20594 4780
rect 21266 4768 21272 4780
rect 21324 4808 21330 4820
rect 21453 4811 21511 4817
rect 21453 4808 21465 4811
rect 21324 4780 21465 4808
rect 21324 4768 21330 4780
rect 21453 4777 21465 4780
rect 21499 4777 21511 4811
rect 21453 4771 21511 4777
rect 19613 4675 19671 4681
rect 19613 4641 19625 4675
rect 19659 4641 19671 4675
rect 20898 4672 20904 4684
rect 20859 4644 20904 4672
rect 19613 4635 19671 4641
rect 20898 4632 20904 4644
rect 20956 4632 20962 4684
rect 18601 4607 18659 4613
rect 18601 4604 18613 4607
rect 18248 4576 18613 4604
rect 18601 4573 18613 4576
rect 18647 4573 18659 4607
rect 18601 4567 18659 4573
rect 19426 4564 19432 4616
rect 19484 4604 19490 4616
rect 20533 4607 20591 4613
rect 20533 4604 20545 4607
rect 19484 4576 20545 4604
rect 19484 4564 19490 4576
rect 20533 4573 20545 4576
rect 20579 4604 20591 4607
rect 20714 4604 20720 4616
rect 20579 4576 20720 4604
rect 20579 4573 20591 4576
rect 20533 4567 20591 4573
rect 20714 4564 20720 4576
rect 20772 4564 20778 4616
rect 16448 4508 17172 4536
rect 16448 4496 16454 4508
rect 17954 4496 17960 4548
rect 18012 4536 18018 4548
rect 18049 4539 18107 4545
rect 18049 4536 18061 4539
rect 18012 4508 18061 4536
rect 18012 4496 18018 4508
rect 18049 4505 18061 4508
rect 18095 4505 18107 4539
rect 18049 4499 18107 4505
rect 20254 4496 20260 4548
rect 20312 4536 20318 4548
rect 21085 4539 21143 4545
rect 21085 4536 21097 4539
rect 20312 4508 21097 4536
rect 20312 4496 20318 4508
rect 21085 4505 21097 4508
rect 21131 4505 21143 4539
rect 21085 4499 21143 4505
rect 6270 4468 6276 4480
rect 5828 4440 6276 4468
rect 6270 4428 6276 4440
rect 6328 4428 6334 4480
rect 7469 4471 7527 4477
rect 7469 4437 7481 4471
rect 7515 4468 7527 4471
rect 7742 4468 7748 4480
rect 7515 4440 7748 4468
rect 7515 4437 7527 4440
rect 7469 4431 7527 4437
rect 7742 4428 7748 4440
rect 7800 4428 7806 4480
rect 10134 4468 10140 4480
rect 10095 4440 10140 4468
rect 10134 4428 10140 4440
rect 10192 4428 10198 4480
rect 12526 4468 12532 4480
rect 12487 4440 12532 4468
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 13814 4428 13820 4480
rect 13872 4468 13878 4480
rect 13909 4471 13967 4477
rect 13909 4468 13921 4471
rect 13872 4440 13921 4468
rect 13872 4428 13878 4440
rect 13909 4437 13921 4440
rect 13955 4437 13967 4471
rect 14274 4468 14280 4480
rect 14235 4440 14280 4468
rect 13909 4431 13967 4437
rect 14274 4428 14280 4440
rect 14332 4428 14338 4480
rect 16482 4468 16488 4480
rect 16443 4440 16488 4468
rect 16482 4428 16488 4440
rect 16540 4428 16546 4480
rect 19794 4468 19800 4480
rect 19755 4440 19800 4468
rect 19794 4428 19800 4440
rect 19852 4428 19858 4480
rect 20070 4428 20076 4480
rect 20128 4468 20134 4480
rect 20165 4471 20223 4477
rect 20165 4468 20177 4471
rect 20128 4440 20177 4468
rect 20128 4428 20134 4440
rect 20165 4437 20177 4440
rect 20211 4437 20223 4471
rect 20165 4431 20223 4437
rect 20714 4428 20720 4480
rect 20772 4468 20778 4480
rect 21821 4471 21879 4477
rect 21821 4468 21833 4471
rect 20772 4440 21833 4468
rect 20772 4428 20778 4440
rect 21821 4437 21833 4440
rect 21867 4437 21879 4471
rect 21821 4431 21879 4437
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 3789 4267 3847 4273
rect 3789 4233 3801 4267
rect 3835 4264 3847 4267
rect 4154 4264 4160 4276
rect 3835 4236 4160 4264
rect 3835 4233 3847 4236
rect 3789 4227 3847 4233
rect 4154 4224 4160 4236
rect 4212 4224 4218 4276
rect 5994 4264 6000 4276
rect 5955 4236 6000 4264
rect 5994 4224 6000 4236
rect 6052 4224 6058 4276
rect 6362 4264 6368 4276
rect 6323 4236 6368 4264
rect 6362 4224 6368 4236
rect 6420 4224 6426 4276
rect 7285 4267 7343 4273
rect 7285 4233 7297 4267
rect 7331 4264 7343 4267
rect 8018 4264 8024 4276
rect 7331 4236 8024 4264
rect 7331 4233 7343 4236
rect 7285 4227 7343 4233
rect 8018 4224 8024 4236
rect 8076 4224 8082 4276
rect 10689 4267 10747 4273
rect 10689 4233 10701 4267
rect 10735 4264 10747 4267
rect 11514 4264 11520 4276
rect 10735 4236 11520 4264
rect 10735 4233 10747 4236
rect 10689 4227 10747 4233
rect 2314 4156 2320 4208
rect 2372 4196 2378 4208
rect 8662 4196 8668 4208
rect 2372 4168 2912 4196
rect 2372 4156 2378 4168
rect 1762 4128 1768 4140
rect 1723 4100 1768 4128
rect 1762 4088 1768 4100
rect 1820 4088 1826 4140
rect 2682 4088 2688 4140
rect 2740 4128 2746 4140
rect 2777 4131 2835 4137
rect 2777 4128 2789 4131
rect 2740 4100 2789 4128
rect 2740 4088 2746 4100
rect 2777 4097 2789 4100
rect 2823 4097 2835 4131
rect 2884 4128 2912 4168
rect 8496 4168 8668 4196
rect 2961 4131 3019 4137
rect 2961 4128 2973 4131
rect 2884 4100 2973 4128
rect 2777 4091 2835 4097
rect 2961 4097 2973 4100
rect 3007 4128 3019 4131
rect 3050 4128 3056 4140
rect 3007 4100 3056 4128
rect 3007 4097 3019 4100
rect 2961 4091 3019 4097
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 8202 4088 8208 4140
rect 8260 4128 8266 4140
rect 8496 4137 8524 4168
rect 8662 4156 8668 4168
rect 8720 4156 8726 4208
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 8260 4100 8309 4128
rect 8260 4088 8266 4100
rect 8297 4097 8309 4100
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 8481 4131 8539 4137
rect 8481 4097 8493 4131
rect 8527 4097 8539 4131
rect 8481 4091 8539 4097
rect 8941 4131 8999 4137
rect 8941 4097 8953 4131
rect 8987 4128 8999 4131
rect 9950 4128 9956 4140
rect 8987 4100 9956 4128
rect 8987 4097 8999 4100
rect 8941 4091 8999 4097
rect 3421 4063 3479 4069
rect 3421 4029 3433 4063
rect 3467 4060 3479 4063
rect 3786 4060 3792 4072
rect 3467 4032 3792 4060
rect 3467 4029 3479 4032
rect 3421 4023 3479 4029
rect 3786 4020 3792 4032
rect 3844 4060 3850 4072
rect 3881 4063 3939 4069
rect 3881 4060 3893 4063
rect 3844 4032 3893 4060
rect 3844 4020 3850 4032
rect 3881 4029 3893 4032
rect 3927 4029 3939 4063
rect 3881 4023 3939 4029
rect 7190 4020 7196 4072
rect 7248 4060 7254 4072
rect 7561 4063 7619 4069
rect 7561 4060 7573 4063
rect 7248 4032 7573 4060
rect 7248 4020 7254 4032
rect 7561 4029 7573 4032
rect 7607 4029 7619 4063
rect 7561 4023 7619 4029
rect 7742 4020 7748 4072
rect 7800 4060 7806 4072
rect 8956 4060 8984 4091
rect 9950 4088 9956 4100
rect 10008 4128 10014 4140
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 10008 4100 10057 4128
rect 10008 4088 10014 4100
rect 10045 4097 10057 4100
rect 10091 4128 10103 4131
rect 10704 4128 10732 4227
rect 11514 4224 11520 4236
rect 11572 4224 11578 4276
rect 11885 4267 11943 4273
rect 11885 4233 11897 4267
rect 11931 4264 11943 4267
rect 11974 4264 11980 4276
rect 11931 4236 11980 4264
rect 11931 4233 11943 4236
rect 11885 4227 11943 4233
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 12618 4224 12624 4276
rect 12676 4264 12682 4276
rect 13909 4267 13967 4273
rect 12676 4236 13860 4264
rect 12676 4224 12682 4236
rect 11057 4199 11115 4205
rect 11057 4165 11069 4199
rect 11103 4196 11115 4199
rect 11790 4196 11796 4208
rect 11103 4168 11796 4196
rect 11103 4165 11115 4168
rect 11057 4159 11115 4165
rect 11790 4156 11796 4168
rect 11848 4156 11854 4208
rect 12526 4156 12532 4208
rect 12584 4196 12590 4208
rect 13832 4196 13860 4236
rect 13909 4233 13921 4267
rect 13955 4264 13967 4267
rect 14090 4264 14096 4276
rect 13955 4236 14096 4264
rect 13955 4233 13967 4236
rect 13909 4227 13967 4233
rect 14090 4224 14096 4236
rect 14148 4224 14154 4276
rect 15378 4264 15384 4276
rect 15339 4236 15384 4264
rect 15378 4224 15384 4236
rect 15436 4224 15442 4276
rect 16117 4267 16175 4273
rect 16117 4233 16129 4267
rect 16163 4264 16175 4267
rect 16850 4264 16856 4276
rect 16163 4236 16856 4264
rect 16163 4233 16175 4236
rect 16117 4227 16175 4233
rect 16850 4224 16856 4236
rect 16908 4224 16914 4276
rect 18046 4264 18052 4276
rect 18007 4236 18052 4264
rect 18046 4224 18052 4236
rect 18104 4224 18110 4276
rect 20898 4264 20904 4276
rect 20859 4236 20904 4264
rect 20898 4224 20904 4236
rect 20956 4224 20962 4276
rect 14001 4199 14059 4205
rect 14001 4196 14013 4199
rect 12584 4168 13768 4196
rect 13832 4168 14013 4196
rect 12584 4156 12590 4168
rect 12710 4128 12716 4140
rect 10091 4100 10732 4128
rect 12176 4100 12716 4128
rect 10091 4097 10103 4100
rect 10045 4091 10103 4097
rect 7800 4032 8984 4060
rect 7800 4020 7806 4032
rect 9214 4020 9220 4072
rect 9272 4060 9278 4072
rect 9769 4063 9827 4069
rect 9769 4060 9781 4063
rect 9272 4032 9781 4060
rect 9272 4020 9278 4032
rect 9769 4029 9781 4032
rect 9815 4060 9827 4063
rect 10686 4060 10692 4072
rect 9815 4032 10692 4060
rect 9815 4029 9827 4032
rect 9769 4023 9827 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 11238 4060 11244 4072
rect 11199 4032 11244 4060
rect 11238 4020 11244 4032
rect 11296 4020 11302 4072
rect 2133 3995 2191 4001
rect 2133 3961 2145 3995
rect 2179 3992 2191 3995
rect 2222 3992 2228 4004
rect 2179 3964 2228 3992
rect 2179 3961 2191 3964
rect 2133 3955 2191 3961
rect 2222 3952 2228 3964
rect 2280 3952 2286 4004
rect 4148 3995 4206 4001
rect 4148 3961 4160 3995
rect 4194 3992 4206 3995
rect 4338 3992 4344 4004
rect 4194 3964 4344 3992
rect 4194 3961 4206 3964
rect 4148 3955 4206 3961
rect 4338 3952 4344 3964
rect 4396 3992 4402 4004
rect 5442 3992 5448 4004
rect 4396 3964 5448 3992
rect 4396 3952 4402 3964
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 8018 3952 8024 4004
rect 8076 3992 8082 4004
rect 8205 3995 8263 4001
rect 8205 3992 8217 3995
rect 8076 3964 8217 3992
rect 8076 3952 8082 3964
rect 8205 3961 8217 3964
rect 8251 3992 8263 3995
rect 8294 3992 8300 4004
rect 8251 3964 8300 3992
rect 8251 3961 8263 3964
rect 8205 3955 8263 3961
rect 8294 3952 8300 3964
rect 8352 3952 8358 4004
rect 9306 3992 9312 4004
rect 9267 3964 9312 3992
rect 9306 3952 9312 3964
rect 9364 3992 9370 4004
rect 9861 3995 9919 4001
rect 9861 3992 9873 3995
rect 9364 3964 9873 3992
rect 9364 3952 9370 3964
rect 9861 3961 9873 3964
rect 9907 3961 9919 3995
rect 9861 3955 9919 3961
rect 11514 3952 11520 4004
rect 11572 3992 11578 4004
rect 12176 4001 12204 4100
rect 12710 4088 12716 4100
rect 12768 4128 12774 4140
rect 12897 4131 12955 4137
rect 12768 4100 12848 4128
rect 12768 4088 12774 4100
rect 12820 4069 12848 4100
rect 12897 4097 12909 4131
rect 12943 4128 12955 4131
rect 12986 4128 12992 4140
rect 12943 4100 12992 4128
rect 12943 4097 12955 4100
rect 12897 4091 12955 4097
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 13081 4131 13139 4137
rect 13081 4097 13093 4131
rect 13127 4128 13139 4131
rect 13262 4128 13268 4140
rect 13127 4100 13268 4128
rect 13127 4097 13139 4100
rect 13081 4091 13139 4097
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 13740 4128 13768 4168
rect 14001 4165 14013 4168
rect 14047 4165 14059 4199
rect 14001 4159 14059 4165
rect 15930 4156 15936 4208
rect 15988 4196 15994 4208
rect 15988 4168 16528 4196
rect 15988 4156 15994 4168
rect 13740 4100 13860 4128
rect 12805 4063 12863 4069
rect 12805 4029 12817 4063
rect 12851 4029 12863 4063
rect 13004 4060 13032 4088
rect 13449 4063 13507 4069
rect 13449 4060 13461 4063
rect 13004 4032 13461 4060
rect 12805 4023 12863 4029
rect 13449 4029 13461 4032
rect 13495 4060 13507 4063
rect 13538 4060 13544 4072
rect 13495 4032 13544 4060
rect 13495 4029 13507 4032
rect 13449 4023 13507 4029
rect 13538 4020 13544 4032
rect 13596 4020 13602 4072
rect 13832 4060 13860 4100
rect 14090 4088 14096 4140
rect 14148 4128 14154 4140
rect 14553 4131 14611 4137
rect 14553 4128 14565 4131
rect 14148 4100 14565 4128
rect 14148 4088 14154 4100
rect 14553 4097 14565 4100
rect 14599 4097 14611 4131
rect 16022 4128 16028 4140
rect 15935 4100 16028 4128
rect 14553 4091 14611 4097
rect 16022 4088 16028 4100
rect 16080 4128 16086 4140
rect 16390 4128 16396 4140
rect 16080 4100 16396 4128
rect 16080 4088 16086 4100
rect 16390 4088 16396 4100
rect 16448 4088 16454 4140
rect 16500 4128 16528 4168
rect 16942 4156 16948 4208
rect 17000 4196 17006 4208
rect 20070 4196 20076 4208
rect 17000 4168 17908 4196
rect 17000 4156 17006 4168
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 16500 4100 16681 4128
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 17880 4128 17908 4168
rect 18616 4168 20076 4196
rect 18046 4128 18052 4140
rect 17880 4100 18052 4128
rect 16669 4091 16727 4097
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 18506 4088 18512 4140
rect 18564 4128 18570 4140
rect 18616 4137 18644 4168
rect 20070 4156 20076 4168
rect 20128 4196 20134 4208
rect 20128 4168 20208 4196
rect 20128 4156 20134 4168
rect 18601 4131 18659 4137
rect 18601 4128 18613 4131
rect 18564 4100 18613 4128
rect 18564 4088 18570 4100
rect 18601 4097 18613 4100
rect 18647 4097 18659 4131
rect 19150 4128 19156 4140
rect 19111 4100 19156 4128
rect 18601 4091 18659 4097
rect 19150 4088 19156 4100
rect 19208 4088 19214 4140
rect 20180 4137 20208 4168
rect 20165 4131 20223 4137
rect 20165 4097 20177 4131
rect 20211 4097 20223 4131
rect 20165 4091 20223 4097
rect 14369 4063 14427 4069
rect 14369 4060 14381 4063
rect 13832 4032 14381 4060
rect 14369 4029 14381 4032
rect 14415 4060 14427 4063
rect 14734 4060 14740 4072
rect 14415 4032 14740 4060
rect 14415 4029 14427 4032
rect 14369 4023 14427 4029
rect 14734 4020 14740 4032
rect 14792 4020 14798 4072
rect 16482 4020 16488 4072
rect 16540 4060 16546 4072
rect 16577 4063 16635 4069
rect 16577 4060 16589 4063
rect 16540 4032 16589 4060
rect 16540 4020 16546 4032
rect 16577 4029 16589 4032
rect 16623 4029 16635 4063
rect 16577 4023 16635 4029
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 19981 4063 20039 4069
rect 19981 4060 19993 4063
rect 19484 4032 19993 4060
rect 19484 4020 19490 4032
rect 19981 4029 19993 4032
rect 20027 4029 20039 4063
rect 19981 4023 20039 4029
rect 21082 4020 21088 4072
rect 21140 4060 21146 4072
rect 21177 4063 21235 4069
rect 21177 4060 21189 4063
rect 21140 4032 21189 4060
rect 21140 4020 21146 4032
rect 21177 4029 21189 4032
rect 21223 4060 21235 4063
rect 21729 4063 21787 4069
rect 21729 4060 21741 4063
rect 21223 4032 21741 4060
rect 21223 4029 21235 4032
rect 21177 4023 21235 4029
rect 21729 4029 21741 4032
rect 21775 4029 21787 4063
rect 22278 4060 22284 4072
rect 22239 4032 22284 4060
rect 21729 4023 21787 4029
rect 22278 4020 22284 4032
rect 22336 4060 22342 4072
rect 22741 4063 22799 4069
rect 22741 4060 22753 4063
rect 22336 4032 22753 4060
rect 22336 4020 22342 4032
rect 22741 4029 22753 4032
rect 22787 4029 22799 4063
rect 22741 4023 22799 4029
rect 12161 3995 12219 4001
rect 12161 3992 12173 3995
rect 11572 3964 12173 3992
rect 11572 3952 11578 3964
rect 12161 3961 12173 3964
rect 12207 3961 12219 3995
rect 13722 3992 13728 4004
rect 12161 3955 12219 3961
rect 12452 3964 13728 3992
rect 12452 3936 12480 3964
rect 13722 3952 13728 3964
rect 13780 3952 13786 4004
rect 14461 3995 14519 4001
rect 14461 3961 14473 3995
rect 14507 3992 14519 3995
rect 14826 3992 14832 4004
rect 14507 3964 14832 3992
rect 14507 3961 14519 3964
rect 14461 3955 14519 3961
rect 14826 3952 14832 3964
rect 14884 3952 14890 4004
rect 18417 3995 18475 4001
rect 18417 3992 18429 3995
rect 17420 3964 18429 3992
rect 17420 3936 17448 3964
rect 18417 3961 18429 3964
rect 18463 3961 18475 3995
rect 18417 3955 18475 3961
rect 19334 3952 19340 4004
rect 19392 3992 19398 4004
rect 20073 3995 20131 4001
rect 19392 3964 19656 3992
rect 19392 3952 19398 3964
rect 2314 3924 2320 3936
rect 2275 3896 2320 3924
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 2682 3924 2688 3936
rect 2643 3896 2688 3924
rect 2682 3884 2688 3896
rect 2740 3884 2746 3936
rect 4614 3884 4620 3936
rect 4672 3924 4678 3936
rect 5261 3927 5319 3933
rect 5261 3924 5273 3927
rect 4672 3896 5273 3924
rect 4672 3884 4678 3896
rect 5261 3893 5273 3896
rect 5307 3893 5319 3927
rect 5261 3887 5319 3893
rect 5350 3884 5356 3936
rect 5408 3924 5414 3936
rect 6546 3924 6552 3936
rect 5408 3896 6552 3924
rect 5408 3884 5414 3896
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 7837 3927 7895 3933
rect 7837 3893 7849 3927
rect 7883 3924 7895 3927
rect 7926 3924 7932 3936
rect 7883 3896 7932 3924
rect 7883 3893 7895 3896
rect 7837 3887 7895 3893
rect 7926 3884 7932 3896
rect 7984 3884 7990 3936
rect 9398 3924 9404 3936
rect 9359 3896 9404 3924
rect 9398 3884 9404 3896
rect 9456 3884 9462 3936
rect 11422 3924 11428 3936
rect 11383 3896 11428 3924
rect 11422 3884 11428 3896
rect 11480 3884 11486 3936
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 12492 3896 12585 3924
rect 12492 3884 12498 3896
rect 12802 3884 12808 3936
rect 12860 3924 12866 3936
rect 13446 3924 13452 3936
rect 12860 3896 13452 3924
rect 12860 3884 12866 3896
rect 13446 3884 13452 3896
rect 13504 3884 13510 3936
rect 16390 3884 16396 3936
rect 16448 3924 16454 3936
rect 16485 3927 16543 3933
rect 16485 3924 16497 3927
rect 16448 3896 16497 3924
rect 16448 3884 16454 3896
rect 16485 3893 16497 3896
rect 16531 3893 16543 3927
rect 17402 3924 17408 3936
rect 17363 3896 17408 3924
rect 16485 3887 16543 3893
rect 17402 3884 17408 3896
rect 17460 3884 17466 3936
rect 17770 3924 17776 3936
rect 17731 3896 17776 3924
rect 17770 3884 17776 3896
rect 17828 3924 17834 3936
rect 18509 3927 18567 3933
rect 18509 3924 18521 3927
rect 17828 3896 18521 3924
rect 17828 3884 17834 3896
rect 18509 3893 18521 3896
rect 18555 3893 18567 3927
rect 19426 3924 19432 3936
rect 19387 3896 19432 3924
rect 18509 3887 18567 3893
rect 19426 3884 19432 3896
rect 19484 3884 19490 3936
rect 19628 3933 19656 3964
rect 20073 3961 20085 3995
rect 20119 3992 20131 3995
rect 20162 3992 20168 4004
rect 20119 3964 20168 3992
rect 20119 3961 20131 3964
rect 20073 3955 20131 3961
rect 20162 3952 20168 3964
rect 20220 3952 20226 4004
rect 22370 3992 22376 4004
rect 21376 3964 22376 3992
rect 21376 3933 21404 3964
rect 22370 3952 22376 3964
rect 22428 3952 22434 4004
rect 19613 3927 19671 3933
rect 19613 3893 19625 3927
rect 19659 3893 19671 3927
rect 19613 3887 19671 3893
rect 21361 3927 21419 3933
rect 21361 3893 21373 3927
rect 21407 3893 21419 3927
rect 22186 3924 22192 3936
rect 22147 3896 22192 3924
rect 21361 3887 21419 3893
rect 22186 3884 22192 3896
rect 22244 3884 22250 3936
rect 22462 3924 22468 3936
rect 22423 3896 22468 3924
rect 22462 3884 22468 3896
rect 22520 3884 22526 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1670 3720 1676 3732
rect 1631 3692 1676 3720
rect 1670 3680 1676 3692
rect 1728 3680 1734 3732
rect 1762 3680 1768 3732
rect 1820 3720 1826 3732
rect 2041 3723 2099 3729
rect 2041 3720 2053 3723
rect 1820 3692 2053 3720
rect 1820 3680 1826 3692
rect 2041 3689 2053 3692
rect 2087 3689 2099 3723
rect 2041 3683 2099 3689
rect 2130 3680 2136 3732
rect 2188 3720 2194 3732
rect 2685 3723 2743 3729
rect 2685 3720 2697 3723
rect 2188 3692 2697 3720
rect 2188 3680 2194 3692
rect 2685 3689 2697 3692
rect 2731 3720 2743 3723
rect 3786 3720 3792 3732
rect 2731 3692 3792 3720
rect 2731 3689 2743 3692
rect 2685 3683 2743 3689
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 5166 3720 5172 3732
rect 3936 3692 3981 3720
rect 5127 3692 5172 3720
rect 3936 3680 3942 3692
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 5994 3680 6000 3732
rect 6052 3720 6058 3732
rect 7006 3720 7012 3732
rect 6052 3692 7012 3720
rect 6052 3680 6058 3692
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 7190 3680 7196 3732
rect 7248 3720 7254 3732
rect 8389 3723 8447 3729
rect 8389 3720 8401 3723
rect 7248 3692 8401 3720
rect 7248 3680 7254 3692
rect 8389 3689 8401 3692
rect 8435 3689 8447 3723
rect 9030 3720 9036 3732
rect 8991 3692 9036 3720
rect 8389 3683 8447 3689
rect 9030 3680 9036 3692
rect 9088 3680 9094 3732
rect 9214 3680 9220 3732
rect 9272 3720 9278 3732
rect 9401 3723 9459 3729
rect 9401 3720 9413 3723
rect 9272 3692 9413 3720
rect 9272 3680 9278 3692
rect 9401 3689 9413 3692
rect 9447 3689 9459 3723
rect 9950 3720 9956 3732
rect 9911 3692 9956 3720
rect 9401 3683 9459 3689
rect 9950 3680 9956 3692
rect 10008 3680 10014 3732
rect 10597 3723 10655 3729
rect 10597 3689 10609 3723
rect 10643 3720 10655 3723
rect 10686 3720 10692 3732
rect 10643 3692 10692 3720
rect 10643 3689 10655 3692
rect 10597 3683 10655 3689
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 10962 3680 10968 3732
rect 11020 3680 11026 3732
rect 11238 3720 11244 3732
rect 11199 3692 11244 3720
rect 11238 3680 11244 3692
rect 11296 3680 11302 3732
rect 11609 3723 11667 3729
rect 11609 3689 11621 3723
rect 11655 3720 11667 3723
rect 11698 3720 11704 3732
rect 11655 3692 11704 3720
rect 11655 3689 11667 3692
rect 11609 3683 11667 3689
rect 11698 3680 11704 3692
rect 11756 3680 11762 3732
rect 14182 3720 14188 3732
rect 14143 3692 14188 3720
rect 14182 3680 14188 3692
rect 14240 3680 14246 3732
rect 15010 3720 15016 3732
rect 14971 3692 15016 3720
rect 15010 3680 15016 3692
rect 15068 3680 15074 3732
rect 15933 3723 15991 3729
rect 15933 3689 15945 3723
rect 15979 3720 15991 3723
rect 16022 3720 16028 3732
rect 15979 3692 16028 3720
rect 15979 3689 15991 3692
rect 15933 3683 15991 3689
rect 16022 3680 16028 3692
rect 16080 3720 16086 3732
rect 16298 3720 16304 3732
rect 16080 3692 16304 3720
rect 16080 3680 16086 3692
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 18049 3723 18107 3729
rect 18049 3689 18061 3723
rect 18095 3720 18107 3723
rect 18138 3720 18144 3732
rect 18095 3692 18144 3720
rect 18095 3689 18107 3692
rect 18049 3683 18107 3689
rect 18138 3680 18144 3692
rect 18196 3680 18202 3732
rect 18506 3680 18512 3732
rect 18564 3720 18570 3732
rect 18601 3723 18659 3729
rect 18601 3720 18613 3723
rect 18564 3692 18613 3720
rect 18564 3680 18570 3692
rect 18601 3689 18613 3692
rect 18647 3689 18659 3723
rect 18966 3720 18972 3732
rect 18927 3692 18972 3720
rect 18601 3683 18659 3689
rect 18966 3680 18972 3692
rect 19024 3720 19030 3732
rect 19613 3723 19671 3729
rect 19613 3720 19625 3723
rect 19024 3692 19625 3720
rect 19024 3680 19030 3692
rect 19613 3689 19625 3692
rect 19659 3689 19671 3723
rect 20162 3720 20168 3732
rect 20123 3692 20168 3720
rect 19613 3683 19671 3689
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 3513 3655 3571 3661
rect 3513 3621 3525 3655
rect 3559 3652 3571 3655
rect 3602 3652 3608 3664
rect 3559 3624 3608 3652
rect 3559 3621 3571 3624
rect 3513 3615 3571 3621
rect 3602 3612 3608 3624
rect 3660 3612 3666 3664
rect 3970 3612 3976 3664
rect 4028 3652 4034 3664
rect 4893 3655 4951 3661
rect 4893 3652 4905 3655
rect 4028 3624 4905 3652
rect 4028 3612 4034 3624
rect 4893 3621 4905 3624
rect 4939 3652 4951 3655
rect 5258 3652 5264 3664
rect 4939 3624 5264 3652
rect 4939 3621 4951 3624
rect 4893 3615 4951 3621
rect 5258 3612 5264 3624
rect 5316 3652 5322 3664
rect 5782 3655 5840 3661
rect 5782 3652 5794 3655
rect 5316 3624 5794 3652
rect 5316 3612 5322 3624
rect 5782 3621 5794 3624
rect 5828 3652 5840 3655
rect 6086 3652 6092 3664
rect 5828 3624 6092 3652
rect 5828 3621 5840 3624
rect 5782 3615 5840 3621
rect 6086 3612 6092 3624
rect 6144 3612 6150 3664
rect 6454 3612 6460 3664
rect 6512 3612 6518 3664
rect 7558 3652 7564 3664
rect 7519 3624 7564 3652
rect 7558 3612 7564 3624
rect 7616 3612 7622 3664
rect 10505 3655 10563 3661
rect 10505 3621 10517 3655
rect 10551 3652 10563 3655
rect 10980 3652 11008 3680
rect 10551 3624 11008 3652
rect 11716 3652 11744 3680
rect 11946 3655 12004 3661
rect 11946 3652 11958 3655
rect 11716 3624 11958 3652
rect 10551 3621 10563 3624
rect 10505 3615 10563 3621
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 2133 3587 2191 3593
rect 2133 3584 2145 3587
rect 1728 3556 2145 3584
rect 1728 3544 1734 3556
rect 2133 3553 2145 3556
rect 2179 3584 2191 3587
rect 2590 3584 2596 3596
rect 2179 3556 2596 3584
rect 2179 3553 2191 3556
rect 2133 3547 2191 3553
rect 2590 3544 2596 3556
rect 2648 3544 2654 3596
rect 5537 3587 5595 3593
rect 5537 3553 5549 3587
rect 5583 3584 5595 3587
rect 6472 3584 6500 3612
rect 11716 3584 11744 3624
rect 11946 3621 11958 3624
rect 11992 3621 12004 3655
rect 11946 3615 12004 3621
rect 12066 3612 12072 3664
rect 12124 3612 12130 3664
rect 14642 3652 14648 3664
rect 14603 3624 14648 3652
rect 14642 3612 14648 3624
rect 14700 3612 14706 3664
rect 12084 3584 12112 3612
rect 5583 3556 6500 3584
rect 10796 3556 11744 3584
rect 11808 3556 12112 3584
rect 15028 3584 15056 3680
rect 17310 3652 17316 3664
rect 16684 3624 17316 3652
rect 16684 3593 16712 3624
rect 17310 3612 17316 3624
rect 17368 3612 17374 3664
rect 21450 3652 21456 3664
rect 21100 3624 21456 3652
rect 16942 3593 16948 3596
rect 15289 3587 15347 3593
rect 15289 3584 15301 3587
rect 15028 3556 15301 3584
rect 5583 3553 5595 3556
rect 5537 3547 5595 3553
rect 10796 3528 10824 3556
rect 2222 3516 2228 3528
rect 2183 3488 2228 3516
rect 2222 3476 2228 3488
rect 2280 3476 2286 3528
rect 7742 3476 7748 3528
rect 7800 3516 7806 3528
rect 8478 3516 8484 3528
rect 7800 3488 8484 3516
rect 7800 3476 7806 3488
rect 8478 3476 8484 3488
rect 8536 3476 8542 3528
rect 8665 3519 8723 3525
rect 8665 3485 8677 3519
rect 8711 3516 8723 3519
rect 8754 3516 8760 3528
rect 8711 3488 8760 3516
rect 8711 3485 8723 3488
rect 8665 3479 8723 3485
rect 8754 3476 8760 3488
rect 8812 3476 8818 3528
rect 10778 3516 10784 3528
rect 10691 3488 10784 3516
rect 10778 3476 10784 3488
rect 10836 3476 10842 3528
rect 11701 3519 11759 3525
rect 11701 3485 11713 3519
rect 11747 3516 11759 3519
rect 11808 3516 11836 3556
rect 15289 3553 15301 3556
rect 15335 3553 15347 3587
rect 15289 3547 15347 3553
rect 16669 3587 16727 3593
rect 16669 3553 16681 3587
rect 16715 3553 16727 3587
rect 16936 3584 16948 3593
rect 16903 3556 16948 3584
rect 16669 3547 16727 3553
rect 16936 3547 16948 3556
rect 16942 3544 16948 3547
rect 17000 3544 17006 3596
rect 19518 3584 19524 3596
rect 19479 3556 19524 3584
rect 19518 3544 19524 3556
rect 19576 3544 19582 3596
rect 21100 3593 21128 3624
rect 21450 3612 21456 3624
rect 21508 3652 21514 3664
rect 22462 3652 22468 3664
rect 21508 3624 22468 3652
rect 21508 3612 21514 3624
rect 22462 3612 22468 3624
rect 22520 3612 22526 3664
rect 21085 3587 21143 3593
rect 21085 3553 21097 3587
rect 21131 3553 21143 3587
rect 21634 3584 21640 3596
rect 21595 3556 21640 3584
rect 21085 3547 21143 3553
rect 21634 3544 21640 3556
rect 21692 3544 21698 3596
rect 22189 3587 22247 3593
rect 22189 3553 22201 3587
rect 22235 3584 22247 3587
rect 22278 3584 22284 3596
rect 22235 3556 22284 3584
rect 22235 3553 22247 3556
rect 22189 3547 22247 3553
rect 22278 3544 22284 3556
rect 22336 3544 22342 3596
rect 19794 3516 19800 3528
rect 11747 3488 11836 3516
rect 19755 3488 19800 3516
rect 11747 3485 11759 3488
rect 11701 3479 11759 3485
rect 19794 3476 19800 3488
rect 19852 3476 19858 3528
rect 6638 3408 6644 3460
rect 6696 3448 6702 3460
rect 6917 3451 6975 3457
rect 6917 3448 6929 3451
rect 6696 3420 6929 3448
rect 6696 3408 6702 3420
rect 6917 3417 6929 3420
rect 6963 3448 6975 3451
rect 7926 3448 7932 3460
rect 6963 3420 7932 3448
rect 6963 3417 6975 3420
rect 6917 3411 6975 3417
rect 7926 3408 7932 3420
rect 7984 3408 7990 3460
rect 13630 3408 13636 3460
rect 13688 3448 13694 3460
rect 15473 3451 15531 3457
rect 13688 3420 14228 3448
rect 13688 3408 13694 3420
rect 3142 3380 3148 3392
rect 3103 3352 3148 3380
rect 3142 3340 3148 3352
rect 3200 3340 3206 3392
rect 4430 3380 4436 3392
rect 4391 3352 4436 3380
rect 4430 3340 4436 3352
rect 4488 3340 4494 3392
rect 8018 3380 8024 3392
rect 7979 3352 8024 3380
rect 8018 3340 8024 3352
rect 8076 3340 8082 3392
rect 10134 3380 10140 3392
rect 10095 3352 10140 3380
rect 10134 3340 10140 3352
rect 10192 3340 10198 3392
rect 10870 3340 10876 3392
rect 10928 3380 10934 3392
rect 11698 3380 11704 3392
rect 10928 3352 11704 3380
rect 10928 3340 10934 3352
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 13081 3383 13139 3389
rect 13081 3349 13093 3383
rect 13127 3380 13139 3383
rect 13170 3380 13176 3392
rect 13127 3352 13176 3380
rect 13127 3349 13139 3352
rect 13081 3343 13139 3349
rect 13170 3340 13176 3352
rect 13228 3380 13234 3392
rect 13722 3380 13728 3392
rect 13228 3352 13728 3380
rect 13228 3340 13234 3352
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 14090 3380 14096 3392
rect 14051 3352 14096 3380
rect 14090 3340 14096 3352
rect 14148 3340 14154 3392
rect 14200 3380 14228 3420
rect 15473 3417 15485 3451
rect 15519 3448 15531 3451
rect 16206 3448 16212 3460
rect 15519 3420 16212 3448
rect 15519 3417 15531 3420
rect 15473 3411 15531 3417
rect 16206 3408 16212 3420
rect 16264 3408 16270 3460
rect 19334 3408 19340 3460
rect 19392 3448 19398 3460
rect 20533 3451 20591 3457
rect 20533 3448 20545 3451
rect 19392 3420 20545 3448
rect 19392 3408 19398 3420
rect 20533 3417 20545 3420
rect 20579 3417 20591 3451
rect 20533 3411 20591 3417
rect 16577 3383 16635 3389
rect 16577 3380 16589 3383
rect 14200 3352 16589 3380
rect 16577 3349 16589 3352
rect 16623 3380 16635 3383
rect 17034 3380 17040 3392
rect 16623 3352 17040 3380
rect 16623 3349 16635 3352
rect 16577 3343 16635 3349
rect 17034 3340 17040 3352
rect 17092 3380 17098 3392
rect 17678 3380 17684 3392
rect 17092 3352 17684 3380
rect 17092 3340 17098 3352
rect 17678 3340 17684 3352
rect 17736 3340 17742 3392
rect 19150 3380 19156 3392
rect 19111 3352 19156 3380
rect 19150 3340 19156 3352
rect 19208 3340 19214 3392
rect 21266 3380 21272 3392
rect 21227 3352 21272 3380
rect 21266 3340 21272 3352
rect 21324 3340 21330 3392
rect 21910 3340 21916 3392
rect 21968 3380 21974 3392
rect 22373 3383 22431 3389
rect 22373 3380 22385 3383
rect 21968 3352 22385 3380
rect 21968 3340 21974 3352
rect 22373 3349 22385 3352
rect 22419 3349 22431 3383
rect 22373 3343 22431 3349
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 4893 3179 4951 3185
rect 4893 3145 4905 3179
rect 4939 3176 4951 3179
rect 5166 3176 5172 3188
rect 4939 3148 5172 3176
rect 4939 3145 4951 3148
rect 4893 3139 4951 3145
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 5997 3179 6055 3185
rect 5997 3145 6009 3179
rect 6043 3176 6055 3179
rect 6454 3176 6460 3188
rect 6043 3148 6460 3176
rect 6043 3145 6055 3148
rect 5997 3139 6055 3145
rect 6454 3136 6460 3148
rect 6512 3136 6518 3188
rect 6917 3179 6975 3185
rect 6917 3145 6929 3179
rect 6963 3176 6975 3179
rect 8202 3176 8208 3188
rect 6963 3148 8208 3176
rect 6963 3145 6975 3148
rect 6917 3139 6975 3145
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 9861 3179 9919 3185
rect 9861 3176 9873 3179
rect 9824 3148 9873 3176
rect 9824 3136 9830 3148
rect 9861 3145 9873 3148
rect 9907 3176 9919 3179
rect 10778 3176 10784 3188
rect 9907 3148 10784 3176
rect 9907 3145 9919 3148
rect 9861 3139 9919 3145
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 11885 3179 11943 3185
rect 11885 3145 11897 3179
rect 11931 3176 11943 3179
rect 12066 3176 12072 3188
rect 11931 3148 12072 3176
rect 11931 3145 11943 3148
rect 11885 3139 11943 3145
rect 12066 3136 12072 3148
rect 12124 3176 12130 3188
rect 12161 3179 12219 3185
rect 12161 3176 12173 3179
rect 12124 3148 12173 3176
rect 12124 3136 12130 3148
rect 12161 3145 12173 3148
rect 12207 3145 12219 3179
rect 12161 3139 12219 3145
rect 17129 3179 17187 3185
rect 17129 3145 17141 3179
rect 17175 3176 17187 3179
rect 17310 3176 17316 3188
rect 17175 3148 17316 3176
rect 17175 3145 17187 3148
rect 17129 3139 17187 3145
rect 3050 3068 3056 3120
rect 3108 3108 3114 3120
rect 3421 3111 3479 3117
rect 3421 3108 3433 3111
rect 3108 3080 3433 3108
rect 3108 3068 3114 3080
rect 3421 3077 3433 3080
rect 3467 3108 3479 3111
rect 4062 3108 4068 3120
rect 3467 3080 4068 3108
rect 3467 3077 3479 3080
rect 3421 3071 3479 3077
rect 4062 3068 4068 3080
rect 4120 3068 4126 3120
rect 7742 3068 7748 3120
rect 7800 3108 7806 3120
rect 8021 3111 8079 3117
rect 8021 3108 8033 3111
rect 7800 3080 8033 3108
rect 7800 3068 7806 3080
rect 8021 3077 8033 3080
rect 8067 3077 8079 3111
rect 8021 3071 8079 3077
rect 9582 3068 9588 3120
rect 9640 3108 9646 3120
rect 9950 3108 9956 3120
rect 9640 3080 9956 3108
rect 9640 3068 9646 3080
rect 9950 3068 9956 3080
rect 10008 3108 10014 3120
rect 10413 3111 10471 3117
rect 10413 3108 10425 3111
rect 10008 3080 10425 3108
rect 10008 3068 10014 3080
rect 10413 3077 10425 3080
rect 10459 3077 10471 3111
rect 10413 3071 10471 3077
rect 3142 3000 3148 3052
rect 3200 3040 3206 3052
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 3200 3012 4445 3040
rect 3200 3000 3206 3012
rect 4433 3009 4445 3012
rect 4479 3040 4491 3043
rect 4706 3040 4712 3052
rect 4479 3012 4712 3040
rect 4479 3009 4491 3012
rect 4433 3003 4491 3009
rect 4706 3000 4712 3012
rect 4764 3040 4770 3052
rect 5537 3043 5595 3049
rect 5537 3040 5549 3043
rect 4764 3012 5549 3040
rect 4764 3000 4770 3012
rect 5537 3009 5549 3012
rect 5583 3040 5595 3043
rect 6638 3040 6644 3052
rect 5583 3012 6644 3040
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 10870 3040 10876 3052
rect 7607 3012 8616 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 2041 2975 2099 2981
rect 2041 2941 2053 2975
rect 2087 2972 2099 2975
rect 2130 2972 2136 2984
rect 2087 2944 2136 2972
rect 2087 2941 2099 2944
rect 2041 2935 2099 2941
rect 2130 2932 2136 2944
rect 2188 2932 2194 2984
rect 2308 2975 2366 2981
rect 2308 2941 2320 2975
rect 2354 2972 2366 2975
rect 3160 2972 3188 3000
rect 2354 2944 3188 2972
rect 2354 2941 2366 2944
rect 2308 2935 2366 2941
rect 2222 2864 2228 2916
rect 2280 2904 2286 2916
rect 2323 2904 2351 2935
rect 4246 2932 4252 2984
rect 4304 2972 4310 2984
rect 4801 2975 4859 2981
rect 4801 2972 4813 2975
rect 4304 2944 4813 2972
rect 4304 2932 4310 2944
rect 4801 2941 4813 2944
rect 4847 2972 4859 2975
rect 5258 2972 5264 2984
rect 4847 2944 5264 2972
rect 4847 2941 4859 2944
rect 4801 2935 4859 2941
rect 5258 2932 5264 2944
rect 5316 2932 5322 2984
rect 7282 2972 7288 2984
rect 7243 2944 7288 2972
rect 7282 2932 7288 2944
rect 7340 2932 7346 2984
rect 8481 2975 8539 2981
rect 8481 2941 8493 2975
rect 8527 2941 8539 2975
rect 8588 2972 8616 3012
rect 9692 3012 10876 3040
rect 8754 2981 8760 2984
rect 8748 2972 8760 2981
rect 8588 2944 8760 2972
rect 8481 2935 8539 2941
rect 8748 2935 8760 2944
rect 8812 2972 8818 2984
rect 9582 2972 9588 2984
rect 8812 2944 9588 2972
rect 2280 2876 2351 2904
rect 2280 2864 2286 2876
rect 2774 2864 2780 2916
rect 2832 2904 2838 2916
rect 4065 2907 4123 2913
rect 4065 2904 4077 2907
rect 2832 2876 4077 2904
rect 2832 2864 2838 2876
rect 4065 2873 4077 2876
rect 4111 2904 4123 2907
rect 5353 2907 5411 2913
rect 5353 2904 5365 2907
rect 4111 2876 5365 2904
rect 4111 2873 4123 2876
rect 4065 2867 4123 2873
rect 5353 2873 5365 2876
rect 5399 2873 5411 2907
rect 5353 2867 5411 2873
rect 6641 2907 6699 2913
rect 6641 2873 6653 2907
rect 6687 2904 6699 2907
rect 7374 2904 7380 2916
rect 6687 2876 7380 2904
rect 6687 2873 6699 2876
rect 6641 2867 6699 2873
rect 7374 2864 7380 2876
rect 7432 2864 7438 2916
rect 8496 2904 8524 2935
rect 8754 2932 8760 2935
rect 8812 2932 8818 2944
rect 9582 2932 9588 2944
rect 9640 2932 9646 2984
rect 9030 2904 9036 2916
rect 8496 2876 9036 2904
rect 9030 2864 9036 2876
rect 9088 2864 9094 2916
rect 1670 2836 1676 2848
rect 1631 2808 1676 2836
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 8386 2796 8392 2848
rect 8444 2836 8450 2848
rect 9306 2836 9312 2848
rect 8444 2808 9312 2836
rect 8444 2796 8450 2808
rect 9306 2796 9312 2808
rect 9364 2836 9370 2848
rect 9692 2836 9720 3012
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 12176 3040 12204 3139
rect 17310 3136 17316 3148
rect 17368 3136 17374 3188
rect 17770 3176 17776 3188
rect 17731 3148 17776 3176
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 18046 3176 18052 3188
rect 18007 3148 18052 3176
rect 18046 3136 18052 3148
rect 18104 3136 18110 3188
rect 19058 3176 19064 3188
rect 19019 3148 19064 3176
rect 19058 3136 19064 3148
rect 19116 3136 19122 3188
rect 19334 3136 19340 3188
rect 19392 3176 19398 3188
rect 19794 3176 19800 3188
rect 19392 3148 19800 3176
rect 19392 3136 19398 3148
rect 19794 3136 19800 3148
rect 19852 3176 19858 3188
rect 20625 3179 20683 3185
rect 20625 3176 20637 3179
rect 19852 3148 20637 3176
rect 19852 3136 19858 3148
rect 20625 3145 20637 3148
rect 20671 3145 20683 3179
rect 21450 3176 21456 3188
rect 21411 3148 21456 3176
rect 20625 3139 20683 3145
rect 21450 3136 21456 3148
rect 21508 3136 21514 3188
rect 22278 3136 22284 3188
rect 22336 3176 22342 3188
rect 22557 3179 22615 3185
rect 22557 3176 22569 3179
rect 22336 3148 22569 3176
rect 22336 3136 22342 3148
rect 22557 3145 22569 3148
rect 22603 3145 22615 3179
rect 23842 3176 23848 3188
rect 23803 3148 23848 3176
rect 22557 3139 22615 3145
rect 23842 3136 23848 3148
rect 23900 3136 23906 3188
rect 13906 3068 13912 3120
rect 13964 3108 13970 3120
rect 14458 3108 14464 3120
rect 13964 3080 14464 3108
rect 13964 3068 13970 3080
rect 14458 3068 14464 3080
rect 14516 3068 14522 3120
rect 16485 3111 16543 3117
rect 16485 3077 16497 3111
rect 16531 3077 16543 3111
rect 16485 3071 16543 3077
rect 12621 3043 12679 3049
rect 12621 3040 12633 3043
rect 12176 3012 12633 3040
rect 12621 3009 12633 3012
rect 12667 3009 12679 3043
rect 16500 3040 16528 3071
rect 16666 3040 16672 3052
rect 16500 3012 16672 3040
rect 12621 3003 12679 3009
rect 11241 2975 11299 2981
rect 11241 2941 11253 2975
rect 11287 2972 11299 2975
rect 12342 2972 12348 2984
rect 11287 2944 12348 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 12342 2932 12348 2944
rect 12400 2932 12406 2984
rect 12636 2972 12664 3003
rect 16666 3000 16672 3012
rect 16724 3040 16730 3052
rect 16942 3040 16948 3052
rect 16724 3012 16948 3040
rect 16724 3000 16730 3012
rect 16942 3000 16948 3012
rect 17000 3040 17006 3052
rect 17497 3043 17555 3049
rect 17497 3040 17509 3043
rect 17000 3012 17509 3040
rect 17000 3000 17006 3012
rect 17497 3009 17509 3012
rect 17543 3040 17555 3043
rect 18601 3043 18659 3049
rect 18601 3040 18613 3043
rect 17543 3012 18613 3040
rect 17543 3009 17555 3012
rect 17497 3003 17555 3009
rect 18601 3009 18613 3012
rect 18647 3009 18659 3043
rect 19076 3040 19104 3136
rect 19518 3068 19524 3120
rect 19576 3108 19582 3120
rect 19613 3111 19671 3117
rect 19613 3108 19625 3111
rect 19576 3080 19625 3108
rect 19576 3068 19582 3080
rect 19613 3077 19625 3080
rect 19659 3108 19671 3111
rect 20993 3111 21051 3117
rect 20993 3108 21005 3111
rect 19659 3080 21005 3108
rect 19659 3077 19671 3080
rect 19613 3071 19671 3077
rect 20993 3077 21005 3080
rect 21039 3077 21051 3111
rect 20993 3071 21051 3077
rect 20165 3043 20223 3049
rect 20165 3040 20177 3043
rect 19076 3012 20177 3040
rect 18601 3003 18659 3009
rect 20165 3009 20177 3012
rect 20211 3009 20223 3043
rect 20165 3003 20223 3009
rect 14921 2975 14979 2981
rect 14921 2972 14933 2975
rect 12636 2944 14933 2972
rect 14921 2941 14933 2944
rect 14967 2972 14979 2975
rect 15105 2975 15163 2981
rect 15105 2972 15117 2975
rect 14967 2944 15117 2972
rect 14967 2941 14979 2944
rect 14921 2935 14979 2941
rect 15105 2941 15117 2944
rect 15151 2941 15163 2975
rect 15105 2935 15163 2941
rect 17770 2932 17776 2984
rect 17828 2972 17834 2984
rect 18417 2975 18475 2981
rect 18417 2972 18429 2975
rect 17828 2944 18429 2972
rect 17828 2932 17834 2944
rect 18417 2941 18429 2944
rect 18463 2972 18475 2975
rect 19426 2972 19432 2984
rect 18463 2944 19432 2972
rect 18463 2941 18475 2944
rect 18417 2935 18475 2941
rect 19426 2932 19432 2944
rect 19484 2932 19490 2984
rect 20073 2975 20131 2981
rect 20073 2941 20085 2975
rect 20119 2972 20131 2975
rect 20346 2972 20352 2984
rect 20119 2944 20352 2972
rect 20119 2941 20131 2944
rect 20073 2935 20131 2941
rect 12888 2907 12946 2913
rect 12888 2873 12900 2907
rect 12934 2904 12946 2907
rect 13722 2904 13728 2916
rect 12934 2876 13728 2904
rect 12934 2873 12946 2876
rect 12888 2867 12946 2873
rect 13722 2864 13728 2876
rect 13780 2864 13786 2916
rect 14090 2904 14096 2916
rect 14003 2876 14096 2904
rect 11422 2836 11428 2848
rect 9364 2808 9720 2836
rect 11383 2808 11428 2836
rect 9364 2796 9370 2808
rect 11422 2796 11428 2808
rect 11480 2796 11486 2848
rect 14016 2845 14044 2876
rect 14090 2864 14096 2876
rect 14148 2904 14154 2916
rect 14645 2907 14703 2913
rect 14645 2904 14657 2907
rect 14148 2876 14657 2904
rect 14148 2864 14154 2876
rect 14645 2873 14657 2876
rect 14691 2904 14703 2907
rect 15350 2907 15408 2913
rect 15350 2904 15362 2907
rect 14691 2876 15362 2904
rect 14691 2873 14703 2876
rect 14645 2867 14703 2873
rect 15350 2873 15362 2876
rect 15396 2873 15408 2907
rect 15350 2867 15408 2873
rect 18230 2864 18236 2916
rect 18288 2904 18294 2916
rect 18509 2907 18567 2913
rect 18509 2904 18521 2907
rect 18288 2876 18521 2904
rect 18288 2864 18294 2876
rect 18509 2873 18521 2876
rect 18555 2873 18567 2907
rect 18509 2867 18567 2873
rect 19518 2864 19524 2916
rect 19576 2904 19582 2916
rect 19981 2907 20039 2913
rect 19981 2904 19993 2907
rect 19576 2876 19993 2904
rect 19576 2864 19582 2876
rect 19981 2873 19993 2876
rect 20027 2873 20039 2907
rect 19981 2867 20039 2873
rect 14001 2839 14059 2845
rect 14001 2805 14013 2839
rect 14047 2805 14059 2839
rect 14001 2799 14059 2805
rect 14734 2796 14740 2848
rect 14792 2836 14798 2848
rect 15194 2836 15200 2848
rect 14792 2808 15200 2836
rect 14792 2796 14798 2808
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 19429 2839 19487 2845
rect 19429 2805 19441 2839
rect 19475 2836 19487 2839
rect 20088 2836 20116 2935
rect 20346 2932 20352 2944
rect 20404 2932 20410 2984
rect 21450 2932 21456 2984
rect 21508 2972 21514 2984
rect 21637 2975 21695 2981
rect 21637 2972 21649 2975
rect 21508 2944 21649 2972
rect 21508 2932 21514 2944
rect 21637 2941 21649 2944
rect 21683 2972 21695 2975
rect 22189 2975 22247 2981
rect 22189 2972 22201 2975
rect 21683 2944 22201 2972
rect 21683 2941 21695 2944
rect 21637 2935 21695 2941
rect 22189 2941 22201 2944
rect 22235 2941 22247 2975
rect 22189 2935 22247 2941
rect 23566 2932 23572 2984
rect 23624 2972 23630 2984
rect 23661 2975 23719 2981
rect 23661 2972 23673 2975
rect 23624 2944 23673 2972
rect 23624 2932 23630 2944
rect 23661 2941 23673 2944
rect 23707 2972 23719 2975
rect 24213 2975 24271 2981
rect 24213 2972 24225 2975
rect 23707 2944 24225 2972
rect 23707 2941 23719 2944
rect 23661 2935 23719 2941
rect 24213 2941 24225 2944
rect 24259 2941 24271 2975
rect 24213 2935 24271 2941
rect 21818 2836 21824 2848
rect 19475 2808 20116 2836
rect 21779 2808 21824 2836
rect 19475 2805 19487 2808
rect 19429 2799 19487 2805
rect 21818 2796 21824 2808
rect 21876 2796 21882 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 2409 2635 2467 2641
rect 2409 2601 2421 2635
rect 2455 2632 2467 2635
rect 2682 2632 2688 2644
rect 2455 2604 2688 2632
rect 2455 2601 2467 2604
rect 2409 2595 2467 2601
rect 2682 2592 2688 2604
rect 2740 2592 2746 2644
rect 3786 2632 3792 2644
rect 3747 2604 3792 2632
rect 3786 2592 3792 2604
rect 3844 2592 3850 2644
rect 4062 2592 4068 2644
rect 4120 2632 4126 2644
rect 6086 2632 6092 2644
rect 4120 2604 4200 2632
rect 6047 2604 6092 2632
rect 4120 2592 4126 2604
rect 1949 2567 2007 2573
rect 1949 2533 1961 2567
rect 1995 2564 2007 2567
rect 2777 2567 2835 2573
rect 2777 2564 2789 2567
rect 1995 2536 2789 2564
rect 1995 2533 2007 2536
rect 1949 2527 2007 2533
rect 2777 2533 2789 2536
rect 2823 2564 2835 2567
rect 2866 2564 2872 2576
rect 2823 2536 2872 2564
rect 2823 2533 2835 2536
rect 2777 2527 2835 2533
rect 2866 2524 2872 2536
rect 2924 2524 2930 2576
rect 3804 2496 3832 2592
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3804 2468 4077 2496
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 4172 2496 4200 2604
rect 6086 2592 6092 2604
rect 6144 2592 6150 2644
rect 7193 2635 7251 2641
rect 7193 2601 7205 2635
rect 7239 2632 7251 2635
rect 7282 2632 7288 2644
rect 7239 2604 7288 2632
rect 7239 2601 7251 2604
rect 7193 2595 7251 2601
rect 7282 2592 7288 2604
rect 7340 2592 7346 2644
rect 8113 2635 8171 2641
rect 8113 2601 8125 2635
rect 8159 2632 8171 2635
rect 8294 2632 8300 2644
rect 8159 2604 8300 2632
rect 8159 2601 8171 2604
rect 8113 2595 8171 2601
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 9582 2632 9588 2644
rect 9543 2604 9588 2632
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 9858 2592 9864 2644
rect 9916 2632 9922 2644
rect 10137 2635 10195 2641
rect 10137 2632 10149 2635
rect 9916 2604 10149 2632
rect 9916 2592 9922 2604
rect 10137 2601 10149 2604
rect 10183 2601 10195 2635
rect 10778 2632 10784 2644
rect 10739 2604 10784 2632
rect 10137 2595 10195 2601
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 11330 2632 11336 2644
rect 11291 2604 11336 2632
rect 11330 2592 11336 2604
rect 11388 2592 11394 2644
rect 12158 2592 12164 2644
rect 12216 2632 12222 2644
rect 12621 2635 12679 2641
rect 12621 2632 12633 2635
rect 12216 2604 12633 2632
rect 12216 2592 12222 2604
rect 12621 2601 12633 2604
rect 12667 2601 12679 2635
rect 12986 2632 12992 2644
rect 12947 2604 12992 2632
rect 12621 2595 12679 2601
rect 12986 2592 12992 2604
rect 13044 2592 13050 2644
rect 13081 2635 13139 2641
rect 13081 2601 13093 2635
rect 13127 2632 13139 2635
rect 13630 2632 13636 2644
rect 13127 2604 13636 2632
rect 13127 2601 13139 2604
rect 13081 2595 13139 2601
rect 6914 2524 6920 2576
rect 6972 2564 6978 2576
rect 7653 2567 7711 2573
rect 7653 2564 7665 2567
rect 6972 2536 7665 2564
rect 6972 2524 6978 2536
rect 7653 2533 7665 2536
rect 7699 2564 7711 2567
rect 8570 2564 8576 2576
rect 7699 2536 8576 2564
rect 7699 2533 7711 2536
rect 7653 2527 7711 2533
rect 8570 2524 8576 2536
rect 8628 2524 8634 2576
rect 9674 2524 9680 2576
rect 9732 2564 9738 2576
rect 10229 2567 10287 2573
rect 10229 2564 10241 2567
rect 9732 2536 10241 2564
rect 9732 2524 9738 2536
rect 10229 2533 10241 2536
rect 10275 2564 10287 2567
rect 10962 2564 10968 2576
rect 10275 2536 10968 2564
rect 10275 2533 10287 2536
rect 10229 2527 10287 2533
rect 10962 2524 10968 2536
rect 11020 2524 11026 2576
rect 4332 2499 4390 2505
rect 4332 2496 4344 2499
rect 4172 2468 4344 2496
rect 4065 2459 4123 2465
rect 4332 2465 4344 2468
rect 4378 2496 4390 2499
rect 6454 2496 6460 2508
rect 4378 2468 6460 2496
rect 4378 2465 4390 2468
rect 4332 2459 4390 2465
rect 6454 2456 6460 2468
rect 6512 2456 6518 2508
rect 8110 2456 8116 2508
rect 8168 2496 8174 2508
rect 8481 2499 8539 2505
rect 8481 2496 8493 2499
rect 8168 2468 8493 2496
rect 8168 2456 8174 2468
rect 8481 2465 8493 2468
rect 8527 2496 8539 2499
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8527 2468 9137 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 9125 2465 9137 2468
rect 9171 2496 9183 2499
rect 9490 2496 9496 2508
rect 9171 2468 9496 2496
rect 9171 2465 9183 2468
rect 9125 2459 9183 2465
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 11348 2496 11376 2592
rect 12437 2567 12495 2573
rect 12437 2533 12449 2567
rect 12483 2564 12495 2567
rect 13004 2564 13032 2592
rect 12483 2536 13032 2564
rect 12483 2533 12495 2536
rect 12437 2527 12495 2533
rect 11425 2499 11483 2505
rect 11425 2496 11437 2499
rect 11348 2468 11437 2496
rect 11425 2465 11437 2468
rect 11471 2465 11483 2499
rect 11425 2459 11483 2465
rect 1394 2428 1400 2440
rect 1355 2400 1400 2428
rect 1394 2388 1400 2400
rect 1452 2388 1458 2440
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 2317 2431 2375 2437
rect 2317 2428 2329 2431
rect 2004 2400 2329 2428
rect 2004 2388 2010 2400
rect 2317 2397 2329 2400
rect 2363 2428 2375 2431
rect 2869 2431 2927 2437
rect 2869 2428 2881 2431
rect 2363 2400 2881 2428
rect 2363 2397 2375 2400
rect 2317 2391 2375 2397
rect 2869 2397 2881 2400
rect 2915 2428 2927 2431
rect 2958 2428 2964 2440
rect 2915 2400 2964 2428
rect 2915 2397 2927 2400
rect 2869 2391 2927 2397
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 3513 2431 3571 2437
rect 3513 2428 3525 2431
rect 3099 2400 3525 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 3513 2397 3525 2400
rect 3559 2428 3571 2431
rect 3970 2428 3976 2440
rect 3559 2400 3976 2428
rect 3559 2397 3571 2400
rect 3513 2391 3571 2397
rect 3970 2388 3976 2400
rect 4028 2388 4034 2440
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 7248 2400 7941 2428
rect 7248 2388 7254 2400
rect 7929 2397 7941 2400
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2428 8815 2431
rect 9582 2428 9588 2440
rect 8803 2400 9588 2428
rect 8803 2397 8815 2400
rect 8757 2391 8815 2397
rect 9582 2388 9588 2400
rect 9640 2388 9646 2440
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2428 10471 2431
rect 10778 2428 10784 2440
rect 10459 2400 10784 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 10778 2388 10784 2400
rect 10836 2388 10842 2440
rect 11974 2428 11980 2440
rect 11935 2400 11980 2428
rect 11974 2388 11980 2400
rect 12032 2428 12038 2440
rect 13096 2428 13124 2595
rect 13630 2592 13636 2604
rect 13688 2592 13694 2644
rect 13998 2592 14004 2644
rect 14056 2632 14062 2644
rect 14185 2635 14243 2641
rect 14185 2632 14197 2635
rect 14056 2604 14197 2632
rect 14056 2592 14062 2604
rect 14185 2601 14197 2604
rect 14231 2632 14243 2635
rect 14734 2632 14740 2644
rect 14231 2604 14740 2632
rect 14231 2601 14243 2604
rect 14185 2595 14243 2601
rect 14292 2505 14320 2604
rect 14734 2592 14740 2604
rect 14792 2592 14798 2644
rect 15473 2635 15531 2641
rect 15473 2601 15485 2635
rect 15519 2632 15531 2635
rect 16390 2632 16396 2644
rect 15519 2604 16396 2632
rect 15519 2601 15531 2604
rect 15473 2595 15531 2601
rect 16390 2592 16396 2604
rect 16448 2592 16454 2644
rect 16666 2632 16672 2644
rect 16627 2604 16672 2632
rect 16666 2592 16672 2604
rect 16724 2592 16730 2644
rect 18138 2632 18144 2644
rect 18099 2604 18144 2632
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 18690 2632 18696 2644
rect 18651 2604 18696 2632
rect 18690 2592 18696 2604
rect 18748 2592 18754 2644
rect 18785 2635 18843 2641
rect 18785 2601 18797 2635
rect 18831 2632 18843 2635
rect 19242 2632 19248 2644
rect 18831 2604 19248 2632
rect 18831 2601 18843 2604
rect 18785 2595 18843 2601
rect 19242 2592 19248 2604
rect 19300 2592 19306 2644
rect 19334 2564 19340 2576
rect 14660 2536 19340 2564
rect 14277 2499 14335 2505
rect 14277 2465 14289 2499
rect 14323 2465 14335 2499
rect 14277 2459 14335 2465
rect 13262 2428 13268 2440
rect 12032 2400 13124 2428
rect 13223 2400 13268 2428
rect 12032 2388 12038 2400
rect 13262 2388 13268 2400
rect 13320 2428 13326 2440
rect 13633 2431 13691 2437
rect 13633 2428 13645 2431
rect 13320 2400 13645 2428
rect 13320 2388 13326 2400
rect 13633 2397 13645 2400
rect 13679 2397 13691 2431
rect 13633 2391 13691 2397
rect 9769 2363 9827 2369
rect 9769 2329 9781 2363
rect 9815 2360 9827 2363
rect 11146 2360 11152 2372
rect 9815 2332 11152 2360
rect 9815 2329 9827 2332
rect 9769 2323 9827 2329
rect 11146 2320 11152 2332
rect 11204 2320 11210 2372
rect 13170 2320 13176 2372
rect 13228 2360 13234 2372
rect 14660 2360 14688 2536
rect 19334 2524 19340 2536
rect 19392 2524 19398 2576
rect 14734 2456 14740 2508
rect 14792 2496 14798 2508
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 14792 2468 14841 2496
rect 14792 2456 14798 2468
rect 14829 2465 14841 2468
rect 14875 2496 14887 2499
rect 15841 2499 15899 2505
rect 15841 2496 15853 2499
rect 14875 2468 15853 2496
rect 14875 2465 14887 2468
rect 14829 2459 14887 2465
rect 15841 2465 15853 2468
rect 15887 2465 15899 2499
rect 17126 2496 17132 2508
rect 17087 2468 17132 2496
rect 15841 2459 15899 2465
rect 17126 2456 17132 2468
rect 17184 2496 17190 2508
rect 17681 2499 17739 2505
rect 17681 2496 17693 2499
rect 17184 2468 17693 2496
rect 17184 2456 17190 2468
rect 17681 2465 17693 2468
rect 17727 2465 17739 2499
rect 17681 2459 17739 2465
rect 19426 2456 19432 2508
rect 19484 2496 19490 2508
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 19484 2468 19901 2496
rect 19484 2456 19490 2468
rect 19889 2465 19901 2468
rect 19935 2496 19947 2499
rect 20441 2499 20499 2505
rect 20441 2496 20453 2499
rect 19935 2468 20453 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 20441 2465 20453 2468
rect 20487 2465 20499 2499
rect 21542 2496 21548 2508
rect 21503 2468 21548 2496
rect 20441 2459 20499 2465
rect 21542 2456 21548 2468
rect 21600 2456 21606 2508
rect 22738 2496 22744 2508
rect 21652 2468 21864 2496
rect 22699 2468 22744 2496
rect 21652 2440 21680 2468
rect 15933 2431 15991 2437
rect 15933 2397 15945 2431
rect 15979 2397 15991 2431
rect 15933 2391 15991 2397
rect 16117 2431 16175 2437
rect 16117 2397 16129 2431
rect 16163 2428 16175 2431
rect 16298 2428 16304 2440
rect 16163 2400 16304 2428
rect 16163 2397 16175 2400
rect 16117 2391 16175 2397
rect 13228 2332 14688 2360
rect 13228 2320 13234 2332
rect 5442 2292 5448 2304
rect 5403 2264 5448 2292
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 6454 2292 6460 2304
rect 6415 2264 6460 2292
rect 6454 2252 6460 2264
rect 6512 2252 6518 2304
rect 11606 2292 11612 2304
rect 11567 2264 11612 2292
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 14458 2292 14464 2304
rect 14419 2264 14464 2292
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 15286 2292 15292 2304
rect 15247 2264 15292 2292
rect 15286 2252 15292 2264
rect 15344 2292 15350 2304
rect 15948 2292 15976 2391
rect 16298 2388 16304 2400
rect 16356 2388 16362 2440
rect 18877 2431 18935 2437
rect 18877 2428 18889 2431
rect 16960 2400 18889 2428
rect 16960 2304 16988 2400
rect 18877 2397 18889 2400
rect 18923 2397 18935 2431
rect 21634 2428 21640 2440
rect 21595 2400 21640 2428
rect 18877 2391 18935 2397
rect 21634 2388 21640 2400
rect 21692 2388 21698 2440
rect 21729 2431 21787 2437
rect 21729 2397 21741 2431
rect 21775 2397 21787 2431
rect 21729 2391 21787 2397
rect 17218 2320 17224 2372
rect 17276 2360 17282 2372
rect 18325 2363 18383 2369
rect 18325 2360 18337 2363
rect 17276 2332 18337 2360
rect 17276 2320 17282 2332
rect 18325 2329 18337 2332
rect 18371 2329 18383 2363
rect 21744 2360 21772 2391
rect 18325 2323 18383 2329
rect 20916 2332 21772 2360
rect 21836 2360 21864 2468
rect 22738 2456 22744 2468
rect 22796 2496 22802 2508
rect 23293 2499 23351 2505
rect 23293 2496 23305 2499
rect 22796 2468 23305 2496
rect 22796 2456 22802 2468
rect 23293 2465 23305 2468
rect 23339 2465 23351 2499
rect 23293 2459 23351 2465
rect 23474 2456 23480 2508
rect 23532 2496 23538 2508
rect 23661 2499 23719 2505
rect 23661 2496 23673 2499
rect 23532 2468 23673 2496
rect 23532 2456 23538 2468
rect 23661 2465 23673 2468
rect 23707 2465 23719 2499
rect 24026 2496 24032 2508
rect 23987 2468 24032 2496
rect 23661 2459 23719 2465
rect 24026 2456 24032 2468
rect 24084 2496 24090 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 24084 2468 24593 2496
rect 24084 2456 24090 2468
rect 24581 2465 24593 2468
rect 24627 2465 24639 2499
rect 24581 2459 24639 2465
rect 22189 2363 22247 2369
rect 22189 2360 22201 2363
rect 21836 2332 22201 2360
rect 20916 2304 20944 2332
rect 22189 2329 22201 2332
rect 22235 2329 22247 2363
rect 22189 2323 22247 2329
rect 22925 2363 22983 2369
rect 22925 2329 22937 2363
rect 22971 2360 22983 2363
rect 24118 2360 24124 2372
rect 22971 2332 24124 2360
rect 22971 2329 22983 2332
rect 22925 2323 22983 2329
rect 24118 2320 24124 2332
rect 24176 2320 24182 2372
rect 16942 2292 16948 2304
rect 15344 2264 15976 2292
rect 16903 2264 16948 2292
rect 15344 2252 15350 2264
rect 16942 2252 16948 2264
rect 17000 2252 17006 2304
rect 17310 2292 17316 2304
rect 17271 2264 17316 2292
rect 17310 2252 17316 2264
rect 17368 2252 17374 2304
rect 19518 2252 19524 2304
rect 19576 2292 19582 2304
rect 19613 2295 19671 2301
rect 19613 2292 19625 2295
rect 19576 2264 19625 2292
rect 19576 2252 19582 2264
rect 19613 2261 19625 2264
rect 19659 2261 19671 2295
rect 20070 2292 20076 2304
rect 20031 2264 20076 2292
rect 19613 2255 19671 2261
rect 20070 2252 20076 2264
rect 20128 2252 20134 2304
rect 20898 2292 20904 2304
rect 20859 2264 20904 2292
rect 20898 2252 20904 2264
rect 20956 2252 20962 2304
rect 21174 2292 21180 2304
rect 21135 2264 21180 2292
rect 21174 2252 21180 2264
rect 21232 2252 21238 2304
rect 21542 2252 21548 2304
rect 21600 2292 21606 2304
rect 22557 2295 22615 2301
rect 22557 2292 22569 2295
rect 21600 2264 22569 2292
rect 21600 2252 21606 2264
rect 22557 2261 22569 2264
rect 22603 2261 22615 2295
rect 24210 2292 24216 2304
rect 24171 2264 24216 2292
rect 22557 2255 22615 2261
rect 24210 2252 24216 2264
rect 24268 2252 24274 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 1394 1708 1400 1760
rect 1452 1748 1458 1760
rect 3510 1748 3516 1760
rect 1452 1720 3516 1748
rect 1452 1708 1458 1720
rect 3510 1708 3516 1720
rect 3568 1748 3574 1760
rect 7190 1748 7196 1760
rect 3568 1720 7196 1748
rect 3568 1708 3574 1720
rect 7190 1708 7196 1720
rect 7248 1708 7254 1760
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 1860 25304 1912 25356
rect 2412 25304 2464 25356
rect 5356 25304 5408 25356
rect 2964 25168 3016 25220
rect 2228 25143 2280 25152
rect 2228 25109 2237 25143
rect 2237 25109 2271 25143
rect 2271 25109 2280 25143
rect 2228 25100 2280 25109
rect 2872 25100 2924 25152
rect 3240 25100 3292 25152
rect 4896 25100 4948 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 2412 24939 2464 24948
rect 2412 24905 2421 24939
rect 2421 24905 2455 24939
rect 2455 24905 2464 24939
rect 2412 24896 2464 24905
rect 4068 24828 4120 24880
rect 6092 24828 6144 24880
rect 2044 24803 2096 24812
rect 2044 24769 2053 24803
rect 2053 24769 2087 24803
rect 2087 24769 2096 24803
rect 2044 24760 2096 24769
rect 4896 24760 4948 24812
rect 2780 24692 2832 24744
rect 4344 24692 4396 24744
rect 7104 24692 7156 24744
rect 16028 24735 16080 24744
rect 16028 24701 16037 24735
rect 16037 24701 16071 24735
rect 16071 24701 16080 24735
rect 16028 24692 16080 24701
rect 5080 24624 5132 24676
rect 1584 24599 1636 24608
rect 1584 24565 1593 24599
rect 1593 24565 1627 24599
rect 1627 24565 1636 24599
rect 1584 24556 1636 24565
rect 2596 24599 2648 24608
rect 2596 24565 2605 24599
rect 2605 24565 2639 24599
rect 2639 24565 2648 24599
rect 2596 24556 2648 24565
rect 3240 24556 3292 24608
rect 4160 24599 4212 24608
rect 4160 24565 4169 24599
rect 4169 24565 4203 24599
rect 4203 24565 4212 24599
rect 4160 24556 4212 24565
rect 7196 24599 7248 24608
rect 7196 24565 7205 24599
rect 7205 24565 7239 24599
rect 7239 24565 7248 24599
rect 7196 24556 7248 24565
rect 7380 24556 7432 24608
rect 7840 24599 7892 24608
rect 7840 24565 7849 24599
rect 7849 24565 7883 24599
rect 7883 24565 7892 24599
rect 7840 24556 7892 24565
rect 16212 24599 16264 24608
rect 16212 24565 16221 24599
rect 16221 24565 16255 24599
rect 16255 24565 16264 24599
rect 16212 24556 16264 24565
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 1860 24395 1912 24404
rect 1860 24361 1869 24395
rect 1869 24361 1903 24395
rect 1903 24361 1912 24395
rect 1860 24352 1912 24361
rect 2228 24352 2280 24404
rect 2780 24352 2832 24404
rect 3516 24352 3568 24404
rect 4804 24352 4856 24404
rect 6184 24352 6236 24404
rect 10784 24395 10836 24404
rect 10784 24361 10793 24395
rect 10793 24361 10827 24395
rect 10827 24361 10836 24395
rect 10784 24352 10836 24361
rect 14280 24395 14332 24404
rect 14280 24361 14289 24395
rect 14289 24361 14323 24395
rect 14323 24361 14332 24395
rect 14280 24352 14332 24361
rect 16488 24352 16540 24404
rect 18512 24352 18564 24404
rect 18972 24395 19024 24404
rect 18972 24361 18981 24395
rect 18981 24361 19015 24395
rect 19015 24361 19024 24395
rect 18972 24352 19024 24361
rect 22468 24352 22520 24404
rect 3056 24284 3108 24336
rect 4252 24284 4304 24336
rect 4712 24284 4764 24336
rect 6000 24284 6052 24336
rect 2044 24216 2096 24268
rect 3700 24216 3752 24268
rect 6920 24216 6972 24268
rect 7840 24259 7892 24268
rect 7840 24225 7849 24259
rect 7849 24225 7883 24259
rect 7883 24225 7892 24259
rect 7840 24216 7892 24225
rect 10600 24259 10652 24268
rect 10600 24225 10609 24259
rect 10609 24225 10643 24259
rect 10643 24225 10652 24259
rect 10600 24216 10652 24225
rect 11980 24216 12032 24268
rect 14096 24259 14148 24268
rect 14096 24225 14105 24259
rect 14105 24225 14139 24259
rect 14139 24225 14148 24259
rect 14096 24216 14148 24225
rect 15476 24216 15528 24268
rect 16764 24216 16816 24268
rect 17684 24216 17736 24268
rect 19064 24216 19116 24268
rect 20812 24216 20864 24268
rect 4252 24148 4304 24200
rect 3332 24080 3384 24132
rect 4896 24148 4948 24200
rect 7196 24148 7248 24200
rect 8116 24191 8168 24200
rect 7380 24080 7432 24132
rect 8116 24157 8125 24191
rect 8125 24157 8159 24191
rect 8159 24157 8168 24191
rect 8116 24148 8168 24157
rect 12256 24123 12308 24132
rect 12256 24089 12265 24123
rect 12265 24089 12299 24123
rect 12299 24089 12308 24123
rect 12256 24080 12308 24089
rect 17776 24123 17828 24132
rect 17776 24089 17785 24123
rect 17785 24089 17819 24123
rect 17819 24089 17828 24123
rect 17776 24080 17828 24089
rect 2504 24012 2556 24064
rect 4988 24012 5040 24064
rect 5448 24012 5500 24064
rect 7104 24055 7156 24064
rect 7104 24021 7113 24055
rect 7113 24021 7147 24055
rect 7147 24021 7156 24055
rect 7104 24012 7156 24021
rect 7472 24055 7524 24064
rect 7472 24021 7481 24055
rect 7481 24021 7515 24055
rect 7515 24021 7524 24055
rect 7472 24012 7524 24021
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2044 23851 2096 23860
rect 2044 23817 2053 23851
rect 2053 23817 2087 23851
rect 2087 23817 2096 23851
rect 2044 23808 2096 23817
rect 3056 23808 3108 23860
rect 3700 23851 3752 23860
rect 1676 23740 1728 23792
rect 2504 23740 2556 23792
rect 3700 23817 3709 23851
rect 3709 23817 3743 23851
rect 3743 23817 3752 23851
rect 3700 23808 3752 23817
rect 4896 23808 4948 23860
rect 6184 23851 6236 23860
rect 6184 23817 6193 23851
rect 6193 23817 6227 23851
rect 6227 23817 6236 23851
rect 6184 23808 6236 23817
rect 2596 23715 2648 23724
rect 2596 23681 2605 23715
rect 2605 23681 2639 23715
rect 2639 23681 2648 23715
rect 2596 23672 2648 23681
rect 3792 23740 3844 23792
rect 4252 23740 4304 23792
rect 6000 23740 6052 23792
rect 6736 23740 6788 23792
rect 2228 23604 2280 23656
rect 4252 23647 4304 23656
rect 4252 23613 4261 23647
rect 4261 23613 4295 23647
rect 4295 23613 4304 23647
rect 4252 23604 4304 23613
rect 6276 23604 6328 23656
rect 7104 23647 7156 23656
rect 7104 23613 7113 23647
rect 7113 23613 7147 23647
rect 7147 23613 7156 23647
rect 7104 23604 7156 23613
rect 9864 23604 9916 23656
rect 10600 23647 10652 23656
rect 10600 23613 10609 23647
rect 10609 23613 10643 23647
rect 10643 23613 10652 23647
rect 10600 23604 10652 23613
rect 11336 23604 11388 23656
rect 13360 23808 13412 23860
rect 14096 23808 14148 23860
rect 15660 23808 15712 23860
rect 18328 23851 18380 23860
rect 18328 23817 18337 23851
rect 18337 23817 18371 23851
rect 18371 23817 18380 23851
rect 18328 23808 18380 23817
rect 19524 23851 19576 23860
rect 19524 23817 19533 23851
rect 19533 23817 19567 23851
rect 19567 23817 19576 23851
rect 19524 23808 19576 23817
rect 21272 23851 21324 23860
rect 21272 23817 21281 23851
rect 21281 23817 21315 23851
rect 21315 23817 21324 23851
rect 21272 23808 21324 23817
rect 25320 23808 25372 23860
rect 15200 23783 15252 23792
rect 15200 23749 15209 23783
rect 15209 23749 15243 23783
rect 15243 23749 15252 23783
rect 15200 23740 15252 23749
rect 19708 23740 19760 23792
rect 3332 23536 3384 23588
rect 4804 23536 4856 23588
rect 7196 23536 7248 23588
rect 7748 23536 7800 23588
rect 1400 23468 1452 23520
rect 1584 23468 1636 23520
rect 2136 23511 2188 23520
rect 2136 23477 2145 23511
rect 2145 23477 2179 23511
rect 2179 23477 2188 23511
rect 2136 23468 2188 23477
rect 6644 23468 6696 23520
rect 8116 23468 8168 23520
rect 11428 23511 11480 23520
rect 11428 23477 11437 23511
rect 11437 23477 11471 23511
rect 11471 23477 11480 23511
rect 11428 23468 11480 23477
rect 11980 23468 12032 23520
rect 12624 23511 12676 23520
rect 12624 23477 12633 23511
rect 12633 23477 12667 23511
rect 12667 23477 12676 23511
rect 12624 23468 12676 23477
rect 13820 23468 13872 23520
rect 14648 23468 14700 23520
rect 16580 23604 16632 23656
rect 19340 23647 19392 23656
rect 19340 23613 19349 23647
rect 19349 23613 19383 23647
rect 19383 23613 19392 23647
rect 19340 23604 19392 23613
rect 21088 23647 21140 23656
rect 21088 23613 21097 23647
rect 21097 23613 21131 23647
rect 21131 23613 21140 23647
rect 21088 23604 21140 23613
rect 23480 23604 23532 23656
rect 15476 23468 15528 23520
rect 16764 23468 16816 23520
rect 17684 23511 17736 23520
rect 17684 23477 17693 23511
rect 17693 23477 17727 23511
rect 17727 23477 17736 23511
rect 17684 23468 17736 23477
rect 18696 23511 18748 23520
rect 18696 23477 18705 23511
rect 18705 23477 18739 23511
rect 18739 23477 18748 23511
rect 18696 23468 18748 23477
rect 19064 23511 19116 23520
rect 19064 23477 19073 23511
rect 19073 23477 19107 23511
rect 19107 23477 19116 23511
rect 19064 23468 19116 23477
rect 20812 23468 20864 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 2780 23264 2832 23316
rect 7196 23264 7248 23316
rect 9864 23307 9916 23316
rect 9864 23273 9873 23307
rect 9873 23273 9907 23307
rect 9907 23273 9916 23307
rect 9864 23264 9916 23273
rect 14096 23264 14148 23316
rect 17224 23307 17276 23316
rect 17224 23273 17233 23307
rect 17233 23273 17267 23307
rect 17267 23273 17276 23307
rect 17224 23264 17276 23273
rect 19064 23264 19116 23316
rect 21088 23307 21140 23316
rect 21088 23273 21097 23307
rect 21097 23273 21131 23307
rect 21131 23273 21140 23307
rect 21088 23264 21140 23273
rect 23480 23264 23532 23316
rect 3332 23196 3384 23248
rect 5172 23196 5224 23248
rect 6644 23196 6696 23248
rect 2136 23171 2188 23180
rect 2136 23137 2145 23171
rect 2145 23137 2179 23171
rect 2179 23137 2188 23171
rect 2136 23128 2188 23137
rect 4252 23128 4304 23180
rect 9680 23171 9732 23180
rect 9680 23137 9689 23171
rect 9689 23137 9723 23171
rect 9723 23137 9732 23171
rect 9680 23128 9732 23137
rect 13084 23128 13136 23180
rect 14280 23128 14332 23180
rect 15292 23171 15344 23180
rect 15292 23137 15301 23171
rect 15301 23137 15335 23171
rect 15335 23137 15344 23171
rect 15292 23128 15344 23137
rect 17040 23171 17092 23180
rect 17040 23137 17049 23171
rect 17049 23137 17083 23171
rect 17083 23137 17092 23171
rect 17040 23128 17092 23137
rect 18144 23171 18196 23180
rect 18144 23137 18153 23171
rect 18153 23137 18187 23171
rect 18187 23137 18196 23171
rect 18144 23128 18196 23137
rect 20904 23171 20956 23180
rect 20904 23137 20913 23171
rect 20913 23137 20947 23171
rect 20947 23137 20956 23171
rect 20904 23128 20956 23137
rect 22376 23171 22428 23180
rect 22376 23137 22385 23171
rect 22385 23137 22419 23171
rect 22419 23137 22428 23171
rect 22376 23128 22428 23137
rect 2228 23103 2280 23112
rect 2228 23069 2237 23103
rect 2237 23069 2271 23103
rect 2271 23069 2280 23103
rect 2228 23060 2280 23069
rect 2688 23060 2740 23112
rect 3976 23060 4028 23112
rect 5264 23060 5316 23112
rect 6276 23103 6328 23112
rect 4804 22992 4856 23044
rect 6276 23069 6285 23103
rect 6285 23069 6319 23103
rect 6319 23069 6328 23103
rect 6276 23060 6328 23069
rect 12900 23035 12952 23044
rect 1768 22967 1820 22976
rect 1768 22933 1777 22967
rect 1777 22933 1811 22967
rect 1811 22933 1820 22967
rect 1768 22924 1820 22933
rect 4436 22924 4488 22976
rect 12900 23001 12909 23035
rect 12909 23001 12943 23035
rect 12943 23001 12952 23035
rect 12900 22992 12952 23001
rect 8484 22967 8536 22976
rect 8484 22933 8493 22967
rect 8493 22933 8527 22967
rect 8527 22933 8536 22967
rect 8484 22924 8536 22933
rect 13636 22967 13688 22976
rect 13636 22933 13645 22967
rect 13645 22933 13679 22967
rect 13679 22933 13688 22967
rect 13636 22924 13688 22933
rect 14280 22967 14332 22976
rect 14280 22933 14289 22967
rect 14289 22933 14323 22967
rect 14323 22933 14332 22967
rect 14280 22924 14332 22933
rect 15568 22924 15620 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 2044 22763 2096 22772
rect 2044 22729 2053 22763
rect 2053 22729 2087 22763
rect 2087 22729 2096 22763
rect 2044 22720 2096 22729
rect 2596 22584 2648 22636
rect 4252 22720 4304 22772
rect 4804 22763 4856 22772
rect 4804 22729 4813 22763
rect 4813 22729 4847 22763
rect 4847 22729 4856 22763
rect 4804 22720 4856 22729
rect 6092 22720 6144 22772
rect 6368 22720 6420 22772
rect 15660 22763 15712 22772
rect 5632 22627 5684 22636
rect 5632 22593 5641 22627
rect 5641 22593 5675 22627
rect 5675 22593 5684 22627
rect 5632 22584 5684 22593
rect 6000 22584 6052 22636
rect 6644 22584 6696 22636
rect 15660 22729 15669 22763
rect 15669 22729 15703 22763
rect 15703 22729 15712 22763
rect 15660 22720 15712 22729
rect 16764 22763 16816 22772
rect 16764 22729 16773 22763
rect 16773 22729 16807 22763
rect 16807 22729 16816 22763
rect 16764 22720 16816 22729
rect 20904 22763 20956 22772
rect 20904 22729 20913 22763
rect 20913 22729 20947 22763
rect 20947 22729 20956 22763
rect 20904 22720 20956 22729
rect 8392 22695 8444 22704
rect 8392 22661 8401 22695
rect 8401 22661 8435 22695
rect 8435 22661 8444 22695
rect 8392 22652 8444 22661
rect 7748 22584 7800 22636
rect 2044 22516 2096 22568
rect 3332 22516 3384 22568
rect 5540 22559 5592 22568
rect 5540 22525 5549 22559
rect 5549 22525 5583 22559
rect 5583 22525 5592 22559
rect 5540 22516 5592 22525
rect 6092 22516 6144 22568
rect 8484 22516 8536 22568
rect 13360 22491 13412 22500
rect 13360 22457 13369 22491
rect 13369 22457 13403 22491
rect 13403 22457 13412 22491
rect 13360 22448 13412 22457
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 4068 22423 4120 22432
rect 4068 22389 4077 22423
rect 4077 22389 4111 22423
rect 4111 22389 4120 22423
rect 4068 22380 4120 22389
rect 5172 22423 5224 22432
rect 5172 22389 5181 22423
rect 5181 22389 5215 22423
rect 5215 22389 5224 22423
rect 5172 22380 5224 22389
rect 8208 22423 8260 22432
rect 8208 22389 8217 22423
rect 8217 22389 8251 22423
rect 8251 22389 8260 22423
rect 8208 22380 8260 22389
rect 9312 22380 9364 22432
rect 9680 22423 9732 22432
rect 9680 22389 9689 22423
rect 9689 22389 9723 22423
rect 9723 22389 9732 22423
rect 9680 22380 9732 22389
rect 10968 22380 11020 22432
rect 13084 22380 13136 22432
rect 13544 22423 13596 22432
rect 13544 22389 13553 22423
rect 13553 22389 13587 22423
rect 13587 22389 13596 22423
rect 13544 22380 13596 22389
rect 13636 22380 13688 22432
rect 15200 22516 15252 22568
rect 15292 22448 15344 22500
rect 15752 22448 15804 22500
rect 15108 22380 15160 22432
rect 17040 22423 17092 22432
rect 17040 22389 17049 22423
rect 17049 22389 17083 22423
rect 17083 22389 17092 22423
rect 17040 22380 17092 22389
rect 17500 22423 17552 22432
rect 17500 22389 17509 22423
rect 17509 22389 17543 22423
rect 17543 22389 17552 22423
rect 17500 22380 17552 22389
rect 18144 22380 18196 22432
rect 22376 22423 22428 22432
rect 22376 22389 22385 22423
rect 22385 22389 22419 22423
rect 22419 22389 22428 22423
rect 22376 22380 22428 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 5172 22176 5224 22228
rect 5632 22219 5684 22228
rect 5632 22185 5641 22219
rect 5641 22185 5675 22219
rect 5675 22185 5684 22219
rect 5632 22176 5684 22185
rect 6000 22219 6052 22228
rect 6000 22185 6009 22219
rect 6009 22185 6043 22219
rect 6043 22185 6052 22219
rect 6000 22176 6052 22185
rect 8484 22176 8536 22228
rect 10876 22219 10928 22228
rect 10876 22185 10885 22219
rect 10885 22185 10919 22219
rect 10919 22185 10928 22219
rect 10876 22176 10928 22185
rect 13084 22176 13136 22228
rect 13544 22176 13596 22228
rect 1676 22083 1728 22092
rect 1676 22049 1710 22083
rect 1710 22049 1728 22083
rect 1676 22040 1728 22049
rect 2228 22040 2280 22092
rect 2504 22040 2556 22092
rect 1308 21972 1360 22024
rect 2412 21972 2464 22024
rect 2688 21972 2740 22024
rect 3976 22040 4028 22092
rect 4988 22108 5040 22160
rect 5540 22108 5592 22160
rect 13636 22108 13688 22160
rect 6644 22040 6696 22092
rect 15108 22040 15160 22092
rect 15568 22083 15620 22092
rect 15568 22049 15591 22083
rect 15591 22049 15620 22083
rect 15568 22040 15620 22049
rect 4160 21972 4212 22024
rect 4528 22015 4580 22024
rect 4528 21981 4537 22015
rect 4537 21981 4571 22015
rect 4571 21981 4580 22015
rect 4528 21972 4580 21981
rect 6552 21972 6604 22024
rect 10968 22015 11020 22024
rect 6828 21904 6880 21956
rect 10968 21981 10977 22015
rect 10977 21981 11011 22015
rect 11011 21981 11020 22015
rect 10968 21972 11020 21981
rect 7748 21904 7800 21956
rect 9588 21904 9640 21956
rect 13636 21972 13688 22024
rect 15292 22015 15344 22024
rect 4160 21836 4212 21888
rect 4344 21836 4396 21888
rect 4620 21836 4672 21888
rect 6276 21836 6328 21888
rect 7104 21836 7156 21888
rect 7656 21836 7708 21888
rect 9036 21879 9088 21888
rect 9036 21845 9045 21879
rect 9045 21845 9079 21879
rect 9079 21845 9088 21879
rect 9036 21836 9088 21845
rect 9956 21836 10008 21888
rect 13728 21904 13780 21956
rect 15292 21981 15301 22015
rect 15301 21981 15335 22015
rect 15335 21981 15344 22015
rect 15292 21972 15344 21981
rect 16672 21947 16724 21956
rect 16672 21913 16681 21947
rect 16681 21913 16715 21947
rect 16715 21913 16724 21947
rect 16672 21904 16724 21913
rect 11520 21879 11572 21888
rect 11520 21845 11529 21879
rect 11529 21845 11563 21879
rect 11563 21845 11572 21879
rect 11520 21836 11572 21845
rect 13360 21879 13412 21888
rect 13360 21845 13369 21879
rect 13369 21845 13403 21879
rect 13403 21845 13412 21879
rect 13360 21836 13412 21845
rect 14464 21879 14516 21888
rect 14464 21845 14473 21879
rect 14473 21845 14507 21879
rect 14507 21845 14516 21879
rect 14464 21836 14516 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1308 21632 1360 21684
rect 2596 21632 2648 21684
rect 3608 21632 3660 21684
rect 8208 21632 8260 21684
rect 10876 21632 10928 21684
rect 13728 21632 13780 21684
rect 15568 21675 15620 21684
rect 15568 21641 15577 21675
rect 15577 21641 15611 21675
rect 15611 21641 15620 21675
rect 15568 21632 15620 21641
rect 5448 21539 5500 21548
rect 5448 21505 5457 21539
rect 5457 21505 5491 21539
rect 5491 21505 5500 21539
rect 5448 21496 5500 21505
rect 8208 21496 8260 21548
rect 9036 21496 9088 21548
rect 11060 21496 11112 21548
rect 12072 21496 12124 21548
rect 13728 21496 13780 21548
rect 13912 21496 13964 21548
rect 1860 21428 1912 21480
rect 6644 21428 6696 21480
rect 11244 21428 11296 21480
rect 14004 21428 14056 21480
rect 14188 21471 14240 21480
rect 14188 21437 14197 21471
rect 14197 21437 14231 21471
rect 14231 21437 14240 21471
rect 14188 21428 14240 21437
rect 2320 21360 2372 21412
rect 7564 21360 7616 21412
rect 8484 21360 8536 21412
rect 10876 21360 10928 21412
rect 3608 21335 3660 21344
rect 3608 21301 3617 21335
rect 3617 21301 3651 21335
rect 3651 21301 3660 21335
rect 3608 21292 3660 21301
rect 5172 21292 5224 21344
rect 5264 21335 5316 21344
rect 5264 21301 5273 21335
rect 5273 21301 5307 21335
rect 5307 21301 5316 21335
rect 6552 21335 6604 21344
rect 5264 21292 5316 21301
rect 6552 21301 6561 21335
rect 6561 21301 6595 21335
rect 6595 21301 6604 21335
rect 6552 21292 6604 21301
rect 7012 21335 7064 21344
rect 7012 21301 7021 21335
rect 7021 21301 7055 21335
rect 7055 21301 7064 21335
rect 7012 21292 7064 21301
rect 7656 21292 7708 21344
rect 8944 21335 8996 21344
rect 8944 21301 8953 21335
rect 8953 21301 8987 21335
rect 8987 21301 8996 21335
rect 8944 21292 8996 21301
rect 9036 21292 9088 21344
rect 10968 21292 11020 21344
rect 11520 21292 11572 21344
rect 12348 21292 12400 21344
rect 13912 21360 13964 21412
rect 14464 21403 14516 21412
rect 14464 21369 14476 21403
rect 14476 21369 14516 21403
rect 14464 21360 14516 21369
rect 26240 21360 26292 21412
rect 27620 21360 27672 21412
rect 13728 21292 13780 21344
rect 14188 21292 14240 21344
rect 15292 21292 15344 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1676 21131 1728 21140
rect 1676 21097 1685 21131
rect 1685 21097 1719 21131
rect 1719 21097 1728 21131
rect 1676 21088 1728 21097
rect 2320 21131 2372 21140
rect 2320 21097 2329 21131
rect 2329 21097 2363 21131
rect 2363 21097 2372 21131
rect 2320 21088 2372 21097
rect 2504 21088 2556 21140
rect 4528 21088 4580 21140
rect 5540 21088 5592 21140
rect 6092 21088 6144 21140
rect 7564 21088 7616 21140
rect 9036 21131 9088 21140
rect 9036 21097 9045 21131
rect 9045 21097 9079 21131
rect 9079 21097 9088 21131
rect 9036 21088 9088 21097
rect 13636 21131 13688 21140
rect 13636 21097 13645 21131
rect 13645 21097 13679 21131
rect 13679 21097 13688 21131
rect 13636 21088 13688 21097
rect 15568 21131 15620 21140
rect 15568 21097 15577 21131
rect 15577 21097 15611 21131
rect 15611 21097 15620 21131
rect 15568 21088 15620 21097
rect 9956 21063 10008 21072
rect 9956 21029 9990 21063
rect 9990 21029 10008 21063
rect 9956 21020 10008 21029
rect 1676 20884 1728 20936
rect 4068 20952 4120 21004
rect 5172 20952 5224 21004
rect 7288 20952 7340 21004
rect 9772 20952 9824 21004
rect 13360 21020 13412 21072
rect 14004 20995 14056 21004
rect 14004 20961 14013 20995
rect 14013 20961 14047 20995
rect 14047 20961 14056 20995
rect 14004 20952 14056 20961
rect 14740 20952 14792 21004
rect 4160 20884 4212 20936
rect 3608 20816 3660 20868
rect 4896 20927 4948 20936
rect 4896 20893 4905 20927
rect 4905 20893 4939 20927
rect 4939 20893 4948 20927
rect 4896 20884 4948 20893
rect 6000 20884 6052 20936
rect 6368 20927 6420 20936
rect 6368 20893 6377 20927
rect 6377 20893 6411 20927
rect 6411 20893 6420 20927
rect 6368 20884 6420 20893
rect 1492 20748 1544 20800
rect 2320 20748 2372 20800
rect 4160 20748 4212 20800
rect 5448 20748 5500 20800
rect 6184 20748 6236 20800
rect 7196 20884 7248 20936
rect 7288 20859 7340 20868
rect 7288 20825 7297 20859
rect 7297 20825 7331 20859
rect 7331 20825 7340 20859
rect 7288 20816 7340 20825
rect 12072 20884 12124 20936
rect 15568 20884 15620 20936
rect 7748 20748 7800 20800
rect 8484 20791 8536 20800
rect 8484 20757 8493 20791
rect 8493 20757 8527 20791
rect 8527 20757 8536 20791
rect 8484 20748 8536 20757
rect 11060 20791 11112 20800
rect 11060 20757 11069 20791
rect 11069 20757 11103 20791
rect 11103 20757 11112 20791
rect 11060 20748 11112 20757
rect 11244 20748 11296 20800
rect 11704 20748 11756 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1492 20544 1544 20596
rect 1952 20544 2004 20596
rect 2136 20544 2188 20596
rect 4896 20544 4948 20596
rect 5540 20587 5592 20596
rect 5540 20553 5549 20587
rect 5549 20553 5583 20587
rect 5583 20553 5592 20587
rect 5540 20544 5592 20553
rect 6092 20544 6144 20596
rect 7196 20587 7248 20596
rect 7196 20553 7205 20587
rect 7205 20553 7239 20587
rect 7239 20553 7248 20587
rect 7196 20544 7248 20553
rect 8300 20544 8352 20596
rect 3424 20451 3476 20460
rect 3424 20417 3433 20451
rect 3433 20417 3467 20451
rect 3467 20417 3476 20451
rect 3424 20408 3476 20417
rect 10048 20544 10100 20596
rect 12072 20544 12124 20596
rect 15568 20544 15620 20596
rect 4068 20340 4120 20392
rect 7104 20340 7156 20392
rect 8024 20340 8076 20392
rect 3608 20272 3660 20324
rect 8484 20272 8536 20324
rect 12440 20383 12492 20392
rect 12440 20349 12449 20383
rect 12449 20349 12483 20383
rect 12483 20349 12492 20383
rect 12440 20340 12492 20349
rect 12072 20272 12124 20324
rect 14004 20272 14056 20324
rect 14648 20272 14700 20324
rect 14832 20272 14884 20324
rect 1676 20247 1728 20256
rect 1676 20213 1685 20247
rect 1685 20213 1719 20247
rect 1719 20213 1728 20247
rect 1676 20204 1728 20213
rect 2044 20247 2096 20256
rect 2044 20213 2053 20247
rect 2053 20213 2087 20247
rect 2087 20213 2096 20247
rect 2044 20204 2096 20213
rect 6000 20247 6052 20256
rect 6000 20213 6009 20247
rect 6009 20213 6043 20247
rect 6043 20213 6052 20247
rect 6000 20204 6052 20213
rect 9772 20247 9824 20256
rect 9772 20213 9781 20247
rect 9781 20213 9815 20247
rect 9815 20213 9824 20247
rect 9772 20204 9824 20213
rect 13636 20204 13688 20256
rect 14740 20247 14792 20256
rect 14740 20213 14749 20247
rect 14749 20213 14783 20247
rect 14783 20213 14792 20247
rect 14740 20204 14792 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 2964 20043 3016 20052
rect 2964 20009 2973 20043
rect 2973 20009 3007 20043
rect 3007 20009 3016 20043
rect 2964 20000 3016 20009
rect 3608 20000 3660 20052
rect 6644 20000 6696 20052
rect 6920 20043 6972 20052
rect 6920 20009 6929 20043
rect 6929 20009 6963 20043
rect 6963 20009 6972 20043
rect 6920 20000 6972 20009
rect 7840 20000 7892 20052
rect 8024 20043 8076 20052
rect 8024 20009 8033 20043
rect 8033 20009 8067 20043
rect 8067 20009 8076 20043
rect 8024 20000 8076 20009
rect 9036 20000 9088 20052
rect 10048 20000 10100 20052
rect 12072 20000 12124 20052
rect 3332 19932 3384 19984
rect 4896 19932 4948 19984
rect 2136 19864 2188 19916
rect 3056 19864 3108 19916
rect 3424 19864 3476 19916
rect 7104 19932 7156 19984
rect 8944 19932 8996 19984
rect 11060 19932 11112 19984
rect 7288 19864 7340 19916
rect 14004 19864 14056 19916
rect 2044 19771 2096 19780
rect 2044 19737 2053 19771
rect 2053 19737 2087 19771
rect 2087 19737 2096 19771
rect 2044 19728 2096 19737
rect 6184 19728 6236 19780
rect 9772 19796 9824 19848
rect 10508 19839 10560 19848
rect 10508 19805 10517 19839
rect 10517 19805 10551 19839
rect 10551 19805 10560 19839
rect 10508 19796 10560 19805
rect 13268 19796 13320 19848
rect 13912 19839 13964 19848
rect 13912 19805 13921 19839
rect 13921 19805 13955 19839
rect 13955 19805 13964 19839
rect 13912 19796 13964 19805
rect 1400 19660 1452 19712
rect 5448 19703 5500 19712
rect 5448 19669 5457 19703
rect 5457 19669 5491 19703
rect 5491 19669 5500 19703
rect 5448 19660 5500 19669
rect 5540 19660 5592 19712
rect 8484 19703 8536 19712
rect 8484 19669 8493 19703
rect 8493 19669 8527 19703
rect 8527 19669 8536 19703
rect 8484 19660 8536 19669
rect 13176 19660 13228 19712
rect 13360 19703 13412 19712
rect 13360 19669 13369 19703
rect 13369 19669 13403 19703
rect 13403 19669 13412 19703
rect 13360 19660 13412 19669
rect 13728 19728 13780 19780
rect 14464 19660 14516 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 3332 19499 3384 19508
rect 3332 19465 3341 19499
rect 3341 19465 3375 19499
rect 3375 19465 3384 19499
rect 3332 19456 3384 19465
rect 6184 19499 6236 19508
rect 6184 19465 6193 19499
rect 6193 19465 6227 19499
rect 6227 19465 6236 19499
rect 6184 19456 6236 19465
rect 7656 19499 7708 19508
rect 7656 19465 7665 19499
rect 7665 19465 7699 19499
rect 7699 19465 7708 19499
rect 7656 19456 7708 19465
rect 10508 19456 10560 19508
rect 12440 19456 12492 19508
rect 12716 19456 12768 19508
rect 1584 19159 1636 19168
rect 1584 19125 1593 19159
rect 1593 19125 1627 19159
rect 1627 19125 1636 19159
rect 1584 19116 1636 19125
rect 2504 19295 2556 19304
rect 2504 19261 2513 19295
rect 2513 19261 2547 19295
rect 2547 19261 2556 19295
rect 2504 19252 2556 19261
rect 4344 19320 4396 19372
rect 5448 19320 5500 19372
rect 4160 19295 4212 19304
rect 4160 19261 4169 19295
rect 4169 19261 4203 19295
rect 4203 19261 4212 19295
rect 4160 19252 4212 19261
rect 5172 19295 5224 19304
rect 5172 19261 5181 19295
rect 5181 19261 5215 19295
rect 5215 19261 5224 19295
rect 5172 19252 5224 19261
rect 5264 19252 5316 19304
rect 7104 19320 7156 19372
rect 7288 19320 7340 19372
rect 7840 19320 7892 19372
rect 8484 19320 8536 19372
rect 11060 19388 11112 19440
rect 13728 19388 13780 19440
rect 13176 19363 13228 19372
rect 8944 19252 8996 19304
rect 11060 19252 11112 19304
rect 13176 19329 13185 19363
rect 13185 19329 13219 19363
rect 13219 19329 13228 19363
rect 13176 19320 13228 19329
rect 13912 19320 13964 19372
rect 13268 19252 13320 19304
rect 13636 19184 13688 19236
rect 14188 19295 14240 19304
rect 14188 19261 14197 19295
rect 14197 19261 14231 19295
rect 14231 19261 14240 19295
rect 14188 19252 14240 19261
rect 14464 19295 14516 19304
rect 14464 19261 14498 19295
rect 14498 19261 14516 19295
rect 14464 19252 14516 19261
rect 3700 19116 3752 19168
rect 4252 19159 4304 19168
rect 4252 19125 4261 19159
rect 4261 19125 4295 19159
rect 4295 19125 4304 19159
rect 4252 19116 4304 19125
rect 4712 19116 4764 19168
rect 6644 19116 6696 19168
rect 6920 19116 6972 19168
rect 7932 19116 7984 19168
rect 8484 19116 8536 19168
rect 9220 19159 9272 19168
rect 9220 19125 9229 19159
rect 9229 19125 9263 19159
rect 9263 19125 9272 19159
rect 9220 19116 9272 19125
rect 9588 19116 9640 19168
rect 10784 19159 10836 19168
rect 10784 19125 10793 19159
rect 10793 19125 10827 19159
rect 10827 19125 10836 19159
rect 10784 19116 10836 19125
rect 11796 19116 11848 19168
rect 12900 19116 12952 19168
rect 13268 19116 13320 19168
rect 14188 19116 14240 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1676 18912 1728 18964
rect 2688 18955 2740 18964
rect 2688 18921 2697 18955
rect 2697 18921 2731 18955
rect 2731 18921 2740 18955
rect 2688 18912 2740 18921
rect 3424 18912 3476 18964
rect 4252 18912 4304 18964
rect 5172 18912 5224 18964
rect 7472 18955 7524 18964
rect 7472 18921 7481 18955
rect 7481 18921 7515 18955
rect 7515 18921 7524 18955
rect 7472 18912 7524 18921
rect 9588 18912 9640 18964
rect 11244 18955 11296 18964
rect 11244 18921 11253 18955
rect 11253 18921 11287 18955
rect 11287 18921 11296 18955
rect 11244 18912 11296 18921
rect 11796 18955 11848 18964
rect 11796 18921 11805 18955
rect 11805 18921 11839 18955
rect 11839 18921 11848 18955
rect 11796 18912 11848 18921
rect 12348 18912 12400 18964
rect 13728 18912 13780 18964
rect 4160 18844 4212 18896
rect 4344 18887 4396 18896
rect 4344 18853 4353 18887
rect 4353 18853 4387 18887
rect 4387 18853 4396 18887
rect 4344 18844 4396 18853
rect 2228 18776 2280 18828
rect 2504 18819 2556 18828
rect 2504 18785 2513 18819
rect 2513 18785 2547 18819
rect 2547 18785 2556 18819
rect 2504 18776 2556 18785
rect 4252 18776 4304 18828
rect 5540 18844 5592 18896
rect 6644 18844 6696 18896
rect 10140 18844 10192 18896
rect 11060 18844 11112 18896
rect 12992 18887 13044 18896
rect 12992 18853 13026 18887
rect 13026 18853 13044 18887
rect 12992 18844 13044 18853
rect 13636 18844 13688 18896
rect 14096 18844 14148 18896
rect 14556 18844 14608 18896
rect 6184 18776 6236 18828
rect 8024 18819 8076 18828
rect 4896 18708 4948 18760
rect 8024 18785 8033 18819
rect 8033 18785 8067 18819
rect 8067 18785 8076 18819
rect 8024 18776 8076 18785
rect 11152 18819 11204 18828
rect 11152 18785 11161 18819
rect 11161 18785 11195 18819
rect 11195 18785 11204 18819
rect 11152 18776 11204 18785
rect 12716 18819 12768 18828
rect 12716 18785 12725 18819
rect 12725 18785 12759 18819
rect 12759 18785 12768 18819
rect 12716 18776 12768 18785
rect 13268 18776 13320 18828
rect 8208 18751 8260 18760
rect 8208 18717 8217 18751
rect 8217 18717 8251 18751
rect 8251 18717 8260 18751
rect 8208 18708 8260 18717
rect 10324 18751 10376 18760
rect 6828 18640 6880 18692
rect 10324 18717 10333 18751
rect 10333 18717 10367 18751
rect 10367 18717 10376 18751
rect 10324 18708 10376 18717
rect 15292 18751 15344 18760
rect 15292 18717 15301 18751
rect 15301 18717 15335 18751
rect 15335 18717 15344 18751
rect 15292 18708 15344 18717
rect 11336 18640 11388 18692
rect 14464 18640 14516 18692
rect 1400 18572 1452 18624
rect 2596 18572 2648 18624
rect 7012 18572 7064 18624
rect 7656 18615 7708 18624
rect 7656 18581 7665 18615
rect 7665 18581 7699 18615
rect 7699 18581 7708 18615
rect 7656 18572 7708 18581
rect 9864 18572 9916 18624
rect 10692 18615 10744 18624
rect 10692 18581 10701 18615
rect 10701 18581 10735 18615
rect 10735 18581 10744 18615
rect 10692 18572 10744 18581
rect 12716 18572 12768 18624
rect 13820 18572 13872 18624
rect 17592 18572 17644 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 2504 18411 2556 18420
rect 2504 18377 2513 18411
rect 2513 18377 2547 18411
rect 2547 18377 2556 18411
rect 2504 18368 2556 18377
rect 4896 18368 4948 18420
rect 8484 18411 8536 18420
rect 8484 18377 8493 18411
rect 8493 18377 8527 18411
rect 8527 18377 8536 18411
rect 8484 18368 8536 18377
rect 10048 18368 10100 18420
rect 10324 18368 10376 18420
rect 14004 18411 14056 18420
rect 14004 18377 14013 18411
rect 14013 18377 14047 18411
rect 14047 18377 14056 18411
rect 14004 18368 14056 18377
rect 9772 18300 9824 18352
rect 10600 18300 10652 18352
rect 3240 18232 3292 18284
rect 3516 18232 3568 18284
rect 9680 18232 9732 18284
rect 10692 18232 10744 18284
rect 12256 18275 12308 18284
rect 12256 18241 12265 18275
rect 12265 18241 12299 18275
rect 12299 18241 12308 18275
rect 12256 18232 12308 18241
rect 1676 18164 1728 18216
rect 3424 18164 3476 18216
rect 4344 18164 4396 18216
rect 7012 18164 7064 18216
rect 11244 18164 11296 18216
rect 13728 18164 13780 18216
rect 4712 18096 4764 18148
rect 6644 18096 6696 18148
rect 7380 18139 7432 18148
rect 7380 18105 7414 18139
rect 7414 18105 7432 18139
rect 7380 18096 7432 18105
rect 10140 18096 10192 18148
rect 10968 18096 11020 18148
rect 1492 18028 1544 18080
rect 2504 18028 2556 18080
rect 4160 18071 4212 18080
rect 4160 18037 4169 18071
rect 4169 18037 4203 18071
rect 4203 18037 4212 18071
rect 4160 18028 4212 18037
rect 4988 18028 5040 18080
rect 6828 18028 6880 18080
rect 9956 18071 10008 18080
rect 9956 18037 9965 18071
rect 9965 18037 9999 18071
rect 9999 18037 10008 18071
rect 9956 18028 10008 18037
rect 10876 18028 10928 18080
rect 11336 18071 11388 18080
rect 11336 18037 11345 18071
rect 11345 18037 11379 18071
rect 11379 18037 11388 18071
rect 11336 18028 11388 18037
rect 11612 18028 11664 18080
rect 12808 18071 12860 18080
rect 12808 18037 12817 18071
rect 12817 18037 12851 18071
rect 12851 18037 12860 18071
rect 12808 18028 12860 18037
rect 13268 18028 13320 18080
rect 14464 18300 14516 18352
rect 14464 18164 14516 18216
rect 15292 18164 15344 18216
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2044 17824 2096 17876
rect 4528 17867 4580 17876
rect 4528 17833 4537 17867
rect 4537 17833 4571 17867
rect 4571 17833 4580 17867
rect 4528 17824 4580 17833
rect 5172 17867 5224 17876
rect 5172 17833 5181 17867
rect 5181 17833 5215 17867
rect 5215 17833 5224 17867
rect 5172 17824 5224 17833
rect 6184 17867 6236 17876
rect 6184 17833 6193 17867
rect 6193 17833 6227 17867
rect 6227 17833 6236 17867
rect 6184 17824 6236 17833
rect 10692 17824 10744 17876
rect 12992 17867 13044 17876
rect 12992 17833 13001 17867
rect 13001 17833 13035 17867
rect 13035 17833 13044 17867
rect 12992 17824 13044 17833
rect 13452 17824 13504 17876
rect 13636 17824 13688 17876
rect 14464 17867 14516 17876
rect 14464 17833 14473 17867
rect 14473 17833 14507 17867
rect 14507 17833 14516 17867
rect 14464 17824 14516 17833
rect 2228 17799 2280 17808
rect 2228 17765 2237 17799
rect 2237 17765 2271 17799
rect 2271 17765 2280 17799
rect 2228 17756 2280 17765
rect 4252 17756 4304 17808
rect 8024 17756 8076 17808
rect 11428 17756 11480 17808
rect 5264 17688 5316 17740
rect 8208 17688 8260 17740
rect 10784 17688 10836 17740
rect 13360 17688 13412 17740
rect 13820 17731 13872 17740
rect 13820 17697 13829 17731
rect 13829 17697 13863 17731
rect 13863 17697 13872 17731
rect 13820 17688 13872 17697
rect 2504 17620 2556 17672
rect 3056 17663 3108 17672
rect 3056 17629 3065 17663
rect 3065 17629 3099 17663
rect 3099 17629 3108 17663
rect 3056 17620 3108 17629
rect 3516 17663 3568 17672
rect 3516 17629 3525 17663
rect 3525 17629 3559 17663
rect 3559 17629 3568 17663
rect 3516 17620 3568 17629
rect 4988 17620 5040 17672
rect 6368 17620 6420 17672
rect 2780 17552 2832 17604
rect 1952 17527 2004 17536
rect 1952 17493 1961 17527
rect 1961 17493 1995 17527
rect 1995 17493 2004 17527
rect 1952 17484 2004 17493
rect 2688 17484 2740 17536
rect 5540 17527 5592 17536
rect 5540 17493 5549 17527
rect 5549 17493 5583 17527
rect 5583 17493 5592 17527
rect 5540 17484 5592 17493
rect 6460 17527 6512 17536
rect 6460 17493 6469 17527
rect 6469 17493 6503 17527
rect 6503 17493 6512 17527
rect 6460 17484 6512 17493
rect 9404 17620 9456 17672
rect 10140 17595 10192 17604
rect 10140 17561 10149 17595
rect 10149 17561 10183 17595
rect 10183 17561 10192 17595
rect 10140 17552 10192 17561
rect 7012 17484 7064 17536
rect 7380 17484 7432 17536
rect 8208 17484 8260 17536
rect 8760 17484 8812 17536
rect 10692 17484 10744 17536
rect 10876 17484 10928 17536
rect 14004 17663 14056 17672
rect 14004 17629 14013 17663
rect 14013 17629 14047 17663
rect 14047 17629 14056 17663
rect 14004 17620 14056 17629
rect 11244 17484 11296 17536
rect 13268 17527 13320 17536
rect 13268 17493 13277 17527
rect 13277 17493 13311 17527
rect 13311 17493 13320 17527
rect 13268 17484 13320 17493
rect 13452 17527 13504 17536
rect 13452 17493 13461 17527
rect 13461 17493 13495 17527
rect 13495 17493 13504 17527
rect 13452 17484 13504 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2688 17280 2740 17332
rect 4528 17280 4580 17332
rect 5264 17323 5316 17332
rect 5264 17289 5273 17323
rect 5273 17289 5307 17323
rect 5307 17289 5316 17323
rect 5264 17280 5316 17289
rect 6460 17280 6512 17332
rect 8024 17280 8076 17332
rect 11244 17280 11296 17332
rect 13912 17280 13964 17332
rect 2320 17212 2372 17264
rect 7380 17187 7432 17196
rect 7380 17153 7389 17187
rect 7389 17153 7423 17187
rect 7423 17153 7432 17187
rect 7380 17144 7432 17153
rect 9404 17187 9456 17196
rect 9404 17153 9413 17187
rect 9413 17153 9447 17187
rect 9447 17153 9456 17187
rect 9404 17144 9456 17153
rect 1952 17076 2004 17128
rect 2964 17119 3016 17128
rect 2964 17085 2973 17119
rect 2973 17085 3007 17119
rect 3007 17085 3016 17119
rect 2964 17076 3016 17085
rect 3516 17076 3568 17128
rect 5724 17076 5776 17128
rect 7656 17076 7708 17128
rect 8668 17076 8720 17128
rect 9220 17076 9272 17128
rect 13268 17119 13320 17128
rect 13268 17085 13277 17119
rect 13277 17085 13311 17119
rect 13311 17085 13320 17119
rect 13268 17076 13320 17085
rect 2780 17008 2832 17060
rect 4068 17008 4120 17060
rect 5540 17008 5592 17060
rect 1584 16983 1636 16992
rect 1584 16949 1593 16983
rect 1593 16949 1627 16983
rect 1627 16949 1636 16983
rect 1584 16940 1636 16949
rect 2412 16940 2464 16992
rect 3056 16940 3108 16992
rect 4804 16940 4856 16992
rect 5632 16983 5684 16992
rect 5632 16949 5641 16983
rect 5641 16949 5675 16983
rect 5675 16949 5684 16983
rect 5632 16940 5684 16949
rect 6368 16940 6420 16992
rect 8760 17008 8812 17060
rect 7288 16983 7340 16992
rect 7288 16949 7297 16983
rect 7297 16949 7331 16983
rect 7331 16949 7340 16983
rect 8576 16983 8628 16992
rect 7288 16940 7340 16949
rect 8576 16949 8585 16983
rect 8585 16949 8619 16983
rect 8619 16949 8628 16983
rect 8576 16940 8628 16949
rect 9220 16983 9272 16992
rect 9220 16949 9229 16983
rect 9229 16949 9263 16983
rect 9263 16949 9272 16983
rect 9220 16940 9272 16949
rect 9588 17008 9640 17060
rect 14004 17008 14056 17060
rect 10140 16940 10192 16992
rect 11428 16940 11480 16992
rect 12072 16940 12124 16992
rect 13360 16940 13412 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1400 16736 1452 16788
rect 2044 16779 2096 16788
rect 2044 16745 2053 16779
rect 2053 16745 2087 16779
rect 2087 16745 2096 16779
rect 2044 16736 2096 16745
rect 2504 16736 2556 16788
rect 2688 16779 2740 16788
rect 2688 16745 2697 16779
rect 2697 16745 2731 16779
rect 2731 16745 2740 16779
rect 2688 16736 2740 16745
rect 3148 16779 3200 16788
rect 3148 16745 3157 16779
rect 3157 16745 3191 16779
rect 3191 16745 3200 16779
rect 3148 16736 3200 16745
rect 3976 16736 4028 16788
rect 6000 16779 6052 16788
rect 6000 16745 6009 16779
rect 6009 16745 6043 16779
rect 6043 16745 6052 16779
rect 6000 16736 6052 16745
rect 1492 16600 1544 16652
rect 4528 16711 4580 16720
rect 4528 16677 4537 16711
rect 4537 16677 4571 16711
rect 4571 16677 4580 16711
rect 7288 16736 7340 16788
rect 8668 16779 8720 16788
rect 4528 16668 4580 16677
rect 7840 16668 7892 16720
rect 8116 16668 8168 16720
rect 8668 16745 8677 16779
rect 8677 16745 8711 16779
rect 8711 16745 8720 16779
rect 8668 16736 8720 16745
rect 9588 16736 9640 16788
rect 9956 16736 10008 16788
rect 10784 16779 10836 16788
rect 10784 16745 10793 16779
rect 10793 16745 10827 16779
rect 10827 16745 10836 16779
rect 10784 16736 10836 16745
rect 14004 16779 14056 16788
rect 14004 16745 14013 16779
rect 14013 16745 14047 16779
rect 14047 16745 14056 16779
rect 14004 16736 14056 16745
rect 13636 16711 13688 16720
rect 13636 16677 13645 16711
rect 13645 16677 13679 16711
rect 13679 16677 13688 16711
rect 13636 16668 13688 16677
rect 3424 16643 3476 16652
rect 3424 16609 3433 16643
rect 3433 16609 3467 16643
rect 3467 16609 3476 16643
rect 3424 16600 3476 16609
rect 4896 16600 4948 16652
rect 5724 16600 5776 16652
rect 4804 16532 4856 16584
rect 6184 16532 6236 16584
rect 7012 16600 7064 16652
rect 11980 16643 12032 16652
rect 11980 16609 12014 16643
rect 12014 16609 12032 16643
rect 4988 16464 5040 16516
rect 5264 16464 5316 16516
rect 7196 16532 7248 16584
rect 8024 16532 8076 16584
rect 9680 16532 9732 16584
rect 11980 16600 12032 16609
rect 10140 16532 10192 16584
rect 11244 16532 11296 16584
rect 11704 16575 11756 16584
rect 11704 16541 11713 16575
rect 11713 16541 11747 16575
rect 11747 16541 11756 16575
rect 11704 16532 11756 16541
rect 4068 16439 4120 16448
rect 4068 16405 4077 16439
rect 4077 16405 4111 16439
rect 4111 16405 4120 16439
rect 4068 16396 4120 16405
rect 6368 16396 6420 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2044 16235 2096 16244
rect 2044 16201 2053 16235
rect 2053 16201 2087 16235
rect 2087 16201 2096 16235
rect 2044 16192 2096 16201
rect 4804 16235 4856 16244
rect 4804 16201 4813 16235
rect 4813 16201 4847 16235
rect 4847 16201 4856 16235
rect 4804 16192 4856 16201
rect 5264 16235 5316 16244
rect 5264 16201 5273 16235
rect 5273 16201 5307 16235
rect 5307 16201 5316 16235
rect 5264 16192 5316 16201
rect 6000 16192 6052 16244
rect 11060 16192 11112 16244
rect 11980 16192 12032 16244
rect 11704 16167 11756 16176
rect 11704 16133 11713 16167
rect 11713 16133 11747 16167
rect 11747 16133 11756 16167
rect 11704 16124 11756 16133
rect 2412 16099 2464 16108
rect 2412 16065 2421 16099
rect 2421 16065 2455 16099
rect 2455 16065 2464 16099
rect 2412 16056 2464 16065
rect 2044 15988 2096 16040
rect 6368 16056 6420 16108
rect 9220 16056 9272 16108
rect 1584 15895 1636 15904
rect 1584 15861 1593 15895
rect 1593 15861 1627 15895
rect 1627 15861 1636 15895
rect 1584 15852 1636 15861
rect 7196 15988 7248 16040
rect 9680 16031 9732 16040
rect 9680 15997 9689 16031
rect 9689 15997 9723 16031
rect 9723 15997 9732 16031
rect 9680 15988 9732 15997
rect 10048 16031 10100 16040
rect 10048 15997 10082 16031
rect 10082 15997 10100 16031
rect 10048 15988 10100 15997
rect 12808 16056 12860 16108
rect 13268 15988 13320 16040
rect 13912 15920 13964 15972
rect 2964 15852 3016 15904
rect 4344 15852 4396 15904
rect 5724 15895 5776 15904
rect 5724 15861 5733 15895
rect 5733 15861 5767 15895
rect 5767 15861 5776 15895
rect 5724 15852 5776 15861
rect 6276 15895 6328 15904
rect 6276 15861 6285 15895
rect 6285 15861 6319 15895
rect 6319 15861 6328 15895
rect 6276 15852 6328 15861
rect 6920 15852 6972 15904
rect 8760 15852 8812 15904
rect 9220 15895 9272 15904
rect 9220 15861 9229 15895
rect 9229 15861 9263 15895
rect 9263 15861 9272 15895
rect 9220 15852 9272 15861
rect 13728 15852 13780 15904
rect 15108 15895 15160 15904
rect 15108 15861 15117 15895
rect 15117 15861 15151 15895
rect 15151 15861 15160 15895
rect 15108 15852 15160 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1492 15648 1544 15700
rect 2320 15691 2372 15700
rect 2320 15657 2329 15691
rect 2329 15657 2363 15691
rect 2363 15657 2372 15691
rect 2320 15648 2372 15657
rect 4068 15648 4120 15700
rect 4252 15691 4304 15700
rect 4252 15657 4261 15691
rect 4261 15657 4295 15691
rect 4295 15657 4304 15691
rect 4252 15648 4304 15657
rect 4528 15691 4580 15700
rect 4528 15657 4537 15691
rect 4537 15657 4571 15691
rect 4571 15657 4580 15691
rect 4528 15648 4580 15657
rect 5540 15648 5592 15700
rect 5724 15648 5776 15700
rect 7196 15648 7248 15700
rect 7840 15648 7892 15700
rect 8024 15691 8076 15700
rect 8024 15657 8033 15691
rect 8033 15657 8067 15691
rect 8067 15657 8076 15691
rect 8024 15648 8076 15657
rect 9956 15648 10008 15700
rect 10140 15648 10192 15700
rect 10784 15691 10836 15700
rect 10784 15657 10793 15691
rect 10793 15657 10827 15691
rect 10827 15657 10836 15691
rect 10784 15648 10836 15657
rect 11244 15691 11296 15700
rect 11244 15657 11253 15691
rect 11253 15657 11287 15691
rect 11287 15657 11296 15691
rect 11244 15648 11296 15657
rect 3976 15580 4028 15632
rect 2044 15512 2096 15564
rect 4160 15512 4212 15564
rect 6184 15580 6236 15632
rect 6368 15580 6420 15632
rect 8484 15580 8536 15632
rect 11612 15580 11664 15632
rect 12808 15580 12860 15632
rect 6000 15555 6052 15564
rect 6000 15521 6034 15555
rect 6034 15521 6052 15555
rect 6000 15512 6052 15521
rect 10048 15512 10100 15564
rect 3056 15487 3108 15496
rect 3056 15453 3065 15487
rect 3065 15453 3099 15487
rect 3099 15453 3108 15487
rect 3056 15444 3108 15453
rect 8576 15487 8628 15496
rect 8576 15453 8585 15487
rect 8585 15453 8619 15487
rect 8619 15453 8628 15487
rect 8576 15444 8628 15453
rect 10968 15444 11020 15496
rect 11428 15487 11480 15496
rect 11428 15453 11437 15487
rect 11437 15453 11471 15487
rect 11471 15453 11480 15487
rect 11428 15444 11480 15453
rect 12440 15444 12492 15496
rect 13452 15512 13504 15564
rect 13176 15444 13228 15496
rect 13912 15648 13964 15700
rect 14372 15691 14424 15700
rect 14372 15657 14381 15691
rect 14381 15657 14415 15691
rect 14415 15657 14424 15691
rect 14372 15648 14424 15657
rect 16304 15580 16356 15632
rect 14188 15555 14240 15564
rect 14188 15521 14197 15555
rect 14197 15521 14231 15555
rect 14231 15521 14240 15555
rect 14188 15512 14240 15521
rect 2504 15376 2556 15428
rect 14648 15419 14700 15428
rect 14648 15385 14657 15419
rect 14657 15385 14691 15419
rect 14691 15385 14700 15419
rect 14648 15376 14700 15385
rect 15844 15376 15896 15428
rect 2780 15308 2832 15360
rect 5448 15308 5500 15360
rect 6828 15308 6880 15360
rect 8300 15308 8352 15360
rect 9036 15351 9088 15360
rect 9036 15317 9045 15351
rect 9045 15317 9079 15351
rect 9079 15317 9088 15351
rect 9036 15308 9088 15317
rect 15476 15308 15528 15360
rect 16488 15351 16540 15360
rect 16488 15317 16497 15351
rect 16497 15317 16531 15351
rect 16531 15317 16540 15351
rect 16488 15308 16540 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2044 15147 2096 15156
rect 2044 15113 2053 15147
rect 2053 15113 2087 15147
rect 2087 15113 2096 15147
rect 2044 15104 2096 15113
rect 4068 15104 4120 15156
rect 5448 15104 5500 15156
rect 7196 15104 7248 15156
rect 8484 15147 8536 15156
rect 8484 15113 8493 15147
rect 8493 15113 8527 15147
rect 8527 15113 8536 15147
rect 8484 15104 8536 15113
rect 10048 15147 10100 15156
rect 10048 15113 10057 15147
rect 10057 15113 10091 15147
rect 10091 15113 10100 15147
rect 10048 15104 10100 15113
rect 10968 15104 11020 15156
rect 11244 15147 11296 15156
rect 11244 15113 11253 15147
rect 11253 15113 11287 15147
rect 11287 15113 11296 15147
rect 11244 15104 11296 15113
rect 11612 15147 11664 15156
rect 11612 15113 11621 15147
rect 11621 15113 11655 15147
rect 11655 15113 11664 15147
rect 11612 15104 11664 15113
rect 12348 15104 12400 15156
rect 13176 15104 13228 15156
rect 16304 15104 16356 15156
rect 4160 15079 4212 15088
rect 4160 15045 4169 15079
rect 4169 15045 4203 15079
rect 4203 15045 4212 15079
rect 4160 15036 4212 15045
rect 5356 15036 5408 15088
rect 2596 14968 2648 15020
rect 2872 14968 2924 15020
rect 6000 14968 6052 15020
rect 2504 14943 2556 14952
rect 2504 14909 2513 14943
rect 2513 14909 2547 14943
rect 2547 14909 2556 14943
rect 2504 14900 2556 14909
rect 2780 14900 2832 14952
rect 3608 14943 3660 14952
rect 3608 14909 3617 14943
rect 3617 14909 3651 14943
rect 3651 14909 3660 14943
rect 3608 14900 3660 14909
rect 5540 14943 5592 14952
rect 5540 14909 5549 14943
rect 5549 14909 5583 14943
rect 5583 14909 5592 14943
rect 5540 14900 5592 14909
rect 6828 14900 6880 14952
rect 7288 14943 7340 14952
rect 7288 14909 7297 14943
rect 7297 14909 7331 14943
rect 7331 14909 7340 14943
rect 7288 14900 7340 14909
rect 8208 14900 8260 14952
rect 16488 14968 16540 15020
rect 17868 14968 17920 15020
rect 9220 14900 9272 14952
rect 13728 14900 13780 14952
rect 3056 14832 3108 14884
rect 4344 14832 4396 14884
rect 6552 14832 6604 14884
rect 8760 14832 8812 14884
rect 13176 14832 13228 14884
rect 14096 14832 14148 14884
rect 1400 14764 1452 14816
rect 2688 14807 2740 14816
rect 2688 14773 2697 14807
rect 2697 14773 2731 14807
rect 2731 14773 2740 14807
rect 2688 14764 2740 14773
rect 4160 14764 4212 14816
rect 6184 14807 6236 14816
rect 6184 14773 6193 14807
rect 6193 14773 6227 14807
rect 6227 14773 6236 14807
rect 6184 14764 6236 14773
rect 6828 14807 6880 14816
rect 6828 14773 6837 14807
rect 6837 14773 6871 14807
rect 6871 14773 6880 14807
rect 6828 14764 6880 14773
rect 7840 14807 7892 14816
rect 7840 14773 7849 14807
rect 7849 14773 7883 14807
rect 7883 14773 7892 14807
rect 7840 14764 7892 14773
rect 12808 14764 12860 14816
rect 14372 14764 14424 14816
rect 15384 14764 15436 14816
rect 15844 14807 15896 14816
rect 15844 14773 15853 14807
rect 15853 14773 15887 14807
rect 15887 14773 15896 14807
rect 15844 14764 15896 14773
rect 16212 14807 16264 14816
rect 16212 14773 16221 14807
rect 16221 14773 16255 14807
rect 16255 14773 16264 14807
rect 16212 14764 16264 14773
rect 16396 14764 16448 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2504 14560 2556 14612
rect 3608 14603 3660 14612
rect 3608 14569 3617 14603
rect 3617 14569 3651 14603
rect 3651 14569 3660 14603
rect 3608 14560 3660 14569
rect 6000 14603 6052 14612
rect 6000 14569 6009 14603
rect 6009 14569 6043 14603
rect 6043 14569 6052 14603
rect 6000 14560 6052 14569
rect 7380 14560 7432 14612
rect 9772 14560 9824 14612
rect 9864 14560 9916 14612
rect 14096 14603 14148 14612
rect 14096 14569 14105 14603
rect 14105 14569 14139 14603
rect 14139 14569 14148 14603
rect 14096 14560 14148 14569
rect 16304 14560 16356 14612
rect 6552 14492 6604 14544
rect 2044 14424 2096 14476
rect 2228 14424 2280 14476
rect 4160 14424 4212 14476
rect 4344 14467 4396 14476
rect 4344 14433 4378 14467
rect 4378 14433 4396 14467
rect 4344 14424 4396 14433
rect 9956 14424 10008 14476
rect 13360 14424 13412 14476
rect 15660 14467 15712 14476
rect 2872 14399 2924 14408
rect 2872 14365 2881 14399
rect 2881 14365 2915 14399
rect 2915 14365 2924 14399
rect 2872 14356 2924 14365
rect 3516 14356 3568 14408
rect 6184 14356 6236 14408
rect 11060 14356 11112 14408
rect 12716 14399 12768 14408
rect 12716 14365 12725 14399
rect 12725 14365 12759 14399
rect 12759 14365 12768 14399
rect 12716 14356 12768 14365
rect 15660 14433 15669 14467
rect 15669 14433 15703 14467
rect 15703 14433 15712 14467
rect 15660 14424 15712 14433
rect 17224 14467 17276 14476
rect 17224 14433 17233 14467
rect 17233 14433 17267 14467
rect 17267 14433 17276 14467
rect 17224 14424 17276 14433
rect 15844 14399 15896 14408
rect 15844 14365 15853 14399
rect 15853 14365 15887 14399
rect 15887 14365 15896 14399
rect 15844 14356 15896 14365
rect 16396 14399 16448 14408
rect 16396 14365 16405 14399
rect 16405 14365 16439 14399
rect 16439 14365 16448 14399
rect 16396 14356 16448 14365
rect 16856 14356 16908 14408
rect 17868 14356 17920 14408
rect 14096 14288 14148 14340
rect 16212 14288 16264 14340
rect 1860 14263 1912 14272
rect 1860 14229 1869 14263
rect 1869 14229 1903 14263
rect 1903 14229 1912 14263
rect 1860 14220 1912 14229
rect 2412 14263 2464 14272
rect 2412 14229 2421 14263
rect 2421 14229 2455 14263
rect 2455 14229 2464 14263
rect 2412 14220 2464 14229
rect 6368 14263 6420 14272
rect 6368 14229 6377 14263
rect 6377 14229 6411 14263
rect 6411 14229 6420 14263
rect 6368 14220 6420 14229
rect 8760 14263 8812 14272
rect 8760 14229 8769 14263
rect 8769 14229 8803 14263
rect 8803 14229 8812 14263
rect 8760 14220 8812 14229
rect 9588 14220 9640 14272
rect 12532 14263 12584 14272
rect 12532 14229 12541 14263
rect 12541 14229 12575 14263
rect 12575 14229 12584 14263
rect 12532 14220 12584 14229
rect 14648 14263 14700 14272
rect 14648 14229 14657 14263
rect 14657 14229 14691 14263
rect 14691 14229 14700 14263
rect 14648 14220 14700 14229
rect 15292 14263 15344 14272
rect 15292 14229 15301 14263
rect 15301 14229 15335 14263
rect 15335 14229 15344 14263
rect 15292 14220 15344 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 4344 14016 4396 14068
rect 4804 14016 4856 14068
rect 5172 14059 5224 14068
rect 1584 13991 1636 14000
rect 1584 13957 1593 13991
rect 1593 13957 1627 13991
rect 1627 13957 1636 13991
rect 1584 13948 1636 13957
rect 3792 13948 3844 14000
rect 3332 13923 3384 13932
rect 3332 13889 3341 13923
rect 3341 13889 3375 13923
rect 3375 13889 3384 13923
rect 3332 13880 3384 13889
rect 3516 13923 3568 13932
rect 3516 13889 3525 13923
rect 3525 13889 3559 13923
rect 3559 13889 3568 13923
rect 3516 13880 3568 13889
rect 5172 14025 5181 14059
rect 5181 14025 5215 14059
rect 5215 14025 5224 14059
rect 5172 14016 5224 14025
rect 6184 14059 6236 14068
rect 6184 14025 6193 14059
rect 6193 14025 6227 14059
rect 6227 14025 6236 14059
rect 6184 14016 6236 14025
rect 7288 14016 7340 14068
rect 8576 14016 8628 14068
rect 9772 14059 9824 14068
rect 6092 13948 6144 14000
rect 6736 13948 6788 14000
rect 8208 13948 8260 14000
rect 5448 13880 5500 13932
rect 6368 13880 6420 13932
rect 7380 13923 7432 13932
rect 7380 13889 7389 13923
rect 7389 13889 7423 13923
rect 7423 13889 7432 13923
rect 7380 13880 7432 13889
rect 9036 13923 9088 13932
rect 9036 13889 9045 13923
rect 9045 13889 9079 13923
rect 9079 13889 9088 13923
rect 9036 13880 9088 13889
rect 1860 13812 1912 13864
rect 2228 13812 2280 13864
rect 2136 13719 2188 13728
rect 2136 13685 2145 13719
rect 2145 13685 2179 13719
rect 2179 13685 2188 13719
rect 2136 13676 2188 13685
rect 2320 13676 2372 13728
rect 2964 13812 3016 13864
rect 4252 13812 4304 13864
rect 3240 13787 3292 13796
rect 3240 13753 3249 13787
rect 3249 13753 3283 13787
rect 3283 13753 3292 13787
rect 3240 13744 3292 13753
rect 4528 13744 4580 13796
rect 4712 13744 4764 13796
rect 7196 13812 7248 13864
rect 7840 13812 7892 13864
rect 8392 13812 8444 13864
rect 8852 13855 8904 13864
rect 8852 13821 8861 13855
rect 8861 13821 8895 13855
rect 8895 13821 8904 13855
rect 8852 13812 8904 13821
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 9956 14059 10008 14068
rect 9956 14025 9965 14059
rect 9965 14025 9999 14059
rect 9999 14025 10008 14059
rect 9956 14016 10008 14025
rect 11060 14059 11112 14068
rect 11060 14025 11069 14059
rect 11069 14025 11103 14059
rect 11103 14025 11112 14059
rect 11060 14016 11112 14025
rect 14188 14016 14240 14068
rect 14648 14016 14700 14068
rect 9864 13948 9916 14000
rect 12716 13948 12768 14000
rect 14372 13948 14424 14000
rect 10048 13880 10100 13932
rect 10692 13880 10744 13932
rect 12256 13923 12308 13932
rect 12256 13889 12265 13923
rect 12265 13889 12299 13923
rect 12299 13889 12308 13923
rect 12256 13880 12308 13889
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 8668 13744 8720 13796
rect 14372 13812 14424 13864
rect 14924 13812 14976 13864
rect 15384 13812 15436 13864
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 17224 13855 17276 13864
rect 17224 13821 17233 13855
rect 17233 13821 17267 13855
rect 17267 13821 17276 13855
rect 17224 13812 17276 13821
rect 15292 13744 15344 13796
rect 8392 13676 8444 13728
rect 13636 13719 13688 13728
rect 13636 13685 13645 13719
rect 13645 13685 13679 13719
rect 13679 13685 13688 13719
rect 13636 13676 13688 13685
rect 13728 13719 13780 13728
rect 13728 13685 13737 13719
rect 13737 13685 13771 13719
rect 13771 13685 13780 13719
rect 13728 13676 13780 13685
rect 15384 13676 15436 13728
rect 15568 13676 15620 13728
rect 16212 13719 16264 13728
rect 16212 13685 16221 13719
rect 16221 13685 16255 13719
rect 16255 13685 16264 13719
rect 16212 13676 16264 13685
rect 17868 13676 17920 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1860 13472 1912 13524
rect 2136 13472 2188 13524
rect 2780 13515 2832 13524
rect 2780 13481 2789 13515
rect 2789 13481 2823 13515
rect 2823 13481 2832 13515
rect 2780 13472 2832 13481
rect 4160 13472 4212 13524
rect 3424 13404 3476 13456
rect 3884 13447 3936 13456
rect 3884 13413 3893 13447
rect 3893 13413 3927 13447
rect 3927 13413 3936 13447
rect 3884 13404 3936 13413
rect 4528 13472 4580 13524
rect 6552 13472 6604 13524
rect 7196 13515 7248 13524
rect 6184 13404 6236 13456
rect 7196 13481 7205 13515
rect 7205 13481 7239 13515
rect 7239 13481 7248 13515
rect 7196 13472 7248 13481
rect 7472 13472 7524 13524
rect 8576 13472 8628 13524
rect 9404 13515 9456 13524
rect 9404 13481 9413 13515
rect 9413 13481 9447 13515
rect 9447 13481 9456 13515
rect 9404 13472 9456 13481
rect 10692 13515 10744 13524
rect 10692 13481 10701 13515
rect 10701 13481 10735 13515
rect 10735 13481 10744 13515
rect 10692 13472 10744 13481
rect 11336 13472 11388 13524
rect 11520 13472 11572 13524
rect 12440 13472 12492 13524
rect 12716 13472 12768 13524
rect 13176 13515 13228 13524
rect 13176 13481 13185 13515
rect 13185 13481 13219 13515
rect 13219 13481 13228 13515
rect 13176 13472 13228 13481
rect 13452 13472 13504 13524
rect 13728 13472 13780 13524
rect 14004 13515 14056 13524
rect 14004 13481 14013 13515
rect 14013 13481 14047 13515
rect 14047 13481 14056 13515
rect 14004 13472 14056 13481
rect 14924 13515 14976 13524
rect 14924 13481 14933 13515
rect 14933 13481 14967 13515
rect 14967 13481 14976 13515
rect 14924 13472 14976 13481
rect 16304 13515 16356 13524
rect 16304 13481 16313 13515
rect 16313 13481 16347 13515
rect 16347 13481 16356 13515
rect 16304 13472 16356 13481
rect 1400 13379 1452 13388
rect 1400 13345 1409 13379
rect 1409 13345 1443 13379
rect 1443 13345 1452 13379
rect 1400 13336 1452 13345
rect 1952 13379 2004 13388
rect 1952 13345 1961 13379
rect 1961 13345 1995 13379
rect 1995 13345 2004 13379
rect 1952 13336 2004 13345
rect 4804 13336 4856 13388
rect 7380 13336 7432 13388
rect 7564 13379 7616 13388
rect 7564 13345 7573 13379
rect 7573 13345 7607 13379
rect 7607 13345 7616 13379
rect 7564 13336 7616 13345
rect 15568 13404 15620 13456
rect 16212 13404 16264 13456
rect 18236 13447 18288 13456
rect 18236 13413 18270 13447
rect 18270 13413 18288 13447
rect 18236 13404 18288 13413
rect 11612 13379 11664 13388
rect 4712 13311 4764 13320
rect 2136 13200 2188 13252
rect 4712 13277 4721 13311
rect 4721 13277 4755 13311
rect 4755 13277 4764 13311
rect 4712 13268 4764 13277
rect 6368 13268 6420 13320
rect 11612 13345 11621 13379
rect 11621 13345 11655 13379
rect 11655 13345 11664 13379
rect 11612 13336 11664 13345
rect 15844 13336 15896 13388
rect 18512 13336 18564 13388
rect 10048 13268 10100 13320
rect 3516 13243 3568 13252
rect 3516 13209 3525 13243
rect 3525 13209 3559 13243
rect 3559 13209 3568 13243
rect 3516 13200 3568 13209
rect 4068 13200 4120 13252
rect 5632 13243 5684 13252
rect 5632 13209 5641 13243
rect 5641 13209 5675 13243
rect 5675 13209 5684 13243
rect 5632 13200 5684 13209
rect 9036 13200 9088 13252
rect 11796 13268 11848 13320
rect 11980 13268 12032 13320
rect 14096 13311 14148 13320
rect 14096 13277 14105 13311
rect 14105 13277 14139 13311
rect 14139 13277 14148 13311
rect 14096 13268 14148 13277
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 15936 13311 15988 13320
rect 15936 13277 15945 13311
rect 15945 13277 15979 13311
rect 15979 13277 15988 13311
rect 15936 13268 15988 13277
rect 16672 13311 16724 13320
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 17408 13200 17460 13252
rect 2596 13132 2648 13184
rect 3148 13132 3200 13184
rect 5540 13132 5592 13184
rect 6828 13132 6880 13184
rect 8392 13175 8444 13184
rect 8392 13141 8401 13175
rect 8401 13141 8435 13175
rect 8435 13141 8444 13175
rect 8392 13132 8444 13141
rect 8484 13132 8536 13184
rect 9864 13132 9916 13184
rect 10876 13132 10928 13184
rect 10968 13132 11020 13184
rect 12440 13175 12492 13184
rect 12440 13141 12449 13175
rect 12449 13141 12483 13175
rect 12483 13141 12492 13175
rect 12440 13132 12492 13141
rect 13360 13132 13412 13184
rect 16028 13132 16080 13184
rect 19340 13175 19392 13184
rect 19340 13141 19349 13175
rect 19349 13141 19383 13175
rect 19383 13141 19392 13175
rect 19340 13132 19392 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2320 12928 2372 12980
rect 4528 12928 4580 12980
rect 5172 12971 5224 12980
rect 4804 12860 4856 12912
rect 5172 12937 5181 12971
rect 5181 12937 5215 12971
rect 5215 12937 5224 12971
rect 5172 12928 5224 12937
rect 6184 12971 6236 12980
rect 6184 12937 6193 12971
rect 6193 12937 6227 12971
rect 6227 12937 6236 12971
rect 6184 12928 6236 12937
rect 6552 12971 6604 12980
rect 6552 12937 6561 12971
rect 6561 12937 6595 12971
rect 6595 12937 6604 12971
rect 6552 12928 6604 12937
rect 7564 12928 7616 12980
rect 7932 12928 7984 12980
rect 8392 12928 8444 12980
rect 6368 12860 6420 12912
rect 5724 12835 5776 12844
rect 5724 12801 5733 12835
rect 5733 12801 5767 12835
rect 5767 12801 5776 12835
rect 5724 12792 5776 12801
rect 6552 12792 6604 12844
rect 6920 12792 6972 12844
rect 7472 12835 7524 12844
rect 7472 12801 7481 12835
rect 7481 12801 7515 12835
rect 7515 12801 7524 12835
rect 7472 12792 7524 12801
rect 9220 12928 9272 12980
rect 11244 12928 11296 12980
rect 11612 12928 11664 12980
rect 11980 12971 12032 12980
rect 11980 12937 11989 12971
rect 11989 12937 12023 12971
rect 12023 12937 12032 12971
rect 11980 12928 12032 12937
rect 13636 12928 13688 12980
rect 14004 12971 14056 12980
rect 14004 12937 14013 12971
rect 14013 12937 14047 12971
rect 14047 12937 14056 12971
rect 14004 12928 14056 12937
rect 14648 12928 14700 12980
rect 15844 12928 15896 12980
rect 17408 12971 17460 12980
rect 17408 12937 17417 12971
rect 17417 12937 17451 12971
rect 17451 12937 17460 12971
rect 17408 12928 17460 12937
rect 18236 12971 18288 12980
rect 18236 12937 18245 12971
rect 18245 12937 18279 12971
rect 18279 12937 18288 12971
rect 18236 12928 18288 12937
rect 18512 12928 18564 12980
rect 12900 12860 12952 12912
rect 11520 12792 11572 12844
rect 13176 12792 13228 12844
rect 2136 12724 2188 12776
rect 4160 12724 4212 12776
rect 7196 12767 7248 12776
rect 7196 12733 7205 12767
rect 7205 12733 7239 12767
rect 7239 12733 7248 12767
rect 7196 12724 7248 12733
rect 12440 12724 12492 12776
rect 12900 12724 12952 12776
rect 2780 12656 2832 12708
rect 2136 12588 2188 12640
rect 3424 12631 3476 12640
rect 3424 12597 3433 12631
rect 3433 12597 3467 12631
rect 3467 12597 3476 12631
rect 3424 12588 3476 12597
rect 5540 12631 5592 12640
rect 5540 12597 5549 12631
rect 5549 12597 5583 12631
rect 5583 12597 5592 12631
rect 5540 12588 5592 12597
rect 5632 12631 5684 12640
rect 5632 12597 5641 12631
rect 5641 12597 5675 12631
rect 5675 12597 5684 12631
rect 9036 12656 9088 12708
rect 12716 12656 12768 12708
rect 13176 12656 13228 12708
rect 14280 12792 14332 12844
rect 17960 12792 18012 12844
rect 18236 12792 18288 12844
rect 13636 12767 13688 12776
rect 13636 12733 13645 12767
rect 13645 12733 13679 12767
rect 13679 12733 13688 12767
rect 13636 12724 13688 12733
rect 14096 12724 14148 12776
rect 15292 12724 15344 12776
rect 15568 12724 15620 12776
rect 15660 12656 15712 12708
rect 5632 12588 5684 12597
rect 7288 12631 7340 12640
rect 7288 12597 7297 12631
rect 7297 12597 7331 12631
rect 7331 12597 7340 12631
rect 7288 12588 7340 12597
rect 9956 12588 10008 12640
rect 12532 12588 12584 12640
rect 13544 12588 13596 12640
rect 13636 12588 13688 12640
rect 16856 12631 16908 12640
rect 16856 12597 16865 12631
rect 16865 12597 16899 12631
rect 16899 12597 16908 12631
rect 16856 12588 16908 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 3700 12427 3752 12436
rect 3700 12393 3709 12427
rect 3709 12393 3743 12427
rect 3743 12393 3752 12427
rect 3700 12384 3752 12393
rect 5724 12384 5776 12436
rect 6184 12384 6236 12436
rect 6460 12384 6512 12436
rect 6552 12384 6604 12436
rect 7380 12427 7432 12436
rect 7380 12393 7389 12427
rect 7389 12393 7423 12427
rect 7423 12393 7432 12427
rect 7380 12384 7432 12393
rect 7472 12384 7524 12436
rect 8484 12384 8536 12436
rect 9036 12427 9088 12436
rect 9036 12393 9045 12427
rect 9045 12393 9079 12427
rect 9079 12393 9088 12427
rect 9036 12384 9088 12393
rect 9404 12427 9456 12436
rect 9404 12393 9413 12427
rect 9413 12393 9447 12427
rect 9447 12393 9456 12427
rect 9404 12384 9456 12393
rect 9864 12384 9916 12436
rect 12348 12384 12400 12436
rect 12532 12427 12584 12436
rect 12532 12393 12541 12427
rect 12541 12393 12575 12427
rect 12575 12393 12584 12427
rect 12532 12384 12584 12393
rect 13176 12427 13228 12436
rect 13176 12393 13185 12427
rect 13185 12393 13219 12427
rect 13219 12393 13228 12427
rect 13176 12384 13228 12393
rect 13360 12384 13412 12436
rect 13912 12384 13964 12436
rect 15568 12427 15620 12436
rect 15568 12393 15577 12427
rect 15577 12393 15611 12427
rect 15611 12393 15620 12427
rect 15568 12384 15620 12393
rect 16488 12384 16540 12436
rect 1952 12316 2004 12368
rect 10876 12316 10928 12368
rect 15476 12316 15528 12368
rect 4804 12248 4856 12300
rect 5448 12248 5500 12300
rect 8208 12291 8260 12300
rect 4252 12180 4304 12232
rect 5356 12223 5408 12232
rect 5356 12189 5365 12223
rect 5365 12189 5399 12223
rect 5399 12189 5408 12223
rect 5356 12180 5408 12189
rect 8208 12257 8217 12291
rect 8217 12257 8251 12291
rect 8251 12257 8260 12291
rect 8208 12248 8260 12257
rect 9956 12248 10008 12300
rect 11612 12291 11664 12300
rect 8760 12180 8812 12232
rect 6920 12112 6972 12164
rect 7288 12112 7340 12164
rect 11612 12257 11621 12291
rect 11621 12257 11655 12291
rect 11655 12257 11664 12291
rect 11612 12248 11664 12257
rect 11704 12291 11756 12300
rect 11704 12257 11713 12291
rect 11713 12257 11747 12291
rect 11747 12257 11756 12291
rect 11704 12248 11756 12257
rect 12348 12248 12400 12300
rect 15568 12248 15620 12300
rect 16212 12291 16264 12300
rect 16212 12257 16221 12291
rect 16221 12257 16255 12291
rect 16255 12257 16264 12291
rect 16212 12248 16264 12257
rect 17500 12248 17552 12300
rect 11888 12223 11940 12232
rect 11888 12189 11897 12223
rect 11897 12189 11931 12223
rect 11931 12189 11940 12223
rect 11888 12180 11940 12189
rect 13360 12223 13412 12232
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 14464 12180 14516 12232
rect 13452 12112 13504 12164
rect 15660 12112 15712 12164
rect 15936 12112 15988 12164
rect 16856 12155 16908 12164
rect 16856 12121 16865 12155
rect 16865 12121 16899 12155
rect 16899 12121 16908 12155
rect 16856 12112 16908 12121
rect 17776 12112 17828 12164
rect 17960 12223 18012 12232
rect 17960 12189 17969 12223
rect 17969 12189 18003 12223
rect 18003 12189 18012 12223
rect 17960 12180 18012 12189
rect 2136 12044 2188 12096
rect 2780 12087 2832 12096
rect 2780 12053 2789 12087
rect 2789 12053 2823 12087
rect 2823 12053 2832 12087
rect 2780 12044 2832 12053
rect 3976 12044 4028 12096
rect 4252 12087 4304 12096
rect 4252 12053 4261 12087
rect 4261 12053 4295 12087
rect 4295 12053 4304 12087
rect 4252 12044 4304 12053
rect 4712 12087 4764 12096
rect 4712 12053 4721 12087
rect 4721 12053 4755 12087
rect 4755 12053 4764 12087
rect 4712 12044 4764 12053
rect 6000 12044 6052 12096
rect 6736 12087 6788 12096
rect 6736 12053 6745 12087
rect 6745 12053 6779 12087
rect 6779 12053 6788 12087
rect 6736 12044 6788 12053
rect 7472 12044 7524 12096
rect 9220 12044 9272 12096
rect 9588 12044 9640 12096
rect 9680 12044 9732 12096
rect 13360 12044 13412 12096
rect 15844 12087 15896 12096
rect 15844 12053 15853 12087
rect 15853 12053 15887 12087
rect 15887 12053 15896 12087
rect 15844 12044 15896 12053
rect 17408 12087 17460 12096
rect 17408 12053 17417 12087
rect 17417 12053 17451 12087
rect 17451 12053 17460 12087
rect 17408 12044 17460 12053
rect 18420 12087 18472 12096
rect 18420 12053 18429 12087
rect 18429 12053 18463 12087
rect 18463 12053 18472 12087
rect 18420 12044 18472 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1584 11883 1636 11892
rect 1584 11849 1593 11883
rect 1593 11849 1627 11883
rect 1627 11849 1636 11883
rect 1584 11840 1636 11849
rect 3976 11840 4028 11892
rect 4804 11883 4856 11892
rect 4804 11849 4813 11883
rect 4813 11849 4847 11883
rect 4847 11849 4856 11883
rect 4804 11840 4856 11849
rect 6184 11883 6236 11892
rect 6184 11849 6193 11883
rect 6193 11849 6227 11883
rect 6227 11849 6236 11883
rect 6184 11840 6236 11849
rect 8760 11883 8812 11892
rect 8760 11849 8769 11883
rect 8769 11849 8803 11883
rect 8803 11849 8812 11883
rect 8760 11840 8812 11849
rect 9312 11883 9364 11892
rect 9312 11849 9321 11883
rect 9321 11849 9355 11883
rect 9355 11849 9364 11883
rect 9312 11840 9364 11849
rect 11704 11840 11756 11892
rect 13912 11883 13964 11892
rect 13912 11849 13921 11883
rect 13921 11849 13955 11883
rect 13955 11849 13964 11883
rect 13912 11840 13964 11849
rect 14464 11883 14516 11892
rect 14464 11849 14473 11883
rect 14473 11849 14507 11883
rect 14507 11849 14516 11883
rect 14464 11840 14516 11849
rect 16488 11883 16540 11892
rect 16488 11849 16497 11883
rect 16497 11849 16531 11883
rect 16531 11849 16540 11883
rect 16488 11840 16540 11849
rect 17776 11883 17828 11892
rect 17776 11849 17785 11883
rect 17785 11849 17819 11883
rect 17819 11849 17828 11883
rect 17776 11840 17828 11849
rect 19156 11883 19208 11892
rect 5356 11772 5408 11824
rect 3424 11636 3476 11688
rect 4436 11636 4488 11688
rect 5264 11636 5316 11688
rect 11888 11772 11940 11824
rect 14556 11772 14608 11824
rect 16212 11772 16264 11824
rect 9864 11747 9916 11756
rect 9864 11713 9873 11747
rect 9873 11713 9907 11747
rect 9907 11713 9916 11747
rect 9864 11704 9916 11713
rect 15568 11747 15620 11756
rect 6184 11636 6236 11688
rect 6920 11636 6972 11688
rect 9680 11636 9732 11688
rect 11612 11636 11664 11688
rect 11888 11636 11940 11688
rect 2136 11500 2188 11552
rect 4252 11543 4304 11552
rect 4252 11509 4261 11543
rect 4261 11509 4295 11543
rect 4295 11509 4304 11543
rect 4252 11500 4304 11509
rect 5448 11500 5500 11552
rect 8208 11543 8260 11552
rect 8208 11509 8217 11543
rect 8217 11509 8251 11543
rect 8251 11509 8260 11543
rect 8208 11500 8260 11509
rect 10048 11568 10100 11620
rect 10968 11568 11020 11620
rect 14004 11636 14056 11688
rect 14740 11636 14792 11688
rect 15568 11713 15577 11747
rect 15577 11713 15611 11747
rect 15611 11713 15620 11747
rect 15568 11704 15620 11713
rect 19156 11849 19165 11883
rect 19165 11849 19199 11883
rect 19199 11849 19208 11883
rect 19156 11840 19208 11849
rect 17960 11636 18012 11688
rect 18420 11679 18472 11688
rect 18420 11645 18429 11679
rect 18429 11645 18463 11679
rect 18463 11645 18472 11679
rect 18420 11636 18472 11645
rect 10876 11500 10928 11552
rect 11336 11543 11388 11552
rect 11336 11509 11345 11543
rect 11345 11509 11379 11543
rect 11379 11509 11388 11543
rect 11336 11500 11388 11509
rect 12532 11500 12584 11552
rect 14740 11500 14792 11552
rect 18696 11568 18748 11620
rect 15016 11543 15068 11552
rect 15016 11509 15025 11543
rect 15025 11509 15059 11543
rect 15059 11509 15068 11543
rect 15016 11500 15068 11509
rect 15108 11500 15160 11552
rect 15752 11500 15804 11552
rect 17500 11543 17552 11552
rect 17500 11509 17509 11543
rect 17509 11509 17543 11543
rect 17543 11509 17552 11543
rect 17500 11500 17552 11509
rect 18052 11543 18104 11552
rect 18052 11509 18061 11543
rect 18061 11509 18095 11543
rect 18095 11509 18104 11543
rect 18052 11500 18104 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 2504 11296 2556 11348
rect 2596 11296 2648 11348
rect 2780 11296 2832 11348
rect 3884 11339 3936 11348
rect 3884 11305 3893 11339
rect 3893 11305 3927 11339
rect 3927 11305 3936 11339
rect 3884 11296 3936 11305
rect 3976 11296 4028 11348
rect 5264 11339 5316 11348
rect 5264 11305 5273 11339
rect 5273 11305 5307 11339
rect 5307 11305 5316 11339
rect 5264 11296 5316 11305
rect 6920 11296 6972 11348
rect 8300 11339 8352 11348
rect 8300 11305 8309 11339
rect 8309 11305 8343 11339
rect 8343 11305 8352 11339
rect 8300 11296 8352 11305
rect 8484 11296 8536 11348
rect 9864 11296 9916 11348
rect 9956 11339 10008 11348
rect 9956 11305 9965 11339
rect 9965 11305 9999 11339
rect 9999 11305 10008 11339
rect 9956 11296 10008 11305
rect 12532 11296 12584 11348
rect 12900 11339 12952 11348
rect 12900 11305 12909 11339
rect 12909 11305 12943 11339
rect 12943 11305 12952 11339
rect 12900 11296 12952 11305
rect 13360 11339 13412 11348
rect 13360 11305 13369 11339
rect 13369 11305 13403 11339
rect 13403 11305 13412 11339
rect 13360 11296 13412 11305
rect 15844 11296 15896 11348
rect 18052 11339 18104 11348
rect 18052 11305 18061 11339
rect 18061 11305 18095 11339
rect 18095 11305 18104 11339
rect 18052 11296 18104 11305
rect 2872 11228 2924 11280
rect 6000 11228 6052 11280
rect 6736 11228 6788 11280
rect 8208 11228 8260 11280
rect 11060 11228 11112 11280
rect 11336 11228 11388 11280
rect 13452 11228 13504 11280
rect 14648 11271 14700 11280
rect 14648 11237 14657 11271
rect 14657 11237 14691 11271
rect 14691 11237 14700 11271
rect 14648 11228 14700 11237
rect 17776 11228 17828 11280
rect 18512 11271 18564 11280
rect 18512 11237 18521 11271
rect 18521 11237 18555 11271
rect 18555 11237 18564 11271
rect 18512 11228 18564 11237
rect 2596 11160 2648 11212
rect 3884 11160 3936 11212
rect 4068 11203 4120 11212
rect 4068 11169 4077 11203
rect 4077 11169 4111 11203
rect 4111 11169 4120 11203
rect 4068 11160 4120 11169
rect 5356 11160 5408 11212
rect 1768 11092 1820 11144
rect 2872 11135 2924 11144
rect 2872 11101 2881 11135
rect 2881 11101 2915 11135
rect 2915 11101 2924 11135
rect 2872 11092 2924 11101
rect 3424 11092 3476 11144
rect 7288 11092 7340 11144
rect 9772 11160 9824 11212
rect 11888 11160 11940 11212
rect 13912 11160 13964 11212
rect 15660 11160 15712 11212
rect 18328 11160 18380 11212
rect 15016 11135 15068 11144
rect 8300 11024 8352 11076
rect 15016 11101 15025 11135
rect 15025 11101 15059 11135
rect 15059 11101 15068 11135
rect 15016 11092 15068 11101
rect 15476 11092 15528 11144
rect 18696 11135 18748 11144
rect 18696 11101 18705 11135
rect 18705 11101 18739 11135
rect 18739 11101 18748 11135
rect 18696 11092 18748 11101
rect 8576 11024 8628 11076
rect 13912 11067 13964 11076
rect 13912 11033 13921 11067
rect 13921 11033 13955 11067
rect 13955 11033 13964 11067
rect 13912 11024 13964 11033
rect 14280 11067 14332 11076
rect 14280 11033 14289 11067
rect 14289 11033 14323 11067
rect 14323 11033 14332 11067
rect 14280 11024 14332 11033
rect 4988 10999 5040 11008
rect 4988 10965 4997 10999
rect 4997 10965 5031 10999
rect 5031 10965 5040 10999
rect 4988 10956 5040 10965
rect 9956 10956 10008 11008
rect 10140 10956 10192 11008
rect 10784 10956 10836 11008
rect 13176 10956 13228 11008
rect 14648 10956 14700 11008
rect 15752 10956 15804 11008
rect 16212 10956 16264 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2596 10752 2648 10804
rect 3148 10795 3200 10804
rect 3148 10761 3157 10795
rect 3157 10761 3191 10795
rect 3191 10761 3200 10795
rect 3148 10752 3200 10761
rect 3332 10752 3384 10804
rect 4896 10752 4948 10804
rect 5448 10752 5500 10804
rect 6184 10795 6236 10804
rect 6184 10761 6193 10795
rect 6193 10761 6227 10795
rect 6227 10761 6236 10795
rect 6184 10752 6236 10761
rect 6828 10752 6880 10804
rect 9772 10795 9824 10804
rect 1860 10659 1912 10668
rect 1860 10625 1869 10659
rect 1869 10625 1903 10659
rect 1903 10625 1912 10659
rect 1860 10616 1912 10625
rect 2688 10616 2740 10668
rect 3884 10659 3936 10668
rect 3884 10625 3893 10659
rect 3893 10625 3927 10659
rect 3927 10625 3936 10659
rect 3884 10616 3936 10625
rect 6000 10616 6052 10668
rect 9772 10761 9781 10795
rect 9781 10761 9815 10795
rect 9815 10761 9824 10795
rect 9772 10752 9824 10761
rect 11060 10752 11112 10804
rect 13452 10795 13504 10804
rect 13452 10761 13461 10795
rect 13461 10761 13495 10795
rect 13495 10761 13504 10795
rect 13452 10752 13504 10761
rect 13544 10752 13596 10804
rect 16120 10752 16172 10804
rect 16672 10795 16724 10804
rect 16672 10761 16681 10795
rect 16681 10761 16715 10795
rect 16715 10761 16724 10795
rect 16672 10752 16724 10761
rect 17408 10752 17460 10804
rect 18604 10752 18656 10804
rect 9680 10684 9732 10736
rect 13820 10727 13872 10736
rect 13820 10693 13829 10727
rect 13829 10693 13863 10727
rect 13863 10693 13872 10727
rect 15476 10727 15528 10736
rect 13820 10684 13872 10693
rect 9312 10616 9364 10668
rect 10784 10616 10836 10668
rect 13176 10616 13228 10668
rect 14464 10659 14516 10668
rect 14464 10625 14473 10659
rect 14473 10625 14507 10659
rect 14507 10625 14516 10659
rect 14464 10616 14516 10625
rect 15476 10693 15485 10727
rect 15485 10693 15519 10727
rect 15519 10693 15528 10727
rect 15476 10684 15528 10693
rect 15936 10684 15988 10736
rect 16028 10659 16080 10668
rect 16028 10625 16037 10659
rect 16037 10625 16071 10659
rect 16071 10625 16080 10659
rect 16028 10616 16080 10625
rect 16120 10659 16172 10668
rect 16120 10625 16129 10659
rect 16129 10625 16163 10659
rect 16163 10625 16172 10659
rect 16120 10616 16172 10625
rect 17408 10616 17460 10668
rect 1400 10548 1452 10600
rect 4528 10548 4580 10600
rect 4988 10548 5040 10600
rect 5448 10548 5500 10600
rect 12164 10591 12216 10600
rect 12164 10557 12173 10591
rect 12173 10557 12207 10591
rect 12207 10557 12216 10591
rect 12164 10548 12216 10557
rect 14372 10591 14424 10600
rect 14372 10557 14381 10591
rect 14381 10557 14415 10591
rect 14415 10557 14424 10591
rect 14372 10548 14424 10557
rect 15844 10548 15896 10600
rect 848 10480 900 10532
rect 7288 10523 7340 10532
rect 7288 10489 7297 10523
rect 7297 10489 7331 10523
rect 7331 10489 7340 10523
rect 7288 10480 7340 10489
rect 8208 10480 8260 10532
rect 10600 10480 10652 10532
rect 13084 10480 13136 10532
rect 3884 10412 3936 10464
rect 4252 10455 4304 10464
rect 4252 10421 4261 10455
rect 4261 10421 4295 10455
rect 4295 10421 4304 10455
rect 4252 10412 4304 10421
rect 5264 10412 5316 10464
rect 9496 10412 9548 10464
rect 12716 10412 12768 10464
rect 15752 10412 15804 10464
rect 17776 10455 17828 10464
rect 17776 10421 17785 10455
rect 17785 10421 17819 10455
rect 17819 10421 17828 10455
rect 17776 10412 17828 10421
rect 18788 10412 18840 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1768 10251 1820 10260
rect 1768 10217 1777 10251
rect 1777 10217 1811 10251
rect 1811 10217 1820 10251
rect 1768 10208 1820 10217
rect 4160 10208 4212 10260
rect 4896 10251 4948 10260
rect 4896 10217 4905 10251
rect 4905 10217 4939 10251
rect 4939 10217 4948 10251
rect 4896 10208 4948 10217
rect 5448 10251 5500 10260
rect 5448 10217 5457 10251
rect 5457 10217 5491 10251
rect 5491 10217 5500 10251
rect 5448 10208 5500 10217
rect 7840 10251 7892 10260
rect 7840 10217 7849 10251
rect 7849 10217 7883 10251
rect 7883 10217 7892 10251
rect 7840 10208 7892 10217
rect 8300 10208 8352 10260
rect 4712 10140 4764 10192
rect 6000 10140 6052 10192
rect 5540 10072 5592 10124
rect 8300 10072 8352 10124
rect 9772 10208 9824 10260
rect 11060 10251 11112 10260
rect 11060 10217 11069 10251
rect 11069 10217 11103 10251
rect 11103 10217 11112 10251
rect 11060 10208 11112 10217
rect 12900 10208 12952 10260
rect 13820 10208 13872 10260
rect 14464 10208 14516 10260
rect 17408 10251 17460 10260
rect 17408 10217 17417 10251
rect 17417 10217 17451 10251
rect 17451 10217 17460 10251
rect 17408 10208 17460 10217
rect 18696 10208 18748 10260
rect 9680 10140 9732 10192
rect 12532 10183 12584 10192
rect 12532 10149 12541 10183
rect 12541 10149 12575 10183
rect 12575 10149 12584 10183
rect 12532 10140 12584 10149
rect 13084 10140 13136 10192
rect 14372 10183 14424 10192
rect 14372 10149 14381 10183
rect 14381 10149 14415 10183
rect 14415 10149 14424 10183
rect 14372 10140 14424 10149
rect 16120 10140 16172 10192
rect 1860 10047 1912 10056
rect 1860 10013 1869 10047
rect 1869 10013 1903 10047
rect 1903 10013 1912 10047
rect 1860 10004 1912 10013
rect 2044 10047 2096 10056
rect 2044 10013 2053 10047
rect 2053 10013 2087 10047
rect 2087 10013 2096 10047
rect 2044 10004 2096 10013
rect 3516 10004 3568 10056
rect 5356 10004 5408 10056
rect 7380 10004 7432 10056
rect 8484 10004 8536 10056
rect 9312 10004 9364 10056
rect 9772 10072 9824 10124
rect 12440 10072 12492 10124
rect 1400 9979 1452 9988
rect 1400 9945 1409 9979
rect 1409 9945 1443 9979
rect 1443 9945 1452 9979
rect 1400 9936 1452 9945
rect 8300 9936 8352 9988
rect 2412 9911 2464 9920
rect 2412 9877 2421 9911
rect 2421 9877 2455 9911
rect 2455 9877 2464 9911
rect 2412 9868 2464 9877
rect 3056 9911 3108 9920
rect 3056 9877 3065 9911
rect 3065 9877 3099 9911
rect 3099 9877 3108 9911
rect 3056 9868 3108 9877
rect 3884 9911 3936 9920
rect 3884 9877 3893 9911
rect 3893 9877 3927 9911
rect 3927 9877 3936 9911
rect 3884 9868 3936 9877
rect 5264 9911 5316 9920
rect 5264 9877 5273 9911
rect 5273 9877 5307 9911
rect 5307 9877 5316 9911
rect 5264 9868 5316 9877
rect 6920 9911 6972 9920
rect 6920 9877 6929 9911
rect 6929 9877 6963 9911
rect 6963 9877 6972 9911
rect 6920 9868 6972 9877
rect 8392 9868 8444 9920
rect 12900 10004 12952 10056
rect 13268 10047 13320 10056
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 13452 10047 13504 10056
rect 13452 10013 13461 10047
rect 13461 10013 13495 10047
rect 13495 10013 13504 10047
rect 13452 10004 13504 10013
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 18328 9936 18380 9988
rect 19248 9936 19300 9988
rect 10324 9868 10376 9920
rect 10968 9868 11020 9920
rect 15660 9911 15712 9920
rect 15660 9877 15669 9911
rect 15669 9877 15703 9911
rect 15703 9877 15712 9911
rect 15660 9868 15712 9877
rect 18788 9911 18840 9920
rect 18788 9877 18797 9911
rect 18797 9877 18831 9911
rect 18831 9877 18840 9911
rect 18788 9868 18840 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1768 9664 1820 9716
rect 5264 9664 5316 9716
rect 8484 9707 8536 9716
rect 8484 9673 8493 9707
rect 8493 9673 8527 9707
rect 8527 9673 8536 9707
rect 8484 9664 8536 9673
rect 10324 9664 10376 9716
rect 1860 9596 1912 9648
rect 5356 9596 5408 9648
rect 6644 9596 6696 9648
rect 8116 9639 8168 9648
rect 8116 9605 8125 9639
rect 8125 9605 8159 9639
rect 8159 9605 8168 9639
rect 8116 9596 8168 9605
rect 9588 9596 9640 9648
rect 10600 9639 10652 9648
rect 10600 9605 10609 9639
rect 10609 9605 10643 9639
rect 10643 9605 10652 9639
rect 10600 9596 10652 9605
rect 12900 9664 12952 9716
rect 15568 9596 15620 9648
rect 16304 9639 16356 9648
rect 16304 9605 16313 9639
rect 16313 9605 16347 9639
rect 16347 9605 16356 9639
rect 16304 9596 16356 9605
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 2136 9528 2188 9580
rect 3056 9571 3108 9580
rect 3056 9537 3065 9571
rect 3065 9537 3099 9571
rect 3099 9537 3108 9571
rect 3056 9528 3108 9537
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 1768 9503 1820 9512
rect 1768 9469 1777 9503
rect 1777 9469 1811 9503
rect 1811 9469 1820 9503
rect 1768 9460 1820 9469
rect 2412 9460 2464 9512
rect 2872 9460 2924 9512
rect 4068 9460 4120 9512
rect 6552 9460 6604 9512
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 8300 9528 8352 9580
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 9772 9528 9824 9580
rect 11888 9528 11940 9580
rect 16120 9528 16172 9580
rect 9680 9460 9732 9512
rect 10600 9460 10652 9512
rect 11980 9460 12032 9512
rect 6368 9392 6420 9444
rect 13452 9392 13504 9444
rect 13912 9392 13964 9444
rect 1584 9324 1636 9376
rect 4620 9324 4672 9376
rect 6000 9367 6052 9376
rect 6000 9333 6009 9367
rect 6009 9333 6043 9367
rect 6043 9333 6052 9367
rect 6000 9324 6052 9333
rect 6920 9324 6972 9376
rect 10784 9367 10836 9376
rect 10784 9333 10793 9367
rect 10793 9333 10827 9367
rect 10827 9333 10836 9367
rect 10784 9324 10836 9333
rect 10876 9324 10928 9376
rect 11704 9324 11756 9376
rect 12348 9324 12400 9376
rect 13360 9367 13412 9376
rect 13360 9333 13369 9367
rect 13369 9333 13403 9367
rect 13403 9333 13412 9367
rect 13360 9324 13412 9333
rect 13820 9324 13872 9376
rect 15752 9460 15804 9512
rect 16028 9324 16080 9376
rect 16672 9324 16724 9376
rect 17684 9367 17736 9376
rect 17684 9333 17693 9367
rect 17693 9333 17727 9367
rect 17727 9333 17736 9367
rect 17684 9324 17736 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2872 9163 2924 9172
rect 2872 9129 2881 9163
rect 2881 9129 2915 9163
rect 2915 9129 2924 9163
rect 2872 9120 2924 9129
rect 3516 9163 3568 9172
rect 3516 9129 3525 9163
rect 3525 9129 3559 9163
rect 3559 9129 3568 9163
rect 3516 9120 3568 9129
rect 4712 9120 4764 9172
rect 6460 9120 6512 9172
rect 6644 9120 6696 9172
rect 7748 9163 7800 9172
rect 7748 9129 7757 9163
rect 7757 9129 7791 9163
rect 7791 9129 7800 9163
rect 7748 9120 7800 9129
rect 8484 9120 8536 9172
rect 10784 9120 10836 9172
rect 12072 9120 12124 9172
rect 16120 9120 16172 9172
rect 4436 9095 4488 9104
rect 4436 9061 4445 9095
rect 4445 9061 4479 9095
rect 4479 9061 4488 9095
rect 4436 9052 4488 9061
rect 9680 9052 9732 9104
rect 10968 9052 11020 9104
rect 14924 9095 14976 9104
rect 14924 9061 14933 9095
rect 14933 9061 14967 9095
rect 14967 9061 14976 9095
rect 14924 9052 14976 9061
rect 17408 9052 17460 9104
rect 6460 8984 6512 9036
rect 7564 8984 7616 9036
rect 9956 8984 10008 9036
rect 11888 8984 11940 9036
rect 12348 8984 12400 9036
rect 16672 8984 16724 9036
rect 3332 8916 3384 8968
rect 3884 8959 3936 8968
rect 3884 8925 3893 8959
rect 3893 8925 3927 8959
rect 3927 8925 3936 8959
rect 4620 8959 4672 8968
rect 3884 8916 3936 8925
rect 4068 8891 4120 8900
rect 4068 8857 4077 8891
rect 4077 8857 4111 8891
rect 4111 8857 4120 8891
rect 4068 8848 4120 8857
rect 4620 8925 4629 8959
rect 4629 8925 4663 8959
rect 4663 8925 4672 8959
rect 4620 8916 4672 8925
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 11796 8959 11848 8968
rect 10232 8916 10284 8925
rect 11796 8925 11805 8959
rect 11805 8925 11839 8959
rect 11839 8925 11848 8959
rect 11796 8916 11848 8925
rect 15292 8916 15344 8968
rect 2136 8780 2188 8832
rect 5540 8780 5592 8832
rect 9312 8848 9364 8900
rect 7380 8780 7432 8832
rect 8392 8823 8444 8832
rect 8392 8789 8401 8823
rect 8401 8789 8435 8823
rect 8435 8789 8444 8823
rect 8392 8780 8444 8789
rect 10048 8780 10100 8832
rect 10876 8823 10928 8832
rect 10876 8789 10885 8823
rect 10885 8789 10919 8823
rect 10919 8789 10928 8823
rect 10876 8780 10928 8789
rect 11612 8823 11664 8832
rect 11612 8789 11621 8823
rect 11621 8789 11655 8823
rect 11655 8789 11664 8823
rect 11612 8780 11664 8789
rect 13176 8823 13228 8832
rect 13176 8789 13185 8823
rect 13185 8789 13219 8823
rect 13219 8789 13228 8823
rect 13176 8780 13228 8789
rect 13912 8823 13964 8832
rect 13912 8789 13921 8823
rect 13921 8789 13955 8823
rect 13955 8789 13964 8823
rect 13912 8780 13964 8789
rect 14188 8823 14240 8832
rect 14188 8789 14197 8823
rect 14197 8789 14231 8823
rect 14231 8789 14240 8823
rect 14188 8780 14240 8789
rect 14556 8823 14608 8832
rect 14556 8789 14565 8823
rect 14565 8789 14599 8823
rect 14599 8789 14608 8823
rect 14556 8780 14608 8789
rect 15660 8780 15712 8832
rect 16488 8780 16540 8832
rect 17960 8823 18012 8832
rect 17960 8789 17969 8823
rect 17969 8789 18003 8823
rect 18003 8789 18012 8823
rect 17960 8780 18012 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2320 8576 2372 8628
rect 6276 8576 6328 8628
rect 7564 8576 7616 8628
rect 10232 8576 10284 8628
rect 13912 8576 13964 8628
rect 15292 8619 15344 8628
rect 15292 8585 15301 8619
rect 15301 8585 15335 8619
rect 15335 8585 15344 8619
rect 15292 8576 15344 8585
rect 15476 8576 15528 8628
rect 15752 8619 15804 8628
rect 2228 8440 2280 8492
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 7380 8483 7432 8492
rect 7380 8449 7389 8483
rect 7389 8449 7423 8483
rect 7423 8449 7432 8483
rect 7380 8440 7432 8449
rect 10876 8440 10928 8492
rect 2136 8347 2188 8356
rect 2136 8313 2145 8347
rect 2145 8313 2179 8347
rect 2179 8313 2188 8347
rect 2136 8304 2188 8313
rect 4620 8304 4672 8356
rect 2596 8279 2648 8288
rect 2596 8245 2605 8279
rect 2605 8245 2639 8279
rect 2639 8245 2648 8279
rect 2596 8236 2648 8245
rect 3148 8279 3200 8288
rect 3148 8245 3157 8279
rect 3157 8245 3191 8279
rect 3191 8245 3200 8279
rect 3148 8236 3200 8245
rect 5540 8236 5592 8288
rect 7196 8415 7248 8424
rect 7196 8381 7205 8415
rect 7205 8381 7239 8415
rect 7239 8381 7248 8415
rect 7196 8372 7248 8381
rect 9404 8372 9456 8424
rect 7104 8304 7156 8356
rect 7472 8304 7524 8356
rect 8484 8304 8536 8356
rect 11428 8304 11480 8356
rect 11796 8304 11848 8356
rect 13820 8372 13872 8424
rect 15752 8585 15761 8619
rect 15761 8585 15795 8619
rect 15795 8585 15804 8619
rect 15752 8576 15804 8585
rect 17408 8576 17460 8628
rect 16212 8483 16264 8492
rect 16212 8449 16221 8483
rect 16221 8449 16255 8483
rect 16255 8449 16264 8483
rect 16212 8440 16264 8449
rect 16488 8440 16540 8492
rect 13176 8304 13228 8356
rect 17500 8347 17552 8356
rect 17500 8313 17509 8347
rect 17509 8313 17543 8347
rect 17543 8313 17552 8347
rect 17500 8304 17552 8313
rect 6460 8236 6512 8288
rect 6828 8236 6880 8288
rect 6920 8236 6972 8288
rect 12440 8236 12492 8288
rect 16672 8236 16724 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1768 8075 1820 8084
rect 1768 8041 1777 8075
rect 1777 8041 1811 8075
rect 1811 8041 1820 8075
rect 1768 8032 1820 8041
rect 2228 8032 2280 8084
rect 3148 8032 3200 8084
rect 7196 8032 7248 8084
rect 9680 8075 9732 8084
rect 9680 8041 9689 8075
rect 9689 8041 9723 8075
rect 9723 8041 9732 8075
rect 9680 8032 9732 8041
rect 11704 8075 11756 8084
rect 11704 8041 11713 8075
rect 11713 8041 11747 8075
rect 11747 8041 11756 8075
rect 11704 8032 11756 8041
rect 12072 8075 12124 8084
rect 12072 8041 12081 8075
rect 12081 8041 12115 8075
rect 12115 8041 12124 8075
rect 12072 8032 12124 8041
rect 13268 8075 13320 8084
rect 13268 8041 13277 8075
rect 13277 8041 13311 8075
rect 13311 8041 13320 8075
rect 13268 8032 13320 8041
rect 13360 8032 13412 8084
rect 16212 8032 16264 8084
rect 16764 8032 16816 8084
rect 17684 8075 17736 8084
rect 17684 8041 17693 8075
rect 17693 8041 17727 8075
rect 17727 8041 17736 8075
rect 17684 8032 17736 8041
rect 4712 8007 4764 8016
rect 4712 7973 4721 8007
rect 4721 7973 4755 8007
rect 4755 7973 4764 8007
rect 4712 7964 4764 7973
rect 1584 7828 1636 7880
rect 2044 7871 2096 7880
rect 2044 7837 2053 7871
rect 2053 7837 2087 7871
rect 2087 7837 2096 7871
rect 2044 7828 2096 7837
rect 4528 7828 4580 7880
rect 4988 7896 5040 7948
rect 5172 7964 5224 8016
rect 12716 7964 12768 8016
rect 6276 7939 6328 7948
rect 6276 7905 6285 7939
rect 6285 7905 6319 7939
rect 6319 7905 6328 7939
rect 6276 7896 6328 7905
rect 8116 7896 8168 7948
rect 8300 7896 8352 7948
rect 1860 7692 1912 7744
rect 3148 7735 3200 7744
rect 3148 7701 3157 7735
rect 3157 7701 3191 7735
rect 3191 7701 3200 7735
rect 3148 7692 3200 7701
rect 3516 7735 3568 7744
rect 3516 7701 3525 7735
rect 3525 7701 3559 7735
rect 3559 7701 3568 7735
rect 3516 7692 3568 7701
rect 4528 7692 4580 7744
rect 4620 7692 4672 7744
rect 9956 7896 10008 7948
rect 16488 7939 16540 7948
rect 16488 7905 16497 7939
rect 16497 7905 16531 7939
rect 16531 7905 16540 7939
rect 16488 7896 16540 7905
rect 18052 7939 18104 7948
rect 18052 7905 18061 7939
rect 18061 7905 18095 7939
rect 18095 7905 18104 7939
rect 18052 7896 18104 7905
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 10140 7871 10192 7880
rect 8576 7828 8628 7837
rect 10140 7837 10149 7871
rect 10149 7837 10183 7871
rect 10183 7837 10192 7871
rect 10140 7828 10192 7837
rect 8024 7803 8076 7812
rect 8024 7769 8033 7803
rect 8033 7769 8067 7803
rect 8067 7769 8076 7803
rect 8024 7760 8076 7769
rect 8484 7760 8536 7812
rect 9864 7760 9916 7812
rect 10784 7828 10836 7880
rect 11612 7828 11664 7880
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 12256 7828 12308 7837
rect 13176 7828 13228 7880
rect 13912 7871 13964 7880
rect 13912 7837 13921 7871
rect 13921 7837 13955 7871
rect 13955 7837 13964 7871
rect 13912 7828 13964 7837
rect 16396 7828 16448 7880
rect 18144 7871 18196 7880
rect 18144 7837 18153 7871
rect 18153 7837 18187 7871
rect 18187 7837 18196 7871
rect 18144 7828 18196 7837
rect 15568 7760 15620 7812
rect 16580 7760 16632 7812
rect 20076 7760 20128 7812
rect 6092 7692 6144 7744
rect 6920 7735 6972 7744
rect 6920 7701 6929 7735
rect 6929 7701 6963 7735
rect 6963 7701 6972 7735
rect 6920 7692 6972 7701
rect 7104 7692 7156 7744
rect 10876 7735 10928 7744
rect 10876 7701 10885 7735
rect 10885 7701 10919 7735
rect 10919 7701 10928 7735
rect 10876 7692 10928 7701
rect 11244 7735 11296 7744
rect 11244 7701 11253 7735
rect 11253 7701 11287 7735
rect 11287 7701 11296 7735
rect 11244 7692 11296 7701
rect 11336 7692 11388 7744
rect 15660 7692 15712 7744
rect 15752 7735 15804 7744
rect 15752 7701 15761 7735
rect 15761 7701 15795 7735
rect 15795 7701 15804 7735
rect 15752 7692 15804 7701
rect 16856 7692 16908 7744
rect 19984 7735 20036 7744
rect 19984 7701 19993 7735
rect 19993 7701 20027 7735
rect 20027 7701 20036 7735
rect 19984 7692 20036 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1400 7531 1452 7540
rect 1400 7497 1409 7531
rect 1409 7497 1443 7531
rect 1443 7497 1452 7531
rect 1400 7488 1452 7497
rect 4160 7488 4212 7540
rect 5172 7531 5224 7540
rect 4436 7420 4488 7472
rect 4712 7463 4764 7472
rect 4712 7429 4721 7463
rect 4721 7429 4755 7463
rect 4755 7429 4764 7463
rect 4712 7420 4764 7429
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 3516 7352 3568 7404
rect 4620 7352 4672 7404
rect 1952 7284 2004 7336
rect 5172 7497 5181 7531
rect 5181 7497 5215 7531
rect 5215 7497 5224 7531
rect 5172 7488 5224 7497
rect 7564 7488 7616 7540
rect 8484 7488 8536 7540
rect 10784 7531 10836 7540
rect 10784 7497 10793 7531
rect 10793 7497 10827 7531
rect 10827 7497 10836 7531
rect 10784 7488 10836 7497
rect 12256 7488 12308 7540
rect 13360 7488 13412 7540
rect 15660 7488 15712 7540
rect 16764 7531 16816 7540
rect 16764 7497 16773 7531
rect 16773 7497 16807 7531
rect 16807 7497 16816 7531
rect 16764 7488 16816 7497
rect 8576 7420 8628 7472
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 6092 7352 6144 7404
rect 10876 7352 10928 7404
rect 12440 7352 12492 7404
rect 13636 7352 13688 7404
rect 6000 7284 6052 7336
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 9680 7284 9732 7336
rect 11796 7284 11848 7336
rect 12808 7284 12860 7336
rect 13360 7284 13412 7336
rect 14096 7395 14148 7404
rect 14096 7361 14105 7395
rect 14105 7361 14139 7395
rect 14139 7361 14148 7395
rect 14280 7395 14332 7404
rect 14096 7352 14148 7361
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 15752 7352 15804 7404
rect 18144 7420 18196 7472
rect 16396 7395 16448 7404
rect 16396 7361 16405 7395
rect 16405 7361 16439 7395
rect 16439 7361 16448 7395
rect 16396 7352 16448 7361
rect 18696 7395 18748 7404
rect 18696 7361 18705 7395
rect 18705 7361 18739 7395
rect 18739 7361 18748 7395
rect 18696 7352 18748 7361
rect 19340 7352 19392 7404
rect 14556 7284 14608 7336
rect 15476 7284 15528 7336
rect 18052 7284 18104 7336
rect 18420 7327 18472 7336
rect 18420 7293 18429 7327
rect 18429 7293 18463 7327
rect 18463 7293 18472 7327
rect 18420 7284 18472 7293
rect 18604 7284 18656 7336
rect 19156 7284 19208 7336
rect 1492 7216 1544 7268
rect 3516 7216 3568 7268
rect 1584 7148 1636 7200
rect 3424 7191 3476 7200
rect 3424 7157 3433 7191
rect 3433 7157 3467 7191
rect 3467 7157 3476 7191
rect 3424 7148 3476 7157
rect 5172 7148 5224 7200
rect 6736 7216 6788 7268
rect 6276 7191 6328 7200
rect 6276 7157 6285 7191
rect 6285 7157 6319 7191
rect 6319 7157 6328 7191
rect 6276 7148 6328 7157
rect 6460 7148 6512 7200
rect 7104 7259 7156 7268
rect 7104 7225 7138 7259
rect 7138 7225 7156 7259
rect 7104 7216 7156 7225
rect 8300 7216 8352 7268
rect 10140 7216 10192 7268
rect 10784 7216 10836 7268
rect 11060 7216 11112 7268
rect 9956 7148 10008 7200
rect 17040 7216 17092 7268
rect 19984 7259 20036 7268
rect 19984 7225 19993 7259
rect 19993 7225 20027 7259
rect 20027 7225 20036 7259
rect 19984 7216 20036 7225
rect 20628 7216 20680 7268
rect 12348 7148 12400 7200
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 12440 7148 12492 7157
rect 16396 7148 16448 7200
rect 18328 7148 18380 7200
rect 19524 7148 19576 7200
rect 20076 7191 20128 7200
rect 20076 7157 20085 7191
rect 20085 7157 20119 7191
rect 20119 7157 20128 7191
rect 20076 7148 20128 7157
rect 20812 7148 20864 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1492 6944 1544 6996
rect 1952 6987 2004 6996
rect 1952 6953 1961 6987
rect 1961 6953 1995 6987
rect 1995 6953 2004 6987
rect 1952 6944 2004 6953
rect 2044 6944 2096 6996
rect 3148 6944 3200 6996
rect 3608 6944 3660 6996
rect 4436 6987 4488 6996
rect 4436 6953 4445 6987
rect 4445 6953 4479 6987
rect 4479 6953 4488 6987
rect 4436 6944 4488 6953
rect 4804 6944 4856 6996
rect 9312 6944 9364 6996
rect 9864 6987 9916 6996
rect 9864 6953 9873 6987
rect 9873 6953 9907 6987
rect 9907 6953 9916 6987
rect 9864 6944 9916 6953
rect 14096 6944 14148 6996
rect 16488 6944 16540 6996
rect 18420 6987 18472 6996
rect 18420 6953 18429 6987
rect 18429 6953 18463 6987
rect 18463 6953 18472 6987
rect 18420 6944 18472 6953
rect 18512 6944 18564 6996
rect 19064 6944 19116 6996
rect 4896 6876 4948 6928
rect 9220 6876 9272 6928
rect 11520 6876 11572 6928
rect 5448 6808 5500 6860
rect 5816 6808 5868 6860
rect 7656 6808 7708 6860
rect 8300 6808 8352 6860
rect 8484 6851 8536 6860
rect 8484 6817 8493 6851
rect 8493 6817 8527 6851
rect 8527 6817 8536 6851
rect 8484 6808 8536 6817
rect 8668 6808 8720 6860
rect 9588 6808 9640 6860
rect 13452 6808 13504 6860
rect 13912 6808 13964 6860
rect 14096 6808 14148 6860
rect 16488 6808 16540 6860
rect 18788 6808 18840 6860
rect 22284 6851 22336 6860
rect 22284 6817 22293 6851
rect 22293 6817 22327 6851
rect 22327 6817 22336 6851
rect 22284 6808 22336 6817
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 4528 6783 4580 6792
rect 4528 6749 4537 6783
rect 4537 6749 4571 6783
rect 4571 6749 4580 6783
rect 4528 6740 4580 6749
rect 6000 6783 6052 6792
rect 4160 6672 4212 6724
rect 5172 6715 5224 6724
rect 5172 6681 5181 6715
rect 5181 6681 5215 6715
rect 5215 6681 5224 6715
rect 5172 6672 5224 6681
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 11060 6740 11112 6792
rect 11612 6783 11664 6792
rect 11612 6749 11621 6783
rect 11621 6749 11655 6783
rect 11655 6749 11664 6783
rect 11612 6740 11664 6749
rect 13084 6783 13136 6792
rect 13084 6749 13093 6783
rect 13093 6749 13127 6783
rect 13127 6749 13136 6783
rect 13084 6740 13136 6749
rect 13636 6740 13688 6792
rect 9680 6672 9732 6724
rect 10876 6672 10928 6724
rect 12900 6672 12952 6724
rect 13820 6672 13872 6724
rect 2228 6647 2280 6656
rect 2228 6613 2237 6647
rect 2237 6613 2271 6647
rect 2271 6613 2280 6647
rect 2228 6604 2280 6613
rect 2688 6604 2740 6656
rect 3516 6604 3568 6656
rect 4068 6647 4120 6656
rect 4068 6613 4077 6647
rect 4077 6613 4111 6647
rect 4111 6613 4120 6647
rect 4068 6604 4120 6613
rect 5264 6604 5316 6656
rect 7104 6604 7156 6656
rect 8944 6647 8996 6656
rect 8944 6613 8953 6647
rect 8953 6613 8987 6647
rect 8987 6613 8996 6647
rect 8944 6604 8996 6613
rect 9312 6647 9364 6656
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 9312 6604 9364 6613
rect 10232 6647 10284 6656
rect 10232 6613 10241 6647
rect 10241 6613 10275 6647
rect 10275 6613 10284 6647
rect 10232 6604 10284 6613
rect 12256 6604 12308 6656
rect 12624 6647 12676 6656
rect 12624 6613 12633 6647
rect 12633 6613 12667 6647
rect 12667 6613 12676 6647
rect 12624 6604 12676 6613
rect 14372 6647 14424 6656
rect 14372 6613 14381 6647
rect 14381 6613 14415 6647
rect 14415 6613 14424 6647
rect 14372 6604 14424 6613
rect 14648 6647 14700 6656
rect 14648 6613 14657 6647
rect 14657 6613 14691 6647
rect 14691 6613 14700 6647
rect 14648 6604 14700 6613
rect 19432 6783 19484 6792
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 21640 6672 21692 6724
rect 16580 6604 16632 6656
rect 17776 6647 17828 6656
rect 17776 6613 17785 6647
rect 17785 6613 17819 6647
rect 17819 6613 17828 6647
rect 17776 6604 17828 6613
rect 18696 6647 18748 6656
rect 18696 6613 18705 6647
rect 18705 6613 18739 6647
rect 18739 6613 18748 6647
rect 18696 6604 18748 6613
rect 20260 6647 20312 6656
rect 20260 6613 20269 6647
rect 20269 6613 20303 6647
rect 20303 6613 20312 6647
rect 20260 6604 20312 6613
rect 21548 6647 21600 6656
rect 21548 6613 21557 6647
rect 21557 6613 21591 6647
rect 21591 6613 21600 6647
rect 21548 6604 21600 6613
rect 22468 6647 22520 6656
rect 22468 6613 22477 6647
rect 22477 6613 22511 6647
rect 22511 6613 22520 6647
rect 22468 6604 22520 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 2044 6400 2096 6452
rect 2136 6443 2188 6452
rect 2136 6409 2145 6443
rect 2145 6409 2179 6443
rect 2179 6409 2188 6443
rect 2136 6400 2188 6409
rect 5448 6400 5500 6452
rect 6000 6400 6052 6452
rect 6460 6400 6512 6452
rect 6828 6443 6880 6452
rect 6828 6409 6837 6443
rect 6837 6409 6871 6443
rect 6871 6409 6880 6443
rect 6828 6400 6880 6409
rect 7564 6400 7616 6452
rect 8300 6443 8352 6452
rect 8300 6409 8309 6443
rect 8309 6409 8343 6443
rect 8343 6409 8352 6443
rect 8300 6400 8352 6409
rect 8576 6443 8628 6452
rect 8576 6409 8585 6443
rect 8585 6409 8619 6443
rect 8619 6409 8628 6443
rect 8576 6400 8628 6409
rect 9404 6443 9456 6452
rect 9404 6409 9413 6443
rect 9413 6409 9447 6443
rect 9447 6409 9456 6443
rect 9404 6400 9456 6409
rect 11888 6400 11940 6452
rect 16672 6400 16724 6452
rect 17684 6400 17736 6452
rect 18052 6443 18104 6452
rect 18052 6409 18061 6443
rect 18061 6409 18095 6443
rect 18095 6409 18104 6443
rect 18052 6400 18104 6409
rect 19064 6443 19116 6452
rect 19064 6409 19073 6443
rect 19073 6409 19107 6443
rect 19107 6409 19116 6443
rect 19064 6400 19116 6409
rect 20720 6400 20772 6452
rect 22284 6443 22336 6452
rect 22284 6409 22293 6443
rect 22293 6409 22327 6443
rect 22327 6409 22336 6443
rect 22284 6400 22336 6409
rect 5264 6307 5316 6316
rect 5264 6273 5273 6307
rect 5273 6273 5307 6307
rect 5307 6273 5316 6307
rect 5264 6264 5316 6273
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 3056 6196 3108 6248
rect 7196 6239 7248 6248
rect 7196 6205 7205 6239
rect 7205 6205 7239 6239
rect 7239 6205 7248 6239
rect 7196 6196 7248 6205
rect 10692 6196 10744 6248
rect 13636 6332 13688 6384
rect 19432 6332 19484 6384
rect 2872 6128 2924 6180
rect 5448 6128 5500 6180
rect 11060 6128 11112 6180
rect 12624 6196 12676 6248
rect 16672 6264 16724 6316
rect 18512 6264 18564 6316
rect 19248 6264 19300 6316
rect 20536 6264 20588 6316
rect 21640 6307 21692 6316
rect 21640 6273 21649 6307
rect 21649 6273 21683 6307
rect 21683 6273 21692 6307
rect 21640 6264 21692 6273
rect 14832 6196 14884 6248
rect 16488 6196 16540 6248
rect 16764 6239 16816 6248
rect 16764 6205 16773 6239
rect 16773 6205 16807 6239
rect 16807 6205 16816 6239
rect 16764 6196 16816 6205
rect 17684 6196 17736 6248
rect 19984 6239 20036 6248
rect 19984 6205 19993 6239
rect 19993 6205 20027 6239
rect 20027 6205 20036 6239
rect 19984 6196 20036 6205
rect 3056 6060 3108 6112
rect 4528 6103 4580 6112
rect 4528 6069 4537 6103
rect 4537 6069 4571 6103
rect 4571 6069 4580 6103
rect 4528 6060 4580 6069
rect 9864 6060 9916 6112
rect 11520 6103 11572 6112
rect 11520 6069 11529 6103
rect 11529 6069 11563 6103
rect 11563 6069 11572 6103
rect 11520 6060 11572 6069
rect 12440 6103 12492 6112
rect 12440 6069 12449 6103
rect 12449 6069 12483 6103
rect 12483 6069 12492 6103
rect 12900 6103 12952 6112
rect 12440 6060 12492 6069
rect 12900 6069 12909 6103
rect 12909 6069 12943 6103
rect 12943 6069 12952 6103
rect 12900 6060 12952 6069
rect 13452 6103 13504 6112
rect 13452 6069 13461 6103
rect 13461 6069 13495 6103
rect 13495 6069 13504 6103
rect 13452 6060 13504 6069
rect 17040 6128 17092 6180
rect 21548 6171 21600 6180
rect 16580 6060 16632 6112
rect 16948 6103 17000 6112
rect 16948 6069 16957 6103
rect 16957 6069 16991 6103
rect 16991 6069 17000 6103
rect 16948 6060 17000 6069
rect 21548 6137 21557 6171
rect 21557 6137 21591 6171
rect 21591 6137 21600 6171
rect 21548 6128 21600 6137
rect 20996 6103 21048 6112
rect 20996 6069 21005 6103
rect 21005 6069 21039 6103
rect 21039 6069 21048 6103
rect 20996 6060 21048 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 3608 5856 3660 5908
rect 5264 5856 5316 5908
rect 7288 5856 7340 5908
rect 7656 5899 7708 5908
rect 7656 5865 7665 5899
rect 7665 5865 7699 5899
rect 7699 5865 7708 5899
rect 7656 5856 7708 5865
rect 8300 5899 8352 5908
rect 8300 5865 8309 5899
rect 8309 5865 8343 5899
rect 8343 5865 8352 5899
rect 8300 5856 8352 5865
rect 11060 5899 11112 5908
rect 11060 5865 11069 5899
rect 11069 5865 11103 5899
rect 11103 5865 11112 5899
rect 11060 5856 11112 5865
rect 11612 5899 11664 5908
rect 11612 5865 11621 5899
rect 11621 5865 11655 5899
rect 11655 5865 11664 5899
rect 11612 5856 11664 5865
rect 12624 5856 12676 5908
rect 14832 5856 14884 5908
rect 15660 5856 15712 5908
rect 16672 5899 16724 5908
rect 16672 5865 16681 5899
rect 16681 5865 16715 5899
rect 16715 5865 16724 5899
rect 16672 5856 16724 5865
rect 19984 5899 20036 5908
rect 19984 5865 19993 5899
rect 19993 5865 20027 5899
rect 20027 5865 20036 5899
rect 19984 5856 20036 5865
rect 20536 5899 20588 5908
rect 20536 5865 20545 5899
rect 20545 5865 20579 5899
rect 20579 5865 20588 5899
rect 20536 5856 20588 5865
rect 20812 5856 20864 5908
rect 21364 5899 21416 5908
rect 21364 5865 21373 5899
rect 21373 5865 21407 5899
rect 21407 5865 21416 5899
rect 21364 5856 21416 5865
rect 2044 5788 2096 5840
rect 6828 5788 6880 5840
rect 9312 5788 9364 5840
rect 2136 5720 2188 5772
rect 4160 5720 4212 5772
rect 4620 5720 4672 5772
rect 7564 5720 7616 5772
rect 8576 5763 8628 5772
rect 8576 5729 8585 5763
rect 8585 5729 8619 5763
rect 8619 5729 8628 5763
rect 8576 5720 8628 5729
rect 9220 5720 9272 5772
rect 9404 5720 9456 5772
rect 9956 5763 10008 5772
rect 9956 5729 9990 5763
rect 9990 5729 10008 5763
rect 9956 5720 10008 5729
rect 12072 5720 12124 5772
rect 12440 5763 12492 5772
rect 12440 5729 12474 5763
rect 12474 5729 12492 5763
rect 12440 5720 12492 5729
rect 15568 5720 15620 5772
rect 17776 5788 17828 5840
rect 16580 5720 16632 5772
rect 17408 5720 17460 5772
rect 19340 5763 19392 5772
rect 19340 5729 19349 5763
rect 19349 5729 19383 5763
rect 19383 5729 19392 5763
rect 19340 5720 19392 5729
rect 21272 5763 21324 5772
rect 21272 5729 21281 5763
rect 21281 5729 21315 5763
rect 21315 5729 21324 5763
rect 21272 5720 21324 5729
rect 22468 5720 22520 5772
rect 23296 5763 23348 5772
rect 23296 5729 23305 5763
rect 23305 5729 23339 5763
rect 23339 5729 23348 5763
rect 23296 5720 23348 5729
rect 7104 5695 7156 5704
rect 7104 5661 7113 5695
rect 7113 5661 7147 5695
rect 7147 5661 7156 5695
rect 15936 5695 15988 5704
rect 7104 5652 7156 5661
rect 15936 5661 15945 5695
rect 15945 5661 15979 5695
rect 15979 5661 15988 5695
rect 15936 5652 15988 5661
rect 20996 5652 21048 5704
rect 2412 5584 2464 5636
rect 2872 5584 2924 5636
rect 9404 5627 9456 5636
rect 3700 5559 3752 5568
rect 3700 5525 3709 5559
rect 3709 5525 3743 5559
rect 3743 5525 3752 5559
rect 3700 5516 3752 5525
rect 3884 5516 3936 5568
rect 9404 5593 9413 5627
rect 9413 5593 9447 5627
rect 9447 5593 9456 5627
rect 9404 5584 9456 5593
rect 13912 5584 13964 5636
rect 14096 5584 14148 5636
rect 16580 5584 16632 5636
rect 20812 5584 20864 5636
rect 7656 5516 7708 5568
rect 13636 5516 13688 5568
rect 14740 5516 14792 5568
rect 16396 5559 16448 5568
rect 16396 5525 16405 5559
rect 16405 5525 16439 5559
rect 16439 5525 16448 5559
rect 16396 5516 16448 5525
rect 18144 5516 18196 5568
rect 18788 5516 18840 5568
rect 23480 5559 23532 5568
rect 23480 5525 23489 5559
rect 23489 5525 23523 5559
rect 23523 5525 23532 5559
rect 23480 5516 23532 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 4160 5312 4212 5364
rect 9956 5312 10008 5364
rect 10692 5355 10744 5364
rect 10692 5321 10701 5355
rect 10701 5321 10735 5355
rect 10735 5321 10744 5355
rect 10692 5312 10744 5321
rect 11060 5312 11112 5364
rect 11244 5312 11296 5364
rect 12072 5312 12124 5364
rect 2872 5244 2924 5296
rect 4068 5244 4120 5296
rect 9220 5287 9272 5296
rect 1860 5219 1912 5228
rect 1860 5185 1869 5219
rect 1869 5185 1903 5219
rect 1903 5185 1912 5219
rect 1860 5176 1912 5185
rect 2412 5176 2464 5228
rect 3700 5176 3752 5228
rect 9220 5253 9229 5287
rect 9229 5253 9263 5287
rect 9263 5253 9272 5287
rect 12440 5312 12492 5364
rect 14832 5312 14884 5364
rect 15936 5355 15988 5364
rect 15936 5321 15945 5355
rect 15945 5321 15979 5355
rect 15979 5321 15988 5355
rect 15936 5312 15988 5321
rect 16488 5312 16540 5364
rect 19432 5355 19484 5364
rect 19432 5321 19441 5355
rect 19441 5321 19475 5355
rect 19475 5321 19484 5355
rect 19432 5312 19484 5321
rect 21364 5312 21416 5364
rect 23296 5355 23348 5364
rect 23296 5321 23305 5355
rect 23305 5321 23339 5355
rect 23339 5321 23348 5355
rect 23296 5312 23348 5321
rect 9220 5244 9272 5253
rect 11244 5219 11296 5228
rect 1400 5108 1452 5160
rect 3056 5108 3108 5160
rect 4620 5108 4672 5160
rect 5356 5108 5408 5160
rect 5540 5108 5592 5160
rect 6460 5108 6512 5160
rect 11244 5185 11253 5219
rect 11253 5185 11287 5219
rect 11287 5185 11296 5219
rect 11244 5176 11296 5185
rect 19340 5244 19392 5296
rect 17868 5176 17920 5228
rect 20536 5176 20588 5228
rect 9404 5108 9456 5160
rect 12348 5108 12400 5160
rect 12624 5108 12676 5160
rect 16856 5151 16908 5160
rect 16856 5117 16865 5151
rect 16865 5117 16899 5151
rect 16899 5117 16908 5151
rect 16856 5108 16908 5117
rect 17408 5151 17460 5160
rect 17408 5117 17417 5151
rect 17417 5117 17451 5151
rect 17451 5117 17460 5151
rect 17408 5108 17460 5117
rect 5632 5083 5684 5092
rect 5632 5049 5641 5083
rect 5641 5049 5675 5083
rect 5675 5049 5684 5083
rect 5632 5040 5684 5049
rect 6276 5083 6328 5092
rect 6276 5049 6285 5083
rect 6285 5049 6319 5083
rect 6319 5049 6328 5083
rect 6276 5040 6328 5049
rect 11612 5083 11664 5092
rect 11612 5049 11621 5083
rect 11621 5049 11655 5083
rect 11655 5049 11664 5083
rect 11612 5040 11664 5049
rect 13636 5040 13688 5092
rect 16580 5040 16632 5092
rect 17500 5040 17552 5092
rect 18144 5108 18196 5160
rect 20996 5108 21048 5160
rect 22192 5108 22244 5160
rect 18420 5040 18472 5092
rect 3700 4972 3752 5024
rect 4160 4972 4212 5024
rect 4712 4972 4764 5024
rect 5172 5015 5224 5024
rect 5172 4981 5181 5015
rect 5181 4981 5215 5015
rect 5215 4981 5224 5015
rect 5172 4972 5224 4981
rect 5540 5015 5592 5024
rect 5540 4981 5549 5015
rect 5549 4981 5583 5015
rect 5583 4981 5592 5015
rect 5540 4972 5592 4981
rect 7748 4972 7800 5024
rect 12440 4972 12492 5024
rect 19432 4972 19484 5024
rect 20536 5015 20588 5024
rect 20536 4981 20545 5015
rect 20545 4981 20579 5015
rect 20579 4981 20588 5015
rect 20536 4972 20588 4981
rect 20720 4972 20772 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 2136 4768 2188 4820
rect 2872 4768 2924 4820
rect 5172 4768 5224 4820
rect 5540 4768 5592 4820
rect 6368 4811 6420 4820
rect 6368 4777 6377 4811
rect 6377 4777 6411 4811
rect 6411 4777 6420 4811
rect 6368 4768 6420 4777
rect 7104 4811 7156 4820
rect 7104 4777 7113 4811
rect 7113 4777 7147 4811
rect 7147 4777 7156 4811
rect 7104 4768 7156 4777
rect 7564 4811 7616 4820
rect 7564 4777 7573 4811
rect 7573 4777 7607 4811
rect 7607 4777 7616 4811
rect 7564 4768 7616 4777
rect 8024 4811 8076 4820
rect 8024 4777 8033 4811
rect 8033 4777 8067 4811
rect 8067 4777 8076 4811
rect 8024 4768 8076 4777
rect 8944 4811 8996 4820
rect 8944 4777 8953 4811
rect 8953 4777 8987 4811
rect 8987 4777 8996 4811
rect 8944 4768 8996 4777
rect 9036 4768 9088 4820
rect 9220 4768 9272 4820
rect 10968 4811 11020 4820
rect 10968 4777 10977 4811
rect 10977 4777 11011 4811
rect 11011 4777 11020 4811
rect 10968 4768 11020 4777
rect 11796 4768 11848 4820
rect 12808 4768 12860 4820
rect 13728 4768 13780 4820
rect 15476 4811 15528 4820
rect 15476 4777 15485 4811
rect 15485 4777 15519 4811
rect 15519 4777 15528 4811
rect 15476 4768 15528 4777
rect 15936 4768 15988 4820
rect 2688 4700 2740 4752
rect 5448 4700 5500 4752
rect 6000 4700 6052 4752
rect 10784 4743 10836 4752
rect 10784 4709 10793 4743
rect 10793 4709 10827 4743
rect 10827 4709 10836 4743
rect 10784 4700 10836 4709
rect 11980 4700 12032 4752
rect 12256 4700 12308 4752
rect 14832 4700 14884 4752
rect 17224 4768 17276 4820
rect 17868 4811 17920 4820
rect 17868 4777 17877 4811
rect 17877 4777 17911 4811
rect 17911 4777 17920 4811
rect 17868 4768 17920 4777
rect 19340 4768 19392 4820
rect 16672 4700 16724 4752
rect 2872 4675 2924 4684
rect 2872 4641 2881 4675
rect 2881 4641 2915 4675
rect 2915 4641 2924 4675
rect 2872 4632 2924 4641
rect 4436 4632 4488 4684
rect 3056 4607 3108 4616
rect 3056 4573 3065 4607
rect 3065 4573 3099 4607
rect 3099 4573 3108 4607
rect 3056 4564 3108 4573
rect 4160 4564 4212 4616
rect 5356 4564 5408 4616
rect 5632 4632 5684 4684
rect 7196 4632 7248 4684
rect 4068 4496 4120 4548
rect 5540 4496 5592 4548
rect 2320 4471 2372 4480
rect 2320 4437 2329 4471
rect 2329 4437 2363 4471
rect 2363 4437 2372 4471
rect 2320 4428 2372 4437
rect 2872 4428 2924 4480
rect 4344 4471 4396 4480
rect 4344 4437 4353 4471
rect 4353 4437 4387 4471
rect 4387 4437 4396 4471
rect 4344 4428 4396 4437
rect 6828 4496 6880 4548
rect 7564 4496 7616 4548
rect 7932 4496 7984 4548
rect 10784 4564 10836 4616
rect 11520 4564 11572 4616
rect 13268 4632 13320 4684
rect 13636 4675 13688 4684
rect 13636 4641 13645 4675
rect 13645 4641 13679 4675
rect 13679 4641 13688 4675
rect 13636 4632 13688 4641
rect 14096 4675 14148 4684
rect 14096 4641 14105 4675
rect 14105 4641 14139 4675
rect 14139 4641 14148 4675
rect 14096 4632 14148 4641
rect 15384 4632 15436 4684
rect 16304 4632 16356 4684
rect 17040 4632 17092 4684
rect 18052 4700 18104 4752
rect 13176 4607 13228 4616
rect 13176 4573 13185 4607
rect 13185 4573 13219 4607
rect 13219 4573 13228 4607
rect 13176 4564 13228 4573
rect 16948 4607 17000 4616
rect 16948 4573 16957 4607
rect 16957 4573 16991 4607
rect 16991 4573 17000 4607
rect 16948 4564 17000 4573
rect 8668 4539 8720 4548
rect 8668 4505 8677 4539
rect 8677 4505 8711 4539
rect 8711 4505 8720 4539
rect 8668 4496 8720 4505
rect 9772 4496 9824 4548
rect 16396 4496 16448 4548
rect 18144 4564 18196 4616
rect 19340 4632 19392 4684
rect 20536 4768 20588 4820
rect 21272 4768 21324 4820
rect 20904 4675 20956 4684
rect 20904 4641 20913 4675
rect 20913 4641 20947 4675
rect 20947 4641 20956 4675
rect 20904 4632 20956 4641
rect 19432 4564 19484 4616
rect 20720 4564 20772 4616
rect 17960 4496 18012 4548
rect 20260 4496 20312 4548
rect 6276 4428 6328 4480
rect 7748 4428 7800 4480
rect 10140 4471 10192 4480
rect 10140 4437 10149 4471
rect 10149 4437 10183 4471
rect 10183 4437 10192 4471
rect 10140 4428 10192 4437
rect 12532 4471 12584 4480
rect 12532 4437 12541 4471
rect 12541 4437 12575 4471
rect 12575 4437 12584 4471
rect 12532 4428 12584 4437
rect 13820 4428 13872 4480
rect 14280 4471 14332 4480
rect 14280 4437 14289 4471
rect 14289 4437 14323 4471
rect 14323 4437 14332 4471
rect 14280 4428 14332 4437
rect 16488 4471 16540 4480
rect 16488 4437 16497 4471
rect 16497 4437 16531 4471
rect 16531 4437 16540 4471
rect 16488 4428 16540 4437
rect 19800 4471 19852 4480
rect 19800 4437 19809 4471
rect 19809 4437 19843 4471
rect 19843 4437 19852 4471
rect 19800 4428 19852 4437
rect 20076 4428 20128 4480
rect 20720 4428 20772 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 4160 4224 4212 4276
rect 6000 4267 6052 4276
rect 6000 4233 6009 4267
rect 6009 4233 6043 4267
rect 6043 4233 6052 4267
rect 6000 4224 6052 4233
rect 6368 4267 6420 4276
rect 6368 4233 6377 4267
rect 6377 4233 6411 4267
rect 6411 4233 6420 4267
rect 6368 4224 6420 4233
rect 8024 4224 8076 4276
rect 2320 4156 2372 4208
rect 1768 4131 1820 4140
rect 1768 4097 1777 4131
rect 1777 4097 1811 4131
rect 1811 4097 1820 4131
rect 1768 4088 1820 4097
rect 2688 4088 2740 4140
rect 3056 4088 3108 4140
rect 8208 4088 8260 4140
rect 8668 4156 8720 4208
rect 3792 4020 3844 4072
rect 7196 4020 7248 4072
rect 7748 4020 7800 4072
rect 9956 4088 10008 4140
rect 11520 4224 11572 4276
rect 11980 4224 12032 4276
rect 12624 4224 12676 4276
rect 11796 4156 11848 4208
rect 12532 4156 12584 4208
rect 14096 4224 14148 4276
rect 15384 4267 15436 4276
rect 15384 4233 15393 4267
rect 15393 4233 15427 4267
rect 15427 4233 15436 4267
rect 15384 4224 15436 4233
rect 16856 4224 16908 4276
rect 18052 4267 18104 4276
rect 18052 4233 18061 4267
rect 18061 4233 18095 4267
rect 18095 4233 18104 4267
rect 18052 4224 18104 4233
rect 20904 4267 20956 4276
rect 20904 4233 20913 4267
rect 20913 4233 20947 4267
rect 20947 4233 20956 4267
rect 20904 4224 20956 4233
rect 9220 4020 9272 4072
rect 10692 4020 10744 4072
rect 11244 4063 11296 4072
rect 11244 4029 11253 4063
rect 11253 4029 11287 4063
rect 11287 4029 11296 4063
rect 11244 4020 11296 4029
rect 2228 3952 2280 4004
rect 4344 3952 4396 4004
rect 5448 3952 5500 4004
rect 8024 3952 8076 4004
rect 8300 3952 8352 4004
rect 9312 3995 9364 4004
rect 9312 3961 9321 3995
rect 9321 3961 9355 3995
rect 9355 3961 9364 3995
rect 9312 3952 9364 3961
rect 11520 3952 11572 4004
rect 12716 4088 12768 4140
rect 12992 4088 13044 4140
rect 13268 4088 13320 4140
rect 15936 4156 15988 4208
rect 13544 4020 13596 4072
rect 14096 4088 14148 4140
rect 16028 4131 16080 4140
rect 16028 4097 16037 4131
rect 16037 4097 16071 4131
rect 16071 4097 16080 4131
rect 16028 4088 16080 4097
rect 16396 4088 16448 4140
rect 16948 4156 17000 4208
rect 18052 4088 18104 4140
rect 18512 4088 18564 4140
rect 20076 4156 20128 4208
rect 19156 4131 19208 4140
rect 19156 4097 19165 4131
rect 19165 4097 19199 4131
rect 19199 4097 19208 4131
rect 19156 4088 19208 4097
rect 14740 4020 14792 4072
rect 16488 4020 16540 4072
rect 19432 4020 19484 4072
rect 21088 4020 21140 4072
rect 22284 4063 22336 4072
rect 22284 4029 22293 4063
rect 22293 4029 22327 4063
rect 22327 4029 22336 4063
rect 22284 4020 22336 4029
rect 13728 3952 13780 4004
rect 14832 3952 14884 4004
rect 19340 3952 19392 4004
rect 2320 3927 2372 3936
rect 2320 3893 2329 3927
rect 2329 3893 2363 3927
rect 2363 3893 2372 3927
rect 2320 3884 2372 3893
rect 2688 3927 2740 3936
rect 2688 3893 2697 3927
rect 2697 3893 2731 3927
rect 2731 3893 2740 3927
rect 2688 3884 2740 3893
rect 4620 3884 4672 3936
rect 5356 3884 5408 3936
rect 6552 3884 6604 3936
rect 7932 3884 7984 3936
rect 9404 3927 9456 3936
rect 9404 3893 9413 3927
rect 9413 3893 9447 3927
rect 9447 3893 9456 3927
rect 9404 3884 9456 3893
rect 11428 3927 11480 3936
rect 11428 3893 11437 3927
rect 11437 3893 11471 3927
rect 11471 3893 11480 3927
rect 11428 3884 11480 3893
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 12440 3884 12492 3893
rect 12808 3884 12860 3936
rect 13452 3884 13504 3936
rect 16396 3884 16448 3936
rect 17408 3927 17460 3936
rect 17408 3893 17417 3927
rect 17417 3893 17451 3927
rect 17451 3893 17460 3927
rect 17408 3884 17460 3893
rect 17776 3927 17828 3936
rect 17776 3893 17785 3927
rect 17785 3893 17819 3927
rect 17819 3893 17828 3927
rect 17776 3884 17828 3893
rect 19432 3927 19484 3936
rect 19432 3893 19441 3927
rect 19441 3893 19475 3927
rect 19475 3893 19484 3927
rect 19432 3884 19484 3893
rect 20168 3952 20220 4004
rect 22376 3952 22428 4004
rect 22192 3927 22244 3936
rect 22192 3893 22201 3927
rect 22201 3893 22235 3927
rect 22235 3893 22244 3927
rect 22192 3884 22244 3893
rect 22468 3927 22520 3936
rect 22468 3893 22477 3927
rect 22477 3893 22511 3927
rect 22511 3893 22520 3927
rect 22468 3884 22520 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1676 3723 1728 3732
rect 1676 3689 1685 3723
rect 1685 3689 1719 3723
rect 1719 3689 1728 3723
rect 1676 3680 1728 3689
rect 1768 3680 1820 3732
rect 2136 3680 2188 3732
rect 3792 3680 3844 3732
rect 3884 3723 3936 3732
rect 3884 3689 3893 3723
rect 3893 3689 3927 3723
rect 3927 3689 3936 3723
rect 5172 3723 5224 3732
rect 3884 3680 3936 3689
rect 5172 3689 5181 3723
rect 5181 3689 5215 3723
rect 5215 3689 5224 3723
rect 5172 3680 5224 3689
rect 6000 3680 6052 3732
rect 7012 3680 7064 3732
rect 7196 3680 7248 3732
rect 9036 3723 9088 3732
rect 9036 3689 9045 3723
rect 9045 3689 9079 3723
rect 9079 3689 9088 3723
rect 9036 3680 9088 3689
rect 9220 3680 9272 3732
rect 9956 3723 10008 3732
rect 9956 3689 9965 3723
rect 9965 3689 9999 3723
rect 9999 3689 10008 3723
rect 9956 3680 10008 3689
rect 10692 3680 10744 3732
rect 10968 3680 11020 3732
rect 11244 3723 11296 3732
rect 11244 3689 11253 3723
rect 11253 3689 11287 3723
rect 11287 3689 11296 3723
rect 11244 3680 11296 3689
rect 11704 3680 11756 3732
rect 14188 3723 14240 3732
rect 14188 3689 14197 3723
rect 14197 3689 14231 3723
rect 14231 3689 14240 3723
rect 14188 3680 14240 3689
rect 15016 3723 15068 3732
rect 15016 3689 15025 3723
rect 15025 3689 15059 3723
rect 15059 3689 15068 3723
rect 15016 3680 15068 3689
rect 16028 3680 16080 3732
rect 16304 3680 16356 3732
rect 18144 3680 18196 3732
rect 18512 3680 18564 3732
rect 18972 3723 19024 3732
rect 18972 3689 18981 3723
rect 18981 3689 19015 3723
rect 19015 3689 19024 3723
rect 18972 3680 19024 3689
rect 20168 3723 20220 3732
rect 20168 3689 20177 3723
rect 20177 3689 20211 3723
rect 20211 3689 20220 3723
rect 20168 3680 20220 3689
rect 3608 3612 3660 3664
rect 3976 3612 4028 3664
rect 5264 3612 5316 3664
rect 6092 3612 6144 3664
rect 6460 3612 6512 3664
rect 7564 3655 7616 3664
rect 7564 3621 7573 3655
rect 7573 3621 7607 3655
rect 7607 3621 7616 3655
rect 7564 3612 7616 3621
rect 1676 3544 1728 3596
rect 2596 3544 2648 3596
rect 12072 3612 12124 3664
rect 14648 3655 14700 3664
rect 14648 3621 14657 3655
rect 14657 3621 14691 3655
rect 14691 3621 14700 3655
rect 14648 3612 14700 3621
rect 17316 3612 17368 3664
rect 2228 3519 2280 3528
rect 2228 3485 2237 3519
rect 2237 3485 2271 3519
rect 2271 3485 2280 3519
rect 2228 3476 2280 3485
rect 7748 3476 7800 3528
rect 8484 3519 8536 3528
rect 8484 3485 8493 3519
rect 8493 3485 8527 3519
rect 8527 3485 8536 3519
rect 8484 3476 8536 3485
rect 8760 3476 8812 3528
rect 10784 3519 10836 3528
rect 10784 3485 10793 3519
rect 10793 3485 10827 3519
rect 10827 3485 10836 3519
rect 10784 3476 10836 3485
rect 16948 3587 17000 3596
rect 16948 3553 16982 3587
rect 16982 3553 17000 3587
rect 16948 3544 17000 3553
rect 19524 3587 19576 3596
rect 19524 3553 19533 3587
rect 19533 3553 19567 3587
rect 19567 3553 19576 3587
rect 19524 3544 19576 3553
rect 21456 3612 21508 3664
rect 22468 3612 22520 3664
rect 21640 3587 21692 3596
rect 21640 3553 21649 3587
rect 21649 3553 21683 3587
rect 21683 3553 21692 3587
rect 21640 3544 21692 3553
rect 22284 3544 22336 3596
rect 19800 3519 19852 3528
rect 19800 3485 19809 3519
rect 19809 3485 19843 3519
rect 19843 3485 19852 3519
rect 19800 3476 19852 3485
rect 6644 3408 6696 3460
rect 7932 3408 7984 3460
rect 13636 3408 13688 3460
rect 3148 3383 3200 3392
rect 3148 3349 3157 3383
rect 3157 3349 3191 3383
rect 3191 3349 3200 3383
rect 3148 3340 3200 3349
rect 4436 3383 4488 3392
rect 4436 3349 4445 3383
rect 4445 3349 4479 3383
rect 4479 3349 4488 3383
rect 4436 3340 4488 3349
rect 8024 3383 8076 3392
rect 8024 3349 8033 3383
rect 8033 3349 8067 3383
rect 8067 3349 8076 3383
rect 8024 3340 8076 3349
rect 10140 3383 10192 3392
rect 10140 3349 10149 3383
rect 10149 3349 10183 3383
rect 10183 3349 10192 3383
rect 10140 3340 10192 3349
rect 10876 3340 10928 3392
rect 11704 3340 11756 3392
rect 13176 3340 13228 3392
rect 13728 3383 13780 3392
rect 13728 3349 13737 3383
rect 13737 3349 13771 3383
rect 13771 3349 13780 3383
rect 13728 3340 13780 3349
rect 14096 3383 14148 3392
rect 14096 3349 14105 3383
rect 14105 3349 14139 3383
rect 14139 3349 14148 3383
rect 14096 3340 14148 3349
rect 16212 3408 16264 3460
rect 19340 3408 19392 3460
rect 17040 3340 17092 3392
rect 17684 3340 17736 3392
rect 19156 3383 19208 3392
rect 19156 3349 19165 3383
rect 19165 3349 19199 3383
rect 19199 3349 19208 3383
rect 19156 3340 19208 3349
rect 21272 3383 21324 3392
rect 21272 3349 21281 3383
rect 21281 3349 21315 3383
rect 21315 3349 21324 3383
rect 21272 3340 21324 3349
rect 21916 3340 21968 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 5172 3136 5224 3188
rect 6460 3136 6512 3188
rect 8208 3136 8260 3188
rect 9772 3136 9824 3188
rect 10784 3179 10836 3188
rect 10784 3145 10793 3179
rect 10793 3145 10827 3179
rect 10827 3145 10836 3179
rect 10784 3136 10836 3145
rect 12072 3136 12124 3188
rect 3056 3068 3108 3120
rect 4068 3068 4120 3120
rect 7748 3068 7800 3120
rect 9588 3068 9640 3120
rect 9956 3068 10008 3120
rect 3148 3000 3200 3052
rect 4712 3000 4764 3052
rect 6644 3000 6696 3052
rect 2136 2932 2188 2984
rect 2228 2864 2280 2916
rect 4252 2932 4304 2984
rect 5264 2975 5316 2984
rect 5264 2941 5273 2975
rect 5273 2941 5307 2975
rect 5307 2941 5316 2975
rect 5264 2932 5316 2941
rect 7288 2975 7340 2984
rect 7288 2941 7297 2975
rect 7297 2941 7331 2975
rect 7331 2941 7340 2975
rect 7288 2932 7340 2941
rect 8760 2975 8812 2984
rect 8760 2941 8794 2975
rect 8794 2941 8812 2975
rect 2780 2864 2832 2916
rect 7380 2907 7432 2916
rect 7380 2873 7389 2907
rect 7389 2873 7423 2907
rect 7423 2873 7432 2907
rect 7380 2864 7432 2873
rect 8760 2932 8812 2941
rect 9588 2932 9640 2984
rect 9036 2864 9088 2916
rect 1676 2839 1728 2848
rect 1676 2805 1685 2839
rect 1685 2805 1719 2839
rect 1719 2805 1728 2839
rect 1676 2796 1728 2805
rect 8392 2796 8444 2848
rect 9312 2796 9364 2848
rect 10876 3000 10928 3052
rect 17316 3136 17368 3188
rect 17776 3179 17828 3188
rect 17776 3145 17785 3179
rect 17785 3145 17819 3179
rect 17819 3145 17828 3179
rect 17776 3136 17828 3145
rect 18052 3179 18104 3188
rect 18052 3145 18061 3179
rect 18061 3145 18095 3179
rect 18095 3145 18104 3179
rect 18052 3136 18104 3145
rect 19064 3179 19116 3188
rect 19064 3145 19073 3179
rect 19073 3145 19107 3179
rect 19107 3145 19116 3179
rect 19064 3136 19116 3145
rect 19340 3136 19392 3188
rect 19800 3136 19852 3188
rect 21456 3179 21508 3188
rect 21456 3145 21465 3179
rect 21465 3145 21499 3179
rect 21499 3145 21508 3179
rect 21456 3136 21508 3145
rect 22284 3136 22336 3188
rect 23848 3179 23900 3188
rect 23848 3145 23857 3179
rect 23857 3145 23891 3179
rect 23891 3145 23900 3179
rect 23848 3136 23900 3145
rect 13912 3068 13964 3120
rect 14464 3068 14516 3120
rect 12348 2932 12400 2984
rect 16672 3000 16724 3052
rect 16948 3000 17000 3052
rect 19524 3068 19576 3120
rect 17776 2932 17828 2984
rect 19432 2932 19484 2984
rect 13728 2864 13780 2916
rect 11428 2839 11480 2848
rect 11428 2805 11437 2839
rect 11437 2805 11471 2839
rect 11471 2805 11480 2839
rect 11428 2796 11480 2805
rect 14096 2864 14148 2916
rect 18236 2864 18288 2916
rect 19524 2864 19576 2916
rect 14740 2796 14792 2848
rect 15200 2796 15252 2848
rect 20352 2932 20404 2984
rect 21456 2932 21508 2984
rect 23572 2932 23624 2984
rect 21824 2839 21876 2848
rect 21824 2805 21833 2839
rect 21833 2805 21867 2839
rect 21867 2805 21876 2839
rect 21824 2796 21876 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 2688 2592 2740 2644
rect 3792 2635 3844 2644
rect 3792 2601 3801 2635
rect 3801 2601 3835 2635
rect 3835 2601 3844 2635
rect 3792 2592 3844 2601
rect 4068 2592 4120 2644
rect 6092 2635 6144 2644
rect 2872 2524 2924 2576
rect 6092 2601 6101 2635
rect 6101 2601 6135 2635
rect 6135 2601 6144 2635
rect 6092 2592 6144 2601
rect 7288 2592 7340 2644
rect 8300 2592 8352 2644
rect 9588 2635 9640 2644
rect 9588 2601 9597 2635
rect 9597 2601 9631 2635
rect 9631 2601 9640 2635
rect 9588 2592 9640 2601
rect 9864 2592 9916 2644
rect 10784 2635 10836 2644
rect 10784 2601 10793 2635
rect 10793 2601 10827 2635
rect 10827 2601 10836 2635
rect 10784 2592 10836 2601
rect 11336 2635 11388 2644
rect 11336 2601 11345 2635
rect 11345 2601 11379 2635
rect 11379 2601 11388 2635
rect 11336 2592 11388 2601
rect 12164 2592 12216 2644
rect 12992 2635 13044 2644
rect 12992 2601 13001 2635
rect 13001 2601 13035 2635
rect 13035 2601 13044 2635
rect 12992 2592 13044 2601
rect 6920 2524 6972 2576
rect 8576 2567 8628 2576
rect 8576 2533 8585 2567
rect 8585 2533 8619 2567
rect 8619 2533 8628 2567
rect 8576 2524 8628 2533
rect 9680 2524 9732 2576
rect 10968 2524 11020 2576
rect 6460 2456 6512 2508
rect 8116 2456 8168 2508
rect 9496 2456 9548 2508
rect 1400 2431 1452 2440
rect 1400 2397 1409 2431
rect 1409 2397 1443 2431
rect 1443 2397 1452 2431
rect 1400 2388 1452 2397
rect 1952 2388 2004 2440
rect 2964 2388 3016 2440
rect 3976 2388 4028 2440
rect 7196 2388 7248 2440
rect 9588 2388 9640 2440
rect 10784 2388 10836 2440
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 13636 2592 13688 2644
rect 14004 2592 14056 2644
rect 14740 2592 14792 2644
rect 16396 2592 16448 2644
rect 16672 2635 16724 2644
rect 16672 2601 16681 2635
rect 16681 2601 16715 2635
rect 16715 2601 16724 2635
rect 16672 2592 16724 2601
rect 18144 2635 18196 2644
rect 18144 2601 18153 2635
rect 18153 2601 18187 2635
rect 18187 2601 18196 2635
rect 18144 2592 18196 2601
rect 18696 2635 18748 2644
rect 18696 2601 18705 2635
rect 18705 2601 18739 2635
rect 18739 2601 18748 2635
rect 18696 2592 18748 2601
rect 19248 2592 19300 2644
rect 13268 2431 13320 2440
rect 11980 2388 12032 2397
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 11152 2320 11204 2372
rect 13176 2320 13228 2372
rect 19340 2524 19392 2576
rect 14740 2456 14792 2508
rect 17132 2499 17184 2508
rect 17132 2465 17141 2499
rect 17141 2465 17175 2499
rect 17175 2465 17184 2499
rect 17132 2456 17184 2465
rect 19432 2456 19484 2508
rect 21548 2499 21600 2508
rect 21548 2465 21557 2499
rect 21557 2465 21591 2499
rect 21591 2465 21600 2499
rect 21548 2456 21600 2465
rect 22744 2499 22796 2508
rect 5448 2295 5500 2304
rect 5448 2261 5457 2295
rect 5457 2261 5491 2295
rect 5491 2261 5500 2295
rect 5448 2252 5500 2261
rect 6460 2295 6512 2304
rect 6460 2261 6469 2295
rect 6469 2261 6503 2295
rect 6503 2261 6512 2295
rect 6460 2252 6512 2261
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 14464 2295 14516 2304
rect 14464 2261 14473 2295
rect 14473 2261 14507 2295
rect 14507 2261 14516 2295
rect 14464 2252 14516 2261
rect 15292 2295 15344 2304
rect 15292 2261 15301 2295
rect 15301 2261 15335 2295
rect 15335 2261 15344 2295
rect 16304 2388 16356 2440
rect 21640 2431 21692 2440
rect 21640 2397 21649 2431
rect 21649 2397 21683 2431
rect 21683 2397 21692 2431
rect 21640 2388 21692 2397
rect 17224 2320 17276 2372
rect 22744 2465 22753 2499
rect 22753 2465 22787 2499
rect 22787 2465 22796 2499
rect 22744 2456 22796 2465
rect 23480 2456 23532 2508
rect 24032 2499 24084 2508
rect 24032 2465 24041 2499
rect 24041 2465 24075 2499
rect 24075 2465 24084 2499
rect 24032 2456 24084 2465
rect 24124 2320 24176 2372
rect 16948 2295 17000 2304
rect 15292 2252 15344 2261
rect 16948 2261 16957 2295
rect 16957 2261 16991 2295
rect 16991 2261 17000 2295
rect 16948 2252 17000 2261
rect 17316 2295 17368 2304
rect 17316 2261 17325 2295
rect 17325 2261 17359 2295
rect 17359 2261 17368 2295
rect 17316 2252 17368 2261
rect 19524 2252 19576 2304
rect 20076 2295 20128 2304
rect 20076 2261 20085 2295
rect 20085 2261 20119 2295
rect 20119 2261 20128 2295
rect 20076 2252 20128 2261
rect 20904 2295 20956 2304
rect 20904 2261 20913 2295
rect 20913 2261 20947 2295
rect 20947 2261 20956 2295
rect 20904 2252 20956 2261
rect 21180 2295 21232 2304
rect 21180 2261 21189 2295
rect 21189 2261 21223 2295
rect 21223 2261 21232 2295
rect 21180 2252 21232 2261
rect 21548 2252 21600 2304
rect 24216 2295 24268 2304
rect 24216 2261 24225 2295
rect 24225 2261 24259 2295
rect 24259 2261 24268 2295
rect 24216 2252 24268 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 1400 1708 1452 1760
rect 3516 1708 3568 1760
rect 7196 1708 7248 1760
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 1950 27520 2006 28000
rect 2502 27520 2558 28000
rect 3054 27704 3110 27713
rect 3054 27639 3110 27648
rect 308 24834 336 27520
rect 32 24806 336 24834
rect 32 12889 60 24806
rect 18 12880 74 12889
rect 18 12815 74 12824
rect 860 10538 888 27520
rect 1412 24834 1440 27520
rect 1860 25356 1912 25362
rect 1860 25298 1912 25304
rect 1412 24806 1532 24834
rect 1400 23520 1452 23526
rect 1400 23462 1452 23468
rect 1308 22024 1360 22030
rect 1308 21966 1360 21972
rect 1320 21690 1348 21966
rect 1308 21684 1360 21690
rect 1308 21626 1360 21632
rect 1412 21321 1440 23462
rect 1398 21312 1454 21321
rect 1398 21247 1454 21256
rect 1504 20806 1532 24806
rect 1872 24721 1900 25298
rect 1858 24712 1914 24721
rect 1858 24647 1914 24656
rect 1584 24608 1636 24614
rect 1584 24550 1636 24556
rect 1596 23526 1624 24550
rect 1872 24410 1900 24647
rect 1860 24404 1912 24410
rect 1860 24346 1912 24352
rect 1676 23792 1728 23798
rect 1676 23734 1728 23740
rect 1584 23520 1636 23526
rect 1584 23462 1636 23468
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1596 21865 1624 22374
rect 1688 22098 1716 23734
rect 1858 23624 1914 23633
rect 1858 23559 1914 23568
rect 1768 22976 1820 22982
rect 1768 22918 1820 22924
rect 1676 22092 1728 22098
rect 1676 22034 1728 22040
rect 1582 21856 1638 21865
rect 1582 21791 1638 21800
rect 1688 21146 1716 22034
rect 1676 21140 1728 21146
rect 1676 21082 1728 21088
rect 1688 20942 1716 21082
rect 1676 20936 1728 20942
rect 1676 20878 1728 20884
rect 1492 20800 1544 20806
rect 1492 20742 1544 20748
rect 1492 20596 1544 20602
rect 1492 20538 1544 20544
rect 1400 19712 1452 19718
rect 1400 19654 1452 19660
rect 1412 19009 1440 19654
rect 1398 19000 1454 19009
rect 1398 18935 1454 18944
rect 1400 18624 1452 18630
rect 1400 18566 1452 18572
rect 1412 17785 1440 18566
rect 1504 18306 1532 20538
rect 1676 20256 1728 20262
rect 1676 20198 1728 20204
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1596 18465 1624 19110
rect 1688 18970 1716 20198
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 1582 18456 1638 18465
rect 1582 18391 1638 18400
rect 1504 18278 1624 18306
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1596 18034 1624 18278
rect 1688 18222 1716 18906
rect 1676 18216 1728 18222
rect 1676 18158 1728 18164
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 1504 16833 1532 18022
rect 1596 18006 1716 18034
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1490 16824 1546 16833
rect 1400 16788 1452 16794
rect 1490 16759 1546 16768
rect 1400 16730 1452 16736
rect 1412 15473 1440 16730
rect 1492 16652 1544 16658
rect 1492 16594 1544 16600
rect 1504 15706 1532 16594
rect 1596 16017 1624 16934
rect 1582 16008 1638 16017
rect 1582 15943 1638 15952
rect 1584 15904 1636 15910
rect 1584 15846 1636 15852
rect 1492 15700 1544 15706
rect 1492 15642 1544 15648
rect 1398 15464 1454 15473
rect 1398 15399 1454 15408
rect 1596 14929 1624 15846
rect 1582 14920 1638 14929
rect 1582 14855 1638 14864
rect 1400 14816 1452 14822
rect 1400 14758 1452 14764
rect 1412 13705 1440 14758
rect 1584 14000 1636 14006
rect 1584 13942 1636 13948
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 1398 13424 1454 13433
rect 1398 13359 1400 13368
rect 1452 13359 1454 13368
rect 1400 13330 1452 13336
rect 1596 13161 1624 13942
rect 1688 13297 1716 18006
rect 1674 13288 1730 13297
rect 1674 13223 1730 13232
rect 1582 13152 1638 13161
rect 1582 13087 1638 13096
rect 1582 12608 1638 12617
rect 1582 12543 1638 12552
rect 1596 11898 1624 12543
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 1780 11529 1808 22918
rect 1872 21486 1900 23559
rect 1860 21480 1912 21486
rect 1860 21422 1912 21428
rect 1964 20602 1992 27520
rect 2412 25356 2464 25362
rect 2412 25298 2464 25304
rect 2228 25152 2280 25158
rect 2228 25094 2280 25100
rect 2042 24848 2098 24857
rect 2042 24783 2044 24792
rect 2096 24783 2098 24792
rect 2044 24754 2096 24760
rect 2240 24410 2268 25094
rect 2424 24954 2452 25298
rect 2412 24948 2464 24954
rect 2412 24890 2464 24896
rect 2516 24834 2544 27520
rect 2778 26616 2834 26625
rect 2778 26551 2834 26560
rect 2332 24806 2544 24834
rect 2228 24404 2280 24410
rect 2228 24346 2280 24352
rect 2044 24268 2096 24274
rect 2044 24210 2096 24216
rect 2056 23866 2084 24210
rect 2044 23860 2096 23866
rect 2044 23802 2096 23808
rect 2240 23662 2268 24346
rect 2228 23656 2280 23662
rect 2042 23624 2098 23633
rect 2228 23598 2280 23604
rect 2042 23559 2098 23568
rect 2056 22778 2084 23559
rect 2136 23520 2188 23526
rect 2136 23462 2188 23468
rect 2148 23186 2176 23462
rect 2136 23180 2188 23186
rect 2136 23122 2188 23128
rect 2044 22772 2096 22778
rect 2044 22714 2096 22720
rect 2056 22574 2084 22714
rect 2044 22568 2096 22574
rect 2044 22510 2096 22516
rect 2148 20602 2176 23122
rect 2228 23112 2280 23118
rect 2228 23054 2280 23060
rect 2240 22098 2268 23054
rect 2228 22092 2280 22098
rect 2228 22034 2280 22040
rect 2332 21978 2360 24806
rect 2792 24750 2820 26551
rect 2964 25220 3016 25226
rect 2964 25162 3016 25168
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 2780 24744 2832 24750
rect 2780 24686 2832 24692
rect 2596 24608 2648 24614
rect 2596 24550 2648 24556
rect 2504 24064 2556 24070
rect 2504 24006 2556 24012
rect 2516 23798 2544 24006
rect 2504 23792 2556 23798
rect 2504 23734 2556 23740
rect 2608 23730 2636 24550
rect 2792 24410 2820 24686
rect 2780 24404 2832 24410
rect 2780 24346 2832 24352
rect 2596 23724 2648 23730
rect 2648 23684 2820 23712
rect 2596 23666 2648 23672
rect 2792 23322 2820 23684
rect 2780 23316 2832 23322
rect 2780 23258 2832 23264
rect 2688 23112 2740 23118
rect 2884 23089 2912 25094
rect 2688 23054 2740 23060
rect 2870 23080 2926 23089
rect 2596 22636 2648 22642
rect 2596 22578 2648 22584
rect 2504 22092 2556 22098
rect 2504 22034 2556 22040
rect 2240 21950 2360 21978
rect 2412 22024 2464 22030
rect 2412 21966 2464 21972
rect 1952 20596 2004 20602
rect 1952 20538 2004 20544
rect 2136 20596 2188 20602
rect 2136 20538 2188 20544
rect 2240 20482 2268 21950
rect 2424 21842 2452 21966
rect 2332 21814 2452 21842
rect 2332 21418 2360 21814
rect 2320 21412 2372 21418
rect 2320 21354 2372 21360
rect 2332 21146 2360 21354
rect 2516 21146 2544 22034
rect 2608 21690 2636 22578
rect 2700 22030 2728 23054
rect 2870 23015 2926 23024
rect 2976 22545 3004 25162
rect 3068 24342 3096 27639
rect 3146 27520 3202 28000
rect 3698 27520 3754 28000
rect 4250 27520 4306 28000
rect 4802 27520 4858 28000
rect 5354 27520 5410 28000
rect 5998 27520 6054 28000
rect 6550 27520 6606 28000
rect 7102 27520 7158 28000
rect 7654 27520 7710 28000
rect 8206 27520 8262 28000
rect 8850 27520 8906 28000
rect 9402 27520 9458 28000
rect 9954 27520 10010 28000
rect 10506 27520 10562 28000
rect 11058 27520 11114 28000
rect 11702 27520 11758 28000
rect 12254 27520 12310 28000
rect 12806 27520 12862 28000
rect 13358 27520 13414 28000
rect 13910 27520 13966 28000
rect 14554 27520 14610 28000
rect 15106 27520 15162 28000
rect 15658 27520 15714 28000
rect 16210 27520 16266 28000
rect 16762 27520 16818 28000
rect 17406 27520 17462 28000
rect 17958 27520 18014 28000
rect 18510 27520 18566 28000
rect 19062 27520 19118 28000
rect 19614 27520 19670 28000
rect 20258 27520 20314 28000
rect 20810 27520 20866 28000
rect 21362 27520 21418 28000
rect 21914 27520 21970 28000
rect 22466 27520 22522 28000
rect 23110 27520 23166 28000
rect 23662 27520 23718 28000
rect 24214 27520 24270 28000
rect 24766 27520 24822 28000
rect 25318 27520 25374 28000
rect 25962 27520 26018 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 3056 24336 3108 24342
rect 3056 24278 3108 24284
rect 3068 23866 3096 24278
rect 3056 23860 3108 23866
rect 3056 23802 3108 23808
rect 3054 23216 3110 23225
rect 3054 23151 3110 23160
rect 2962 22536 3018 22545
rect 2962 22471 3018 22480
rect 2688 22024 2740 22030
rect 2688 21966 2740 21972
rect 2596 21684 2648 21690
rect 2596 21626 2648 21632
rect 2320 21140 2372 21146
rect 2320 21082 2372 21088
rect 2504 21140 2556 21146
rect 2504 21082 2556 21088
rect 2962 20904 3018 20913
rect 2962 20839 3018 20848
rect 2320 20800 2372 20806
rect 2320 20742 2372 20748
rect 1872 20454 2268 20482
rect 1872 14521 1900 20454
rect 2044 20256 2096 20262
rect 2044 20198 2096 20204
rect 2056 19961 2084 20198
rect 2042 19952 2098 19961
rect 2042 19887 2098 19896
rect 2136 19916 2188 19922
rect 2136 19858 2188 19864
rect 2042 19816 2098 19825
rect 2042 19751 2044 19760
rect 2096 19751 2098 19760
rect 2044 19722 2096 19728
rect 2044 17876 2096 17882
rect 2044 17818 2096 17824
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 17134 1992 17478
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1964 15745 1992 17070
rect 2056 16794 2084 17818
rect 2044 16788 2096 16794
rect 2044 16730 2096 16736
rect 2042 16552 2098 16561
rect 2042 16487 2098 16496
rect 2056 16250 2084 16487
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 2056 16046 2084 16186
rect 2044 16040 2096 16046
rect 2044 15982 2096 15988
rect 1950 15736 2006 15745
rect 1950 15671 2006 15680
rect 2042 15600 2098 15609
rect 2042 15535 2044 15544
rect 2096 15535 2098 15544
rect 2044 15506 2096 15512
rect 2056 15162 2084 15506
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 2148 14634 2176 19858
rect 2228 18828 2280 18834
rect 2228 18770 2280 18776
rect 2240 17814 2268 18770
rect 2228 17808 2280 17814
rect 2228 17750 2280 17756
rect 2240 17649 2268 17750
rect 2226 17640 2282 17649
rect 2226 17575 2282 17584
rect 2332 17490 2360 20742
rect 2870 20360 2926 20369
rect 2700 20318 2870 20346
rect 2700 20097 2728 20318
rect 2870 20295 2926 20304
rect 2686 20088 2742 20097
rect 2976 20058 3004 20839
rect 2686 20023 2742 20032
rect 2964 20052 3016 20058
rect 2964 19994 3016 20000
rect 3068 19922 3096 23151
rect 3056 19916 3108 19922
rect 3056 19858 3108 19864
rect 2686 19544 2742 19553
rect 2686 19479 2742 19488
rect 2504 19304 2556 19310
rect 2502 19272 2504 19281
rect 2556 19272 2558 19281
rect 2502 19207 2558 19216
rect 2700 18970 2728 19479
rect 2688 18964 2740 18970
rect 2688 18906 2740 18912
rect 2502 18864 2558 18873
rect 2502 18799 2504 18808
rect 2556 18799 2558 18808
rect 2504 18770 2556 18776
rect 2516 18426 2544 18770
rect 2596 18624 2648 18630
rect 2596 18566 2648 18572
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 2504 18080 2556 18086
rect 2504 18022 2556 18028
rect 2516 17678 2544 18022
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 2240 17462 2360 17490
rect 2240 15337 2268 17462
rect 2320 17264 2372 17270
rect 2320 17206 2372 17212
rect 2332 15706 2360 17206
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 2424 16114 2452 16934
rect 2516 16794 2544 17614
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2412 16108 2464 16114
rect 2412 16050 2464 16056
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 2504 15428 2556 15434
rect 2504 15370 2556 15376
rect 2226 15328 2282 15337
rect 2226 15263 2282 15272
rect 2516 14958 2544 15370
rect 2608 15026 2636 18566
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 2780 17604 2832 17610
rect 2780 17546 2832 17552
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2700 17338 2728 17478
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 2686 17232 2742 17241
rect 2686 17167 2742 17176
rect 2700 16794 2728 17167
rect 2792 17066 2820 17546
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 2780 17060 2832 17066
rect 2780 17002 2832 17008
rect 2688 16788 2740 16794
rect 2688 16730 2740 16736
rect 2976 15910 3004 17070
rect 3068 16998 3096 17614
rect 3160 17252 3188 27520
rect 3606 27160 3662 27169
rect 3606 27095 3662 27104
rect 3238 25392 3294 25401
rect 3238 25327 3294 25336
rect 3252 25158 3280 25327
rect 3240 25152 3292 25158
rect 3240 25094 3292 25100
rect 3252 24614 3280 25094
rect 3240 24608 3292 24614
rect 3240 24550 3292 24556
rect 3252 19009 3280 24550
rect 3516 24404 3568 24410
rect 3516 24346 3568 24352
rect 3332 24132 3384 24138
rect 3332 24074 3384 24080
rect 3344 23594 3372 24074
rect 3332 23588 3384 23594
rect 3332 23530 3384 23536
rect 3344 23254 3372 23530
rect 3332 23248 3384 23254
rect 3332 23190 3384 23196
rect 3344 22574 3372 23190
rect 3332 22568 3384 22574
rect 3332 22510 3384 22516
rect 3528 21457 3556 24346
rect 3620 21690 3648 27095
rect 3712 24834 3740 27520
rect 4066 25936 4122 25945
rect 4066 25871 4122 25880
rect 4080 24886 4108 25871
rect 4068 24880 4120 24886
rect 3712 24806 3924 24834
rect 4068 24822 4120 24828
rect 3700 24268 3752 24274
rect 3700 24210 3752 24216
rect 3712 24177 3740 24210
rect 3698 24168 3754 24177
rect 3698 24103 3754 24112
rect 3712 23866 3740 24103
rect 3700 23860 3752 23866
rect 3700 23802 3752 23808
rect 3608 21684 3660 21690
rect 3608 21626 3660 21632
rect 3514 21448 3570 21457
rect 3514 21383 3570 21392
rect 3424 20460 3476 20466
rect 3424 20402 3476 20408
rect 3332 19984 3384 19990
rect 3332 19926 3384 19932
rect 3344 19514 3372 19926
rect 3436 19922 3464 20402
rect 3424 19916 3476 19922
rect 3424 19858 3476 19864
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 3238 19000 3294 19009
rect 3238 18935 3294 18944
rect 3424 18964 3476 18970
rect 3252 18290 3280 18935
rect 3528 18952 3556 21383
rect 3608 21344 3660 21350
rect 3608 21286 3660 21292
rect 3620 20874 3648 21286
rect 3608 20868 3660 20874
rect 3608 20810 3660 20816
rect 3620 20330 3648 20810
rect 3608 20324 3660 20330
rect 3608 20266 3660 20272
rect 3620 20058 3648 20266
rect 3608 20052 3660 20058
rect 3608 19994 3660 20000
rect 3712 19258 3740 23802
rect 3792 23792 3844 23798
rect 3792 23734 3844 23740
rect 3476 18924 3556 18952
rect 3620 19230 3740 19258
rect 3424 18906 3476 18912
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 3436 18222 3464 18906
rect 3620 18873 3648 19230
rect 3700 19168 3752 19174
rect 3700 19110 3752 19116
rect 3606 18864 3662 18873
rect 3606 18799 3662 18808
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 3424 18216 3476 18222
rect 3424 18158 3476 18164
rect 3528 17678 3556 18226
rect 3516 17672 3568 17678
rect 3516 17614 3568 17620
rect 3160 17224 3280 17252
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 3146 16824 3202 16833
rect 3146 16759 3148 16768
rect 3200 16759 3202 16768
rect 3148 16730 3200 16736
rect 3252 16017 3280 17224
rect 3330 17232 3386 17241
rect 3330 17167 3386 17176
rect 3238 16008 3294 16017
rect 3238 15943 3294 15952
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2792 14958 2820 15302
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2504 14952 2556 14958
rect 2504 14894 2556 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2148 14606 2452 14634
rect 2516 14618 2544 14894
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 1858 14512 1914 14521
rect 2424 14498 2452 14606
rect 2504 14612 2556 14618
rect 2504 14554 2556 14560
rect 1858 14447 1914 14456
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 2228 14476 2280 14482
rect 2424 14470 2544 14498
rect 2228 14418 2280 14424
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 1872 13870 1900 14214
rect 1860 13864 1912 13870
rect 2056 13841 2084 14418
rect 2240 13870 2268 14418
rect 2412 14272 2464 14278
rect 2412 14214 2464 14220
rect 2228 13864 2280 13870
rect 1860 13806 1912 13812
rect 2042 13832 2098 13841
rect 1872 13530 1900 13806
rect 2228 13806 2280 13812
rect 2042 13767 2098 13776
rect 2136 13728 2188 13734
rect 2136 13670 2188 13676
rect 2148 13530 2176 13670
rect 1860 13524 1912 13530
rect 1860 13466 1912 13472
rect 2136 13524 2188 13530
rect 2136 13466 2188 13472
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 1964 12374 1992 13330
rect 2148 13258 2176 13466
rect 2136 13252 2188 13258
rect 2136 13194 2188 13200
rect 2148 12782 2176 13194
rect 2136 12776 2188 12782
rect 2136 12718 2188 12724
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 1952 12368 2004 12374
rect 1952 12310 2004 12316
rect 2148 12102 2176 12582
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 2148 11558 2176 12038
rect 2136 11552 2188 11558
rect 1766 11520 1822 11529
rect 2136 11494 2188 11500
rect 1766 11455 1822 11464
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 848 10532 900 10538
rect 848 10474 900 10480
rect 1412 10033 1440 10542
rect 1780 10266 1808 11086
rect 1858 10976 1914 10985
rect 1858 10911 1914 10920
rect 1872 10674 1900 10911
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1872 10146 1900 10610
rect 1780 10118 1900 10146
rect 1398 10024 1454 10033
rect 1398 9959 1400 9968
rect 1452 9959 1454 9968
rect 1400 9930 1452 9936
rect 1780 9722 1808 10118
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 1768 9716 1820 9722
rect 1768 9658 1820 9664
rect 1872 9654 1900 9998
rect 1860 9648 1912 9654
rect 1858 9616 1860 9625
rect 1912 9616 1914 9625
rect 1914 9574 1992 9602
rect 2056 9586 2084 9998
rect 2148 9586 2176 11494
rect 1858 9551 1914 9560
rect 1872 9525 1900 9551
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1398 8392 1454 8401
rect 1398 8327 1454 8336
rect 1412 7546 1440 8327
rect 1596 7886 1624 9318
rect 1780 8090 1808 9454
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 1412 5166 1440 7482
rect 1492 7268 1544 7274
rect 1492 7210 1544 7216
rect 1504 7002 1532 7210
rect 1596 7206 1624 7822
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1492 6996 1544 7002
rect 1492 6938 1544 6944
rect 1400 5160 1452 5166
rect 1400 5102 1452 5108
rect 294 4176 350 4185
rect 294 4111 350 4120
rect 308 480 336 4111
rect 846 3360 902 3369
rect 846 3295 902 3304
rect 860 480 888 3295
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 1412 1873 1440 2382
rect 1398 1864 1454 1873
rect 1398 1799 1454 1808
rect 1400 1760 1452 1766
rect 1400 1702 1452 1708
rect 1412 480 1440 1702
rect 1596 1465 1624 7142
rect 1872 5273 1900 7686
rect 1964 7342 1992 9574
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2148 8838 2176 9522
rect 2136 8832 2188 8838
rect 2136 8774 2188 8780
rect 2148 8362 2176 8774
rect 2240 8498 2268 13806
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2332 12986 2360 13670
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2318 12608 2374 12617
rect 2318 12543 2374 12552
rect 2332 8634 2360 12543
rect 2424 10010 2452 14214
rect 2516 11354 2544 14470
rect 2700 14385 2728 14758
rect 2884 14414 2912 14962
rect 2872 14408 2924 14414
rect 2686 14376 2742 14385
rect 2872 14350 2924 14356
rect 2686 14311 2742 14320
rect 2884 13705 2912 14350
rect 2976 13870 3004 15846
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 3068 14890 3096 15438
rect 3056 14884 3108 14890
rect 3056 14826 3108 14832
rect 3238 14376 3294 14385
rect 3238 14311 3294 14320
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 3252 13802 3280 14311
rect 3344 13938 3372 17167
rect 3528 17134 3556 17614
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 3424 16652 3476 16658
rect 3424 16594 3476 16600
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3240 13796 3292 13802
rect 3240 13738 3292 13744
rect 2870 13696 2926 13705
rect 2870 13631 2926 13640
rect 2778 13560 2834 13569
rect 2778 13495 2780 13504
rect 2832 13495 2834 13504
rect 2780 13466 2832 13472
rect 3146 13288 3202 13297
rect 3146 13223 3202 13232
rect 3160 13190 3188 13223
rect 2596 13184 2648 13190
rect 2596 13126 2648 13132
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 2608 11354 2636 13126
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2792 12102 2820 12650
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2792 11354 2820 12038
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2596 11348 2648 11354
rect 2780 11348 2832 11354
rect 2596 11290 2648 11296
rect 2700 11308 2780 11336
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2608 10810 2636 11154
rect 2596 10804 2648 10810
rect 2596 10746 2648 10752
rect 2700 10674 2728 11308
rect 2780 11290 2832 11296
rect 2872 11280 2924 11286
rect 2872 11222 2924 11228
rect 2884 11150 2912 11222
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 2884 10169 2912 11086
rect 3160 10810 3188 13126
rect 3252 12617 3280 13738
rect 3238 12608 3294 12617
rect 3238 12543 3294 12552
rect 3344 10810 3372 13874
rect 3436 13462 3464 16594
rect 3608 14952 3660 14958
rect 3608 14894 3660 14900
rect 3620 14618 3648 14894
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 3528 13938 3556 14350
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3424 13456 3476 13462
rect 3424 13398 3476 13404
rect 3528 13258 3556 13874
rect 3712 13433 3740 19110
rect 3804 18193 3832 23734
rect 3790 18184 3846 18193
rect 3790 18119 3846 18128
rect 3792 14000 3844 14006
rect 3792 13942 3844 13948
rect 3896 13954 3924 24806
rect 4160 24608 4212 24614
rect 4066 24576 4122 24585
rect 4160 24550 4212 24556
rect 4066 24511 4122 24520
rect 3976 23112 4028 23118
rect 4080 23089 4108 24511
rect 3976 23054 4028 23060
rect 4066 23080 4122 23089
rect 3988 22098 4016 23054
rect 4066 23015 4122 23024
rect 4068 22432 4120 22438
rect 4068 22374 4120 22380
rect 3976 22092 4028 22098
rect 3976 22034 4028 22040
rect 4080 21876 4108 22374
rect 4172 22030 4200 24550
rect 4264 24342 4292 27520
rect 4344 24744 4396 24750
rect 4344 24686 4396 24692
rect 4252 24336 4304 24342
rect 4252 24278 4304 24284
rect 4252 24200 4304 24206
rect 4252 24142 4304 24148
rect 4264 23798 4292 24142
rect 4252 23792 4304 23798
rect 4250 23760 4252 23769
rect 4304 23760 4306 23769
rect 4250 23695 4306 23704
rect 4252 23656 4304 23662
rect 4252 23598 4304 23604
rect 4264 23186 4292 23598
rect 4252 23180 4304 23186
rect 4252 23122 4304 23128
rect 4264 22778 4292 23122
rect 4252 22772 4304 22778
rect 4252 22714 4304 22720
rect 4160 22024 4212 22030
rect 4160 21966 4212 21972
rect 4356 21894 4384 24686
rect 4816 24410 4844 27520
rect 5368 25362 5396 27520
rect 5356 25356 5408 25362
rect 5356 25298 5408 25304
rect 4896 25152 4948 25158
rect 4896 25094 4948 25100
rect 4908 24818 4936 25094
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 4896 24812 4948 24818
rect 4896 24754 4948 24760
rect 4804 24404 4856 24410
rect 4804 24346 4856 24352
rect 4712 24336 4764 24342
rect 4712 24278 4764 24284
rect 4436 22976 4488 22982
rect 4436 22918 4488 22924
rect 4160 21888 4212 21894
rect 4080 21848 4160 21876
rect 4080 21010 4108 21848
rect 4160 21830 4212 21836
rect 4344 21888 4396 21894
rect 4344 21830 4396 21836
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 4160 20936 4212 20942
rect 4080 20884 4160 20890
rect 4080 20878 4212 20884
rect 4080 20862 4200 20878
rect 4080 20398 4108 20862
rect 4160 20800 4212 20806
rect 4160 20742 4212 20748
rect 4068 20392 4120 20398
rect 4068 20334 4120 20340
rect 4172 19310 4200 20742
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 4172 18902 4200 19246
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4264 18970 4292 19110
rect 4252 18964 4304 18970
rect 4252 18906 4304 18912
rect 4356 18902 4384 19314
rect 4160 18896 4212 18902
rect 4160 18838 4212 18844
rect 4344 18896 4396 18902
rect 4344 18838 4396 18844
rect 4252 18828 4304 18834
rect 4252 18770 4304 18776
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4172 17898 4200 18022
rect 4080 17870 4200 17898
rect 4080 17066 4108 17870
rect 4264 17814 4292 18770
rect 4356 18222 4384 18838
rect 4344 18216 4396 18222
rect 4344 18158 4396 18164
rect 4252 17808 4304 17814
rect 4252 17750 4304 17756
rect 4068 17060 4120 17066
rect 4068 17002 4120 17008
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 3988 15638 4016 16730
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4080 15706 4108 16390
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4250 15736 4306 15745
rect 4068 15700 4120 15706
rect 4250 15671 4252 15680
rect 4068 15642 4120 15648
rect 4304 15671 4306 15680
rect 4252 15642 4304 15648
rect 3976 15632 4028 15638
rect 3976 15574 4028 15580
rect 4080 15162 4108 15642
rect 4160 15564 4212 15570
rect 4160 15506 4212 15512
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4172 15094 4200 15506
rect 4160 15088 4212 15094
rect 4160 15030 4212 15036
rect 4356 14890 4384 15846
rect 4344 14884 4396 14890
rect 4344 14826 4396 14832
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4172 14482 4200 14758
rect 4356 14482 4384 14826
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4344 14476 4396 14482
rect 4344 14418 4396 14424
rect 4172 14362 4200 14418
rect 4172 14334 4292 14362
rect 3698 13424 3754 13433
rect 3698 13359 3754 13368
rect 3516 13252 3568 13258
rect 3516 13194 3568 13200
rect 3606 12880 3662 12889
rect 3606 12815 3662 12824
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 3436 11694 3464 12582
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3436 11150 3464 11630
rect 3620 11393 3648 12815
rect 3712 12442 3740 13359
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3606 11384 3662 11393
rect 3606 11319 3662 11328
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3422 10432 3478 10441
rect 3422 10367 3478 10376
rect 2870 10160 2926 10169
rect 2870 10095 2926 10104
rect 2424 9982 2544 10010
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 2424 9518 2452 9862
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2516 9217 2544 9982
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 3068 9586 3096 9862
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2502 9208 2558 9217
rect 2884 9178 2912 9454
rect 2502 9143 2558 9152
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 3344 8498 3372 8910
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2056 7410 2084 7822
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 1952 7336 2004 7342
rect 1952 7278 2004 7284
rect 1964 7002 1992 7278
rect 2056 7002 2084 7346
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 2044 6996 2096 7002
rect 2044 6938 2096 6944
rect 2056 6458 2084 6938
rect 2148 6458 2176 8298
rect 2596 8288 2648 8294
rect 3148 8288 3200 8294
rect 2596 8230 2648 8236
rect 3146 8256 3148 8265
rect 3200 8256 3202 8265
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2240 6662 2268 8026
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2056 5846 2084 6394
rect 2044 5840 2096 5846
rect 2044 5782 2096 5788
rect 2148 5778 2176 6394
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 1858 5264 1914 5273
rect 1858 5199 1860 5208
rect 1912 5199 1914 5208
rect 1860 5170 1912 5176
rect 1766 4992 1822 5001
rect 1766 4927 1822 4936
rect 1780 4146 1808 4927
rect 2148 4826 2176 5714
rect 2240 5545 2268 6598
rect 2412 5636 2464 5642
rect 2412 5578 2464 5584
rect 2226 5536 2282 5545
rect 2226 5471 2282 5480
rect 2424 5234 2452 5578
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1674 3768 1730 3777
rect 1780 3738 1808 4082
rect 2148 3738 2176 4762
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2332 4214 2360 4422
rect 2320 4208 2372 4214
rect 2320 4150 2372 4156
rect 2228 4004 2280 4010
rect 2228 3946 2280 3952
rect 1674 3703 1676 3712
rect 1728 3703 1730 3712
rect 1768 3732 1820 3738
rect 1676 3674 1728 3680
rect 1768 3674 1820 3680
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1688 2854 1716 3538
rect 2148 2990 2176 3674
rect 2240 3534 2268 3946
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 2240 2922 2268 3470
rect 2228 2916 2280 2922
rect 2228 2858 2280 2864
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1582 1456 1638 1465
rect 1582 1391 1638 1400
rect 1688 921 1716 2790
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 1674 912 1730 921
rect 1674 847 1730 856
rect 1964 480 1992 2382
rect 2332 1601 2360 3878
rect 2502 3632 2558 3641
rect 2608 3602 2636 8230
rect 3146 8191 3202 8200
rect 3160 8090 3188 8191
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 3160 7002 3188 7686
rect 3436 7313 3464 10367
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3528 9178 3556 9998
rect 3804 9489 3832 13942
rect 3896 13926 4016 13954
rect 3882 13832 3938 13841
rect 3882 13767 3938 13776
rect 3896 13462 3924 13767
rect 3988 13512 4016 13926
rect 4264 13870 4292 14334
rect 4356 14074 4384 14418
rect 4344 14068 4396 14074
rect 4344 14010 4396 14016
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4160 13524 4212 13530
rect 3988 13484 4160 13512
rect 4160 13466 4212 13472
rect 3884 13456 3936 13462
rect 3884 13398 3936 13404
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 3882 12608 3938 12617
rect 3882 12543 3938 12552
rect 3896 11354 3924 12543
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3988 11898 4016 12038
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3988 11354 4016 11834
rect 4080 11642 4108 13194
rect 4172 12782 4200 13466
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4264 12238 4292 13806
rect 4342 13560 4398 13569
rect 4342 13495 4398 13504
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 4264 11937 4292 12038
rect 4250 11928 4306 11937
rect 4250 11863 4306 11872
rect 4356 11665 4384 13495
rect 4448 11694 4476 22918
rect 4724 22148 4752 24278
rect 4908 24206 4936 24754
rect 5080 24676 5132 24682
rect 5080 24618 5132 24624
rect 4896 24200 4948 24206
rect 4896 24142 4948 24148
rect 4908 23866 4936 24142
rect 4988 24064 5040 24070
rect 4988 24006 5040 24012
rect 4896 23860 4948 23866
rect 4896 23802 4948 23808
rect 4804 23588 4856 23594
rect 4804 23530 4856 23536
rect 4816 23050 4844 23530
rect 4804 23044 4856 23050
rect 4804 22986 4856 22992
rect 4816 22778 4844 22986
rect 4804 22772 4856 22778
rect 4804 22714 4856 22720
rect 5000 22166 5028 24006
rect 4988 22160 5040 22166
rect 4724 22120 4936 22148
rect 4528 22024 4580 22030
rect 4908 21978 4936 22120
rect 4988 22102 5040 22108
rect 4528 21966 4580 21972
rect 4540 21146 4568 21966
rect 4816 21950 4936 21978
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 4528 21140 4580 21146
rect 4528 21082 4580 21088
rect 4526 18184 4582 18193
rect 4526 18119 4582 18128
rect 4540 17882 4568 18119
rect 4528 17876 4580 17882
rect 4528 17818 4580 17824
rect 4540 17338 4568 17818
rect 4528 17332 4580 17338
rect 4528 17274 4580 17280
rect 4528 16720 4580 16726
rect 4528 16662 4580 16668
rect 4540 15706 4568 16662
rect 4528 15700 4580 15706
rect 4528 15642 4580 15648
rect 4528 13796 4580 13802
rect 4528 13738 4580 13744
rect 4540 13530 4568 13738
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4540 12986 4568 13466
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4436 11688 4488 11694
rect 4342 11656 4398 11665
rect 4080 11614 4200 11642
rect 4066 11520 4122 11529
rect 4066 11455 4122 11464
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 3882 11248 3938 11257
rect 4080 11218 4108 11455
rect 3882 11183 3884 11192
rect 3936 11183 3938 11192
rect 4068 11212 4120 11218
rect 3884 11154 3936 11160
rect 4068 11154 4120 11160
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3896 10470 3924 10610
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 3896 9926 3924 10406
rect 4172 10266 4200 11614
rect 4436 11630 4488 11636
rect 4342 11591 4398 11600
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4264 10470 4292 11494
rect 4540 10606 4568 12922
rect 4528 10600 4580 10606
rect 4528 10542 4580 10548
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3974 9888 4030 9897
rect 3790 9480 3846 9489
rect 3790 9415 3846 9424
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3896 8974 3924 9862
rect 3974 9823 4030 9832
rect 3988 9625 4016 9823
rect 4172 9738 4200 10202
rect 4080 9710 4200 9738
rect 3974 9616 4030 9625
rect 3974 9551 4030 9560
rect 4080 9518 4108 9710
rect 4068 9512 4120 9518
rect 4632 9466 4660 21830
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4724 18154 4752 19110
rect 4712 18148 4764 18154
rect 4712 18090 4764 18096
rect 4816 17082 4844 21950
rect 4896 20936 4948 20942
rect 4896 20878 4948 20884
rect 4908 20602 4936 20878
rect 4896 20596 4948 20602
rect 4896 20538 4948 20544
rect 4908 19990 4936 20538
rect 4896 19984 4948 19990
rect 4896 19926 4948 19932
rect 4908 18766 4936 19926
rect 4896 18760 4948 18766
rect 4896 18702 4948 18708
rect 4908 18426 4936 18702
rect 4896 18420 4948 18426
rect 4896 18362 4948 18368
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 5000 17678 5028 18022
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 4724 17054 4844 17082
rect 4724 13802 4752 17054
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4816 16590 4844 16934
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4816 16250 4844 16526
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4802 15328 4858 15337
rect 4802 15263 4858 15272
rect 4816 14074 4844 15263
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4712 13796 4764 13802
rect 4712 13738 4764 13744
rect 4816 13394 4844 14010
rect 4908 13569 4936 16594
rect 5000 16522 5028 17614
rect 4988 16516 5040 16522
rect 4988 16458 5040 16464
rect 4894 13560 4950 13569
rect 4894 13495 4950 13504
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4724 12102 4752 13262
rect 4816 12918 4844 13330
rect 4804 12912 4856 12918
rect 4804 12854 4856 12860
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4724 10198 4752 12038
rect 4816 11898 4844 12242
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4908 10266 4936 10746
rect 5000 10606 5028 10950
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 4712 10192 4764 10198
rect 4712 10134 4764 10140
rect 4068 9454 4120 9460
rect 4540 9438 4660 9466
rect 4710 9480 4766 9489
rect 4436 9104 4488 9110
rect 4434 9072 4436 9081
rect 4488 9072 4490 9081
rect 4434 9007 4490 9016
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 4066 8936 4122 8945
rect 4066 8871 4068 8880
rect 4120 8871 4122 8880
rect 4068 8842 4120 8848
rect 3790 8528 3846 8537
rect 3846 8486 4200 8514
rect 3790 8463 3846 8472
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3528 7410 3556 7686
rect 4172 7546 4200 8486
rect 4540 7886 4568 9438
rect 4710 9415 4766 9424
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4632 8974 4660 9318
rect 4724 9178 4752 9415
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4632 8362 4660 8910
rect 4620 8356 4672 8362
rect 4620 8298 4672 8304
rect 4712 8016 4764 8022
rect 4712 7958 4764 7964
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4436 7472 4488 7478
rect 4436 7414 4488 7420
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3422 7304 3478 7313
rect 3422 7239 3478 7248
rect 3516 7268 3568 7274
rect 3516 7210 3568 7216
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 4758 2728 6598
rect 3068 6254 3096 6734
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 2872 6180 2924 6186
rect 2872 6122 2924 6128
rect 2884 5642 2912 6122
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 2872 5636 2924 5642
rect 2872 5578 2924 5584
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 2884 4826 2912 5238
rect 3068 5166 3096 6054
rect 3330 5944 3386 5953
rect 3330 5879 3386 5888
rect 3056 5160 3108 5166
rect 3054 5128 3056 5137
rect 3108 5128 3110 5137
rect 3054 5063 3110 5072
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2688 4752 2740 4758
rect 2688 4694 2740 4700
rect 2870 4720 2926 4729
rect 2870 4655 2872 4664
rect 2924 4655 2926 4664
rect 2872 4626 2924 4632
rect 3068 4622 3096 5063
rect 3056 4616 3108 4622
rect 2686 4584 2742 4593
rect 3056 4558 3108 4564
rect 2686 4519 2742 4528
rect 2700 4146 2728 4519
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2502 3567 2558 3576
rect 2596 3596 2648 3602
rect 2318 1592 2374 1601
rect 2318 1527 2374 1536
rect 2516 480 2544 3567
rect 2596 3538 2648 3544
rect 2700 3233 2728 3878
rect 2884 3505 2912 4422
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 2870 3496 2926 3505
rect 2870 3431 2926 3440
rect 2686 3224 2742 3233
rect 2686 3159 2742 3168
rect 3068 3126 3096 4082
rect 3344 3913 3372 5879
rect 3436 4185 3464 7142
rect 3528 6662 3556 7210
rect 4448 7041 4476 7414
rect 4434 7032 4490 7041
rect 3608 6996 3660 7002
rect 4434 6967 4436 6976
rect 3608 6938 3660 6944
rect 4488 6967 4490 6976
rect 4436 6938 4488 6944
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3422 4176 3478 4185
rect 3422 4111 3478 4120
rect 3330 3904 3386 3913
rect 3330 3839 3386 3848
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 3056 3120 3108 3126
rect 3056 3062 3108 3068
rect 3160 3058 3188 3334
rect 3422 3088 3478 3097
rect 3148 3052 3200 3058
rect 3422 3023 3478 3032
rect 3148 2994 3200 3000
rect 2870 2952 2926 2961
rect 2780 2916 2832 2922
rect 2870 2887 2926 2896
rect 2780 2858 2832 2864
rect 2792 2802 2820 2858
rect 2700 2774 2820 2802
rect 2700 2650 2728 2774
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 2884 2582 2912 2887
rect 2872 2576 2924 2582
rect 2872 2518 2924 2524
rect 2962 2544 3018 2553
rect 2884 1306 2912 2518
rect 2962 2479 3018 2488
rect 2976 2446 3004 2479
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2884 1278 3188 1306
rect 3160 480 3188 1278
rect 3436 1057 3464 3023
rect 3528 1766 3556 6598
rect 3620 5914 3648 6938
rect 4540 6798 4568 7686
rect 4632 7410 4660 7686
rect 4724 7478 4752 7958
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4528 6792 4580 6798
rect 4526 6760 4528 6769
rect 4580 6760 4582 6769
rect 3804 6730 4200 6746
rect 3804 6724 4212 6730
rect 3804 6718 4160 6724
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3620 3670 3648 5850
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3712 5234 3740 5510
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3712 4865 3740 4966
rect 3698 4856 3754 4865
rect 3698 4791 3754 4800
rect 3804 4457 3832 6718
rect 4526 6695 4582 6704
rect 4160 6666 4212 6672
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3974 6352 4030 6361
rect 3974 6287 4030 6296
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3790 4448 3846 4457
rect 3790 4383 3846 4392
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3698 3904 3754 3913
rect 3698 3839 3754 3848
rect 3608 3664 3660 3670
rect 3608 3606 3660 3612
rect 3516 1760 3568 1766
rect 3516 1702 3568 1708
rect 3422 1048 3478 1057
rect 3422 983 3478 992
rect 3712 480 3740 3839
rect 3804 3738 3832 4014
rect 3896 3738 3924 5510
rect 3988 5001 4016 6287
rect 4080 6225 4108 6598
rect 4066 6216 4122 6225
rect 4066 6151 4122 6160
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4066 5672 4122 5681
rect 4066 5607 4122 5616
rect 4080 5302 4108 5607
rect 4172 5370 4200 5714
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 4160 5024 4212 5030
rect 3974 4992 4030 5001
rect 3974 4927 4030 4936
rect 4080 4984 4160 5012
rect 4080 4554 4108 4984
rect 4160 4966 4212 4972
rect 4436 4684 4488 4690
rect 4436 4626 4488 4632
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 4172 4282 4200 4558
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4356 4010 4384 4422
rect 4344 4004 4396 4010
rect 4344 3946 4396 3952
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3804 2650 3832 3674
rect 3976 3664 4028 3670
rect 3976 3606 4028 3612
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3988 2446 4016 3606
rect 4448 3398 4476 4626
rect 4540 3641 4568 6054
rect 4632 5778 4660 7346
rect 4804 6996 4856 7002
rect 4804 6938 4856 6944
rect 4816 6905 4844 6938
rect 4896 6928 4948 6934
rect 4802 6896 4858 6905
rect 4896 6870 4948 6876
rect 4802 6831 4858 6840
rect 4908 6089 4936 6870
rect 4894 6080 4950 6089
rect 4894 6015 4950 6024
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4632 5166 4660 5714
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4632 3942 4660 5102
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4526 3632 4582 3641
rect 4526 3567 4582 3576
rect 4436 3392 4488 3398
rect 4434 3360 4436 3369
rect 4488 3360 4490 3369
rect 4434 3295 4490 3304
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 4080 2650 4108 3062
rect 4724 3058 4752 4966
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 4264 480 4292 2926
rect 5000 2417 5028 7890
rect 4986 2408 5042 2417
rect 4986 2343 5042 2352
rect 5092 1034 5120 24618
rect 6012 24342 6040 27520
rect 6092 24880 6144 24886
rect 6092 24822 6144 24828
rect 6000 24336 6052 24342
rect 6000 24278 6052 24284
rect 5448 24064 5500 24070
rect 5448 24006 5500 24012
rect 5262 23488 5318 23497
rect 5262 23423 5318 23432
rect 5172 23248 5224 23254
rect 5172 23190 5224 23196
rect 5184 22438 5212 23190
rect 5276 23118 5304 23423
rect 5264 23112 5316 23118
rect 5264 23054 5316 23060
rect 5460 22930 5488 24006
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 6012 23798 6040 24278
rect 6000 23792 6052 23798
rect 6000 23734 6052 23740
rect 5460 22902 5580 22930
rect 5552 22681 5580 22902
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 6104 22778 6132 24822
rect 6564 24721 6592 27520
rect 7116 24750 7144 27520
rect 7104 24744 7156 24750
rect 6550 24712 6606 24721
rect 7104 24686 7156 24692
rect 6550 24647 6606 24656
rect 7196 24608 7248 24614
rect 7196 24550 7248 24556
rect 7380 24608 7432 24614
rect 7380 24550 7432 24556
rect 6184 24404 6236 24410
rect 6184 24346 6236 24352
rect 6196 23866 6224 24346
rect 6920 24268 6972 24274
rect 6920 24210 6972 24216
rect 6932 24154 6960 24210
rect 7208 24206 7236 24550
rect 6840 24126 6960 24154
rect 7196 24200 7248 24206
rect 7196 24142 7248 24148
rect 6184 23860 6236 23866
rect 6184 23802 6236 23808
rect 6736 23792 6788 23798
rect 6736 23734 6788 23740
rect 6276 23656 6328 23662
rect 6276 23598 6328 23604
rect 6288 23118 6316 23598
rect 6644 23520 6696 23526
rect 6644 23462 6696 23468
rect 6656 23254 6684 23462
rect 6644 23248 6696 23254
rect 6644 23190 6696 23196
rect 6276 23112 6328 23118
rect 6276 23054 6328 23060
rect 6366 23080 6422 23089
rect 6092 22772 6144 22778
rect 6092 22714 6144 22720
rect 5538 22672 5594 22681
rect 5538 22607 5594 22616
rect 5632 22636 5684 22642
rect 5552 22574 5580 22607
rect 5632 22578 5684 22584
rect 6000 22636 6052 22642
rect 6000 22578 6052 22584
rect 5540 22568 5592 22574
rect 5540 22510 5592 22516
rect 5172 22432 5224 22438
rect 5172 22374 5224 22380
rect 5184 22234 5212 22374
rect 5644 22234 5672 22578
rect 6012 22234 6040 22578
rect 6104 22574 6132 22714
rect 6092 22568 6144 22574
rect 6092 22510 6144 22516
rect 5172 22228 5224 22234
rect 5172 22170 5224 22176
rect 5632 22228 5684 22234
rect 5632 22170 5684 22176
rect 6000 22228 6052 22234
rect 6000 22170 6052 22176
rect 5540 22160 5592 22166
rect 5540 22102 5592 22108
rect 5448 21548 5500 21554
rect 5448 21490 5500 21496
rect 5172 21344 5224 21350
rect 5172 21286 5224 21292
rect 5264 21344 5316 21350
rect 5264 21286 5316 21292
rect 5184 21010 5212 21286
rect 5172 21004 5224 21010
rect 5172 20946 5224 20952
rect 5184 19310 5212 20946
rect 5276 19310 5304 21286
rect 5460 20806 5488 21490
rect 5552 21146 5580 22102
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6104 21146 6132 22510
rect 6288 21894 6316 23054
rect 6366 23015 6422 23024
rect 6380 22778 6408 23015
rect 6368 22772 6420 22778
rect 6368 22714 6420 22720
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 5540 21140 5592 21146
rect 5540 21082 5592 21088
rect 6092 21140 6144 21146
rect 6092 21082 6144 21088
rect 6000 20936 6052 20942
rect 6000 20878 6052 20884
rect 5448 20800 5500 20806
rect 5500 20760 5580 20788
rect 5448 20742 5500 20748
rect 5552 20602 5580 20760
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 6012 20262 6040 20878
rect 6104 20602 6132 21082
rect 6380 20942 6408 22714
rect 6656 22642 6684 23190
rect 6644 22636 6696 22642
rect 6644 22578 6696 22584
rect 6642 22536 6698 22545
rect 6642 22471 6698 22480
rect 6656 22098 6684 22471
rect 6644 22092 6696 22098
rect 6644 22034 6696 22040
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6564 21350 6592 21966
rect 6656 21486 6684 22034
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6552 21344 6604 21350
rect 6550 21312 6552 21321
rect 6604 21312 6606 21321
rect 6550 21247 6606 21256
rect 6368 20936 6420 20942
rect 6368 20878 6420 20884
rect 6184 20800 6236 20806
rect 6184 20742 6236 20748
rect 6092 20596 6144 20602
rect 6092 20538 6144 20544
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 5448 19712 5500 19718
rect 5448 19654 5500 19660
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5460 19378 5488 19654
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 5184 17882 5212 18906
rect 5552 18902 5580 19654
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5540 18896 5592 18902
rect 6012 18873 6040 20198
rect 6196 19786 6224 20742
rect 6656 20058 6684 21422
rect 6644 20052 6696 20058
rect 6644 19994 6696 20000
rect 6184 19780 6236 19786
rect 6184 19722 6236 19728
rect 6196 19514 6224 19722
rect 6184 19508 6236 19514
rect 6184 19450 6236 19456
rect 5540 18838 5592 18844
rect 5998 18864 6054 18873
rect 6196 18834 6224 19450
rect 6644 19168 6696 19174
rect 6564 19116 6644 19122
rect 6564 19110 6696 19116
rect 6564 19094 6684 19110
rect 5998 18799 6054 18808
rect 6184 18828 6236 18834
rect 6184 18770 6236 18776
rect 5998 18728 6054 18737
rect 5998 18663 6054 18672
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 5264 17740 5316 17746
rect 5264 17682 5316 17688
rect 5276 17338 5304 17682
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5552 17241 5580 17478
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5538 17232 5594 17241
rect 5538 17167 5594 17176
rect 5724 17128 5776 17134
rect 5724 17070 5776 17076
rect 5540 17060 5592 17066
rect 5540 17002 5592 17008
rect 5264 16516 5316 16522
rect 5264 16458 5316 16464
rect 5276 16250 5304 16458
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5552 15858 5580 17002
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5644 16561 5672 16934
rect 5736 16697 5764 17070
rect 6012 16794 6040 18663
rect 6196 17882 6224 18770
rect 6184 17876 6236 17882
rect 6184 17818 6236 17824
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 6380 16998 6408 17614
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6472 17338 6500 17478
rect 6460 17332 6512 17338
rect 6460 17274 6512 17280
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 5722 16688 5778 16697
rect 5722 16623 5724 16632
rect 5776 16623 5778 16632
rect 5724 16594 5776 16600
rect 5630 16552 5686 16561
rect 5630 16487 5686 16496
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6012 16250 6040 16730
rect 6184 16584 6236 16590
rect 6236 16532 6316 16538
rect 6184 16526 6316 16532
rect 6196 16510 6316 16526
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5368 15830 5580 15858
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 5170 15464 5226 15473
rect 5170 15399 5226 15408
rect 5184 14074 5212 15399
rect 5368 15094 5396 15830
rect 5736 15706 5764 15846
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5724 15700 5776 15706
rect 6012 15688 6040 16186
rect 6288 15910 6316 16510
rect 6380 16454 6408 16934
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6380 16114 6408 16390
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 6012 15660 6132 15688
rect 5724 15642 5776 15648
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5460 15162 5488 15302
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5356 15088 5408 15094
rect 5356 15030 5408 15036
rect 5552 14958 5580 15642
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6012 15026 6040 15506
rect 6000 15020 6052 15026
rect 6000 14962 6052 14968
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 6012 14618 6040 14962
rect 6000 14612 6052 14618
rect 6000 14554 6052 14560
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6104 14113 6132 15660
rect 6184 15632 6236 15638
rect 6184 15574 6236 15580
rect 6196 14822 6224 15574
rect 6288 15337 6316 15846
rect 6380 15638 6408 16050
rect 6368 15632 6420 15638
rect 6368 15574 6420 15580
rect 6274 15328 6330 15337
rect 6274 15263 6330 15272
rect 6564 14890 6592 19094
rect 6644 18896 6696 18902
rect 6644 18838 6696 18844
rect 6656 18154 6684 18838
rect 6644 18148 6696 18154
rect 6644 18090 6696 18096
rect 6552 14884 6604 14890
rect 6552 14826 6604 14832
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6196 14414 6224 14758
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6090 14104 6146 14113
rect 5172 14068 5224 14074
rect 6196 14074 6224 14350
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6090 14039 6146 14048
rect 6184 14068 6236 14074
rect 5172 14010 5224 14016
rect 6184 14010 6236 14016
rect 6092 14000 6144 14006
rect 6092 13942 6144 13948
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5460 13569 5488 13874
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5446 13560 5502 13569
rect 5446 13495 5502 13504
rect 5170 13424 5226 13433
rect 5170 13359 5226 13368
rect 5184 12986 5212 13359
rect 5552 13190 5580 13670
rect 5630 13288 5686 13297
rect 5630 13223 5632 13232
rect 5684 13223 5686 13232
rect 5632 13194 5684 13200
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5540 12640 5592 12646
rect 5632 12640 5684 12646
rect 5540 12582 5592 12588
rect 5630 12608 5632 12617
rect 5684 12608 5686 12617
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 5368 11830 5396 12174
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 5276 11354 5304 11630
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5368 11218 5396 11766
rect 5460 11558 5488 12242
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 5460 11098 5488 11494
rect 5368 11070 5488 11098
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5276 9926 5304 10406
rect 5368 10062 5396 11070
rect 5448 10804 5500 10810
rect 5552 10792 5580 12582
rect 5630 12543 5686 12552
rect 5736 12442 5764 12786
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 6000 12096 6052 12102
rect 5998 12064 6000 12073
rect 6052 12064 6054 12073
rect 5622 11996 5918 12016
rect 5998 11999 6054 12008
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6000 11280 6052 11286
rect 6000 11222 6052 11228
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5500 10764 5580 10792
rect 5448 10746 5500 10752
rect 6012 10674 6040 11222
rect 6104 10690 6132 13942
rect 6380 13938 6408 14214
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6274 13696 6330 13705
rect 6274 13631 6330 13640
rect 6184 13456 6236 13462
rect 6184 13398 6236 13404
rect 6196 13161 6224 13398
rect 6182 13152 6238 13161
rect 6182 13087 6238 13096
rect 6196 12986 6224 13087
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6184 12436 6236 12442
rect 6184 12378 6236 12384
rect 6196 11898 6224 12378
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 6196 10810 6224 11630
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6000 10668 6052 10674
rect 6104 10662 6224 10690
rect 6000 10610 6052 10616
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 6090 10568 6146 10577
rect 5460 10266 5488 10542
rect 6090 10503 6146 10512
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 6000 10192 6052 10198
rect 6000 10134 6052 10140
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5276 9722 5304 9862
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5368 9654 5396 9998
rect 5356 9648 5408 9654
rect 5356 9590 5408 9596
rect 5552 9586 5580 10066
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 6012 9382 6040 10134
rect 6104 9897 6132 10503
rect 6090 9888 6146 9897
rect 6090 9823 6146 9832
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5540 8968 5592 8974
rect 5460 8916 5540 8922
rect 5460 8910 5592 8916
rect 5460 8894 5580 8910
rect 5172 8016 5224 8022
rect 5172 7958 5224 7964
rect 5184 7546 5212 7958
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5184 6730 5212 7142
rect 5460 6866 5488 8894
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5552 8401 5580 8774
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5538 8392 5594 8401
rect 5538 8327 5594 8336
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5276 6322 5304 6598
rect 5460 6458 5488 6802
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5276 5914 5304 6258
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5172 5024 5224 5030
rect 5170 4992 5172 5001
rect 5224 4992 5226 5001
rect 5226 4950 5304 4978
rect 5170 4927 5226 4936
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5184 3738 5212 4762
rect 5276 4593 5304 4950
rect 5368 4622 5396 5102
rect 5460 4758 5488 6122
rect 5552 5166 5580 8230
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5828 6866 5856 7346
rect 6012 7342 6040 9318
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6104 7410 6132 7686
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6012 6458 6040 6734
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5552 4826 5580 4966
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5448 4752 5500 4758
rect 5448 4694 5500 4700
rect 5644 4690 5672 5034
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5356 4616 5408 4622
rect 5262 4584 5318 4593
rect 5356 4558 5408 4564
rect 5262 4519 5318 4528
rect 5368 4128 5396 4558
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5552 4185 5580 4490
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6012 4282 6040 4694
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 5276 4100 5396 4128
rect 5538 4176 5594 4185
rect 5538 4111 5594 4120
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5276 3670 5304 4100
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5264 3664 5316 3670
rect 5170 3632 5226 3641
rect 5264 3606 5316 3612
rect 5170 3567 5226 3576
rect 5184 3233 5212 3567
rect 5170 3224 5226 3233
rect 5170 3159 5172 3168
rect 5224 3159 5226 3168
rect 5172 3130 5224 3136
rect 5184 3099 5212 3130
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 5276 2689 5304 2926
rect 5262 2680 5318 2689
rect 5262 2615 5318 2624
rect 4816 1006 5120 1034
rect 4816 480 4844 1006
rect 5368 480 5396 3878
rect 5460 2310 5488 3946
rect 6012 3913 6040 4218
rect 6196 4185 6224 10662
rect 6288 8634 6316 13631
rect 6380 13326 6408 13874
rect 6564 13530 6592 14486
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6380 13025 6408 13262
rect 6366 13016 6422 13025
rect 6564 12986 6592 13466
rect 6366 12951 6422 12960
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6368 12912 6420 12918
rect 6368 12854 6420 12860
rect 6380 10849 6408 12854
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6564 12442 6592 12786
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6366 10840 6422 10849
rect 6366 10775 6422 10784
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6380 8514 6408 9386
rect 6472 9178 6500 12378
rect 6656 9654 6684 18090
rect 6748 14006 6776 23734
rect 6840 21962 6868 24126
rect 7104 24064 7156 24070
rect 7104 24006 7156 24012
rect 7116 23662 7144 24006
rect 7104 23656 7156 23662
rect 7104 23598 7156 23604
rect 7208 23594 7236 24142
rect 7392 24138 7420 24550
rect 7380 24132 7432 24138
rect 7380 24074 7432 24080
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 7196 23588 7248 23594
rect 7196 23530 7248 23536
rect 7208 23322 7236 23530
rect 7484 23497 7512 24006
rect 7470 23488 7526 23497
rect 7470 23423 7526 23432
rect 7668 23338 7696 27520
rect 7840 24608 7892 24614
rect 7840 24550 7892 24556
rect 7852 24274 7880 24550
rect 7840 24268 7892 24274
rect 7840 24210 7892 24216
rect 8116 24200 8168 24206
rect 8116 24142 8168 24148
rect 7748 23588 7800 23594
rect 7748 23530 7800 23536
rect 7196 23316 7248 23322
rect 7196 23258 7248 23264
rect 7484 23310 7696 23338
rect 6828 21956 6880 21962
rect 6828 21898 6880 21904
rect 7104 21888 7156 21894
rect 7104 21830 7156 21836
rect 7012 21344 7064 21350
rect 7012 21286 7064 21292
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6932 19174 6960 19994
rect 7024 19961 7052 21286
rect 7116 20398 7144 21830
rect 7484 21026 7512 23310
rect 7760 22642 7788 23530
rect 8128 23526 8156 24142
rect 8116 23520 8168 23526
rect 8116 23462 8168 23468
rect 8220 23338 8248 27520
rect 8864 24834 8892 27520
rect 8772 24806 8892 24834
rect 8772 23633 8800 24806
rect 9416 24698 9444 27520
rect 9968 24857 9996 27520
rect 10520 25786 10548 27520
rect 10520 25758 10732 25786
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 9954 24848 10010 24857
rect 9954 24783 10010 24792
rect 8864 24670 9444 24698
rect 8758 23624 8814 23633
rect 8758 23559 8814 23568
rect 8128 23310 8248 23338
rect 7748 22636 7800 22642
rect 7748 22578 7800 22584
rect 7760 21962 7788 22578
rect 7748 21956 7800 21962
rect 7748 21898 7800 21904
rect 7656 21888 7708 21894
rect 7656 21830 7708 21836
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7576 21146 7604 21354
rect 7668 21350 7696 21830
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7564 21140 7616 21146
rect 7564 21082 7616 21088
rect 7288 21004 7340 21010
rect 7484 20998 7604 21026
rect 7288 20946 7340 20952
rect 7196 20936 7248 20942
rect 7300 20913 7328 20946
rect 7196 20878 7248 20884
rect 7286 20904 7342 20913
rect 7208 20602 7236 20878
rect 7286 20839 7288 20848
rect 7340 20839 7342 20848
rect 7288 20810 7340 20816
rect 7196 20596 7248 20602
rect 7196 20538 7248 20544
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 7116 19990 7144 20334
rect 7104 19984 7156 19990
rect 7010 19952 7066 19961
rect 7104 19926 7156 19932
rect 7286 19952 7342 19961
rect 7010 19887 7066 19896
rect 7116 19836 7144 19926
rect 7286 19887 7288 19896
rect 7340 19887 7342 19896
rect 7288 19858 7340 19864
rect 7024 19808 7144 19836
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 6828 18692 6880 18698
rect 6828 18634 6880 18640
rect 6840 18086 6868 18634
rect 7024 18630 7052 19808
rect 7300 19378 7328 19858
rect 7104 19372 7156 19378
rect 7104 19314 7156 19320
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 7024 18222 7052 18566
rect 7012 18216 7064 18222
rect 7012 18158 7064 18164
rect 6828 18080 6880 18086
rect 6826 18048 6828 18057
rect 6880 18048 6882 18057
rect 6826 17983 6882 17992
rect 7024 17542 7052 18158
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 6920 15904 6972 15910
rect 7024 15892 7052 16594
rect 6972 15864 7052 15892
rect 6920 15846 6972 15852
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6840 14958 6868 15302
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6736 14000 6788 14006
rect 6736 13942 6788 13948
rect 6840 13841 6868 14758
rect 6826 13832 6882 13841
rect 6826 13767 6882 13776
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6840 12594 6868 13126
rect 6932 12850 6960 15846
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6840 12566 7052 12594
rect 6920 12164 6972 12170
rect 6920 12106 6972 12112
rect 6736 12096 6788 12102
rect 6932 12050 6960 12106
rect 6736 12038 6788 12044
rect 6748 11286 6776 12038
rect 6840 12022 6960 12050
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6840 10810 6868 12022
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6932 11354 6960 11630
rect 7024 11393 7052 12566
rect 7116 11937 7144 19314
rect 7470 19000 7526 19009
rect 7470 18935 7472 18944
rect 7524 18935 7526 18944
rect 7472 18906 7524 18912
rect 7380 18148 7432 18154
rect 7380 18090 7432 18096
rect 7392 17542 7420 18090
rect 7576 18057 7604 20998
rect 7668 19514 7696 21286
rect 7760 20806 7788 21898
rect 7748 20800 7800 20806
rect 7748 20742 7800 20748
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7562 18048 7618 18057
rect 7562 17983 7618 17992
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7392 17202 7420 17478
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7668 17134 7696 18566
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 7300 16794 7328 16934
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7196 16584 7248 16590
rect 7196 16526 7248 16532
rect 7208 16046 7236 16526
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7208 15706 7236 15982
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7208 15162 7236 15642
rect 7654 15328 7710 15337
rect 7654 15263 7710 15272
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7300 14074 7328 14894
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7392 13938 7420 14554
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7208 13530 7236 13806
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7392 13394 7420 13874
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7484 13274 7512 13466
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7392 13246 7512 13274
rect 7196 12776 7248 12782
rect 7194 12744 7196 12753
rect 7248 12744 7250 12753
rect 7194 12679 7250 12688
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7300 12170 7328 12582
rect 7392 12442 7420 13246
rect 7576 12986 7604 13330
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7484 12442 7512 12786
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7484 12102 7512 12378
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7102 11928 7158 11937
rect 7102 11863 7158 11872
rect 7010 11384 7066 11393
rect 6920 11348 6972 11354
rect 7010 11319 7066 11328
rect 6920 11290 6972 11296
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6288 8486 6408 8514
rect 6288 8106 6316 8486
rect 6472 8294 6500 8978
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6288 8078 6408 8106
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6288 7206 6316 7890
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6288 6905 6316 7142
rect 6274 6896 6330 6905
rect 6274 6831 6330 6840
rect 6274 5128 6330 5137
rect 6274 5063 6276 5072
rect 6328 5063 6330 5072
rect 6276 5034 6328 5040
rect 6380 4826 6408 8078
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6472 6458 6500 7142
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6472 5166 6500 6394
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 6182 4176 6238 4185
rect 6182 4111 6238 4120
rect 5998 3904 6054 3913
rect 5998 3839 6054 3848
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 5460 1465 5488 2246
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5446 1456 5502 1465
rect 5446 1391 5502 1400
rect 6012 480 6040 3674
rect 6092 3664 6144 3670
rect 6092 3606 6144 3612
rect 6104 2650 6132 3606
rect 6092 2644 6144 2650
rect 6092 2586 6144 2592
rect 6288 2417 6316 4422
rect 6380 4282 6408 4762
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6274 2408 6330 2417
rect 6274 2343 6330 2352
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 1950 0 2006 480
rect 2502 0 2558 480
rect 3146 0 3202 480
rect 3698 0 3754 480
rect 4250 0 4306 480
rect 4802 0 4858 480
rect 5354 0 5410 480
rect 5998 0 6054 480
rect 6380 377 6408 4218
rect 6472 3670 6500 5102
rect 6564 3942 6592 9454
rect 6932 9382 6960 9862
rect 6920 9376 6972 9382
rect 6748 9324 6920 9330
rect 6748 9318 6972 9324
rect 7010 9344 7066 9353
rect 6748 9302 6960 9318
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6656 3754 6684 9114
rect 6748 7274 6776 9302
rect 7010 9279 7066 9288
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6840 7342 6868 8230
rect 6932 7750 6960 8230
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 6826 6488 6882 6497
rect 6826 6423 6828 6432
rect 6880 6423 6882 6432
rect 6828 6394 6880 6400
rect 6932 6361 6960 7686
rect 6918 6352 6974 6361
rect 6918 6287 6974 6296
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 6840 4554 6868 5782
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 6564 3726 6684 3754
rect 7024 3738 7052 9279
rect 7116 8362 7144 11863
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7300 10538 7328 11086
rect 7288 10532 7340 10538
rect 7288 10474 7340 10480
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7392 9586 7420 9998
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7668 9058 7696 15263
rect 7760 9178 7788 20742
rect 7838 20496 7894 20505
rect 7838 20431 7894 20440
rect 7852 20058 7880 20431
rect 8024 20392 8076 20398
rect 8024 20334 8076 20340
rect 8036 20058 8064 20334
rect 7840 20052 7892 20058
rect 7840 19994 7892 20000
rect 8024 20052 8076 20058
rect 8024 19994 8076 20000
rect 7852 19378 7880 19994
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 7852 16810 7880 19314
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 7944 18737 7972 19110
rect 8024 18828 8076 18834
rect 8024 18770 8076 18776
rect 7930 18728 7986 18737
rect 7930 18663 7986 18672
rect 8036 17814 8064 18770
rect 8024 17808 8076 17814
rect 8024 17750 8076 17756
rect 8036 17338 8064 17750
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 7852 16782 7972 16810
rect 7840 16720 7892 16726
rect 7840 16662 7892 16668
rect 7852 16153 7880 16662
rect 7838 16144 7894 16153
rect 7838 16079 7894 16088
rect 7852 15706 7880 16079
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7944 15586 7972 16782
rect 8128 16726 8156 23310
rect 8484 22976 8536 22982
rect 8484 22918 8536 22924
rect 8392 22704 8444 22710
rect 8390 22672 8392 22681
rect 8444 22672 8446 22681
rect 8390 22607 8446 22616
rect 8496 22574 8524 22918
rect 8484 22568 8536 22574
rect 8484 22510 8536 22516
rect 8208 22432 8260 22438
rect 8208 22374 8260 22380
rect 8220 22001 8248 22374
rect 8496 22234 8524 22510
rect 8484 22228 8536 22234
rect 8484 22170 8536 22176
rect 8206 21992 8262 22001
rect 8206 21927 8262 21936
rect 8220 21690 8248 21927
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 8220 20618 8248 21490
rect 8482 21448 8538 21457
rect 8482 21383 8484 21392
rect 8536 21383 8538 21392
rect 8484 21354 8536 21360
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 8220 20602 8340 20618
rect 8220 20596 8352 20602
rect 8220 20590 8300 20596
rect 8300 20538 8352 20544
rect 8496 20330 8524 20742
rect 8484 20324 8536 20330
rect 8484 20266 8536 20272
rect 8496 19718 8524 20266
rect 8484 19712 8536 19718
rect 8484 19654 8536 19660
rect 8496 19378 8524 19654
rect 8484 19372 8536 19378
rect 8484 19314 8536 19320
rect 8496 19174 8524 19314
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8220 17746 8248 18702
rect 8496 18426 8524 19110
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8208 17740 8260 17746
rect 8208 17682 8260 17688
rect 8220 17542 8248 17682
rect 8208 17536 8260 17542
rect 8208 17478 8260 17484
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8588 16833 8616 16934
rect 8574 16824 8630 16833
rect 8680 16794 8708 17070
rect 8772 17066 8800 17478
rect 8760 17060 8812 17066
rect 8760 17002 8812 17008
rect 8574 16759 8630 16768
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8116 16720 8168 16726
rect 8116 16662 8168 16668
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 8036 15706 8064 16526
rect 8114 16008 8170 16017
rect 8864 15994 8892 24670
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10600 24268 10652 24274
rect 10600 24210 10652 24216
rect 9494 23760 9550 23769
rect 9494 23695 9550 23704
rect 9312 22432 9364 22438
rect 9312 22374 9364 22380
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 9048 21554 9076 21830
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 9036 21344 9088 21350
rect 9036 21286 9088 21292
rect 9126 21312 9182 21321
rect 8956 19990 8984 21286
rect 9048 21146 9076 21286
rect 9126 21247 9182 21256
rect 9036 21140 9088 21146
rect 9036 21082 9088 21088
rect 9048 20058 9076 21082
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 8944 19984 8996 19990
rect 8944 19926 8996 19932
rect 8956 19310 8984 19926
rect 8944 19304 8996 19310
rect 8944 19246 8996 19252
rect 8114 15943 8170 15952
rect 8680 15966 8892 15994
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 7944 15558 8064 15586
rect 7840 14816 7892 14822
rect 7840 14758 7892 14764
rect 7852 13870 7880 14758
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 7838 11384 7894 11393
rect 7838 11319 7894 11328
rect 7852 10266 7880 11319
rect 7944 11121 7972 12922
rect 7930 11112 7986 11121
rect 7930 11047 7986 11056
rect 7840 10260 7892 10266
rect 7840 10202 7892 10208
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7564 9036 7616 9042
rect 7668 9030 7880 9058
rect 7564 8978 7616 8984
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7194 8528 7250 8537
rect 7392 8498 7420 8774
rect 7576 8634 7604 8978
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7194 8463 7250 8472
rect 7380 8492 7432 8498
rect 7208 8430 7236 8463
rect 7380 8434 7432 8440
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7116 7274 7144 7686
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 7116 6662 7144 7210
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7116 5710 7144 6598
rect 7208 6254 7236 8026
rect 7286 6352 7342 6361
rect 7286 6287 7288 6296
rect 7340 6287 7342 6296
rect 7288 6258 7340 6264
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7300 5914 7328 6258
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7116 4826 7144 5646
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7208 4078 7236 4626
rect 7196 4072 7248 4078
rect 7102 4040 7158 4049
rect 7196 4014 7248 4020
rect 7102 3975 7158 3984
rect 7012 3732 7064 3738
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6472 3194 6500 3606
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6460 2508 6512 2514
rect 6460 2450 6512 2456
rect 6472 2310 6500 2450
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 6472 2145 6500 2246
rect 6458 2136 6514 2145
rect 6458 2071 6514 2080
rect 6564 480 6592 3726
rect 7012 3674 7064 3680
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6656 3058 6684 3402
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6918 2680 6974 2689
rect 6918 2615 6974 2624
rect 6932 2582 6960 2615
rect 6920 2576 6972 2582
rect 6920 2518 6972 2524
rect 7116 480 7144 3975
rect 7208 3738 7236 4014
rect 7286 3904 7342 3913
rect 7286 3839 7342 3848
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7208 2446 7236 3674
rect 7300 2990 7328 3839
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 7378 2952 7434 2961
rect 7300 2650 7328 2926
rect 7378 2887 7380 2896
rect 7432 2887 7434 2896
rect 7380 2858 7432 2864
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7208 1766 7236 2382
rect 7196 1760 7248 1766
rect 7196 1702 7248 1708
rect 7484 1306 7512 8298
rect 7576 7546 7604 8570
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7576 6458 7604 7482
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7668 5953 7696 6802
rect 7654 5944 7710 5953
rect 7654 5879 7656 5888
rect 7708 5879 7710 5888
rect 7656 5850 7708 5856
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7576 5137 7604 5714
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7562 5128 7618 5137
rect 7562 5063 7618 5072
rect 7576 4826 7604 5063
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7576 3670 7604 4490
rect 7564 3664 7616 3670
rect 7668 3641 7696 5510
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7760 4486 7788 4966
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 7760 4078 7788 4422
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7564 3606 7616 3612
rect 7654 3632 7710 3641
rect 7654 3567 7710 3576
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7760 3126 7788 3470
rect 7748 3120 7800 3126
rect 7746 3088 7748 3097
rect 7800 3088 7802 3097
rect 7746 3023 7802 3032
rect 7852 1442 7880 9030
rect 8036 8888 8064 15558
rect 8128 10112 8156 15943
rect 8484 15632 8536 15638
rect 8484 15574 8536 15580
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8208 14952 8260 14958
rect 8312 14940 8340 15302
rect 8496 15162 8524 15574
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8260 14912 8340 14940
rect 8208 14894 8260 14900
rect 8390 14512 8446 14521
rect 8390 14447 8446 14456
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8220 12306 8248 13942
rect 8404 13870 8432 14447
rect 8588 14074 8616 15438
rect 8576 14068 8628 14074
rect 8576 14010 8628 14016
rect 8680 13954 8708 15966
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8772 14890 8800 15846
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 8772 14278 8800 14826
rect 9048 14385 9076 15302
rect 9034 14376 9090 14385
rect 9034 14311 9090 14320
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8588 13926 8708 13954
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8404 13190 8432 13670
rect 8588 13530 8616 13926
rect 8668 13796 8720 13802
rect 8668 13738 8720 13744
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8392 13184 8444 13190
rect 8390 13152 8392 13161
rect 8484 13184 8536 13190
rect 8444 13152 8446 13161
rect 8484 13126 8536 13132
rect 8390 13087 8446 13096
rect 8390 13016 8446 13025
rect 8390 12951 8392 12960
rect 8444 12951 8446 12960
rect 8392 12922 8444 12928
rect 8496 12442 8524 13126
rect 8588 12481 8616 13466
rect 8574 12472 8630 12481
rect 8484 12436 8536 12442
rect 8574 12407 8630 12416
rect 8484 12378 8536 12384
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8220 12209 8248 12242
rect 8206 12200 8262 12209
rect 8206 12135 8262 12144
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8220 11286 8248 11494
rect 8298 11384 8354 11393
rect 8496 11354 8524 12378
rect 8298 11319 8300 11328
rect 8352 11319 8354 11328
rect 8484 11348 8536 11354
rect 8300 11290 8352 11296
rect 8484 11290 8536 11296
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 8220 10538 8248 11222
rect 8300 11076 8352 11082
rect 8300 11018 8352 11024
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 8312 10266 8340 11018
rect 8588 10577 8616 11018
rect 8574 10568 8630 10577
rect 8574 10503 8630 10512
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8300 10124 8352 10130
rect 8128 10084 8300 10112
rect 8114 9752 8170 9761
rect 8220 9738 8248 10084
rect 8300 10066 8352 10072
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8170 9710 8248 9738
rect 8114 9687 8170 9696
rect 8128 9654 8156 9687
rect 8116 9648 8168 9654
rect 8116 9590 8168 9596
rect 8312 9586 8340 9930
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8404 8922 8432 9862
rect 8496 9722 8524 9998
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8496 9178 8524 9658
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8220 8894 8432 8922
rect 8036 8860 8156 8888
rect 8022 8800 8078 8809
rect 8022 8735 8078 8744
rect 8036 7818 8064 8735
rect 8128 7954 8156 8860
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8024 7812 8076 7818
rect 8024 7754 8076 7760
rect 8128 7585 8156 7890
rect 8114 7576 8170 7585
rect 8114 7511 8170 7520
rect 7930 5944 7986 5953
rect 7930 5879 7986 5888
rect 7944 4554 7972 5879
rect 8220 5692 8248 8894
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8312 7274 8340 7890
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 8312 6866 8340 7210
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8298 6760 8354 6769
rect 8298 6695 8354 6704
rect 8312 6458 8340 6695
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8298 6216 8354 6225
rect 8298 6151 8354 6160
rect 8312 5914 8340 6151
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8128 5664 8248 5692
rect 8022 5400 8078 5409
rect 8022 5335 8078 5344
rect 8036 4826 8064 5335
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 7932 4548 7984 4554
rect 7932 4490 7984 4496
rect 7930 4448 7986 4457
rect 7930 4383 7986 4392
rect 7944 3942 7972 4383
rect 8036 4282 8064 4762
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 8128 4162 8156 5664
rect 8404 5624 8432 8774
rect 8496 8362 8524 9114
rect 8484 8356 8536 8362
rect 8536 8316 8616 8344
rect 8484 8298 8536 8304
rect 8588 7886 8616 8316
rect 8576 7880 8628 7886
rect 8482 7848 8538 7857
rect 8576 7822 8628 7828
rect 8482 7783 8484 7792
rect 8536 7783 8538 7792
rect 8484 7754 8536 7760
rect 8496 7546 8524 7754
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8588 7478 8616 7822
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 8574 7032 8630 7041
rect 8574 6967 8630 6976
rect 8482 6896 8538 6905
rect 8482 6831 8484 6840
rect 8536 6831 8538 6840
rect 8484 6802 8536 6808
rect 8588 6458 8616 6967
rect 8680 6866 8708 13738
rect 8772 13161 8800 14214
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 8852 13864 8904 13870
rect 8850 13832 8852 13841
rect 8904 13832 8906 13841
rect 8850 13767 8906 13776
rect 9048 13258 9076 13874
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 8758 13152 8814 13161
rect 8758 13087 8814 13096
rect 9048 12714 9076 13194
rect 9140 12832 9168 21247
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9232 17134 9260 19110
rect 9220 17128 9272 17134
rect 9220 17070 9272 17076
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 9232 16114 9260 16934
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9232 15910 9260 16050
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 9232 14958 9260 15846
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 9232 12986 9260 14894
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9140 12804 9260 12832
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 9048 12442 9076 12650
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8772 11898 8800 12174
rect 9232 12102 9260 12804
rect 9220 12096 9272 12102
rect 9140 12056 9220 12084
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8850 11112 8906 11121
rect 8850 11047 8906 11056
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8574 5808 8630 5817
rect 8574 5743 8576 5752
rect 8628 5743 8630 5752
rect 8576 5714 8628 5720
rect 8036 4134 8156 4162
rect 8220 5596 8432 5624
rect 8220 4146 8248 5596
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8680 4214 8708 4490
rect 8668 4208 8720 4214
rect 8668 4150 8720 4156
rect 8208 4140 8260 4146
rect 8036 4010 8064 4134
rect 8208 4082 8260 4088
rect 8024 4004 8076 4010
rect 8024 3946 8076 3952
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7930 3632 7986 3641
rect 7930 3567 7986 3576
rect 7944 3466 7972 3567
rect 7932 3460 7984 3466
rect 7932 3402 7984 3408
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 8036 3097 8064 3334
rect 8220 3194 8248 4082
rect 8300 4004 8352 4010
rect 8300 3946 8352 3952
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8022 3088 8078 3097
rect 8022 3023 8078 3032
rect 8312 2650 8340 3946
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8404 2553 8432 2790
rect 8390 2544 8446 2553
rect 8116 2508 8168 2514
rect 8390 2479 8446 2488
rect 8116 2450 8168 2456
rect 8128 2009 8156 2450
rect 8496 2145 8524 3470
rect 8772 2990 8800 3470
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8576 2576 8628 2582
rect 8574 2544 8576 2553
rect 8628 2544 8630 2553
rect 8574 2479 8630 2488
rect 8482 2136 8538 2145
rect 8482 2071 8538 2080
rect 8114 2000 8170 2009
rect 8114 1935 8170 1944
rect 7852 1414 8248 1442
rect 7484 1278 7696 1306
rect 7668 480 7696 1278
rect 8220 480 8248 1414
rect 8864 480 8892 11047
rect 9140 9704 9168 12056
rect 9220 12038 9272 12044
rect 9324 11898 9352 22374
rect 9508 22137 9536 23695
rect 10612 23662 10640 24210
rect 9864 23656 9916 23662
rect 9864 23598 9916 23604
rect 10600 23656 10652 23662
rect 10600 23598 10652 23604
rect 9876 23322 9904 23598
rect 10704 23497 10732 25758
rect 11072 24993 11100 27520
rect 11058 24984 11114 24993
rect 11058 24919 11114 24928
rect 11518 24848 11574 24857
rect 11716 24834 11744 27520
rect 12268 24834 12296 27520
rect 11518 24783 11574 24792
rect 11624 24806 11744 24834
rect 12176 24806 12296 24834
rect 10782 24712 10838 24721
rect 10782 24647 10838 24656
rect 10796 24410 10824 24647
rect 10784 24404 10836 24410
rect 10784 24346 10836 24352
rect 11336 23656 11388 23662
rect 11336 23598 11388 23604
rect 11426 23624 11482 23633
rect 10690 23488 10746 23497
rect 10289 23420 10585 23440
rect 10690 23423 10746 23432
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 9864 23316 9916 23322
rect 9864 23258 9916 23264
rect 9680 23180 9732 23186
rect 9680 23122 9732 23128
rect 9692 22438 9720 23122
rect 9680 22432 9732 22438
rect 9680 22374 9732 22380
rect 10968 22432 11020 22438
rect 10968 22374 11020 22380
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10876 22228 10928 22234
rect 10876 22170 10928 22176
rect 9494 22128 9550 22137
rect 9494 22063 9550 22072
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 9416 17202 9444 17614
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 9402 13560 9458 13569
rect 9402 13495 9404 13504
rect 9456 13495 9458 13504
rect 9404 13466 9456 13472
rect 9402 12608 9458 12617
rect 9402 12543 9458 12552
rect 9416 12442 9444 12543
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9324 10062 9352 10610
rect 9508 10470 9536 22063
rect 9588 21956 9640 21962
rect 9588 21898 9640 21904
rect 9600 19174 9628 21898
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9968 21078 9996 21830
rect 10888 21690 10916 22170
rect 10980 22114 11008 22374
rect 10980 22086 11100 22114
rect 10968 22024 11020 22030
rect 10968 21966 11020 21972
rect 10876 21684 10928 21690
rect 10876 21626 10928 21632
rect 10980 21434 11008 21966
rect 11072 21554 11100 22086
rect 11060 21548 11112 21554
rect 11060 21490 11112 21496
rect 10888 21418 11008 21434
rect 11244 21480 11296 21486
rect 11244 21422 11296 21428
rect 10876 21412 11008 21418
rect 10928 21406 11008 21412
rect 10876 21354 10928 21360
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 9956 21072 10008 21078
rect 9956 21014 10008 21020
rect 9772 21004 9824 21010
rect 9772 20946 9824 20952
rect 9784 20262 9812 20946
rect 9968 20618 9996 21014
rect 10888 20913 10916 21354
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 10874 20904 10930 20913
rect 10874 20839 10930 20848
rect 9968 20602 10088 20618
rect 9968 20596 10100 20602
rect 9968 20590 10048 20596
rect 10048 20538 10100 20544
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9784 19854 9812 20198
rect 10060 20058 10088 20538
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 10508 19848 10560 19854
rect 10508 19790 10560 19796
rect 10520 19514 10548 19790
rect 10508 19508 10560 19514
rect 10508 19450 10560 19456
rect 10980 19292 11008 21286
rect 11256 20806 11284 21422
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 11244 20800 11296 20806
rect 11244 20742 11296 20748
rect 11072 19990 11100 20742
rect 11060 19984 11112 19990
rect 11060 19926 11112 19932
rect 11072 19530 11100 19926
rect 11072 19502 11192 19530
rect 11072 19446 11100 19502
rect 11060 19440 11112 19446
rect 11060 19382 11112 19388
rect 11060 19304 11112 19310
rect 10980 19264 11060 19292
rect 11060 19246 11112 19252
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 9600 18970 9628 19110
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 10140 18896 10192 18902
rect 10140 18838 10192 18844
rect 9864 18624 9916 18630
rect 9864 18566 9916 18572
rect 9772 18352 9824 18358
rect 9772 18294 9824 18300
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9692 17898 9720 18226
rect 9600 17870 9720 17898
rect 9600 17066 9628 17870
rect 9784 17762 9812 18294
rect 9692 17734 9812 17762
rect 9588 17060 9640 17066
rect 9588 17002 9640 17008
rect 9600 16794 9628 17002
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9692 16674 9720 17734
rect 9600 16646 9720 16674
rect 9770 16688 9826 16697
rect 9600 15858 9628 16646
rect 9770 16623 9826 16632
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9692 16046 9720 16526
rect 9680 16040 9732 16046
rect 9678 16008 9680 16017
rect 9732 16008 9734 16017
rect 9678 15943 9734 15952
rect 9600 15830 9720 15858
rect 9588 14272 9640 14278
rect 9588 14214 9640 14220
rect 9600 13716 9628 14214
rect 9692 13818 9720 15830
rect 9784 14618 9812 16623
rect 9876 14618 9904 18566
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 9968 16794 9996 18022
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9968 15706 9996 16730
rect 10060 16046 10088 18362
rect 10152 18154 10180 18838
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10336 18426 10364 18702
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10600 18352 10652 18358
rect 10600 18294 10652 18300
rect 10612 18193 10640 18294
rect 10704 18290 10732 18566
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10598 18184 10654 18193
rect 10140 18148 10192 18154
rect 10598 18119 10654 18128
rect 10140 18090 10192 18096
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10704 17882 10732 18226
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10796 17746 10824 19110
rect 11072 18902 11100 19246
rect 11060 18896 11112 18902
rect 11060 18838 11112 18844
rect 11164 18834 11192 19502
rect 11256 18970 11284 20742
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11348 18850 11376 23598
rect 11426 23559 11482 23568
rect 11440 23526 11468 23559
rect 11428 23520 11480 23526
rect 11428 23462 11480 23468
rect 11532 23338 11560 24783
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 11256 18822 11376 18850
rect 11440 23310 11560 23338
rect 11256 18222 11284 18822
rect 11336 18692 11388 18698
rect 11336 18634 11388 18640
rect 11244 18216 11296 18222
rect 10874 18184 10930 18193
rect 11244 18158 11296 18164
rect 10874 18119 10930 18128
rect 10968 18148 11020 18154
rect 10888 18086 10916 18119
rect 10968 18090 11020 18096
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10138 17640 10194 17649
rect 10138 17575 10140 17584
rect 10192 17575 10194 17584
rect 10140 17546 10192 17552
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10152 16590 10180 16934
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 10060 15570 10088 15982
rect 10152 15706 10180 16526
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10704 15586 10732 17478
rect 10796 16794 10824 17682
rect 10888 17542 10916 18022
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10980 16561 11008 18090
rect 11348 18086 11376 18634
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11244 17536 11296 17542
rect 11244 17478 11296 17484
rect 11256 17338 11284 17478
rect 11244 17332 11296 17338
rect 11244 17274 11296 17280
rect 11256 16590 11284 17274
rect 11244 16584 11296 16590
rect 10966 16552 11022 16561
rect 10966 16487 11022 16496
rect 11150 16552 11206 16561
rect 11244 16526 11296 16532
rect 11150 16487 11206 16496
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10796 15609 10824 15642
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 10152 15558 10732 15586
rect 10782 15600 10838 15609
rect 10060 15162 10088 15506
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9770 14104 9826 14113
rect 9770 14039 9772 14048
rect 9824 14039 9826 14048
rect 9772 14010 9824 14016
rect 9876 14006 9904 14554
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9968 14074 9996 14418
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 10060 13938 10088 15098
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9692 13790 9904 13818
rect 9600 13688 9812 13716
rect 9784 13002 9812 13688
rect 9876 13190 9904 13790
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9784 12974 9904 13002
rect 9876 12753 9904 12974
rect 9862 12744 9918 12753
rect 9862 12679 9918 12688
rect 9876 12442 9904 12679
rect 9956 12640 10008 12646
rect 10060 12617 10088 13262
rect 9956 12582 10008 12588
rect 10046 12608 10102 12617
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9968 12306 9996 12582
rect 10046 12543 10102 12552
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9954 12200 10010 12209
rect 9954 12135 10010 12144
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9600 11937 9628 12038
rect 9586 11928 9642 11937
rect 9586 11863 9642 11872
rect 9692 11694 9720 12038
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9680 11688 9732 11694
rect 9600 11636 9680 11642
rect 9600 11630 9732 11636
rect 9600 11614 9720 11630
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9048 9676 9168 9704
rect 9048 9353 9076 9676
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9034 9344 9090 9353
rect 9034 9279 9090 9288
rect 9324 8906 9352 9522
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9310 7440 9366 7449
rect 9140 7398 9310 7426
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8956 5681 8984 6598
rect 8942 5672 8998 5681
rect 8942 5607 8998 5616
rect 8942 4992 8998 5001
rect 8942 4927 8998 4936
rect 8956 4826 8984 4927
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 9048 3738 9076 4762
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9048 2922 9076 3674
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 9140 2825 9168 7398
rect 9310 7375 9366 7384
rect 9310 7304 9366 7313
rect 9310 7239 9366 7248
rect 9218 7168 9274 7177
rect 9218 7103 9274 7112
rect 9232 6934 9260 7103
rect 9324 7002 9352 7239
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9220 6928 9272 6934
rect 9220 6870 9272 6876
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9324 5846 9352 6598
rect 9416 6458 9444 8366
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9416 5778 9444 6394
rect 9220 5772 9272 5778
rect 9220 5714 9272 5720
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 9232 5302 9260 5714
rect 9402 5672 9458 5681
rect 9402 5607 9404 5616
rect 9456 5607 9458 5616
rect 9404 5578 9456 5584
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 9232 4826 9260 5238
rect 9416 5166 9444 5578
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9220 4072 9272 4078
rect 9508 4049 9536 10406
rect 9600 9654 9628 11614
rect 9876 11354 9904 11698
rect 9968 11354 9996 12135
rect 10048 11620 10100 11626
rect 10048 11562 10100 11568
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9784 10810 9812 11154
rect 9862 11112 9918 11121
rect 9862 11047 9918 11056
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9692 10198 9720 10678
rect 9784 10266 9812 10746
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9692 9518 9720 10134
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9784 9586 9812 10066
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9876 9330 9904 11047
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9784 9302 9904 9330
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 9692 8090 9720 9046
rect 9680 8084 9732 8090
rect 9784 8072 9812 9302
rect 9968 9217 9996 10950
rect 9954 9208 10010 9217
rect 9954 9143 10010 9152
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9968 8809 9996 8978
rect 10060 8838 10088 11562
rect 10152 11014 10180 15558
rect 10782 15535 10838 15544
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10980 15162 11008 15438
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 11072 14414 11100 16186
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 11072 14074 11100 14350
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 13530 10732 13874
rect 10782 13560 10838 13569
rect 10692 13524 10744 13530
rect 10782 13495 10838 13504
rect 10692 13466 10744 13472
rect 10796 12889 10824 13495
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10782 12880 10838 12889
rect 10782 12815 10838 12824
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10888 12374 10916 13126
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10888 11558 10916 12310
rect 10980 11626 11008 13126
rect 10968 11620 11020 11626
rect 10968 11562 11020 11568
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10598 10840 10654 10849
rect 10598 10775 10654 10784
rect 10612 10538 10640 10775
rect 10796 10674 10824 10950
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10138 10296 10194 10305
rect 10289 10288 10585 10308
rect 10138 10231 10194 10240
rect 10048 8832 10100 8838
rect 9954 8800 10010 8809
rect 10048 8774 10100 8780
rect 9954 8735 10010 8744
rect 9784 8044 10088 8072
rect 9680 8026 9732 8032
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9864 7812 9916 7818
rect 9864 7754 9916 7760
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9692 7177 9720 7278
rect 9678 7168 9734 7177
rect 9678 7103 9734 7112
rect 9586 7032 9642 7041
rect 9580 6976 9586 7018
rect 9876 7002 9904 7754
rect 9968 7206 9996 7890
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9580 6967 9642 6976
rect 9864 6996 9916 7002
rect 9580 6882 9608 6967
rect 9864 6938 9916 6944
rect 9580 6866 9628 6882
rect 9580 6860 9640 6866
rect 9580 6854 9588 6860
rect 9588 6802 9640 6808
rect 9220 4014 9272 4020
rect 9494 4040 9550 4049
rect 9232 3777 9260 4014
rect 9312 4004 9364 4010
rect 9494 3975 9550 3984
rect 9312 3946 9364 3952
rect 9218 3768 9274 3777
rect 9218 3703 9220 3712
rect 9272 3703 9274 3712
rect 9220 3674 9272 3680
rect 9324 2854 9352 3946
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9416 3505 9444 3878
rect 9402 3496 9458 3505
rect 9402 3431 9458 3440
rect 9600 3380 9628 6802
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9416 3352 9628 3380
rect 9312 2848 9364 2854
rect 9126 2816 9182 2825
rect 9312 2790 9364 2796
rect 9126 2751 9182 2760
rect 9416 480 9444 3352
rect 9692 3210 9720 6666
rect 9864 6112 9916 6118
rect 9968 6089 9996 7142
rect 9864 6054 9916 6060
rect 9954 6080 10010 6089
rect 9876 5953 9904 6054
rect 9954 6015 10010 6024
rect 9862 5944 9918 5953
rect 9862 5879 9918 5888
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9968 5370 9996 5714
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9508 3182 9720 3210
rect 9784 3194 9812 4490
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9968 3738 9996 4082
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 9862 3496 9918 3505
rect 9862 3431 9918 3440
rect 9772 3188 9824 3194
rect 9508 2514 9536 3182
rect 9772 3130 9824 3136
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 9678 3088 9734 3097
rect 9600 2990 9628 3062
rect 9678 3023 9734 3032
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9600 2650 9628 2926
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9600 2446 9628 2586
rect 9692 2582 9720 3023
rect 9876 2650 9904 3431
rect 9968 3126 9996 3674
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 10060 2972 10088 8044
rect 10152 7886 10180 10231
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10336 9722 10364 9862
rect 10888 9738 10916 11494
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 11072 10810 11100 11222
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11072 10266 11100 10746
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10704 9710 10916 9738
rect 10600 9648 10652 9654
rect 10598 9616 10600 9625
rect 10652 9616 10654 9625
rect 10598 9551 10654 9560
rect 10612 9518 10640 9551
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10244 8634 10272 8910
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10152 7274 10180 7822
rect 10140 7268 10192 7274
rect 10140 7210 10192 7216
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10704 6610 10732 9710
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10796 9178 10824 9318
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10888 8838 10916 9318
rect 10980 9110 11008 9862
rect 11058 9480 11114 9489
rect 11058 9415 11114 9424
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10876 8832 10928 8838
rect 11072 8809 11100 9415
rect 10876 8774 10928 8780
rect 11058 8800 11114 8809
rect 10888 8498 10916 8774
rect 11058 8735 11114 8744
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10796 7546 10824 7822
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10888 7410 10916 7686
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10784 7268 10836 7274
rect 10784 7210 10836 7216
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 10796 7177 10824 7210
rect 10782 7168 10838 7177
rect 11072 7154 11100 7210
rect 10782 7103 10838 7112
rect 10888 7126 11100 7154
rect 10888 6730 10916 7126
rect 11060 6792 11112 6798
rect 10980 6740 11060 6746
rect 10980 6734 11112 6740
rect 10876 6724 10928 6730
rect 10876 6666 10928 6672
rect 10980 6718 11100 6734
rect 10980 6633 11008 6718
rect 10966 6624 11022 6633
rect 10244 6361 10272 6598
rect 10704 6582 10916 6610
rect 10230 6352 10286 6361
rect 10230 6287 10286 6296
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10704 5370 10732 6190
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10690 4856 10746 4865
rect 10690 4791 10746 4800
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 10152 4049 10180 4422
rect 10704 4078 10732 4791
rect 10784 4752 10836 4758
rect 10782 4720 10784 4729
rect 10836 4720 10838 4729
rect 10782 4655 10838 4664
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10692 4072 10744 4078
rect 10138 4040 10194 4049
rect 10692 4014 10744 4020
rect 10138 3975 10194 3984
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10690 3768 10746 3777
rect 10690 3703 10692 3712
rect 10744 3703 10746 3712
rect 10692 3674 10744 3680
rect 10796 3618 10824 4558
rect 10704 3590 10824 3618
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 10152 3097 10180 3334
rect 10138 3088 10194 3097
rect 10138 3023 10194 3032
rect 9968 2944 10088 2972
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 9968 480 9996 2944
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10506 2272 10562 2281
rect 10506 2207 10562 2216
rect 10520 480 10548 2207
rect 10704 1737 10732 3590
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10796 3194 10824 3470
rect 10888 3398 10916 6582
rect 10966 6559 11022 6568
rect 10980 4826 11008 6559
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 11072 5914 11100 6122
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10966 4720 11022 4729
rect 10966 4655 11022 4664
rect 10980 4185 11008 4655
rect 10966 4176 11022 4185
rect 10966 4111 11022 4120
rect 11072 3754 11100 5306
rect 10980 3738 11100 3754
rect 10968 3732 11100 3738
rect 11020 3726 11100 3732
rect 10968 3674 11020 3680
rect 10876 3392 10928 3398
rect 11072 3369 11100 3726
rect 10876 3334 10928 3340
rect 11058 3360 11114 3369
rect 11058 3295 11114 3304
rect 11164 3210 11192 16487
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11256 15162 11284 15642
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11348 13530 11376 18022
rect 11440 17898 11468 23310
rect 11518 21992 11574 22001
rect 11518 21927 11574 21936
rect 11532 21894 11560 21927
rect 11520 21888 11572 21894
rect 11520 21830 11572 21836
rect 11532 21350 11560 21830
rect 11520 21344 11572 21350
rect 11520 21286 11572 21292
rect 11624 18193 11652 24806
rect 11980 24268 12032 24274
rect 11980 24210 12032 24216
rect 11992 23526 12020 24210
rect 11980 23520 12032 23526
rect 11980 23462 12032 23468
rect 11704 20800 11756 20806
rect 11704 20742 11756 20748
rect 11716 19825 11744 20742
rect 11702 19816 11758 19825
rect 11702 19751 11758 19760
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11808 18970 11836 19110
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 11992 18737 12020 23462
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 12084 20942 12112 21490
rect 12072 20936 12124 20942
rect 12072 20878 12124 20884
rect 12084 20602 12112 20878
rect 12072 20596 12124 20602
rect 12072 20538 12124 20544
rect 12084 20330 12112 20538
rect 12176 20505 12204 24806
rect 12254 24168 12310 24177
rect 12254 24103 12256 24112
rect 12308 24103 12310 24112
rect 12256 24074 12308 24080
rect 12624 23520 12676 23526
rect 12624 23462 12676 23468
rect 12348 21344 12400 21350
rect 12348 21286 12400 21292
rect 12162 20496 12218 20505
rect 12162 20431 12218 20440
rect 12072 20324 12124 20330
rect 12072 20266 12124 20272
rect 12084 20058 12112 20266
rect 12072 20052 12124 20058
rect 12072 19994 12124 20000
rect 12360 18970 12388 21286
rect 12636 21049 12664 23462
rect 12622 21040 12678 21049
rect 12622 20975 12678 20984
rect 12622 20904 12678 20913
rect 12820 20890 12848 27520
rect 13372 23866 13400 27520
rect 13924 27418 13952 27520
rect 13924 27390 14044 27418
rect 13360 23860 13412 23866
rect 13360 23802 13412 23808
rect 13820 23520 13872 23526
rect 13450 23488 13506 23497
rect 13820 23462 13872 23468
rect 13450 23423 13506 23432
rect 13084 23180 13136 23186
rect 13084 23122 13136 23128
rect 12898 23080 12954 23089
rect 12898 23015 12900 23024
rect 12952 23015 12954 23024
rect 12900 22986 12952 22992
rect 13096 22438 13124 23122
rect 13358 22536 13414 22545
rect 13358 22471 13360 22480
rect 13412 22471 13414 22480
rect 13360 22442 13412 22448
rect 13084 22432 13136 22438
rect 13084 22374 13136 22380
rect 13096 22234 13124 22374
rect 13084 22228 13136 22234
rect 13084 22170 13136 22176
rect 12678 20862 12848 20890
rect 12622 20839 12678 20848
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 12452 19514 12480 20334
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12348 18964 12400 18970
rect 12348 18906 12400 18912
rect 12254 18864 12310 18873
rect 12254 18799 12310 18808
rect 11978 18728 12034 18737
rect 11978 18663 12034 18672
rect 12268 18290 12296 18799
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 11610 18184 11666 18193
rect 11610 18119 11666 18128
rect 11612 18080 11664 18086
rect 11612 18022 11664 18028
rect 11440 17870 11560 17898
rect 11428 17808 11480 17814
rect 11428 17750 11480 17756
rect 11440 16998 11468 17750
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11440 15609 11468 16934
rect 11426 15600 11482 15609
rect 11426 15535 11482 15544
rect 11440 15502 11468 15535
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11532 13530 11560 17870
rect 11624 15638 11652 18022
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11716 16182 11744 16526
rect 11992 16250 12020 16594
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11704 16176 11756 16182
rect 11704 16118 11756 16124
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11624 15162 11652 15574
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11256 11121 11284 12922
rect 11532 12850 11560 13466
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11624 12986 11652 13330
rect 11796 13320 11848 13326
rect 11980 13320 12032 13326
rect 11848 13280 11928 13308
rect 11796 13262 11848 13268
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11900 12889 11928 13280
rect 11980 13262 12032 13268
rect 11992 13161 12020 13262
rect 11978 13152 12034 13161
rect 11978 13087 12034 13096
rect 11992 12986 12020 13087
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11886 12880 11942 12889
rect 11520 12844 11572 12850
rect 11886 12815 11942 12824
rect 11520 12786 11572 12792
rect 11532 12481 11560 12786
rect 11702 12608 11758 12617
rect 11702 12543 11758 12552
rect 11518 12472 11574 12481
rect 11518 12407 11574 12416
rect 11716 12306 11744 12543
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11624 11937 11652 12242
rect 11610 11928 11666 11937
rect 11716 11898 11744 12242
rect 11900 12238 11928 12815
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11610 11863 11666 11872
rect 11704 11892 11756 11898
rect 11624 11694 11652 11863
rect 11704 11834 11756 11840
rect 11900 11830 11928 12174
rect 11888 11824 11940 11830
rect 11888 11766 11940 11772
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11348 11286 11376 11494
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11900 11218 11928 11630
rect 11888 11212 11940 11218
rect 11808 11172 11888 11200
rect 11242 11112 11298 11121
rect 11242 11047 11298 11056
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11612 8832 11664 8838
rect 11612 8774 11664 8780
rect 11428 8356 11480 8362
rect 11428 8298 11480 8304
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11256 5370 11284 7686
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 11242 5264 11298 5273
rect 11242 5199 11244 5208
rect 11296 5199 11298 5208
rect 11244 5170 11296 5176
rect 11242 4992 11298 5001
rect 11242 4927 11298 4936
rect 11256 4593 11284 4927
rect 11242 4584 11298 4593
rect 11242 4519 11298 4528
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11256 3913 11284 4014
rect 11242 3904 11298 3913
rect 11242 3839 11298 3848
rect 11256 3738 11284 3839
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11348 3618 11376 7686
rect 11440 4740 11468 8298
rect 11624 7886 11652 8774
rect 11716 8090 11744 9318
rect 11808 8974 11836 11172
rect 11888 11154 11940 11160
rect 12084 10452 12112 16934
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 12452 15314 12480 15438
rect 12360 15286 12480 15314
rect 12360 15162 12388 15286
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12162 14376 12218 14385
rect 12162 14311 12218 14320
rect 12176 10606 12204 14311
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12254 13968 12310 13977
rect 12254 13903 12256 13912
rect 12308 13903 12310 13912
rect 12438 13968 12494 13977
rect 12438 13903 12494 13912
rect 12256 13874 12308 13880
rect 12452 13530 12480 13903
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12346 13016 12402 13025
rect 12346 12951 12402 12960
rect 12360 12442 12388 12951
rect 12452 12782 12480 13126
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12544 12646 12572 14214
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12438 12336 12494 12345
rect 12348 12300 12400 12306
rect 12438 12271 12494 12280
rect 12348 12242 12400 12248
rect 12360 12073 12388 12242
rect 12346 12064 12402 12073
rect 12346 11999 12402 12008
rect 12452 10849 12480 12271
rect 12544 11558 12572 12378
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12544 11354 12572 11494
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12438 10840 12494 10849
rect 12438 10775 12494 10784
rect 12164 10600 12216 10606
rect 12162 10568 12164 10577
rect 12216 10568 12218 10577
rect 12162 10503 12218 10512
rect 12084 10424 12204 10452
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11900 9042 11928 9522
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11808 8362 11836 8910
rect 11796 8356 11848 8362
rect 11796 8298 11848 8304
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11520 6928 11572 6934
rect 11520 6870 11572 6876
rect 11532 6118 11560 6870
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11520 6112 11572 6118
rect 11518 6080 11520 6089
rect 11572 6080 11574 6089
rect 11518 6015 11574 6024
rect 11624 5914 11652 6734
rect 11612 5908 11664 5914
rect 11664 5868 11744 5896
rect 11612 5850 11664 5856
rect 11610 5128 11666 5137
rect 11610 5063 11612 5072
rect 11664 5063 11666 5072
rect 11612 5034 11664 5040
rect 11440 4712 11652 4740
rect 11520 4616 11572 4622
rect 11426 4584 11482 4593
rect 11520 4558 11572 4564
rect 11426 4519 11482 4528
rect 11440 3942 11468 4519
rect 11532 4282 11560 4558
rect 11520 4276 11572 4282
rect 11520 4218 11572 4224
rect 11520 4004 11572 4010
rect 11520 3946 11572 3952
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 11072 3182 11192 3210
rect 11256 3590 11376 3618
rect 10796 2650 10824 3130
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10796 2446 10824 2586
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 10690 1728 10746 1737
rect 10690 1663 10746 1672
rect 10888 1329 10916 2994
rect 10966 2816 11022 2825
rect 10966 2751 11022 2760
rect 10980 2582 11008 2751
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 10874 1320 10930 1329
rect 10874 1255 10930 1264
rect 11072 480 11100 3182
rect 11256 2825 11284 3590
rect 11532 3482 11560 3946
rect 11624 3505 11652 4712
rect 11716 3738 11744 5868
rect 11808 4826 11836 7278
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11900 5681 11928 6394
rect 11886 5672 11942 5681
rect 11886 5607 11942 5616
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11808 4214 11836 4762
rect 11992 4758 12020 9454
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 12084 8090 12112 9114
rect 12176 8401 12204 10424
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12452 9568 12480 10066
rect 12544 9761 12572 10134
rect 12530 9752 12586 9761
rect 12530 9687 12586 9696
rect 12360 9540 12480 9568
rect 12360 9382 12388 9540
rect 12438 9480 12494 9489
rect 12438 9415 12494 9424
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12360 8922 12388 8978
rect 12452 8922 12480 9415
rect 12360 8894 12480 8922
rect 12162 8392 12218 8401
rect 12162 8327 12218 8336
rect 12452 8294 12480 8894
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12268 7546 12296 7822
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12452 7410 12480 8230
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12348 7200 12400 7206
rect 12162 7168 12218 7177
rect 12348 7142 12400 7148
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12162 7103 12218 7112
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 12084 5370 12112 5714
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 11980 4752 12032 4758
rect 11980 4694 12032 4700
rect 11992 4282 12020 4694
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 12084 3670 12112 5306
rect 12176 4570 12204 7103
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12268 4758 12296 6598
rect 12360 5166 12388 7142
rect 12452 6905 12480 7142
rect 12438 6896 12494 6905
rect 12438 6831 12494 6840
rect 12636 6746 12664 20839
rect 12716 19508 12768 19514
rect 12716 19450 12768 19456
rect 12728 18834 12756 19450
rect 12900 19168 12952 19174
rect 12898 19136 12900 19145
rect 12952 19136 12954 19145
rect 12898 19071 12954 19080
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12716 18624 12768 18630
rect 12768 18572 12848 18578
rect 12716 18566 12848 18572
rect 12728 18550 12848 18566
rect 12820 18086 12848 18550
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12820 16114 12848 18022
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12808 15632 12860 15638
rect 12808 15574 12860 15580
rect 12820 14822 12848 15574
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12716 14408 12768 14414
rect 12716 14350 12768 14356
rect 12728 14006 12756 14350
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12728 12714 12756 13466
rect 12716 12708 12768 12714
rect 12716 12650 12768 12656
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12728 8022 12756 10406
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12820 7342 12848 14758
rect 12912 12918 12940 19071
rect 12992 18896 13044 18902
rect 12992 18838 13044 18844
rect 13004 17882 13032 18838
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 12990 17776 13046 17785
rect 12990 17711 13046 17720
rect 12900 12912 12952 12918
rect 12900 12854 12952 12860
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12912 11354 12940 12718
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12898 10296 12954 10305
rect 12898 10231 12900 10240
rect 12952 10231 12954 10240
rect 12900 10202 12952 10208
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12912 9722 12940 9998
rect 12900 9716 12952 9722
rect 12900 9658 12952 9664
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12636 6718 12756 6746
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12636 6254 12664 6598
rect 12624 6248 12676 6254
rect 12530 6216 12586 6225
rect 12624 6190 12676 6196
rect 12530 6151 12586 6160
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12452 5953 12480 6054
rect 12438 5944 12494 5953
rect 12438 5879 12494 5888
rect 12544 5794 12572 6151
rect 12636 5914 12664 6190
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12452 5778 12572 5794
rect 12440 5772 12572 5778
rect 12492 5766 12572 5772
rect 12440 5714 12492 5720
rect 12452 5370 12480 5714
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12256 4752 12308 4758
rect 12256 4694 12308 4700
rect 12176 4542 12296 4570
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 11348 3454 11560 3482
rect 11610 3496 11666 3505
rect 11242 2816 11298 2825
rect 11242 2751 11298 2760
rect 11150 2680 11206 2689
rect 11348 2650 11376 3454
rect 11610 3431 11666 3440
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11428 2848 11480 2854
rect 11426 2816 11428 2825
rect 11480 2816 11482 2825
rect 11426 2751 11482 2760
rect 11150 2615 11206 2624
rect 11336 2644 11388 2650
rect 11164 2378 11192 2615
rect 11336 2586 11388 2592
rect 11152 2372 11204 2378
rect 11152 2314 11204 2320
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 6366 368 6422 377
rect 6366 303 6422 312
rect 6550 0 6606 480
rect 7102 0 7158 480
rect 7654 0 7710 480
rect 8206 0 8262 480
rect 8850 0 8906 480
rect 9402 0 9458 480
rect 9954 0 10010 480
rect 10506 0 10562 480
rect 11058 0 11114 480
rect 11624 105 11652 2246
rect 11716 480 11744 3334
rect 12084 3194 12112 3606
rect 12162 3360 12218 3369
rect 12162 3295 12218 3304
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12176 2650 12204 3295
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 11980 2440 12032 2446
rect 11978 2408 11980 2417
rect 12032 2408 12034 2417
rect 11978 2343 12034 2352
rect 12162 2408 12218 2417
rect 12162 2343 12218 2352
rect 12176 2009 12204 2343
rect 12162 2000 12218 2009
rect 12162 1935 12218 1944
rect 12268 480 12296 4542
rect 12452 4026 12480 4966
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12544 4214 12572 4422
rect 12636 4282 12664 5102
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12728 4146 12756 6718
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 12912 6118 12940 6666
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12912 5681 12940 6054
rect 12898 5672 12954 5681
rect 12898 5607 12954 5616
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12820 4457 12848 4762
rect 12806 4448 12862 4457
rect 12806 4383 12862 4392
rect 13004 4146 13032 17711
rect 13096 12345 13124 22170
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 13372 21078 13400 21830
rect 13360 21072 13412 21078
rect 13360 21014 13412 21020
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 13188 19378 13216 19654
rect 13280 19417 13308 19790
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13266 19408 13322 19417
rect 13176 19372 13228 19378
rect 13266 19343 13322 19352
rect 13176 19314 13228 19320
rect 13280 19310 13308 19343
rect 13268 19304 13320 19310
rect 13372 19281 13400 19654
rect 13268 19246 13320 19252
rect 13358 19272 13414 19281
rect 13358 19207 13414 19216
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13280 18834 13308 19110
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 13280 18086 13308 18770
rect 13268 18080 13320 18086
rect 13268 18022 13320 18028
rect 13280 17542 13308 18022
rect 13464 17882 13492 23423
rect 13636 22976 13688 22982
rect 13636 22918 13688 22924
rect 13648 22438 13676 22918
rect 13544 22432 13596 22438
rect 13544 22374 13596 22380
rect 13636 22432 13688 22438
rect 13636 22374 13688 22380
rect 13556 22234 13584 22374
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13648 22166 13676 22374
rect 13636 22160 13688 22166
rect 13636 22102 13688 22108
rect 13636 22024 13688 22030
rect 13636 21966 13688 21972
rect 13726 21992 13782 22001
rect 13648 21146 13676 21966
rect 13726 21927 13728 21936
rect 13780 21927 13782 21936
rect 13728 21898 13780 21904
rect 13740 21690 13768 21898
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13740 21350 13768 21490
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13636 20256 13688 20262
rect 13636 20198 13688 20204
rect 13740 20210 13768 21286
rect 13832 20369 13860 23462
rect 14016 21570 14044 27390
rect 14278 24440 14334 24449
rect 14278 24375 14280 24384
rect 14332 24375 14334 24384
rect 14280 24346 14332 24352
rect 14096 24268 14148 24274
rect 14096 24210 14148 24216
rect 14108 23866 14136 24210
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 14108 23322 14136 23802
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 14280 23180 14332 23186
rect 14280 23122 14332 23128
rect 14292 22982 14320 23122
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 13924 21554 14044 21570
rect 13912 21548 14044 21554
rect 13964 21542 14044 21548
rect 14094 21584 14150 21593
rect 14094 21519 14150 21528
rect 13912 21490 13964 21496
rect 14004 21480 14056 21486
rect 14108 21434 14136 21519
rect 14056 21428 14136 21434
rect 14004 21422 14136 21428
rect 14188 21480 14240 21486
rect 14188 21422 14240 21428
rect 13912 21412 13964 21418
rect 14016 21406 14136 21422
rect 13912 21354 13964 21360
rect 13818 20360 13874 20369
rect 13818 20295 13874 20304
rect 13648 19242 13676 20198
rect 13740 20182 13860 20210
rect 13728 19780 13780 19786
rect 13728 19722 13780 19728
rect 13740 19446 13768 19722
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13636 19236 13688 19242
rect 13636 19178 13688 19184
rect 13648 18902 13676 19178
rect 13740 18970 13768 19382
rect 13728 18964 13780 18970
rect 13728 18906 13780 18912
rect 13636 18896 13688 18902
rect 13636 18838 13688 18844
rect 13832 18630 13860 20182
rect 13924 19854 13952 21354
rect 14004 21004 14056 21010
rect 14004 20946 14056 20952
rect 14016 20330 14044 20946
rect 14004 20324 14056 20330
rect 14004 20266 14056 20272
rect 14004 19916 14056 19922
rect 14004 19858 14056 19864
rect 13912 19848 13964 19854
rect 13912 19790 13964 19796
rect 13924 19378 13952 19790
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 14016 18426 14044 19858
rect 14108 18902 14136 21406
rect 14200 21350 14228 21422
rect 14188 21344 14240 21350
rect 14188 21286 14240 21292
rect 14200 19310 14228 21286
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14200 19174 14228 19246
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 14004 18420 14056 18426
rect 14004 18362 14056 18368
rect 13728 18216 13780 18222
rect 13728 18158 13780 18164
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13636 17876 13688 17882
rect 13636 17818 13688 17824
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13280 17134 13308 17478
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 13280 16046 13308 17070
rect 13372 16998 13400 17682
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13360 16992 13412 16998
rect 13360 16934 13412 16940
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 13464 15570 13492 17478
rect 13648 16726 13676 17818
rect 13740 17354 13768 18158
rect 13818 17776 13874 17785
rect 13818 17711 13820 17720
rect 13872 17711 13874 17720
rect 13820 17682 13872 17688
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 13740 17338 13952 17354
rect 13740 17332 13964 17338
rect 13740 17326 13912 17332
rect 13912 17274 13964 17280
rect 13636 16720 13688 16726
rect 13636 16662 13688 16668
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 13188 15162 13216 15438
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 13188 13530 13216 14826
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13188 12866 13216 13466
rect 13372 13190 13400 14418
rect 13648 13818 13676 16662
rect 13924 15978 13952 17274
rect 14016 17066 14044 17614
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 14016 16794 14044 17002
rect 14004 16788 14056 16794
rect 14004 16730 14056 16736
rect 13912 15972 13964 15978
rect 13912 15914 13964 15920
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13740 14958 13768 15846
rect 13924 15706 13952 15914
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 14108 14618 14136 14826
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 14096 14340 14148 14346
rect 14096 14282 14148 14288
rect 13556 13790 13676 13818
rect 14002 13832 14058 13841
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13188 12850 13308 12866
rect 13176 12844 13308 12850
rect 13228 12838 13308 12844
rect 13176 12786 13228 12792
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 13188 12442 13216 12650
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 13082 12336 13138 12345
rect 13280 12322 13308 12838
rect 13372 12442 13400 13126
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 13280 12294 13400 12322
rect 13082 12271 13138 12280
rect 13096 11098 13124 12271
rect 13372 12238 13400 12294
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13464 12170 13492 13466
rect 13556 12866 13584 13790
rect 14002 13767 14058 13776
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 13648 12986 13676 13670
rect 13740 13530 13768 13670
rect 14016 13530 14044 13767
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14016 12986 14044 13466
rect 14108 13326 14136 14282
rect 14200 14074 14228 15506
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14292 13433 14320 22918
rect 14370 22400 14426 22409
rect 14370 22335 14426 22344
rect 14384 15706 14412 22335
rect 14464 21888 14516 21894
rect 14464 21830 14516 21836
rect 14476 21418 14504 21830
rect 14464 21412 14516 21418
rect 14464 21354 14516 21360
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 14476 19310 14504 19654
rect 14568 19417 14596 27520
rect 15120 25242 15148 27520
rect 14844 25214 15148 25242
rect 14648 23520 14700 23526
rect 14648 23462 14700 23468
rect 14660 20330 14688 23462
rect 14844 21026 14872 25214
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15476 24268 15528 24274
rect 15476 24210 15528 24216
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15200 23792 15252 23798
rect 15198 23760 15200 23769
rect 15252 23760 15254 23769
rect 15198 23695 15254 23704
rect 15488 23526 15516 24210
rect 15672 23866 15700 27520
rect 16224 24970 16252 27520
rect 16132 24942 16252 24970
rect 16028 24744 16080 24750
rect 16028 24686 16080 24692
rect 15660 23860 15712 23866
rect 15660 23802 15712 23808
rect 15476 23520 15528 23526
rect 15476 23462 15528 23468
rect 15658 23488 15714 23497
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15200 22568 15252 22574
rect 15200 22510 15252 22516
rect 15108 22432 15160 22438
rect 15212 22409 15240 22510
rect 15304 22506 15332 23122
rect 15292 22500 15344 22506
rect 15292 22442 15344 22448
rect 15108 22374 15160 22380
rect 15198 22400 15254 22409
rect 15120 22098 15148 22374
rect 15198 22335 15254 22344
rect 15108 22092 15160 22098
rect 15108 22034 15160 22040
rect 15292 22024 15344 22030
rect 15292 21966 15344 21972
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15304 21350 15332 21966
rect 15292 21344 15344 21350
rect 15292 21286 15344 21292
rect 14752 21010 14872 21026
rect 14740 21004 14872 21010
rect 14792 20998 14872 21004
rect 14740 20946 14792 20952
rect 14648 20324 14700 20330
rect 14648 20266 14700 20272
rect 14752 20262 14780 20946
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14832 20324 14884 20330
rect 14832 20266 14884 20272
rect 14740 20256 14792 20262
rect 14740 20198 14792 20204
rect 14554 19408 14610 19417
rect 14554 19343 14610 19352
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14476 18698 14504 19246
rect 14556 18896 14608 18902
rect 14556 18838 14608 18844
rect 14464 18692 14516 18698
rect 14464 18634 14516 18640
rect 14476 18358 14504 18634
rect 14464 18352 14516 18358
rect 14464 18294 14516 18300
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14476 17882 14504 18158
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14462 17232 14518 17241
rect 14462 17167 14518 17176
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14384 14006 14412 14758
rect 14372 14000 14424 14006
rect 14372 13942 14424 13948
rect 14384 13870 14412 13942
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14278 13424 14334 13433
rect 14278 13359 14334 13368
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 13556 12838 13768 12866
rect 13636 12776 13688 12782
rect 13634 12744 13636 12753
rect 13688 12744 13690 12753
rect 13634 12679 13690 12688
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13372 11393 13400 12038
rect 13358 11384 13414 11393
rect 13358 11319 13360 11328
rect 13412 11319 13414 11328
rect 13360 11290 13412 11296
rect 13452 11280 13504 11286
rect 13452 11222 13504 11228
rect 13096 11070 13308 11098
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 13188 10674 13216 10950
rect 13280 10690 13308 11070
rect 13464 10810 13492 11222
rect 13556 10810 13584 12582
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 13176 10668 13228 10674
rect 13280 10662 13584 10690
rect 13176 10610 13228 10616
rect 13082 10568 13138 10577
rect 13082 10503 13084 10512
rect 13136 10503 13138 10512
rect 13084 10474 13136 10480
rect 13096 10198 13124 10474
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 13188 9489 13216 10610
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13174 9480 13230 9489
rect 13174 9415 13230 9424
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13188 8362 13216 8774
rect 13176 8356 13228 8362
rect 13176 8298 13228 8304
rect 13188 7886 13216 8298
rect 13280 8090 13308 9998
rect 13464 9450 13492 9998
rect 13452 9444 13504 9450
rect 13452 9386 13504 9392
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13372 8090 13400 9318
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13372 7546 13400 8026
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 13084 6792 13136 6798
rect 13082 6760 13084 6769
rect 13136 6760 13138 6769
rect 13082 6695 13138 6704
rect 13082 4992 13138 5001
rect 13082 4927 13138 4936
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12360 3998 12480 4026
rect 12360 3641 12388 3998
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12452 3777 12480 3878
rect 12438 3768 12494 3777
rect 12438 3703 12494 3712
rect 12346 3632 12402 3641
rect 12346 3567 12402 3576
rect 12360 2990 12388 3567
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12820 480 12848 3878
rect 12992 2644 13044 2650
rect 13096 2632 13124 4927
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 13188 3398 13216 4558
rect 13280 4146 13308 4626
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13044 2604 13124 2632
rect 12992 2586 13044 2592
rect 13280 2446 13308 4082
rect 13268 2440 13320 2446
rect 13174 2408 13230 2417
rect 13268 2382 13320 2388
rect 13174 2343 13176 2352
rect 13228 2343 13230 2352
rect 13176 2314 13228 2320
rect 13372 480 13400 7278
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 13464 6118 13492 6802
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13464 5817 13492 6054
rect 13450 5808 13506 5817
rect 13450 5743 13506 5752
rect 13556 5692 13584 10662
rect 13648 7410 13676 12582
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13648 6390 13676 6734
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13648 5817 13676 6326
rect 13634 5808 13690 5817
rect 13634 5743 13690 5752
rect 13464 5664 13584 5692
rect 13464 3942 13492 5664
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13648 5273 13676 5510
rect 13740 5409 13768 12838
rect 14108 12782 14136 13262
rect 14292 12850 14320 13262
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14476 12594 14504 17167
rect 14108 12566 14504 12594
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 13924 11898 13952 12378
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13924 11218 13952 11834
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 13912 11212 13964 11218
rect 13832 11172 13912 11200
rect 13832 10742 13860 11172
rect 13912 11154 13964 11160
rect 13912 11076 13964 11082
rect 13912 11018 13964 11024
rect 13820 10736 13872 10742
rect 13924 10713 13952 11018
rect 13820 10678 13872 10684
rect 13910 10704 13966 10713
rect 13832 10266 13860 10678
rect 13910 10639 13966 10648
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13912 9444 13964 9450
rect 13912 9386 13964 9392
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13832 8430 13860 9318
rect 13924 8838 13952 9386
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13924 8634 13952 8774
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13924 6866 13952 7822
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13726 5400 13782 5409
rect 13726 5335 13782 5344
rect 13634 5264 13690 5273
rect 13634 5199 13690 5208
rect 13648 5098 13676 5199
rect 13740 5137 13768 5335
rect 13726 5128 13782 5137
rect 13636 5092 13688 5098
rect 13726 5063 13782 5072
rect 13636 5034 13688 5040
rect 13648 4690 13676 5034
rect 13728 4820 13780 4826
rect 13832 4808 13860 6666
rect 13912 5636 13964 5642
rect 13912 5578 13964 5584
rect 13780 4780 13860 4808
rect 13728 4762 13780 4768
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13556 2417 13584 4014
rect 13728 4004 13780 4010
rect 13832 3992 13860 4422
rect 13780 3964 13860 3992
rect 13728 3946 13780 3952
rect 13818 3904 13874 3913
rect 13818 3839 13874 3848
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 13648 2650 13676 3402
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13740 2922 13768 3334
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 13542 2408 13598 2417
rect 13542 2343 13598 2352
rect 13740 2009 13768 2858
rect 13832 2145 13860 3839
rect 13924 3233 13952 5578
rect 13910 3224 13966 3233
rect 13910 3159 13966 3168
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 13818 2136 13874 2145
rect 13818 2071 13874 2080
rect 13726 2000 13782 2009
rect 13726 1935 13782 1944
rect 13924 480 13952 3062
rect 14016 2650 14044 11630
rect 14108 7410 14136 12566
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14476 11898 14504 12174
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14568 11830 14596 18838
rect 14646 15464 14702 15473
rect 14646 15399 14648 15408
rect 14700 15399 14702 15408
rect 14648 15370 14700 15376
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14660 14074 14688 14214
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 14660 12617 14688 12922
rect 14646 12608 14702 12617
rect 14646 12543 14702 12552
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 14462 11520 14518 11529
rect 14462 11455 14518 11464
rect 14280 11076 14332 11082
rect 14280 11018 14332 11024
rect 14292 10033 14320 11018
rect 14370 10704 14426 10713
rect 14476 10674 14504 11455
rect 14370 10639 14426 10648
rect 14464 10668 14516 10674
rect 14384 10606 14412 10639
rect 14464 10610 14516 10616
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14476 10266 14504 10610
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14372 10192 14424 10198
rect 14370 10160 14372 10169
rect 14424 10160 14426 10169
rect 14370 10095 14426 10104
rect 14278 10024 14334 10033
rect 14278 9959 14334 9968
rect 14568 9738 14596 11766
rect 14752 11694 14780 20198
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14740 11552 14792 11558
rect 14844 11540 14872 20266
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15488 19145 15516 23462
rect 15658 23423 15714 23432
rect 15568 22976 15620 22982
rect 15566 22944 15568 22953
rect 15620 22944 15622 22953
rect 15566 22879 15622 22888
rect 15672 22778 15700 23423
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15752 22500 15804 22506
rect 15752 22442 15804 22448
rect 15568 22092 15620 22098
rect 15568 22034 15620 22040
rect 15580 21690 15608 22034
rect 15568 21684 15620 21690
rect 15568 21626 15620 21632
rect 15580 21146 15608 21626
rect 15568 21140 15620 21146
rect 15568 21082 15620 21088
rect 15580 20942 15608 21082
rect 15568 20936 15620 20942
rect 15568 20878 15620 20884
rect 15580 20602 15608 20878
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15474 19136 15530 19145
rect 15474 19071 15530 19080
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15304 18222 15332 18702
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15566 16008 15622 16017
rect 15566 15943 15622 15952
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 15120 15609 15148 15846
rect 15106 15600 15162 15609
rect 15106 15535 15162 15544
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15304 13977 15332 14214
rect 15290 13968 15346 13977
rect 15290 13903 15346 13912
rect 15396 13870 15424 14758
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 14936 13530 14964 13806
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 14924 13524 14976 13530
rect 14924 13466 14976 13472
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15304 12782 15332 13738
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15014 11656 15070 11665
rect 15014 11591 15070 11600
rect 15028 11558 15056 11591
rect 14792 11512 14872 11540
rect 15016 11552 15068 11558
rect 14740 11494 14792 11500
rect 15016 11494 15068 11500
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 14648 11280 14700 11286
rect 14646 11248 14648 11257
rect 14700 11248 14702 11257
rect 14646 11183 14702 11192
rect 14648 11008 14700 11014
rect 14646 10976 14648 10985
rect 14700 10976 14702 10985
rect 14646 10911 14702 10920
rect 14646 10840 14702 10849
rect 14646 10775 14702 10784
rect 14660 10169 14688 10775
rect 14646 10160 14702 10169
rect 14646 10095 14702 10104
rect 14476 9710 14596 9738
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14200 8673 14228 8774
rect 14186 8664 14242 8673
rect 14186 8599 14242 8608
rect 14278 8392 14334 8401
rect 14278 8327 14334 8336
rect 14292 7410 14320 8327
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14108 7041 14136 7346
rect 14094 7032 14150 7041
rect 14094 6967 14096 6976
rect 14148 6967 14150 6976
rect 14096 6938 14148 6944
rect 14108 6907 14136 6938
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14108 5642 14136 6802
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14186 6080 14242 6089
rect 14186 6015 14242 6024
rect 14096 5636 14148 5642
rect 14096 5578 14148 5584
rect 14094 4720 14150 4729
rect 14094 4655 14096 4664
rect 14148 4655 14150 4664
rect 14096 4626 14148 4632
rect 14108 4282 14136 4626
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14108 3398 14136 4082
rect 14200 3738 14228 6015
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 14292 4185 14320 4422
rect 14278 4176 14334 4185
rect 14278 4111 14334 4120
rect 14384 3777 14412 6598
rect 14370 3768 14426 3777
rect 14188 3732 14240 3738
rect 14370 3703 14426 3712
rect 14188 3674 14240 3680
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14108 2922 14136 3334
rect 14476 3126 14504 9710
rect 14556 8832 14608 8838
rect 14554 8800 14556 8809
rect 14608 8800 14610 8809
rect 14554 8735 14610 8744
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 14464 3120 14516 3126
rect 14464 3062 14516 3068
rect 14096 2916 14148 2922
rect 14096 2858 14148 2864
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14476 921 14504 2246
rect 14462 912 14518 921
rect 14462 847 14518 856
rect 14568 480 14596 7278
rect 14648 6656 14700 6662
rect 14646 6624 14648 6633
rect 14700 6624 14702 6633
rect 14646 6559 14702 6568
rect 14752 6474 14780 11494
rect 15120 11370 15148 11494
rect 15028 11342 15148 11370
rect 15028 11150 15056 11342
rect 15016 11144 15068 11150
rect 15014 11112 15016 11121
rect 15068 11112 15070 11121
rect 15014 11047 15070 11056
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14924 9104 14976 9110
rect 14922 9072 14924 9081
rect 14976 9072 14978 9081
rect 14922 9007 14978 9016
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15304 8634 15332 8910
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14830 7032 14886 7041
rect 14830 6967 14886 6976
rect 14660 6446 14780 6474
rect 14660 3924 14688 6446
rect 14844 6254 14872 6967
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14832 6248 14884 6254
rect 14832 6190 14884 6196
rect 14844 5914 14872 6190
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14752 4078 14780 5510
rect 14844 5370 14872 5850
rect 15396 5658 15424 13670
rect 15488 12374 15516 15302
rect 15580 13734 15608 15943
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15568 13728 15620 13734
rect 15568 13670 15620 13676
rect 15568 13456 15620 13462
rect 15672 13433 15700 14418
rect 15568 13398 15620 13404
rect 15658 13424 15714 13433
rect 15580 12782 15608 13398
rect 15658 13359 15714 13368
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15658 12744 15714 12753
rect 15580 12442 15608 12718
rect 15658 12679 15660 12688
rect 15712 12679 15714 12688
rect 15660 12650 15712 12656
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15580 11762 15608 12242
rect 15660 12164 15712 12170
rect 15660 12106 15712 12112
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15488 10742 15516 11086
rect 15476 10736 15528 10742
rect 15476 10678 15528 10684
rect 15474 10024 15530 10033
rect 15474 9959 15530 9968
rect 15488 8634 15516 9959
rect 15580 9654 15608 11698
rect 15672 11218 15700 12106
rect 15764 11558 15792 22442
rect 16040 21457 16068 24686
rect 16132 24449 16160 24942
rect 16210 24848 16266 24857
rect 16210 24783 16266 24792
rect 16224 24614 16252 24783
rect 16776 24721 16804 27520
rect 16762 24712 16818 24721
rect 16762 24647 16818 24656
rect 16212 24608 16264 24614
rect 16212 24550 16264 24556
rect 16118 24440 16174 24449
rect 17222 24440 17278 24449
rect 16118 24375 16174 24384
rect 16488 24404 16540 24410
rect 17222 24375 17278 24384
rect 16488 24346 16540 24352
rect 16500 24313 16528 24346
rect 16486 24304 16542 24313
rect 16486 24239 16542 24248
rect 16764 24268 16816 24274
rect 16764 24210 16816 24216
rect 16580 23656 16632 23662
rect 16580 23598 16632 23604
rect 16592 21593 16620 23598
rect 16776 23526 16804 24210
rect 16764 23520 16816 23526
rect 16764 23462 16816 23468
rect 16776 22778 16804 23462
rect 17236 23322 17264 24375
rect 17420 23497 17448 27520
rect 17972 24857 18000 27520
rect 17958 24848 18014 24857
rect 17958 24783 18014 24792
rect 18524 24410 18552 27520
rect 18970 24712 19026 24721
rect 18970 24647 19026 24656
rect 18984 24410 19012 24647
rect 19076 24449 19104 27520
rect 19628 25786 19656 27520
rect 19536 25758 19656 25786
rect 19062 24440 19118 24449
rect 18512 24404 18564 24410
rect 18512 24346 18564 24352
rect 18972 24404 19024 24410
rect 19062 24375 19118 24384
rect 18972 24346 19024 24352
rect 17684 24268 17736 24274
rect 17684 24210 17736 24216
rect 19064 24268 19116 24274
rect 19064 24210 19116 24216
rect 17696 23526 17724 24210
rect 17774 24168 17830 24177
rect 17774 24103 17776 24112
rect 17828 24103 17830 24112
rect 17776 24074 17828 24080
rect 18326 23896 18382 23905
rect 18326 23831 18328 23840
rect 18380 23831 18382 23840
rect 18328 23802 18380 23808
rect 19076 23526 19104 24210
rect 19536 24177 19564 25758
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19522 24168 19578 24177
rect 19522 24103 19578 24112
rect 19706 24168 19762 24177
rect 19706 24103 19762 24112
rect 19522 24032 19578 24041
rect 19522 23967 19578 23976
rect 19536 23866 19564 23967
rect 19524 23860 19576 23866
rect 19524 23802 19576 23808
rect 19720 23798 19748 24103
rect 20272 23905 20300 27520
rect 20824 24721 20852 27520
rect 20810 24712 20866 24721
rect 20810 24647 20866 24656
rect 20812 24268 20864 24274
rect 20812 24210 20864 24216
rect 20258 23896 20314 23905
rect 20258 23831 20314 23840
rect 19708 23792 19760 23798
rect 19708 23734 19760 23740
rect 19340 23656 19392 23662
rect 19340 23598 19392 23604
rect 17684 23520 17736 23526
rect 17406 23488 17462 23497
rect 17684 23462 17736 23468
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 19064 23520 19116 23526
rect 19064 23462 19116 23468
rect 17406 23423 17462 23432
rect 17224 23316 17276 23322
rect 17224 23258 17276 23264
rect 17040 23180 17092 23186
rect 17040 23122 17092 23128
rect 16764 22772 16816 22778
rect 16764 22714 16816 22720
rect 17052 22438 17080 23122
rect 17040 22432 17092 22438
rect 17500 22432 17552 22438
rect 17040 22374 17092 22380
rect 17498 22400 17500 22409
rect 17552 22400 17554 22409
rect 17052 22137 17080 22374
rect 17498 22335 17554 22344
rect 17038 22128 17094 22137
rect 17038 22063 17094 22072
rect 16670 21992 16726 22001
rect 16670 21927 16672 21936
rect 16724 21927 16726 21936
rect 16672 21898 16724 21904
rect 16578 21584 16634 21593
rect 16578 21519 16634 21528
rect 16026 21448 16082 21457
rect 16026 21383 16082 21392
rect 17696 19961 17724 23462
rect 18144 23180 18196 23186
rect 18144 23122 18196 23128
rect 18156 22438 18184 23122
rect 18144 22432 18196 22438
rect 18144 22374 18196 22380
rect 18602 22400 18658 22409
rect 17682 19952 17738 19961
rect 17682 19887 17738 19896
rect 16118 19408 16174 19417
rect 16118 19343 16174 19352
rect 15844 15428 15896 15434
rect 15844 15370 15896 15376
rect 15856 14822 15884 15370
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15856 14414 15884 14758
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15842 13424 15898 13433
rect 15842 13359 15844 13368
rect 15896 13359 15898 13368
rect 15844 13330 15896 13336
rect 15856 12986 15884 13330
rect 15936 13320 15988 13326
rect 16132 13308 16160 19343
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 16394 16552 16450 16561
rect 16394 16487 16450 16496
rect 16304 15632 16356 15638
rect 16304 15574 16356 15580
rect 16316 15162 16344 15574
rect 16408 15473 16436 16487
rect 16394 15464 16450 15473
rect 16394 15399 16450 15408
rect 16304 15156 16356 15162
rect 16304 15098 16356 15104
rect 16408 14906 16436 15399
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16500 15026 16528 15302
rect 16488 15020 16540 15026
rect 16488 14962 16540 14968
rect 16408 14878 16528 14906
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16224 14346 16252 14758
rect 16304 14612 16356 14618
rect 16304 14554 16356 14560
rect 16212 14340 16264 14346
rect 16212 14282 16264 14288
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16224 13462 16252 13670
rect 16316 13530 16344 14554
rect 16408 14414 16436 14758
rect 16396 14408 16448 14414
rect 16394 14376 16396 14385
rect 16448 14376 16450 14385
rect 16394 14311 16450 14320
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 16132 13280 16436 13308
rect 15936 13262 15988 13268
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15948 12170 15976 13262
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 15936 12164 15988 12170
rect 15936 12106 15988 12112
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15856 11354 15884 12038
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15672 9926 15700 11154
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15764 10470 15792 10950
rect 15856 10606 15884 11290
rect 15936 10736 15988 10742
rect 15936 10678 15988 10684
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15948 10418 15976 10678
rect 16040 10674 16068 13126
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16224 11830 16252 12242
rect 16212 11824 16264 11830
rect 16212 11766 16264 11772
rect 16212 11008 16264 11014
rect 16132 10956 16212 10962
rect 16132 10950 16264 10956
rect 16132 10934 16252 10950
rect 16132 10810 16160 10934
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16132 10674 16160 10746
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 15948 10390 16068 10418
rect 16040 10062 16068 10390
rect 16132 10198 16160 10610
rect 16120 10192 16172 10198
rect 16120 10134 16172 10140
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15672 8838 15700 9862
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15660 8832 15712 8838
rect 15660 8774 15712 8780
rect 15764 8634 15792 9454
rect 16040 9382 16068 9998
rect 16132 9586 16160 10134
rect 16302 9888 16358 9897
rect 16302 9823 16358 9832
rect 16316 9654 16344 9823
rect 16304 9648 16356 9654
rect 16304 9590 16356 9596
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 16132 9178 16160 9522
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 16224 8090 16252 8434
rect 16408 8129 16436 13280
rect 16500 12442 16528 14878
rect 17224 14476 17276 14482
rect 17224 14418 17276 14424
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16868 13870 16896 14350
rect 17236 13870 17264 14418
rect 16856 13864 16908 13870
rect 16854 13832 16856 13841
rect 17224 13864 17276 13870
rect 16908 13832 16910 13841
rect 17224 13806 17276 13812
rect 16854 13767 16910 13776
rect 16672 13320 16724 13326
rect 16670 13288 16672 13297
rect 16724 13288 16726 13297
rect 16670 13223 16726 13232
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16500 11898 16528 12378
rect 16868 12170 16896 12582
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16684 10713 16712 10746
rect 16670 10704 16726 10713
rect 16670 10639 16726 10648
rect 17236 10577 17264 13806
rect 17408 13252 17460 13258
rect 17408 13194 17460 13200
rect 17420 12986 17448 13194
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17420 10810 17448 12038
rect 17512 11558 17540 12242
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17512 11257 17540 11494
rect 17498 11248 17554 11257
rect 17498 11183 17554 11192
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17222 10568 17278 10577
rect 17222 10503 17278 10512
rect 17420 10266 17448 10610
rect 17408 10260 17460 10266
rect 17408 10202 17460 10208
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16684 9042 16712 9318
rect 17420 9110 17448 10202
rect 17408 9104 17460 9110
rect 17408 9046 17460 9052
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16500 8498 16528 8774
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16500 8242 16528 8434
rect 16684 8294 16712 8978
rect 17420 8634 17448 9046
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17500 8356 17552 8362
rect 17500 8298 17552 8304
rect 16672 8288 16724 8294
rect 16500 8214 16620 8242
rect 16672 8230 16724 8236
rect 16394 8120 16450 8129
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16316 8078 16394 8106
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15476 7336 15528 7342
rect 15474 7304 15476 7313
rect 15528 7304 15530 7313
rect 15474 7239 15530 7248
rect 15580 5778 15608 7754
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15672 7546 15700 7686
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15672 5914 15700 7482
rect 15764 7449 15792 7686
rect 15750 7440 15806 7449
rect 15750 7375 15752 7384
rect 15804 7375 15806 7384
rect 15752 7346 15804 7352
rect 15764 7315 15792 7346
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15936 5704 15988 5710
rect 15396 5630 15700 5658
rect 15936 5646 15988 5652
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 15290 5128 15346 5137
rect 15290 5063 15346 5072
rect 15474 5128 15530 5137
rect 15474 5063 15530 5072
rect 14832 4752 14884 4758
rect 14832 4694 14884 4700
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14844 4010 14872 4694
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15304 4162 15332 5063
rect 15488 4826 15516 5063
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15396 4282 15424 4626
rect 15384 4276 15436 4282
rect 15384 4218 15436 4224
rect 15304 4134 15516 4162
rect 15014 4040 15070 4049
rect 14832 4004 14884 4010
rect 15014 3975 15070 3984
rect 14832 3946 14884 3952
rect 14660 3896 14780 3924
rect 14648 3664 14700 3670
rect 14646 3632 14648 3641
rect 14700 3632 14702 3641
rect 14646 3567 14702 3576
rect 14752 3074 14780 3896
rect 15028 3738 15056 3975
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15198 3088 15254 3097
rect 14752 3046 14872 3074
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 14752 2650 14780 2790
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 14738 2544 14794 2553
rect 14738 2479 14740 2488
rect 14792 2479 14794 2488
rect 14740 2450 14792 2456
rect 14844 1442 14872 3046
rect 15198 3023 15254 3032
rect 15212 2854 15240 3023
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14844 1414 15148 1442
rect 15120 480 15148 1414
rect 15304 1329 15332 2246
rect 15488 1329 15516 4134
rect 15290 1320 15346 1329
rect 15290 1255 15346 1264
rect 15474 1320 15530 1329
rect 15474 1255 15530 1264
rect 15672 480 15700 5630
rect 15948 5370 15976 5646
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 15948 4826 15976 5306
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 15948 4214 15976 4762
rect 16316 4690 16344 8078
rect 16394 8055 16450 8064
rect 16488 7948 16540 7954
rect 16488 7890 16540 7896
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16408 7410 16436 7822
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16408 7206 16436 7346
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16408 6848 16436 7142
rect 16500 7002 16528 7890
rect 16592 7818 16620 8214
rect 16580 7812 16632 7818
rect 16580 7754 16632 7760
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16488 6860 16540 6866
rect 16408 6820 16488 6848
rect 16408 5574 16436 6820
rect 16488 6802 16540 6808
rect 16580 6656 16632 6662
rect 16684 6644 16712 8230
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16776 7546 16804 8026
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16632 6616 16712 6644
rect 16580 6598 16632 6604
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 16408 4554 16436 5510
rect 16500 5370 16528 6190
rect 16592 6118 16620 6598
rect 16762 6488 16818 6497
rect 16672 6452 16724 6458
rect 16762 6423 16818 6432
rect 16672 6394 16724 6400
rect 16684 6322 16712 6394
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16592 5778 16620 6054
rect 16684 5914 16712 6258
rect 16776 6254 16804 6423
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16670 5808 16726 5817
rect 16580 5772 16632 5778
rect 16670 5743 16726 5752
rect 16580 5714 16632 5720
rect 16580 5636 16632 5642
rect 16580 5578 16632 5584
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16592 5098 16620 5578
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16684 4758 16712 5743
rect 16868 5166 16896 7686
rect 17040 7268 17092 7274
rect 17040 7210 17092 7216
rect 17052 6186 17080 7210
rect 17040 6180 17092 6186
rect 17040 6122 17092 6128
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16960 5273 16988 6054
rect 17408 5772 17460 5778
rect 17408 5714 17460 5720
rect 16946 5264 17002 5273
rect 16946 5199 17002 5208
rect 17420 5166 17448 5714
rect 16856 5160 16908 5166
rect 17408 5160 17460 5166
rect 16856 5102 16908 5108
rect 17328 5120 17408 5148
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 16762 4584 16818 4593
rect 16396 4548 16448 4554
rect 16762 4519 16818 4528
rect 16396 4490 16448 4496
rect 15936 4208 15988 4214
rect 15936 4150 15988 4156
rect 16408 4146 16436 4490
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16028 4140 16080 4146
rect 16028 4082 16080 4088
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16040 3738 16068 4082
rect 16500 4078 16528 4422
rect 16488 4072 16540 4078
rect 16394 4040 16450 4049
rect 16488 4014 16540 4020
rect 16394 3975 16450 3984
rect 16408 3942 16436 3975
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 16224 480 16252 3402
rect 16316 2446 16344 3674
rect 16408 2650 16436 3878
rect 16500 3641 16528 4014
rect 16486 3632 16542 3641
rect 16486 3567 16542 3576
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16684 2650 16712 2994
rect 16396 2644 16448 2650
rect 16396 2586 16448 2592
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16776 480 16804 4519
rect 16868 4282 16896 5102
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16960 4214 16988 4558
rect 16948 4208 17000 4214
rect 16948 4150 17000 4156
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16960 3058 16988 3538
rect 17052 3398 17080 4626
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 17130 2544 17186 2553
rect 17130 2479 17132 2488
rect 17184 2479 17186 2488
rect 17132 2450 17184 2456
rect 17236 2378 17264 4762
rect 17328 3670 17356 5120
rect 17408 5102 17460 5108
rect 17512 5098 17540 8298
rect 17500 5092 17552 5098
rect 17500 5034 17552 5040
rect 17604 4434 17632 18566
rect 17866 16144 17922 16153
rect 17866 16079 17922 16088
rect 17880 15178 17908 16079
rect 17880 15150 18000 15178
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 17880 14414 17908 14962
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17880 13734 17908 14350
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 17774 12336 17830 12345
rect 17774 12271 17830 12280
rect 17788 12170 17816 12271
rect 17880 12220 17908 13670
rect 17972 12850 18000 15150
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 17960 12232 18012 12238
rect 17880 12192 17960 12220
rect 17960 12174 18012 12180
rect 17776 12164 17828 12170
rect 17776 12106 17828 12112
rect 17788 11898 17816 12106
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17972 11694 18000 12174
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 18052 11552 18104 11558
rect 18050 11520 18052 11529
rect 18104 11520 18106 11529
rect 18050 11455 18106 11464
rect 18050 11384 18106 11393
rect 18050 11319 18052 11328
rect 18104 11319 18106 11328
rect 18052 11290 18104 11296
rect 17776 11280 17828 11286
rect 17776 11222 17828 11228
rect 17788 10470 17816 11222
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 18156 10305 18184 22374
rect 18602 22335 18658 22344
rect 18234 13968 18290 13977
rect 18234 13903 18290 13912
rect 18248 13462 18276 13903
rect 18326 13560 18382 13569
rect 18326 13495 18382 13504
rect 18236 13456 18288 13462
rect 18236 13398 18288 13404
rect 18248 12986 18276 13398
rect 18236 12980 18288 12986
rect 18236 12922 18288 12928
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18142 10296 18198 10305
rect 18142 10231 18198 10240
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17696 8090 17724 9318
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17972 8401 18000 8774
rect 17958 8392 18014 8401
rect 17958 8327 18014 8336
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17682 7984 17738 7993
rect 17682 7919 17738 7928
rect 18052 7948 18104 7954
rect 17696 6458 17724 7919
rect 18052 7890 18104 7896
rect 18064 7342 18092 7890
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18156 7478 18184 7822
rect 18144 7472 18196 7478
rect 18144 7414 18196 7420
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18050 6760 18106 6769
rect 18050 6695 18106 6704
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17696 6254 17724 6394
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 17788 5846 17816 6598
rect 18064 6458 18092 6695
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 17776 5840 17828 5846
rect 17776 5782 17828 5788
rect 17958 5672 18014 5681
rect 17958 5607 18014 5616
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 17880 4826 17908 5170
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17972 4554 18000 5607
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18156 5166 18184 5510
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18052 4752 18104 4758
rect 18248 4729 18276 12786
rect 18340 11218 18368 13495
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18524 12986 18552 13330
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18524 12753 18552 12922
rect 18510 12744 18566 12753
rect 18510 12679 18566 12688
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18432 11937 18460 12038
rect 18418 11928 18474 11937
rect 18418 11863 18474 11872
rect 18432 11694 18460 11863
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18512 11280 18564 11286
rect 18512 11222 18564 11228
rect 18328 11212 18380 11218
rect 18328 11154 18380 11160
rect 18340 9994 18368 11154
rect 18328 9988 18380 9994
rect 18328 9930 18380 9936
rect 18418 8120 18474 8129
rect 18418 8055 18474 8064
rect 18432 7342 18460 8055
rect 18420 7336 18472 7342
rect 18326 7304 18382 7313
rect 18420 7278 18472 7284
rect 18326 7239 18382 7248
rect 18340 7206 18368 7239
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 18432 7002 18460 7278
rect 18524 7002 18552 11222
rect 18616 10810 18644 22335
rect 18708 16561 18736 23462
rect 19076 23322 19104 23462
rect 19064 23316 19116 23322
rect 19064 23258 19116 23264
rect 19352 17241 19380 23598
rect 20824 23526 20852 24210
rect 21376 24041 21404 27520
rect 21362 24032 21418 24041
rect 21362 23967 21418 23976
rect 21270 23896 21326 23905
rect 21270 23831 21272 23840
rect 21324 23831 21326 23840
rect 21272 23802 21324 23808
rect 21088 23656 21140 23662
rect 21088 23598 21140 23604
rect 20812 23520 20864 23526
rect 20812 23462 20864 23468
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 20824 17785 20852 23462
rect 21100 23322 21128 23598
rect 21088 23316 21140 23322
rect 21088 23258 21140 23264
rect 20902 23216 20958 23225
rect 20902 23151 20904 23160
rect 20956 23151 20958 23160
rect 20904 23122 20956 23128
rect 20916 22778 20944 23122
rect 21928 22953 21956 27520
rect 22480 24410 22508 27520
rect 22468 24404 22520 24410
rect 22468 24346 22520 24352
rect 23124 23905 23152 27520
rect 23110 23896 23166 23905
rect 23110 23831 23166 23840
rect 23480 23656 23532 23662
rect 23676 23633 23704 27520
rect 24228 24857 24256 27520
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24214 24848 24270 24857
rect 24214 24783 24270 24792
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 23480 23598 23532 23604
rect 23662 23624 23718 23633
rect 23492 23322 23520 23598
rect 23662 23559 23718 23568
rect 23570 23352 23626 23361
rect 23480 23316 23532 23322
rect 23570 23287 23626 23296
rect 23480 23258 23532 23264
rect 22376 23180 22428 23186
rect 22376 23122 22428 23128
rect 21914 22944 21970 22953
rect 21914 22879 21970 22888
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 22388 22438 22416 23122
rect 22376 22432 22428 22438
rect 22376 22374 22428 22380
rect 20810 17776 20866 17785
rect 20810 17711 20866 17720
rect 19338 17232 19394 17241
rect 19338 17167 19394 17176
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 18694 16552 18750 16561
rect 18694 16487 18750 16496
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19154 13288 19210 13297
rect 19154 13223 19210 13232
rect 19168 11898 19196 13223
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19352 12889 19380 13126
rect 19338 12880 19394 12889
rect 19338 12815 19394 12824
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 20166 12336 20222 12345
rect 20166 12271 20222 12280
rect 19156 11892 19208 11898
rect 19156 11834 19208 11840
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 18708 11150 18736 11562
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18604 10804 18656 10810
rect 18604 10746 18656 10752
rect 18708 10266 18736 11086
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18602 10160 18658 10169
rect 18602 10095 18658 10104
rect 18616 7342 18644 10095
rect 18800 9926 18828 10406
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 18788 9920 18840 9926
rect 18786 9888 18788 9897
rect 18840 9888 18842 9897
rect 18786 9823 18842 9832
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 18604 7336 18656 7342
rect 18604 7278 18656 7284
rect 18420 6996 18472 7002
rect 18420 6938 18472 6944
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18708 6662 18736 7346
rect 19156 7336 19208 7342
rect 19156 7278 19208 7284
rect 18786 7168 18842 7177
rect 18786 7103 18842 7112
rect 18800 6866 18828 7103
rect 19064 6996 19116 7002
rect 19064 6938 19116 6944
rect 18788 6860 18840 6866
rect 18788 6802 18840 6808
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18420 5092 18472 5098
rect 18420 5034 18472 5040
rect 18052 4694 18104 4700
rect 18234 4720 18290 4729
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 17604 4406 17724 4434
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17316 3664 17368 3670
rect 17316 3606 17368 3612
rect 17328 3194 17356 3606
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 17420 2961 17448 3878
rect 17696 3754 17724 4406
rect 18064 4282 18092 4694
rect 18234 4655 18290 4664
rect 18144 4616 18196 4622
rect 18144 4558 18196 4564
rect 18052 4276 18104 4282
rect 18052 4218 18104 4224
rect 17958 4176 18014 4185
rect 17958 4111 18014 4120
rect 18052 4140 18104 4146
rect 17776 3936 17828 3942
rect 17774 3904 17776 3913
rect 17828 3904 17830 3913
rect 17774 3839 17830 3848
rect 17696 3726 17816 3754
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 17696 2961 17724 3334
rect 17788 3194 17816 3726
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17788 2990 17816 3130
rect 17776 2984 17828 2990
rect 17406 2952 17462 2961
rect 17406 2887 17462 2896
rect 17682 2952 17738 2961
rect 17776 2926 17828 2932
rect 17682 2887 17738 2896
rect 17406 2816 17462 2825
rect 17406 2751 17462 2760
rect 17224 2372 17276 2378
rect 17224 2314 17276 2320
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 16854 2136 16910 2145
rect 16854 2071 16910 2080
rect 16868 1873 16896 2071
rect 16960 2009 16988 2246
rect 16946 2000 17002 2009
rect 16946 1935 17002 1944
rect 16854 1864 16910 1873
rect 16854 1799 16910 1808
rect 17130 1864 17186 1873
rect 17130 1799 17186 1808
rect 17144 1465 17172 1799
rect 17328 1465 17356 2246
rect 17130 1456 17186 1465
rect 17130 1391 17186 1400
rect 17314 1456 17370 1465
rect 17314 1391 17370 1400
rect 17420 480 17448 2751
rect 17972 480 18000 4111
rect 18052 4082 18104 4088
rect 18064 3369 18092 4082
rect 18156 3738 18184 4558
rect 18144 3732 18196 3738
rect 18144 3674 18196 3680
rect 18050 3360 18106 3369
rect 18050 3295 18106 3304
rect 18064 3194 18092 3295
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 18248 2922 18276 4655
rect 18432 4593 18460 5034
rect 18418 4584 18474 4593
rect 18418 4519 18474 4528
rect 18524 4146 18552 6258
rect 18708 6225 18736 6598
rect 18694 6216 18750 6225
rect 18694 6151 18750 6160
rect 18800 5574 18828 6802
rect 19076 6458 19104 6938
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 18788 5568 18840 5574
rect 18788 5510 18840 5516
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18524 3738 18552 4082
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 18510 3224 18566 3233
rect 18510 3159 18566 3168
rect 18236 2916 18288 2922
rect 18156 2876 18236 2904
rect 18156 2650 18184 2876
rect 18236 2858 18288 2864
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18524 480 18552 3159
rect 18694 2680 18750 2689
rect 18694 2615 18696 2624
rect 18748 2615 18750 2624
rect 18696 2586 18748 2592
rect 18800 1057 18828 5510
rect 19168 4808 19196 7278
rect 19260 6322 19288 9930
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 20076 7812 20128 7818
rect 20076 7754 20128 7760
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 19352 7041 19380 7346
rect 19996 7274 20024 7686
rect 19984 7268 20036 7274
rect 19984 7210 20036 7216
rect 20088 7206 20116 7754
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 19338 7032 19394 7041
rect 19338 6967 19394 6976
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 19444 6390 19472 6734
rect 19432 6384 19484 6390
rect 19432 6326 19484 6332
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 19338 6216 19394 6225
rect 19444 6202 19472 6326
rect 19536 6225 19564 7142
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19982 6896 20038 6905
rect 19982 6831 20038 6840
rect 19996 6254 20024 6831
rect 19984 6248 20036 6254
rect 19394 6174 19472 6202
rect 19338 6151 19394 6160
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19352 5302 19380 5714
rect 19444 5370 19472 6174
rect 19522 6216 19578 6225
rect 19984 6190 20036 6196
rect 19522 6151 19578 6160
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19996 5914 20024 6190
rect 19984 5908 20036 5914
rect 19984 5850 20036 5856
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19432 5024 19484 5030
rect 19430 4992 19432 5001
rect 19484 4992 19486 5001
rect 19430 4927 19486 4936
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19430 4856 19486 4865
rect 19340 4820 19392 4826
rect 19168 4780 19340 4808
rect 19168 4146 19196 4780
rect 19622 4848 19918 4868
rect 19430 4791 19486 4800
rect 19340 4762 19392 4768
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 19352 4010 19380 4626
rect 19444 4622 19472 4791
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19800 4480 19852 4486
rect 19800 4422 19852 4428
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 19432 4072 19484 4078
rect 19812 4049 19840 4422
rect 20088 4214 20116 4422
rect 20076 4208 20128 4214
rect 20076 4150 20128 4156
rect 19432 4014 19484 4020
rect 19798 4040 19854 4049
rect 19340 4004 19392 4010
rect 19340 3946 19392 3952
rect 19444 3942 19472 4014
rect 20180 4010 20208 12271
rect 22388 8945 22416 22374
rect 23584 22001 23612 23287
rect 24780 23089 24808 27520
rect 25332 23866 25360 27520
rect 25976 24177 26004 27520
rect 26528 24313 26556 27520
rect 26514 24304 26570 24313
rect 26514 24239 26570 24248
rect 25962 24168 26018 24177
rect 25962 24103 26018 24112
rect 25320 23860 25372 23866
rect 25320 23802 25372 23808
rect 27080 23769 27108 27520
rect 27066 23760 27122 23769
rect 27066 23695 27122 23704
rect 24766 23080 24822 23089
rect 24766 23015 24822 23024
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 23570 21992 23626 22001
rect 23570 21927 23626 21936
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 27632 21418 27660 27520
rect 26240 21412 26292 21418
rect 26240 21354 26292 21360
rect 27620 21412 27672 21418
rect 27620 21354 27672 21360
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 26252 13297 26280 21354
rect 26238 13288 26294 13297
rect 26238 13223 26294 13232
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 22374 8936 22430 8945
rect 22374 8871 22430 8880
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 20350 8528 20406 8537
rect 20350 8463 20406 8472
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20272 6497 20300 6598
rect 20258 6488 20314 6497
rect 20258 6423 20314 6432
rect 20260 4548 20312 4554
rect 20260 4490 20312 4496
rect 19798 3975 19854 3984
rect 20168 4004 20220 4010
rect 20168 3946 20220 3952
rect 19432 3936 19484 3942
rect 19246 3904 19302 3913
rect 19432 3878 19484 3884
rect 19246 3839 19302 3848
rect 18970 3768 19026 3777
rect 18970 3703 18972 3712
rect 19024 3703 19026 3712
rect 18972 3674 19024 3680
rect 19062 3496 19118 3505
rect 19062 3431 19118 3440
rect 19260 3482 19288 3839
rect 19260 3466 19380 3482
rect 19260 3460 19392 3466
rect 19260 3454 19340 3460
rect 19076 3194 19104 3431
rect 19156 3392 19208 3398
rect 19156 3334 19208 3340
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 19168 2417 19196 3334
rect 19260 2650 19288 3454
rect 19340 3402 19392 3408
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 19352 2582 19380 3130
rect 19444 3097 19472 3878
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 20180 3777 20208 3946
rect 20166 3768 20222 3777
rect 20166 3703 20168 3712
rect 20220 3703 20222 3712
rect 20168 3674 20220 3680
rect 20180 3643 20208 3674
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 19536 3126 19564 3538
rect 19800 3528 19852 3534
rect 19800 3470 19852 3476
rect 19812 3194 19840 3470
rect 19800 3188 19852 3194
rect 19800 3130 19852 3136
rect 19524 3120 19576 3126
rect 19430 3088 19486 3097
rect 19524 3062 19576 3068
rect 19430 3023 19486 3032
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19340 2576 19392 2582
rect 19340 2518 19392 2524
rect 19444 2514 19472 2926
rect 19524 2916 19576 2922
rect 19524 2858 19576 2864
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 19154 2408 19210 2417
rect 19154 2343 19210 2352
rect 19536 2310 19564 2858
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19524 2304 19576 2310
rect 19524 2246 19576 2252
rect 20076 2304 20128 2310
rect 20076 2246 20128 2252
rect 19536 2145 19564 2246
rect 19522 2136 19578 2145
rect 19522 2071 19578 2080
rect 18878 2000 18934 2009
rect 18878 1935 18934 1944
rect 18892 1601 18920 1935
rect 18878 1592 18934 1601
rect 18878 1527 18934 1536
rect 19062 1592 19118 1601
rect 19062 1527 19118 1536
rect 18786 1048 18842 1057
rect 18786 983 18842 992
rect 19076 480 19104 1527
rect 20088 1465 20116 2246
rect 19614 1456 19670 1465
rect 19614 1391 19670 1400
rect 20074 1456 20130 1465
rect 20074 1391 20130 1400
rect 19628 480 19656 1391
rect 20272 480 20300 4490
rect 20364 2990 20392 8463
rect 22742 7848 22798 7857
rect 22742 7783 22798 7792
rect 21362 7304 21418 7313
rect 20628 7268 20680 7274
rect 20680 7228 20760 7256
rect 21362 7239 21418 7248
rect 20628 7210 20680 7216
rect 20732 6458 20760 7228
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20548 5914 20576 6258
rect 20824 5914 20852 7142
rect 20996 6112 21048 6118
rect 20996 6054 21048 6060
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20548 5234 20576 5850
rect 21008 5710 21036 6054
rect 21376 5914 21404 7239
rect 22284 6860 22336 6866
rect 22284 6802 22336 6808
rect 21640 6724 21692 6730
rect 21640 6666 21692 6672
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21560 6186 21588 6598
rect 21652 6322 21680 6666
rect 22296 6497 22324 6802
rect 22468 6656 22520 6662
rect 22468 6598 22520 6604
rect 22282 6488 22338 6497
rect 22282 6423 22284 6432
rect 22336 6423 22338 6432
rect 22284 6394 22336 6400
rect 21640 6316 21692 6322
rect 21640 6258 21692 6264
rect 22190 6216 22246 6225
rect 21548 6180 21600 6186
rect 22190 6151 22246 6160
rect 21548 6122 21600 6128
rect 21364 5908 21416 5914
rect 21364 5850 21416 5856
rect 21272 5772 21324 5778
rect 21272 5714 21324 5720
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 20812 5636 20864 5642
rect 20812 5578 20864 5584
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20548 4826 20576 4966
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 20732 4622 20760 4966
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20720 4480 20772 4486
rect 20720 4422 20772 4428
rect 20732 4185 20760 4422
rect 20718 4176 20774 4185
rect 20718 4111 20774 4120
rect 20352 2984 20404 2990
rect 20352 2926 20404 2932
rect 20824 480 20852 5578
rect 21008 5409 21036 5646
rect 20994 5400 21050 5409
rect 20994 5335 21050 5344
rect 21008 5166 21036 5335
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 21284 4826 21312 5714
rect 21376 5370 21404 5850
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 22204 5166 22232 6151
rect 22282 5808 22338 5817
rect 22480 5778 22508 6598
rect 22282 5743 22338 5752
rect 22468 5772 22520 5778
rect 22192 5160 22244 5166
rect 22192 5102 22244 5108
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 20902 4720 20958 4729
rect 20902 4655 20904 4664
rect 20956 4655 20958 4664
rect 20904 4626 20956 4632
rect 20916 4282 20944 4626
rect 20904 4276 20956 4282
rect 20904 4218 20956 4224
rect 22296 4078 22324 5743
rect 22468 5714 22520 5720
rect 21088 4072 21140 4078
rect 22284 4072 22336 4078
rect 21088 4014 21140 4020
rect 21362 4040 21418 4049
rect 20904 2304 20956 2310
rect 20904 2246 20956 2252
rect 20916 1873 20944 2246
rect 20902 1864 20958 1873
rect 20902 1799 20958 1808
rect 21100 1329 21128 4014
rect 22284 4014 22336 4020
rect 21362 3975 21418 3984
rect 22376 4004 22428 4010
rect 21272 3392 21324 3398
rect 21272 3334 21324 3340
rect 21284 2825 21312 3334
rect 21270 2816 21326 2825
rect 21270 2751 21326 2760
rect 21180 2304 21232 2310
rect 21180 2246 21232 2252
rect 21192 1737 21220 2246
rect 21178 1728 21234 1737
rect 21178 1663 21234 1672
rect 21086 1320 21142 1329
rect 21086 1255 21142 1264
rect 21376 480 21404 3975
rect 22376 3946 22428 3952
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 21456 3664 21508 3670
rect 21456 3606 21508 3612
rect 21638 3632 21694 3641
rect 21468 3194 21496 3606
rect 21638 3567 21640 3576
rect 21692 3567 21694 3576
rect 21640 3538 21692 3544
rect 21916 3392 21968 3398
rect 22204 3369 22232 3878
rect 22282 3768 22338 3777
rect 22282 3703 22338 3712
rect 22296 3602 22324 3703
rect 22284 3596 22336 3602
rect 22284 3538 22336 3544
rect 21916 3334 21968 3340
rect 22190 3360 22246 3369
rect 21456 3188 21508 3194
rect 21456 3130 21508 3136
rect 21456 2984 21508 2990
rect 21456 2926 21508 2932
rect 21822 2952 21878 2961
rect 21468 1193 21496 2926
rect 21822 2887 21878 2896
rect 21836 2854 21864 2887
rect 21824 2848 21876 2854
rect 21824 2790 21876 2796
rect 21548 2508 21600 2514
rect 21548 2450 21600 2456
rect 21560 2417 21588 2450
rect 21640 2440 21692 2446
rect 21546 2408 21602 2417
rect 21640 2382 21692 2388
rect 21546 2343 21602 2352
rect 21560 2310 21588 2343
rect 21548 2304 21600 2310
rect 21548 2246 21600 2252
rect 21652 2009 21680 2382
rect 21638 2000 21694 2009
rect 21638 1935 21694 1944
rect 21454 1184 21510 1193
rect 21454 1119 21510 1128
rect 21928 480 21956 3334
rect 22190 3295 22246 3304
rect 22296 3194 22324 3538
rect 22284 3188 22336 3194
rect 22284 3130 22336 3136
rect 22388 1986 22416 3946
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 22480 3670 22508 3878
rect 22468 3664 22520 3670
rect 22468 3606 22520 3612
rect 22756 2514 22784 7783
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 23296 5772 23348 5778
rect 23296 5714 23348 5720
rect 23308 5370 23336 5714
rect 23480 5568 23532 5574
rect 23480 5510 23532 5516
rect 23296 5364 23348 5370
rect 23296 5306 23348 5312
rect 23492 2825 23520 5510
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 23570 5264 23626 5273
rect 23570 5199 23626 5208
rect 23584 2990 23612 5199
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 26514 4040 26570 4049
rect 26514 3975 26570 3984
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 23846 3224 23902 3233
rect 24289 3216 24585 3236
rect 23846 3159 23848 3168
rect 23900 3159 23902 3168
rect 23848 3130 23900 3136
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 23662 2952 23718 2961
rect 23662 2887 23718 2896
rect 23110 2816 23166 2825
rect 23110 2751 23166 2760
rect 23478 2816 23534 2825
rect 23478 2751 23534 2760
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 22388 1958 22508 1986
rect 22480 480 22508 1958
rect 23124 480 23152 2751
rect 23478 2544 23534 2553
rect 23478 2479 23480 2488
rect 23532 2479 23534 2488
rect 23480 2450 23532 2456
rect 23676 480 23704 2887
rect 25318 2816 25374 2825
rect 25318 2751 25374 2760
rect 24032 2508 24084 2514
rect 24032 2450 24084 2456
rect 24044 2417 24072 2450
rect 24030 2408 24086 2417
rect 24030 2343 24086 2352
rect 24124 2372 24176 2378
rect 24124 2314 24176 2320
rect 24136 1170 24164 2314
rect 24216 2304 24268 2310
rect 24216 2246 24268 2252
rect 24228 1601 24256 2246
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24214 1592 24270 1601
rect 24214 1527 24270 1536
rect 24136 1142 24256 1170
rect 24228 480 24256 1142
rect 24688 598 24808 626
rect 11610 96 11666 105
rect 11610 31 11666 40
rect 11702 0 11758 480
rect 12254 0 12310 480
rect 12806 0 12862 480
rect 13358 0 13414 480
rect 13910 0 13966 480
rect 14554 0 14610 480
rect 15106 0 15162 480
rect 15658 0 15714 480
rect 16210 0 16266 480
rect 16762 0 16818 480
rect 17406 0 17462 480
rect 17958 0 18014 480
rect 18510 0 18566 480
rect 19062 0 19118 480
rect 19614 0 19670 480
rect 20258 0 20314 480
rect 20810 0 20866 480
rect 21362 0 21418 480
rect 21914 0 21970 480
rect 22466 0 22522 480
rect 23110 0 23166 480
rect 23662 0 23718 480
rect 24214 0 24270 480
rect 24688 105 24716 598
rect 24780 480 24808 598
rect 25332 480 25360 2751
rect 25962 1456 26018 1465
rect 25962 1391 26018 1400
rect 25976 480 26004 1391
rect 26528 480 26556 3975
rect 27618 3496 27674 3505
rect 27618 3431 27674 3440
rect 27066 912 27122 921
rect 27066 847 27122 856
rect 27080 480 27108 847
rect 27632 480 27660 3431
rect 24674 96 24730 105
rect 24674 31 24730 40
rect 24766 0 24822 480
rect 25318 0 25374 480
rect 25962 0 26018 480
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 3054 27648 3110 27704
rect 18 12824 74 12880
rect 1398 21256 1454 21312
rect 1858 24656 1914 24712
rect 1858 23568 1914 23624
rect 1582 21800 1638 21856
rect 1398 18944 1454 19000
rect 1582 18400 1638 18456
rect 1398 17720 1454 17776
rect 1490 16768 1546 16824
rect 1582 15952 1638 16008
rect 1398 15408 1454 15464
rect 1582 14864 1638 14920
rect 1398 13640 1454 13696
rect 1398 13388 1454 13424
rect 1398 13368 1400 13388
rect 1400 13368 1452 13388
rect 1452 13368 1454 13388
rect 1674 13232 1730 13288
rect 1582 13096 1638 13152
rect 1582 12552 1638 12608
rect 2042 24812 2098 24848
rect 2042 24792 2044 24812
rect 2044 24792 2096 24812
rect 2096 24792 2098 24812
rect 2778 26560 2834 26616
rect 2042 23568 2098 23624
rect 2870 23024 2926 23080
rect 3054 23160 3110 23216
rect 2962 22480 3018 22536
rect 2962 20848 3018 20904
rect 2042 19896 2098 19952
rect 2042 19780 2098 19816
rect 2042 19760 2044 19780
rect 2044 19760 2096 19780
rect 2096 19760 2098 19780
rect 2042 16496 2098 16552
rect 1950 15680 2006 15736
rect 2042 15564 2098 15600
rect 2042 15544 2044 15564
rect 2044 15544 2096 15564
rect 2096 15544 2098 15564
rect 2226 17584 2282 17640
rect 2870 20304 2926 20360
rect 2686 20032 2742 20088
rect 2686 19488 2742 19544
rect 2502 19252 2504 19272
rect 2504 19252 2556 19272
rect 2556 19252 2558 19272
rect 2502 19216 2558 19252
rect 2502 18828 2558 18864
rect 2502 18808 2504 18828
rect 2504 18808 2556 18828
rect 2556 18808 2558 18828
rect 2226 15272 2282 15328
rect 2686 17176 2742 17232
rect 3606 27104 3662 27160
rect 3238 25336 3294 25392
rect 4066 25880 4122 25936
rect 3698 24112 3754 24168
rect 3514 21392 3570 21448
rect 3238 18944 3294 19000
rect 3606 18808 3662 18864
rect 3146 16788 3202 16824
rect 3146 16768 3148 16788
rect 3148 16768 3200 16788
rect 3200 16768 3202 16788
rect 3330 17176 3386 17232
rect 3238 15952 3294 16008
rect 1858 14456 1914 14512
rect 2042 13776 2098 13832
rect 1766 11464 1822 11520
rect 1858 10920 1914 10976
rect 1398 9988 1454 10024
rect 1398 9968 1400 9988
rect 1400 9968 1452 9988
rect 1452 9968 1454 9988
rect 1858 9596 1860 9616
rect 1860 9596 1912 9616
rect 1912 9596 1914 9616
rect 1858 9560 1914 9596
rect 1398 8336 1454 8392
rect 294 4120 350 4176
rect 846 3304 902 3360
rect 1398 1808 1454 1864
rect 2318 12552 2374 12608
rect 2686 14320 2742 14376
rect 3238 14320 3294 14376
rect 2870 13640 2926 13696
rect 2778 13524 2834 13560
rect 2778 13504 2780 13524
rect 2780 13504 2832 13524
rect 2832 13504 2834 13524
rect 3146 13232 3202 13288
rect 3238 12552 3294 12608
rect 3790 18128 3846 18184
rect 4066 24520 4122 24576
rect 4066 23024 4122 23080
rect 4250 23740 4252 23760
rect 4252 23740 4304 23760
rect 4304 23740 4306 23760
rect 4250 23704 4306 23740
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 4250 15700 4306 15736
rect 4250 15680 4252 15700
rect 4252 15680 4304 15700
rect 4304 15680 4306 15700
rect 3698 13368 3754 13424
rect 3606 12824 3662 12880
rect 3606 11328 3662 11384
rect 3422 10376 3478 10432
rect 2870 10104 2926 10160
rect 2502 9152 2558 9208
rect 3146 8236 3148 8256
rect 3148 8236 3200 8256
rect 3200 8236 3202 8256
rect 1858 5228 1914 5264
rect 1858 5208 1860 5228
rect 1860 5208 1912 5228
rect 1912 5208 1914 5228
rect 1766 4936 1822 4992
rect 2226 5480 2282 5536
rect 1674 3732 1730 3768
rect 1674 3712 1676 3732
rect 1676 3712 1728 3732
rect 1728 3712 1730 3732
rect 1582 1400 1638 1456
rect 1674 856 1730 912
rect 2502 3576 2558 3632
rect 3146 8200 3202 8236
rect 3882 13776 3938 13832
rect 3882 12552 3938 12608
rect 4342 13504 4398 13560
rect 4250 11872 4306 11928
rect 4526 18128 4582 18184
rect 4066 11464 4122 11520
rect 3882 11212 3938 11248
rect 3882 11192 3884 11212
rect 3884 11192 3936 11212
rect 3936 11192 3938 11212
rect 4342 11600 4398 11656
rect 3790 9424 3846 9480
rect 3974 9832 4030 9888
rect 3974 9560 4030 9616
rect 4802 15272 4858 15328
rect 4894 13504 4950 13560
rect 4434 9052 4436 9072
rect 4436 9052 4488 9072
rect 4488 9052 4490 9072
rect 4434 9016 4490 9052
rect 4066 8900 4122 8936
rect 4066 8880 4068 8900
rect 4068 8880 4120 8900
rect 4120 8880 4122 8900
rect 3790 8472 3846 8528
rect 4710 9424 4766 9480
rect 3422 7248 3478 7304
rect 3330 5888 3386 5944
rect 3054 5108 3056 5128
rect 3056 5108 3108 5128
rect 3108 5108 3110 5128
rect 3054 5072 3110 5108
rect 2870 4684 2926 4720
rect 2870 4664 2872 4684
rect 2872 4664 2924 4684
rect 2924 4664 2926 4684
rect 2686 4528 2742 4584
rect 2318 1536 2374 1592
rect 2870 3440 2926 3496
rect 2686 3168 2742 3224
rect 4434 6996 4490 7032
rect 4434 6976 4436 6996
rect 4436 6976 4488 6996
rect 4488 6976 4490 6996
rect 3422 4120 3478 4176
rect 3330 3848 3386 3904
rect 3422 3032 3478 3088
rect 2870 2896 2926 2952
rect 2962 2488 3018 2544
rect 4526 6740 4528 6760
rect 4528 6740 4580 6760
rect 4580 6740 4582 6760
rect 3698 4800 3754 4856
rect 4526 6704 4582 6740
rect 3974 6296 4030 6352
rect 3790 4392 3846 4448
rect 3698 3848 3754 3904
rect 3422 992 3478 1048
rect 4066 6160 4122 6216
rect 4066 5616 4122 5672
rect 3974 4936 4030 4992
rect 4802 6840 4858 6896
rect 4894 6024 4950 6080
rect 4526 3576 4582 3632
rect 4434 3340 4436 3360
rect 4436 3340 4488 3360
rect 4488 3340 4490 3360
rect 4434 3304 4490 3340
rect 4986 2352 5042 2408
rect 5262 23432 5318 23488
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 6550 24656 6606 24712
rect 5538 22616 5594 22672
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 6366 23024 6422 23080
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 6642 22480 6698 22536
rect 6550 21292 6552 21312
rect 6552 21292 6604 21312
rect 6604 21292 6606 21312
rect 6550 21256 6606 21292
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5998 18808 6054 18864
rect 5998 18672 6054 18728
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5538 17176 5594 17232
rect 5722 16652 5778 16688
rect 5722 16632 5724 16652
rect 5724 16632 5776 16652
rect 5776 16632 5778 16652
rect 5630 16496 5686 16552
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5170 15408 5226 15464
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 6274 15272 6330 15328
rect 6090 14048 6146 14104
rect 5446 13504 5502 13560
rect 5170 13368 5226 13424
rect 5630 13252 5686 13288
rect 5630 13232 5632 13252
rect 5632 13232 5684 13252
rect 5684 13232 5686 13252
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5630 12588 5632 12608
rect 5632 12588 5684 12608
rect 5684 12588 5686 12608
rect 5630 12552 5686 12588
rect 5998 12044 6000 12064
rect 6000 12044 6052 12064
rect 6052 12044 6054 12064
rect 5998 12008 6054 12044
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 6274 13640 6330 13696
rect 6182 13096 6238 13152
rect 6090 10512 6146 10568
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 6090 9832 6146 9888
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5538 8336 5594 8392
rect 5170 4972 5172 4992
rect 5172 4972 5224 4992
rect 5224 4972 5226 4992
rect 5170 4936 5226 4972
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5262 4528 5318 4584
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5538 4120 5594 4176
rect 5170 3576 5226 3632
rect 5170 3188 5226 3224
rect 5170 3168 5172 3188
rect 5172 3168 5224 3188
rect 5224 3168 5226 3188
rect 5262 2624 5318 2680
rect 6366 12960 6422 13016
rect 6366 10784 6422 10840
rect 7470 23432 7526 23488
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 9954 24792 10010 24848
rect 8758 23568 8814 23624
rect 7286 20868 7342 20904
rect 7286 20848 7288 20868
rect 7288 20848 7340 20868
rect 7340 20848 7342 20868
rect 7010 19896 7066 19952
rect 7286 19916 7342 19952
rect 7286 19896 7288 19916
rect 7288 19896 7340 19916
rect 7340 19896 7342 19916
rect 6826 18028 6828 18048
rect 6828 18028 6880 18048
rect 6880 18028 6882 18048
rect 6826 17992 6882 18028
rect 6826 13776 6882 13832
rect 7470 18964 7526 19000
rect 7470 18944 7472 18964
rect 7472 18944 7524 18964
rect 7524 18944 7526 18964
rect 7562 17992 7618 18048
rect 7654 15272 7710 15328
rect 7194 12724 7196 12744
rect 7196 12724 7248 12744
rect 7248 12724 7250 12744
rect 7194 12688 7250 12724
rect 7102 11872 7158 11928
rect 7010 11328 7066 11384
rect 6274 6840 6330 6896
rect 6274 5092 6330 5128
rect 6274 5072 6276 5092
rect 6276 5072 6328 5092
rect 6328 5072 6330 5092
rect 6182 4120 6238 4176
rect 5998 3848 6054 3904
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 5446 1400 5502 1456
rect 6274 2352 6330 2408
rect 7010 9288 7066 9344
rect 6826 6452 6882 6488
rect 6826 6432 6828 6452
rect 6828 6432 6880 6452
rect 6880 6432 6882 6452
rect 6918 6296 6974 6352
rect 7838 20440 7894 20496
rect 7930 18672 7986 18728
rect 7838 16088 7894 16144
rect 8390 22652 8392 22672
rect 8392 22652 8444 22672
rect 8444 22652 8446 22672
rect 8390 22616 8446 22652
rect 8206 21936 8262 21992
rect 8482 21412 8538 21448
rect 8482 21392 8484 21412
rect 8484 21392 8536 21412
rect 8536 21392 8538 21412
rect 8574 16768 8630 16824
rect 8114 15952 8170 16008
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 9494 23704 9550 23760
rect 9126 21256 9182 21312
rect 7838 11328 7894 11384
rect 7930 11056 7986 11112
rect 7194 8472 7250 8528
rect 7286 6316 7342 6352
rect 7286 6296 7288 6316
rect 7288 6296 7340 6316
rect 7340 6296 7342 6316
rect 7102 3984 7158 4040
rect 6458 2080 6514 2136
rect 6918 2624 6974 2680
rect 7286 3848 7342 3904
rect 7378 2916 7434 2952
rect 7378 2896 7380 2916
rect 7380 2896 7432 2916
rect 7432 2896 7434 2916
rect 7654 5908 7710 5944
rect 7654 5888 7656 5908
rect 7656 5888 7708 5908
rect 7708 5888 7710 5908
rect 7562 5072 7618 5128
rect 7654 3576 7710 3632
rect 7746 3068 7748 3088
rect 7748 3068 7800 3088
rect 7800 3068 7802 3088
rect 7746 3032 7802 3068
rect 8390 14456 8446 14512
rect 9034 14320 9090 14376
rect 8390 13132 8392 13152
rect 8392 13132 8444 13152
rect 8444 13132 8446 13152
rect 8390 13096 8446 13132
rect 8390 12980 8446 13016
rect 8390 12960 8392 12980
rect 8392 12960 8444 12980
rect 8444 12960 8446 12980
rect 8574 12416 8630 12472
rect 8206 12144 8262 12200
rect 8298 11348 8354 11384
rect 8298 11328 8300 11348
rect 8300 11328 8352 11348
rect 8352 11328 8354 11348
rect 8574 10512 8630 10568
rect 8114 9696 8170 9752
rect 8022 8744 8078 8800
rect 8114 7520 8170 7576
rect 7930 5888 7986 5944
rect 8298 6704 8354 6760
rect 8298 6160 8354 6216
rect 8022 5344 8078 5400
rect 7930 4392 7986 4448
rect 8482 7812 8538 7848
rect 8482 7792 8484 7812
rect 8484 7792 8536 7812
rect 8536 7792 8538 7812
rect 8574 6976 8630 7032
rect 8482 6860 8538 6896
rect 8482 6840 8484 6860
rect 8484 6840 8536 6860
rect 8536 6840 8538 6860
rect 8850 13812 8852 13832
rect 8852 13812 8904 13832
rect 8904 13812 8906 13832
rect 8850 13776 8906 13812
rect 8758 13096 8814 13152
rect 8850 11056 8906 11112
rect 8574 5772 8630 5808
rect 8574 5752 8576 5772
rect 8576 5752 8628 5772
rect 8628 5752 8630 5772
rect 7930 3576 7986 3632
rect 8022 3032 8078 3088
rect 8390 2488 8446 2544
rect 8574 2524 8576 2544
rect 8576 2524 8628 2544
rect 8628 2524 8630 2544
rect 8574 2488 8630 2524
rect 8482 2080 8538 2136
rect 8114 1944 8170 2000
rect 11058 24928 11114 24984
rect 11518 24792 11574 24848
rect 10782 24656 10838 24712
rect 10690 23432 10746 23488
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 9494 22072 9550 22128
rect 9402 13524 9458 13560
rect 9402 13504 9404 13524
rect 9404 13504 9456 13524
rect 9456 13504 9458 13524
rect 9402 12552 9458 12608
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10874 20848 10930 20904
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 9770 16632 9826 16688
rect 9678 15988 9680 16008
rect 9680 15988 9732 16008
rect 9732 15988 9734 16008
rect 9678 15952 9734 15988
rect 10598 18128 10654 18184
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 11426 23568 11482 23624
rect 10874 18128 10930 18184
rect 10138 17604 10194 17640
rect 10138 17584 10140 17604
rect 10140 17584 10192 17604
rect 10192 17584 10194 17604
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10966 16496 11022 16552
rect 11150 16496 11206 16552
rect 9770 14068 9826 14104
rect 9770 14048 9772 14068
rect 9772 14048 9824 14068
rect 9824 14048 9826 14068
rect 9862 12688 9918 12744
rect 10046 12552 10102 12608
rect 9954 12144 10010 12200
rect 9586 11872 9642 11928
rect 9034 9288 9090 9344
rect 8942 5616 8998 5672
rect 8942 4936 8998 4992
rect 9310 7384 9366 7440
rect 9310 7248 9366 7304
rect 9218 7112 9274 7168
rect 9402 5636 9458 5672
rect 9402 5616 9404 5636
rect 9404 5616 9456 5636
rect 9456 5616 9458 5636
rect 9862 11056 9918 11112
rect 9954 9152 10010 9208
rect 10782 15544 10838 15600
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10782 13504 10838 13560
rect 10782 12824 10838 12880
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10598 10784 10654 10840
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10138 10240 10194 10296
rect 9954 8744 10010 8800
rect 9678 7112 9734 7168
rect 9586 6976 9642 7032
rect 9494 3984 9550 4040
rect 9218 3732 9274 3768
rect 9218 3712 9220 3732
rect 9220 3712 9272 3732
rect 9272 3712 9274 3732
rect 9402 3440 9458 3496
rect 9126 2760 9182 2816
rect 9954 6024 10010 6080
rect 9862 5888 9918 5944
rect 9862 3440 9918 3496
rect 9678 3032 9734 3088
rect 10598 9596 10600 9616
rect 10600 9596 10652 9616
rect 10652 9596 10654 9616
rect 10598 9560 10654 9596
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 11058 9424 11114 9480
rect 11058 8744 11114 8800
rect 10782 7112 10838 7168
rect 10230 6296 10286 6352
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10690 4800 10746 4856
rect 10782 4700 10784 4720
rect 10784 4700 10836 4720
rect 10836 4700 10838 4720
rect 10782 4664 10838 4700
rect 10138 3984 10194 4040
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10690 3732 10746 3768
rect 10690 3712 10692 3732
rect 10692 3712 10744 3732
rect 10744 3712 10746 3732
rect 10138 3032 10194 3088
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10506 2216 10562 2272
rect 10966 6568 11022 6624
rect 10966 4664 11022 4720
rect 10966 4120 11022 4176
rect 11058 3304 11114 3360
rect 11518 21936 11574 21992
rect 11702 19760 11758 19816
rect 12254 24132 12310 24168
rect 12254 24112 12256 24132
rect 12256 24112 12308 24132
rect 12308 24112 12310 24132
rect 12162 20440 12218 20496
rect 12622 20984 12678 21040
rect 12622 20848 12678 20904
rect 13450 23432 13506 23488
rect 12898 23044 12954 23080
rect 12898 23024 12900 23044
rect 12900 23024 12952 23044
rect 12952 23024 12954 23044
rect 13358 22500 13414 22536
rect 13358 22480 13360 22500
rect 13360 22480 13412 22500
rect 13412 22480 13414 22500
rect 12254 18808 12310 18864
rect 11978 18672 12034 18728
rect 11610 18128 11666 18184
rect 11426 15544 11482 15600
rect 11978 13096 12034 13152
rect 11886 12824 11942 12880
rect 11702 12552 11758 12608
rect 11518 12416 11574 12472
rect 11610 11872 11666 11928
rect 11242 11056 11298 11112
rect 11242 5228 11298 5264
rect 11242 5208 11244 5228
rect 11244 5208 11296 5228
rect 11296 5208 11298 5228
rect 11242 4936 11298 4992
rect 11242 4528 11298 4584
rect 11242 3848 11298 3904
rect 12162 14320 12218 14376
rect 12254 13932 12310 13968
rect 12254 13912 12256 13932
rect 12256 13912 12308 13932
rect 12308 13912 12310 13932
rect 12438 13912 12494 13968
rect 12346 12960 12402 13016
rect 12438 12280 12494 12336
rect 12346 12008 12402 12064
rect 12438 10784 12494 10840
rect 12162 10548 12164 10568
rect 12164 10548 12216 10568
rect 12216 10548 12218 10568
rect 12162 10512 12218 10548
rect 11518 6060 11520 6080
rect 11520 6060 11572 6080
rect 11572 6060 11574 6080
rect 11518 6024 11574 6060
rect 11610 5092 11666 5128
rect 11610 5072 11612 5092
rect 11612 5072 11664 5092
rect 11664 5072 11666 5092
rect 11426 4528 11482 4584
rect 10690 1672 10746 1728
rect 10966 2760 11022 2816
rect 10874 1264 10930 1320
rect 11886 5616 11942 5672
rect 12530 9696 12586 9752
rect 12438 9424 12494 9480
rect 12162 8336 12218 8392
rect 12162 7112 12218 7168
rect 12438 6840 12494 6896
rect 12898 19116 12900 19136
rect 12900 19116 12952 19136
rect 12952 19116 12954 19136
rect 12898 19080 12954 19116
rect 12990 17720 13046 17776
rect 12898 10260 12954 10296
rect 12898 10240 12900 10260
rect 12900 10240 12952 10260
rect 12952 10240 12954 10260
rect 12530 6160 12586 6216
rect 12438 5888 12494 5944
rect 11242 2760 11298 2816
rect 11150 2624 11206 2680
rect 11610 3440 11666 3496
rect 11426 2796 11428 2816
rect 11428 2796 11480 2816
rect 11480 2796 11482 2816
rect 11426 2760 11482 2796
rect 6366 312 6422 368
rect 12162 3304 12218 3360
rect 11978 2388 11980 2408
rect 11980 2388 12032 2408
rect 12032 2388 12034 2408
rect 11978 2352 12034 2388
rect 12162 2352 12218 2408
rect 12162 1944 12218 2000
rect 12898 5616 12954 5672
rect 12806 4392 12862 4448
rect 13266 19352 13322 19408
rect 13358 19216 13414 19272
rect 13726 21956 13782 21992
rect 13726 21936 13728 21956
rect 13728 21936 13780 21956
rect 13780 21936 13782 21956
rect 14278 24404 14334 24440
rect 14278 24384 14280 24404
rect 14280 24384 14332 24404
rect 14332 24384 14334 24404
rect 14094 21528 14150 21584
rect 13818 20304 13874 20360
rect 13818 17740 13874 17776
rect 13818 17720 13820 17740
rect 13820 17720 13872 17740
rect 13872 17720 13874 17740
rect 13082 12280 13138 12336
rect 14002 13776 14058 13832
rect 14370 22344 14426 22400
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15198 23740 15200 23760
rect 15200 23740 15252 23760
rect 15252 23740 15254 23760
rect 15198 23704 15254 23740
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 15198 22344 15254 22400
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14554 19352 14610 19408
rect 14462 17176 14518 17232
rect 14278 13368 14334 13424
rect 13634 12724 13636 12744
rect 13636 12724 13688 12744
rect 13688 12724 13690 12744
rect 13634 12688 13690 12724
rect 13358 11348 13414 11384
rect 13358 11328 13360 11348
rect 13360 11328 13412 11348
rect 13412 11328 13414 11348
rect 13082 10532 13138 10568
rect 13082 10512 13084 10532
rect 13084 10512 13136 10532
rect 13136 10512 13138 10532
rect 13174 9424 13230 9480
rect 13082 6740 13084 6760
rect 13084 6740 13136 6760
rect 13136 6740 13138 6760
rect 13082 6704 13138 6740
rect 13082 4936 13138 4992
rect 12438 3712 12494 3768
rect 12346 3576 12402 3632
rect 13174 2372 13230 2408
rect 13174 2352 13176 2372
rect 13176 2352 13228 2372
rect 13228 2352 13230 2372
rect 13450 5752 13506 5808
rect 13634 5752 13690 5808
rect 13910 10648 13966 10704
rect 13726 5344 13782 5400
rect 13634 5208 13690 5264
rect 13726 5072 13782 5128
rect 13818 3848 13874 3904
rect 13542 2352 13598 2408
rect 13910 3168 13966 3224
rect 13818 2080 13874 2136
rect 13726 1944 13782 2000
rect 14646 15428 14702 15464
rect 14646 15408 14648 15428
rect 14648 15408 14700 15428
rect 14700 15408 14702 15428
rect 14646 12552 14702 12608
rect 14462 11464 14518 11520
rect 14370 10648 14426 10704
rect 14370 10140 14372 10160
rect 14372 10140 14424 10160
rect 14424 10140 14426 10160
rect 14370 10104 14426 10140
rect 14278 9968 14334 10024
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 15658 23432 15714 23488
rect 15566 22924 15568 22944
rect 15568 22924 15620 22944
rect 15620 22924 15622 22944
rect 15566 22888 15622 22924
rect 15474 19080 15530 19136
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 15566 15952 15622 16008
rect 15106 15544 15162 15600
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 15290 13912 15346 13968
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 15014 11600 15070 11656
rect 14646 11228 14648 11248
rect 14648 11228 14700 11248
rect 14700 11228 14702 11248
rect 14646 11192 14702 11228
rect 14646 10956 14648 10976
rect 14648 10956 14700 10976
rect 14700 10956 14702 10976
rect 14646 10920 14702 10956
rect 14646 10784 14702 10840
rect 14646 10104 14702 10160
rect 14186 8608 14242 8664
rect 14278 8336 14334 8392
rect 14094 6996 14150 7032
rect 14094 6976 14096 6996
rect 14096 6976 14148 6996
rect 14148 6976 14150 6996
rect 14186 6024 14242 6080
rect 14094 4684 14150 4720
rect 14094 4664 14096 4684
rect 14096 4664 14148 4684
rect 14148 4664 14150 4684
rect 14278 4120 14334 4176
rect 14370 3712 14426 3768
rect 14554 8780 14556 8800
rect 14556 8780 14608 8800
rect 14608 8780 14610 8800
rect 14554 8744 14610 8780
rect 14462 856 14518 912
rect 14646 6604 14648 6624
rect 14648 6604 14700 6624
rect 14700 6604 14702 6624
rect 14646 6568 14702 6604
rect 15014 11092 15016 11112
rect 15016 11092 15068 11112
rect 15068 11092 15070 11112
rect 15014 11056 15070 11092
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14922 9052 14924 9072
rect 14924 9052 14976 9072
rect 14976 9052 14978 9072
rect 14922 9016 14978 9052
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14830 6976 14886 7032
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15658 13368 15714 13424
rect 15658 12708 15714 12744
rect 15658 12688 15660 12708
rect 15660 12688 15712 12708
rect 15712 12688 15714 12708
rect 15474 9968 15530 10024
rect 16210 24792 16266 24848
rect 16762 24656 16818 24712
rect 16118 24384 16174 24440
rect 17222 24384 17278 24440
rect 16486 24248 16542 24304
rect 17958 24792 18014 24848
rect 18970 24656 19026 24712
rect 19062 24384 19118 24440
rect 17774 24132 17830 24168
rect 17774 24112 17776 24132
rect 17776 24112 17828 24132
rect 17828 24112 17830 24132
rect 18326 23860 18382 23896
rect 18326 23840 18328 23860
rect 18328 23840 18380 23860
rect 18380 23840 18382 23860
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19522 24112 19578 24168
rect 19706 24112 19762 24168
rect 19522 23976 19578 24032
rect 20810 24656 20866 24712
rect 20258 23840 20314 23896
rect 17406 23432 17462 23488
rect 17498 22380 17500 22400
rect 17500 22380 17552 22400
rect 17552 22380 17554 22400
rect 17498 22344 17554 22380
rect 17038 22072 17094 22128
rect 16670 21956 16726 21992
rect 16670 21936 16672 21956
rect 16672 21936 16724 21956
rect 16724 21936 16726 21956
rect 16578 21528 16634 21584
rect 16026 21392 16082 21448
rect 17682 19896 17738 19952
rect 16118 19352 16174 19408
rect 15842 13388 15898 13424
rect 15842 13368 15844 13388
rect 15844 13368 15896 13388
rect 15896 13368 15898 13388
rect 16394 16496 16450 16552
rect 16394 15408 16450 15464
rect 16394 14356 16396 14376
rect 16396 14356 16448 14376
rect 16448 14356 16450 14376
rect 16394 14320 16450 14356
rect 16302 9832 16358 9888
rect 16854 13812 16856 13832
rect 16856 13812 16908 13832
rect 16908 13812 16910 13832
rect 16854 13776 16910 13812
rect 16670 13268 16672 13288
rect 16672 13268 16724 13288
rect 16724 13268 16726 13288
rect 16670 13232 16726 13268
rect 16670 10648 16726 10704
rect 17498 11192 17554 11248
rect 17222 10512 17278 10568
rect 15474 7284 15476 7304
rect 15476 7284 15528 7304
rect 15528 7284 15530 7304
rect 15474 7248 15530 7284
rect 15750 7404 15806 7440
rect 15750 7384 15752 7404
rect 15752 7384 15804 7404
rect 15804 7384 15806 7404
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15290 5072 15346 5128
rect 15474 5072 15530 5128
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15014 3984 15070 4040
rect 14646 3612 14648 3632
rect 14648 3612 14700 3632
rect 14700 3612 14702 3632
rect 14646 3576 14702 3612
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14738 2508 14794 2544
rect 14738 2488 14740 2508
rect 14740 2488 14792 2508
rect 14792 2488 14794 2508
rect 15198 3032 15254 3088
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15290 1264 15346 1320
rect 15474 1264 15530 1320
rect 16394 8064 16450 8120
rect 16762 6432 16818 6488
rect 16670 5752 16726 5808
rect 16946 5208 17002 5264
rect 16762 4528 16818 4584
rect 16394 3984 16450 4040
rect 16486 3576 16542 3632
rect 17130 2508 17186 2544
rect 17130 2488 17132 2508
rect 17132 2488 17184 2508
rect 17184 2488 17186 2508
rect 17866 16088 17922 16144
rect 17774 12280 17830 12336
rect 18050 11500 18052 11520
rect 18052 11500 18104 11520
rect 18104 11500 18106 11520
rect 18050 11464 18106 11500
rect 18050 11348 18106 11384
rect 18050 11328 18052 11348
rect 18052 11328 18104 11348
rect 18104 11328 18106 11348
rect 18602 22344 18658 22400
rect 18234 13912 18290 13968
rect 18326 13504 18382 13560
rect 18142 10240 18198 10296
rect 17958 8336 18014 8392
rect 17682 7928 17738 7984
rect 18050 6704 18106 6760
rect 17958 5616 18014 5672
rect 18510 12688 18566 12744
rect 18418 11872 18474 11928
rect 18418 8064 18474 8120
rect 18326 7248 18382 7304
rect 21362 23976 21418 24032
rect 21270 23860 21326 23896
rect 21270 23840 21272 23860
rect 21272 23840 21324 23860
rect 21324 23840 21326 23860
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 20902 23180 20958 23216
rect 20902 23160 20904 23180
rect 20904 23160 20956 23180
rect 20956 23160 20958 23180
rect 23110 23840 23166 23896
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24214 24792 24270 24848
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 23662 23568 23718 23624
rect 23570 23296 23626 23352
rect 21914 22888 21970 22944
rect 20810 17720 20866 17776
rect 19338 17176 19394 17232
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 18694 16496 18750 16552
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19154 13232 19210 13288
rect 19338 12824 19394 12880
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 20166 12280 20222 12336
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 18602 10104 18658 10160
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 18786 9868 18788 9888
rect 18788 9868 18840 9888
rect 18840 9868 18842 9888
rect 18786 9832 18842 9868
rect 18786 7112 18842 7168
rect 18234 4664 18290 4720
rect 17958 4120 18014 4176
rect 17774 3884 17776 3904
rect 17776 3884 17828 3904
rect 17828 3884 17830 3904
rect 17774 3848 17830 3884
rect 17406 2896 17462 2952
rect 17682 2896 17738 2952
rect 17406 2760 17462 2816
rect 16854 2080 16910 2136
rect 16946 1944 17002 2000
rect 16854 1808 16910 1864
rect 17130 1808 17186 1864
rect 17130 1400 17186 1456
rect 17314 1400 17370 1456
rect 18050 3304 18106 3360
rect 18418 4528 18474 4584
rect 18694 6160 18750 6216
rect 18510 3168 18566 3224
rect 18694 2644 18750 2680
rect 18694 2624 18696 2644
rect 18696 2624 18748 2644
rect 18748 2624 18750 2644
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19338 6976 19394 7032
rect 19338 6160 19394 6216
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19982 6840 20038 6896
rect 19522 6160 19578 6216
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19430 4972 19432 4992
rect 19432 4972 19484 4992
rect 19484 4972 19486 4992
rect 19430 4936 19486 4972
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19430 4800 19486 4856
rect 19798 3984 19854 4040
rect 26514 24248 26570 24304
rect 25962 24112 26018 24168
rect 27066 23704 27122 23760
rect 24766 23024 24822 23080
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 23570 21936 23626 21992
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 26238 13232 26294 13288
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 22374 8880 22430 8936
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 20350 8472 20406 8528
rect 20258 6432 20314 6488
rect 19246 3848 19302 3904
rect 18970 3732 19026 3768
rect 18970 3712 18972 3732
rect 18972 3712 19024 3732
rect 19024 3712 19026 3732
rect 19062 3440 19118 3496
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20166 3732 20222 3768
rect 20166 3712 20168 3732
rect 20168 3712 20220 3732
rect 20220 3712 20222 3732
rect 19430 3032 19486 3088
rect 19154 2352 19210 2408
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 19522 2080 19578 2136
rect 18878 1944 18934 2000
rect 18878 1536 18934 1592
rect 19062 1536 19118 1592
rect 18786 992 18842 1048
rect 19614 1400 19670 1456
rect 20074 1400 20130 1456
rect 22742 7792 22798 7848
rect 21362 7248 21418 7304
rect 22282 6452 22338 6488
rect 22282 6432 22284 6452
rect 22284 6432 22336 6452
rect 22336 6432 22338 6452
rect 22190 6160 22246 6216
rect 20718 4120 20774 4176
rect 20994 5344 21050 5400
rect 22282 5752 22338 5808
rect 20902 4684 20958 4720
rect 20902 4664 20904 4684
rect 20904 4664 20956 4684
rect 20956 4664 20958 4684
rect 20902 1808 20958 1864
rect 21362 3984 21418 4040
rect 21270 2760 21326 2816
rect 21178 1672 21234 1728
rect 21086 1264 21142 1320
rect 21638 3596 21694 3632
rect 21638 3576 21640 3596
rect 21640 3576 21692 3596
rect 21692 3576 21694 3596
rect 22282 3712 22338 3768
rect 21822 2896 21878 2952
rect 21546 2352 21602 2408
rect 21638 1944 21694 2000
rect 21454 1128 21510 1184
rect 22190 3304 22246 3360
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 23570 5208 23626 5264
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 26514 3984 26570 4040
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 23846 3188 23902 3224
rect 23846 3168 23848 3188
rect 23848 3168 23900 3188
rect 23900 3168 23902 3188
rect 23662 2896 23718 2952
rect 23110 2760 23166 2816
rect 23478 2760 23534 2816
rect 23478 2508 23534 2544
rect 23478 2488 23480 2508
rect 23480 2488 23532 2508
rect 23532 2488 23534 2508
rect 25318 2760 25374 2816
rect 24030 2352 24086 2408
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24214 1536 24270 1592
rect 11610 40 11666 96
rect 25962 1400 26018 1456
rect 27618 3440 27674 3496
rect 27066 856 27122 912
rect 24674 40 24730 96
<< metal3 >>
rect 0 27706 480 27736
rect 3049 27706 3115 27709
rect 0 27704 3115 27706
rect 0 27648 3054 27704
rect 3110 27648 3115 27704
rect 0 27646 3115 27648
rect 0 27616 480 27646
rect 3049 27643 3115 27646
rect 0 27162 480 27192
rect 3601 27162 3667 27165
rect 0 27160 3667 27162
rect 0 27104 3606 27160
rect 3662 27104 3667 27160
rect 0 27102 3667 27104
rect 0 27072 480 27102
rect 3601 27099 3667 27102
rect 0 26618 480 26648
rect 2773 26618 2839 26621
rect 0 26616 2839 26618
rect 0 26560 2778 26616
rect 2834 26560 2839 26616
rect 0 26558 2839 26560
rect 0 26528 480 26558
rect 2773 26555 2839 26558
rect 0 25938 480 25968
rect 4061 25938 4127 25941
rect 0 25936 4127 25938
rect 0 25880 4066 25936
rect 4122 25880 4127 25936
rect 0 25878 4127 25880
rect 0 25848 480 25878
rect 4061 25875 4127 25878
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25394 480 25424
rect 3233 25394 3299 25397
rect 0 25392 3299 25394
rect 0 25336 3238 25392
rect 3294 25336 3299 25392
rect 0 25334 3299 25336
rect 0 25304 480 25334
rect 3233 25331 3299 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 11053 24986 11119 24989
rect 9814 24984 11119 24986
rect 9814 24928 11058 24984
rect 11114 24928 11119 24984
rect 9814 24926 11119 24928
rect 0 24850 480 24880
rect 2037 24850 2103 24853
rect 9814 24850 9874 24926
rect 11053 24923 11119 24926
rect 0 24790 1226 24850
rect 0 24760 480 24790
rect 1166 24578 1226 24790
rect 2037 24848 9874 24850
rect 2037 24792 2042 24848
rect 2098 24792 9874 24848
rect 2037 24790 9874 24792
rect 9949 24850 10015 24853
rect 11513 24850 11579 24853
rect 9949 24848 11579 24850
rect 9949 24792 9954 24848
rect 10010 24792 11518 24848
rect 11574 24792 11579 24848
rect 9949 24790 11579 24792
rect 2037 24787 2103 24790
rect 9949 24787 10015 24790
rect 11513 24787 11579 24790
rect 16205 24850 16271 24853
rect 17953 24850 18019 24853
rect 24209 24850 24275 24853
rect 16205 24848 18019 24850
rect 16205 24792 16210 24848
rect 16266 24792 17958 24848
rect 18014 24792 18019 24848
rect 16205 24790 18019 24792
rect 16205 24787 16271 24790
rect 17953 24787 18019 24790
rect 18094 24848 24275 24850
rect 18094 24792 24214 24848
rect 24270 24792 24275 24848
rect 18094 24790 24275 24792
rect 1853 24714 1919 24717
rect 6545 24714 6611 24717
rect 1853 24712 6611 24714
rect 1853 24656 1858 24712
rect 1914 24656 6550 24712
rect 6606 24656 6611 24712
rect 1853 24654 6611 24656
rect 1853 24651 1919 24654
rect 6545 24651 6611 24654
rect 10777 24714 10843 24717
rect 16757 24714 16823 24717
rect 18094 24714 18154 24790
rect 24209 24787 24275 24790
rect 10777 24712 16823 24714
rect 10777 24656 10782 24712
rect 10838 24656 16762 24712
rect 16818 24656 16823 24712
rect 10777 24654 16823 24656
rect 10777 24651 10843 24654
rect 16757 24651 16823 24654
rect 16990 24654 18154 24714
rect 18965 24714 19031 24717
rect 20805 24714 20871 24717
rect 18965 24712 20871 24714
rect 18965 24656 18970 24712
rect 19026 24656 20810 24712
rect 20866 24656 20871 24712
rect 18965 24654 20871 24656
rect 4061 24578 4127 24581
rect 1166 24576 4127 24578
rect 1166 24520 4066 24576
rect 4122 24520 4127 24576
rect 1166 24518 4127 24520
rect 4061 24515 4127 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 14273 24442 14339 24445
rect 16113 24442 16179 24445
rect 16990 24442 17050 24654
rect 18965 24651 19031 24654
rect 20805 24651 20871 24654
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 14273 24440 16179 24442
rect 14273 24384 14278 24440
rect 14334 24384 16118 24440
rect 16174 24384 16179 24440
rect 14273 24382 16179 24384
rect 14273 24379 14339 24382
rect 16113 24379 16179 24382
rect 16254 24382 17050 24442
rect 17217 24442 17283 24445
rect 19057 24442 19123 24445
rect 17217 24440 19123 24442
rect 17217 24384 17222 24440
rect 17278 24384 19062 24440
rect 19118 24384 19123 24440
rect 17217 24382 19123 24384
rect 0 24170 480 24200
rect 3693 24170 3759 24173
rect 0 24168 3759 24170
rect 0 24112 3698 24168
rect 3754 24112 3759 24168
rect 0 24110 3759 24112
rect 0 24080 480 24110
rect 3693 24107 3759 24110
rect 12249 24170 12315 24173
rect 16254 24170 16314 24382
rect 17217 24379 17283 24382
rect 19057 24379 19123 24382
rect 16481 24306 16547 24309
rect 26509 24306 26575 24309
rect 16481 24304 26575 24306
rect 16481 24248 16486 24304
rect 16542 24248 26514 24304
rect 26570 24248 26575 24304
rect 16481 24246 26575 24248
rect 16481 24243 16547 24246
rect 26509 24243 26575 24246
rect 12249 24168 16314 24170
rect 12249 24112 12254 24168
rect 12310 24112 16314 24168
rect 12249 24110 16314 24112
rect 17769 24170 17835 24173
rect 19517 24170 19583 24173
rect 17769 24168 19583 24170
rect 17769 24112 17774 24168
rect 17830 24112 19522 24168
rect 19578 24112 19583 24168
rect 17769 24110 19583 24112
rect 12249 24107 12315 24110
rect 17769 24107 17835 24110
rect 19517 24107 19583 24110
rect 19701 24170 19767 24173
rect 25957 24170 26023 24173
rect 19701 24168 26023 24170
rect 19701 24112 19706 24168
rect 19762 24112 25962 24168
rect 26018 24112 26023 24168
rect 19701 24110 26023 24112
rect 19701 24107 19767 24110
rect 25957 24107 26023 24110
rect 19517 24034 19583 24037
rect 21357 24034 21423 24037
rect 19517 24032 21423 24034
rect 19517 23976 19522 24032
rect 19578 23976 21362 24032
rect 21418 23976 21423 24032
rect 19517 23974 21423 23976
rect 19517 23971 19583 23974
rect 21357 23971 21423 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 18321 23898 18387 23901
rect 20253 23898 20319 23901
rect 18321 23896 20319 23898
rect 18321 23840 18326 23896
rect 18382 23840 20258 23896
rect 20314 23840 20319 23896
rect 18321 23838 20319 23840
rect 18321 23835 18387 23838
rect 20253 23835 20319 23838
rect 21265 23898 21331 23901
rect 23105 23898 23171 23901
rect 21265 23896 23171 23898
rect 21265 23840 21270 23896
rect 21326 23840 23110 23896
rect 23166 23840 23171 23896
rect 21265 23838 23171 23840
rect 21265 23835 21331 23838
rect 23105 23835 23171 23838
rect 4245 23762 4311 23765
rect 9489 23762 9555 23765
rect 4245 23760 9555 23762
rect 4245 23704 4250 23760
rect 4306 23704 9494 23760
rect 9550 23704 9555 23760
rect 4245 23702 9555 23704
rect 4245 23699 4311 23702
rect 9489 23699 9555 23702
rect 15193 23762 15259 23765
rect 27061 23762 27127 23765
rect 15193 23760 27127 23762
rect 15193 23704 15198 23760
rect 15254 23704 27066 23760
rect 27122 23704 27127 23760
rect 15193 23702 27127 23704
rect 15193 23699 15259 23702
rect 27061 23699 27127 23702
rect 0 23626 480 23656
rect 1853 23626 1919 23629
rect 0 23624 1919 23626
rect 0 23568 1858 23624
rect 1914 23568 1919 23624
rect 0 23566 1919 23568
rect 0 23536 480 23566
rect 1853 23563 1919 23566
rect 2037 23626 2103 23629
rect 8753 23626 8819 23629
rect 2037 23624 8819 23626
rect 2037 23568 2042 23624
rect 2098 23568 8758 23624
rect 8814 23568 8819 23624
rect 2037 23566 8819 23568
rect 2037 23563 2103 23566
rect 8753 23563 8819 23566
rect 11421 23626 11487 23629
rect 23657 23626 23723 23629
rect 11421 23624 23723 23626
rect 11421 23568 11426 23624
rect 11482 23568 23662 23624
rect 23718 23568 23723 23624
rect 11421 23566 23723 23568
rect 11421 23563 11487 23566
rect 23657 23563 23723 23566
rect 5257 23490 5323 23493
rect 7465 23490 7531 23493
rect 5257 23488 7531 23490
rect 5257 23432 5262 23488
rect 5318 23432 7470 23488
rect 7526 23432 7531 23488
rect 5257 23430 7531 23432
rect 5257 23427 5323 23430
rect 7465 23427 7531 23430
rect 10685 23490 10751 23493
rect 13445 23490 13511 23493
rect 10685 23488 13511 23490
rect 10685 23432 10690 23488
rect 10746 23432 13450 23488
rect 13506 23432 13511 23488
rect 10685 23430 13511 23432
rect 10685 23427 10751 23430
rect 13445 23427 13511 23430
rect 15653 23490 15719 23493
rect 17401 23490 17467 23493
rect 15653 23488 17467 23490
rect 15653 23432 15658 23488
rect 15714 23432 17406 23488
rect 17462 23432 17467 23488
rect 15653 23430 17467 23432
rect 15653 23427 15719 23430
rect 17401 23427 17467 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 23565 23354 23631 23357
rect 27520 23354 28000 23384
rect 23565 23352 28000 23354
rect 23565 23296 23570 23352
rect 23626 23296 28000 23352
rect 23565 23294 28000 23296
rect 23565 23291 23631 23294
rect 27520 23264 28000 23294
rect 3049 23218 3115 23221
rect 20897 23218 20963 23221
rect 3049 23216 20963 23218
rect 3049 23160 3054 23216
rect 3110 23160 20902 23216
rect 20958 23160 20963 23216
rect 3049 23158 20963 23160
rect 3049 23155 3115 23158
rect 20897 23155 20963 23158
rect 0 23082 480 23112
rect 2865 23082 2931 23085
rect 0 23080 2931 23082
rect 0 23024 2870 23080
rect 2926 23024 2931 23080
rect 0 23022 2931 23024
rect 0 22992 480 23022
rect 2865 23019 2931 23022
rect 4061 23082 4127 23085
rect 6361 23082 6427 23085
rect 4061 23080 6427 23082
rect 4061 23024 4066 23080
rect 4122 23024 6366 23080
rect 6422 23024 6427 23080
rect 4061 23022 6427 23024
rect 4061 23019 4127 23022
rect 6361 23019 6427 23022
rect 12893 23082 12959 23085
rect 24761 23082 24827 23085
rect 12893 23080 24827 23082
rect 12893 23024 12898 23080
rect 12954 23024 24766 23080
rect 24822 23024 24827 23080
rect 12893 23022 24827 23024
rect 12893 23019 12959 23022
rect 24761 23019 24827 23022
rect 15561 22946 15627 22949
rect 21909 22946 21975 22949
rect 15561 22944 21975 22946
rect 15561 22888 15566 22944
rect 15622 22888 21914 22944
rect 21970 22888 21975 22944
rect 15561 22886 21975 22888
rect 15561 22883 15627 22886
rect 21909 22883 21975 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 5533 22674 5599 22677
rect 8385 22674 8451 22677
rect 5533 22672 8451 22674
rect 5533 22616 5538 22672
rect 5594 22616 8390 22672
rect 8446 22616 8451 22672
rect 5533 22614 8451 22616
rect 5533 22611 5599 22614
rect 8385 22611 8451 22614
rect 0 22538 480 22568
rect 2957 22538 3023 22541
rect 0 22536 3023 22538
rect 0 22480 2962 22536
rect 3018 22480 3023 22536
rect 0 22478 3023 22480
rect 0 22448 480 22478
rect 2957 22475 3023 22478
rect 6637 22538 6703 22541
rect 13353 22538 13419 22541
rect 6637 22536 13419 22538
rect 6637 22480 6642 22536
rect 6698 22480 13358 22536
rect 13414 22480 13419 22536
rect 6637 22478 13419 22480
rect 6637 22475 6703 22478
rect 13353 22475 13419 22478
rect 14365 22402 14431 22405
rect 15193 22402 15259 22405
rect 14365 22400 15259 22402
rect 14365 22344 14370 22400
rect 14426 22344 15198 22400
rect 15254 22344 15259 22400
rect 14365 22342 15259 22344
rect 14365 22339 14431 22342
rect 15193 22339 15259 22342
rect 17493 22402 17559 22405
rect 18597 22402 18663 22405
rect 17493 22400 18663 22402
rect 17493 22344 17498 22400
rect 17554 22344 18602 22400
rect 18658 22344 18663 22400
rect 17493 22342 18663 22344
rect 17493 22339 17559 22342
rect 18597 22339 18663 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 9489 22130 9555 22133
rect 17033 22130 17099 22133
rect 9489 22128 17099 22130
rect 9489 22072 9494 22128
rect 9550 22072 17038 22128
rect 17094 22072 17099 22128
rect 9489 22070 17099 22072
rect 9489 22067 9555 22070
rect 17033 22067 17099 22070
rect 8201 21994 8267 21997
rect 11513 21994 11579 21997
rect 8201 21992 11579 21994
rect 8201 21936 8206 21992
rect 8262 21936 11518 21992
rect 11574 21936 11579 21992
rect 8201 21934 11579 21936
rect 8201 21931 8267 21934
rect 11513 21931 11579 21934
rect 13721 21994 13787 21997
rect 16665 21994 16731 21997
rect 23565 21994 23631 21997
rect 13721 21992 23631 21994
rect 13721 21936 13726 21992
rect 13782 21936 16670 21992
rect 16726 21936 23570 21992
rect 23626 21936 23631 21992
rect 13721 21934 23631 21936
rect 13721 21931 13787 21934
rect 16665 21931 16731 21934
rect 23565 21931 23631 21934
rect 0 21858 480 21888
rect 1577 21858 1643 21861
rect 0 21856 1643 21858
rect 0 21800 1582 21856
rect 1638 21800 1643 21856
rect 0 21798 1643 21800
rect 0 21768 480 21798
rect 1577 21795 1643 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 14089 21586 14155 21589
rect 16573 21586 16639 21589
rect 14089 21584 16639 21586
rect 14089 21528 14094 21584
rect 14150 21528 16578 21584
rect 16634 21528 16639 21584
rect 14089 21526 16639 21528
rect 14089 21523 14155 21526
rect 16573 21523 16639 21526
rect 3509 21450 3575 21453
rect 8477 21450 8543 21453
rect 16021 21450 16087 21453
rect 3509 21448 8543 21450
rect 3509 21392 3514 21448
rect 3570 21392 8482 21448
rect 8538 21392 8543 21448
rect 3509 21390 8543 21392
rect 3509 21387 3575 21390
rect 8477 21387 8543 21390
rect 9262 21448 16087 21450
rect 9262 21392 16026 21448
rect 16082 21392 16087 21448
rect 9262 21390 16087 21392
rect 0 21314 480 21344
rect 1393 21314 1459 21317
rect 0 21312 1459 21314
rect 0 21256 1398 21312
rect 1454 21256 1459 21312
rect 0 21254 1459 21256
rect 0 21224 480 21254
rect 1393 21251 1459 21254
rect 6545 21314 6611 21317
rect 9121 21314 9187 21317
rect 9262 21314 9322 21390
rect 16021 21387 16087 21390
rect 6545 21312 9322 21314
rect 6545 21256 6550 21312
rect 6606 21256 9126 21312
rect 9182 21256 9322 21312
rect 6545 21254 9322 21256
rect 6545 21251 6611 21254
rect 9121 21251 9187 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 12617 21042 12683 21045
rect 2822 21040 12683 21042
rect 2822 20984 12622 21040
rect 12678 20984 12683 21040
rect 2822 20982 12683 20984
rect 2822 20906 2882 20982
rect 12617 20979 12683 20982
rect 2638 20846 2882 20906
rect 2957 20906 3023 20909
rect 7281 20906 7347 20909
rect 2957 20904 7347 20906
rect 2957 20848 2962 20904
rect 3018 20848 7286 20904
rect 7342 20848 7347 20904
rect 2957 20846 7347 20848
rect 0 20770 480 20800
rect 2638 20770 2698 20846
rect 2957 20843 3023 20846
rect 7281 20843 7347 20846
rect 10869 20906 10935 20909
rect 12617 20906 12683 20909
rect 10869 20904 12683 20906
rect 10869 20848 10874 20904
rect 10930 20848 12622 20904
rect 12678 20848 12683 20904
rect 10869 20846 12683 20848
rect 10869 20843 10935 20846
rect 12617 20843 12683 20846
rect 0 20710 2698 20770
rect 0 20680 480 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 7833 20498 7899 20501
rect 12157 20498 12223 20501
rect 7833 20496 12223 20498
rect 7833 20440 7838 20496
rect 7894 20440 12162 20496
rect 12218 20440 12223 20496
rect 7833 20438 12223 20440
rect 7833 20435 7899 20438
rect 12157 20435 12223 20438
rect 2865 20362 2931 20365
rect 13813 20362 13879 20365
rect 2865 20360 13879 20362
rect 2865 20304 2870 20360
rect 2926 20304 13818 20360
rect 13874 20304 13879 20360
rect 2865 20302 13879 20304
rect 2865 20299 2931 20302
rect 13813 20299 13879 20302
rect 10277 20160 10597 20161
rect 0 20090 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 2681 20090 2747 20093
rect 0 20088 2747 20090
rect 0 20032 2686 20088
rect 2742 20032 2747 20088
rect 0 20030 2747 20032
rect 0 20000 480 20030
rect 2681 20027 2747 20030
rect 2037 19954 2103 19957
rect 7005 19954 7071 19957
rect 2037 19952 7071 19954
rect 2037 19896 2042 19952
rect 2098 19896 7010 19952
rect 7066 19896 7071 19952
rect 2037 19894 7071 19896
rect 2037 19891 2103 19894
rect 7005 19891 7071 19894
rect 7281 19954 7347 19957
rect 17677 19954 17743 19957
rect 7281 19952 17743 19954
rect 7281 19896 7286 19952
rect 7342 19896 17682 19952
rect 17738 19896 17743 19952
rect 7281 19894 17743 19896
rect 7281 19891 7347 19894
rect 17677 19891 17743 19894
rect 2037 19818 2103 19821
rect 11697 19818 11763 19821
rect 2037 19816 11763 19818
rect 2037 19760 2042 19816
rect 2098 19760 11702 19816
rect 11758 19760 11763 19816
rect 2037 19758 11763 19760
rect 2037 19755 2103 19758
rect 11697 19755 11763 19758
rect 5610 19616 5930 19617
rect 0 19546 480 19576
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 2681 19546 2747 19549
rect 0 19544 2747 19546
rect 0 19488 2686 19544
rect 2742 19488 2747 19544
rect 0 19486 2747 19488
rect 0 19456 480 19486
rect 2681 19483 2747 19486
rect 13261 19410 13327 19413
rect 14549 19410 14615 19413
rect 16113 19410 16179 19413
rect 13261 19408 16179 19410
rect 13261 19352 13266 19408
rect 13322 19352 14554 19408
rect 14610 19352 16118 19408
rect 16174 19352 16179 19408
rect 13261 19350 16179 19352
rect 13261 19347 13327 19350
rect 14549 19347 14615 19350
rect 16113 19347 16179 19350
rect 2497 19274 2563 19277
rect 13353 19274 13419 19277
rect 2497 19272 13419 19274
rect 2497 19216 2502 19272
rect 2558 19216 13358 19272
rect 13414 19216 13419 19272
rect 2497 19214 13419 19216
rect 2497 19211 2563 19214
rect 13353 19211 13419 19214
rect 12893 19138 12959 19141
rect 15469 19138 15535 19141
rect 12893 19136 15535 19138
rect 12893 19080 12898 19136
rect 12954 19080 15474 19136
rect 15530 19080 15535 19136
rect 12893 19078 15535 19080
rect 12893 19075 12959 19078
rect 15469 19075 15535 19078
rect 10277 19072 10597 19073
rect 0 19002 480 19032
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 1393 19002 1459 19005
rect 0 19000 1459 19002
rect 0 18944 1398 19000
rect 1454 18944 1459 19000
rect 0 18942 1459 18944
rect 0 18912 480 18942
rect 1393 18939 1459 18942
rect 3233 19002 3299 19005
rect 7465 19002 7531 19005
rect 3233 19000 7531 19002
rect 3233 18944 3238 19000
rect 3294 18944 7470 19000
rect 7526 18944 7531 19000
rect 3233 18942 7531 18944
rect 3233 18939 3299 18942
rect 7465 18939 7531 18942
rect 2497 18866 2563 18869
rect 3601 18866 3667 18869
rect 5993 18866 6059 18869
rect 12249 18866 12315 18869
rect 2497 18864 5826 18866
rect 2497 18808 2502 18864
rect 2558 18808 3606 18864
rect 3662 18808 5826 18864
rect 2497 18806 5826 18808
rect 2497 18803 2563 18806
rect 3601 18803 3667 18806
rect 5766 18730 5826 18806
rect 5993 18864 12315 18866
rect 5993 18808 5998 18864
rect 6054 18808 12254 18864
rect 12310 18808 12315 18864
rect 5993 18806 12315 18808
rect 5993 18803 6059 18806
rect 12249 18803 12315 18806
rect 5993 18730 6059 18733
rect 5766 18728 6059 18730
rect 5766 18672 5998 18728
rect 6054 18672 6059 18728
rect 5766 18670 6059 18672
rect 5993 18667 6059 18670
rect 7925 18730 7991 18733
rect 9806 18730 9812 18732
rect 7925 18728 9812 18730
rect 7925 18672 7930 18728
rect 7986 18672 9812 18728
rect 7925 18670 9812 18672
rect 7925 18667 7991 18670
rect 9806 18668 9812 18670
rect 9876 18730 9882 18732
rect 11973 18730 12039 18733
rect 9876 18728 12039 18730
rect 9876 18672 11978 18728
rect 12034 18672 12039 18728
rect 9876 18670 12039 18672
rect 9876 18668 9882 18670
rect 11973 18667 12039 18670
rect 5610 18528 5930 18529
rect 0 18458 480 18488
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 1577 18458 1643 18461
rect 0 18456 1643 18458
rect 0 18400 1582 18456
rect 1638 18400 1643 18456
rect 0 18398 1643 18400
rect 0 18368 480 18398
rect 1577 18395 1643 18398
rect 3785 18186 3851 18189
rect 4521 18186 4587 18189
rect 10593 18186 10659 18189
rect 3785 18184 10659 18186
rect 3785 18128 3790 18184
rect 3846 18128 4526 18184
rect 4582 18128 10598 18184
rect 10654 18128 10659 18184
rect 3785 18126 10659 18128
rect 3785 18123 3851 18126
rect 4521 18123 4587 18126
rect 10593 18123 10659 18126
rect 10869 18186 10935 18189
rect 11605 18186 11671 18189
rect 10869 18184 11671 18186
rect 10869 18128 10874 18184
rect 10930 18128 11610 18184
rect 11666 18128 11671 18184
rect 10869 18126 11671 18128
rect 10869 18123 10935 18126
rect 11605 18123 11671 18126
rect 6821 18050 6887 18053
rect 7557 18050 7623 18053
rect 6821 18048 9874 18050
rect 6821 17992 6826 18048
rect 6882 17992 7562 18048
rect 7618 17992 9874 18048
rect 6821 17990 9874 17992
rect 6821 17987 6887 17990
rect 7557 17987 7623 17990
rect 0 17778 480 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 9814 17778 9874 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 12985 17778 13051 17781
rect 9814 17776 13051 17778
rect 9814 17720 12990 17776
rect 13046 17720 13051 17776
rect 9814 17718 13051 17720
rect 0 17688 480 17718
rect 1393 17715 1459 17718
rect 12985 17715 13051 17718
rect 13813 17778 13879 17781
rect 20805 17778 20871 17781
rect 13813 17776 20871 17778
rect 13813 17720 13818 17776
rect 13874 17720 20810 17776
rect 20866 17720 20871 17776
rect 13813 17718 20871 17720
rect 13813 17715 13879 17718
rect 20805 17715 20871 17718
rect 2221 17642 2287 17645
rect 10133 17642 10199 17645
rect 2221 17640 10199 17642
rect 2221 17584 2226 17640
rect 2282 17584 10138 17640
rect 10194 17584 10199 17640
rect 2221 17582 10199 17584
rect 2221 17579 2287 17582
rect 10133 17579 10199 17582
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 0 17234 480 17264
rect 2681 17234 2747 17237
rect 0 17232 2747 17234
rect 0 17176 2686 17232
rect 2742 17176 2747 17232
rect 0 17174 2747 17176
rect 0 17144 480 17174
rect 2681 17171 2747 17174
rect 3325 17234 3391 17237
rect 5533 17234 5599 17237
rect 3325 17232 5599 17234
rect 3325 17176 3330 17232
rect 3386 17176 5538 17232
rect 5594 17176 5599 17232
rect 3325 17174 5599 17176
rect 3325 17171 3391 17174
rect 5533 17171 5599 17174
rect 14457 17234 14523 17237
rect 19333 17234 19399 17237
rect 14457 17232 19399 17234
rect 14457 17176 14462 17232
rect 14518 17176 19338 17232
rect 19394 17176 19399 17232
rect 14457 17174 19399 17176
rect 14457 17171 14523 17174
rect 19333 17171 19399 17174
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 1485 16826 1551 16829
rect 798 16824 1551 16826
rect 798 16768 1490 16824
rect 1546 16768 1551 16824
rect 798 16766 1551 16768
rect 0 16690 480 16720
rect 798 16690 858 16766
rect 1485 16763 1551 16766
rect 3141 16826 3207 16829
rect 8569 16826 8635 16829
rect 3141 16824 8635 16826
rect 3141 16768 3146 16824
rect 3202 16768 8574 16824
rect 8630 16768 8635 16824
rect 3141 16766 8635 16768
rect 3141 16763 3207 16766
rect 8569 16763 8635 16766
rect 0 16630 858 16690
rect 5717 16690 5783 16693
rect 9765 16690 9831 16693
rect 5717 16688 9831 16690
rect 5717 16632 5722 16688
rect 5778 16632 9770 16688
rect 9826 16632 9831 16688
rect 5717 16630 9831 16632
rect 0 16600 480 16630
rect 5717 16627 5783 16630
rect 9765 16627 9831 16630
rect 2037 16554 2103 16557
rect 5625 16554 5691 16557
rect 2037 16552 5691 16554
rect 2037 16496 2042 16552
rect 2098 16496 5630 16552
rect 5686 16496 5691 16552
rect 2037 16494 5691 16496
rect 2037 16491 2103 16494
rect 5625 16491 5691 16494
rect 10961 16554 11027 16557
rect 11145 16554 11211 16557
rect 10961 16552 11211 16554
rect 10961 16496 10966 16552
rect 11022 16496 11150 16552
rect 11206 16496 11211 16552
rect 10961 16494 11211 16496
rect 10961 16491 11027 16494
rect 11145 16491 11211 16494
rect 16389 16554 16455 16557
rect 18689 16554 18755 16557
rect 16389 16552 18755 16554
rect 16389 16496 16394 16552
rect 16450 16496 18694 16552
rect 18750 16496 18755 16552
rect 16389 16494 18755 16496
rect 16389 16491 16455 16494
rect 18689 16491 18755 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 7833 16146 7899 16149
rect 17861 16146 17927 16149
rect 7833 16144 17927 16146
rect 7833 16088 7838 16144
rect 7894 16088 17866 16144
rect 17922 16088 17927 16144
rect 7833 16086 17927 16088
rect 7833 16083 7899 16086
rect 17861 16083 17927 16086
rect 0 16010 480 16040
rect 1577 16010 1643 16013
rect 0 16008 1643 16010
rect 0 15952 1582 16008
rect 1638 15952 1643 16008
rect 0 15950 1643 15952
rect 0 15920 480 15950
rect 1577 15947 1643 15950
rect 3233 16010 3299 16013
rect 8109 16010 8175 16013
rect 3233 16008 8175 16010
rect 3233 15952 3238 16008
rect 3294 15952 8114 16008
rect 8170 15952 8175 16008
rect 3233 15950 8175 15952
rect 3233 15947 3299 15950
rect 8109 15947 8175 15950
rect 9673 16010 9739 16013
rect 15561 16010 15627 16013
rect 9673 16008 15627 16010
rect 9673 15952 9678 16008
rect 9734 15952 15566 16008
rect 15622 15952 15627 16008
rect 9673 15950 15627 15952
rect 9673 15947 9739 15950
rect 15561 15947 15627 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 1945 15738 2011 15741
rect 4245 15738 4311 15741
rect 1945 15736 4311 15738
rect 1945 15680 1950 15736
rect 2006 15680 4250 15736
rect 4306 15680 4311 15736
rect 1945 15678 4311 15680
rect 1945 15675 2011 15678
rect 4245 15675 4311 15678
rect 2037 15602 2103 15605
rect 10777 15602 10843 15605
rect 2037 15600 10843 15602
rect 2037 15544 2042 15600
rect 2098 15544 10782 15600
rect 10838 15544 10843 15600
rect 2037 15542 10843 15544
rect 2037 15539 2103 15542
rect 10777 15539 10843 15542
rect 11421 15602 11487 15605
rect 15101 15602 15167 15605
rect 11421 15600 15167 15602
rect 11421 15544 11426 15600
rect 11482 15544 15106 15600
rect 15162 15544 15167 15600
rect 11421 15542 15167 15544
rect 11421 15539 11487 15542
rect 15101 15539 15167 15542
rect 0 15466 480 15496
rect 1393 15466 1459 15469
rect 0 15464 1459 15466
rect 0 15408 1398 15464
rect 1454 15408 1459 15464
rect 0 15406 1459 15408
rect 0 15376 480 15406
rect 1393 15403 1459 15406
rect 5165 15466 5231 15469
rect 14641 15466 14707 15469
rect 16389 15466 16455 15469
rect 5165 15464 14707 15466
rect 5165 15408 5170 15464
rect 5226 15408 14646 15464
rect 14702 15408 14707 15464
rect 5165 15406 14707 15408
rect 5165 15403 5231 15406
rect 14641 15403 14707 15406
rect 14782 15464 16455 15466
rect 14782 15408 16394 15464
rect 16450 15408 16455 15464
rect 14782 15406 16455 15408
rect 2221 15330 2287 15333
rect 4797 15330 4863 15333
rect 2221 15328 4863 15330
rect 2221 15272 2226 15328
rect 2282 15272 4802 15328
rect 4858 15272 4863 15328
rect 2221 15270 4863 15272
rect 2221 15267 2287 15270
rect 4797 15267 4863 15270
rect 6269 15330 6335 15333
rect 7649 15330 7715 15333
rect 14782 15330 14842 15406
rect 16389 15403 16455 15406
rect 6269 15328 14842 15330
rect 6269 15272 6274 15328
rect 6330 15272 7654 15328
rect 7710 15272 14842 15328
rect 6269 15270 14842 15272
rect 6269 15267 6335 15270
rect 7649 15267 7715 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 0 14922 480 14952
rect 1577 14922 1643 14925
rect 0 14920 1643 14922
rect 0 14864 1582 14920
rect 1638 14864 1643 14920
rect 0 14862 1643 14864
rect 0 14832 480 14862
rect 1577 14859 1643 14862
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 1853 14514 1919 14517
rect 8385 14514 8451 14517
rect 1853 14512 8451 14514
rect 1853 14456 1858 14512
rect 1914 14456 8390 14512
rect 8446 14456 8451 14512
rect 1853 14454 8451 14456
rect 1853 14451 1919 14454
rect 8385 14451 8451 14454
rect 0 14378 480 14408
rect 2681 14378 2747 14381
rect 0 14376 2747 14378
rect 0 14320 2686 14376
rect 2742 14320 2747 14376
rect 0 14318 2747 14320
rect 0 14288 480 14318
rect 2681 14315 2747 14318
rect 3233 14378 3299 14381
rect 9029 14378 9095 14381
rect 3233 14376 9095 14378
rect 3233 14320 3238 14376
rect 3294 14320 9034 14376
rect 9090 14320 9095 14376
rect 3233 14318 9095 14320
rect 3233 14315 3299 14318
rect 9029 14315 9095 14318
rect 12157 14378 12223 14381
rect 16389 14378 16455 14381
rect 12157 14376 16455 14378
rect 12157 14320 12162 14376
rect 12218 14320 16394 14376
rect 16450 14320 16455 14376
rect 12157 14318 16455 14320
rect 12157 14315 12223 14318
rect 16389 14315 16455 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 6085 14106 6151 14109
rect 9765 14106 9831 14109
rect 6085 14104 9831 14106
rect 6085 14048 6090 14104
rect 6146 14048 9770 14104
rect 9826 14048 9831 14104
rect 6085 14046 9831 14048
rect 6085 14043 6151 14046
rect 9765 14043 9831 14046
rect 12249 13970 12315 13973
rect 12433 13970 12499 13973
rect 15285 13970 15351 13973
rect 12249 13968 15351 13970
rect 12249 13912 12254 13968
rect 12310 13912 12438 13968
rect 12494 13912 15290 13968
rect 15346 13912 15351 13968
rect 12249 13910 15351 13912
rect 12249 13907 12315 13910
rect 12433 13907 12499 13910
rect 15285 13907 15351 13910
rect 18229 13970 18295 13973
rect 27520 13970 28000 14000
rect 18229 13968 28000 13970
rect 18229 13912 18234 13968
rect 18290 13912 28000 13968
rect 18229 13910 28000 13912
rect 18229 13907 18295 13910
rect 27520 13880 28000 13910
rect 2037 13834 2103 13837
rect 3877 13834 3943 13837
rect 6821 13834 6887 13837
rect 2037 13832 6887 13834
rect 2037 13776 2042 13832
rect 2098 13776 3882 13832
rect 3938 13776 6826 13832
rect 6882 13776 6887 13832
rect 2037 13774 6887 13776
rect 2037 13771 2103 13774
rect 3877 13771 3943 13774
rect 6821 13771 6887 13774
rect 8845 13834 8911 13837
rect 13997 13834 14063 13837
rect 16849 13834 16915 13837
rect 8845 13832 16915 13834
rect 8845 13776 8850 13832
rect 8906 13776 14002 13832
rect 14058 13776 16854 13832
rect 16910 13776 16915 13832
rect 8845 13774 16915 13776
rect 8845 13771 8911 13774
rect 13997 13771 14063 13774
rect 16849 13771 16915 13774
rect 0 13698 480 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 480 13638
rect 1393 13635 1459 13638
rect 2865 13698 2931 13701
rect 6269 13698 6335 13701
rect 2865 13696 6335 13698
rect 2865 13640 2870 13696
rect 2926 13640 6274 13696
rect 6330 13640 6335 13696
rect 2865 13638 6335 13640
rect 2865 13635 2931 13638
rect 6269 13635 6335 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 2773 13562 2839 13565
rect 4337 13562 4403 13565
rect 4889 13562 4955 13565
rect 2773 13560 4955 13562
rect 2773 13504 2778 13560
rect 2834 13504 4342 13560
rect 4398 13504 4894 13560
rect 4950 13504 4955 13560
rect 2773 13502 4955 13504
rect 2773 13499 2839 13502
rect 4337 13499 4403 13502
rect 4889 13499 4955 13502
rect 5441 13562 5507 13565
rect 9397 13562 9463 13565
rect 5441 13560 9463 13562
rect 5441 13504 5446 13560
rect 5502 13504 9402 13560
rect 9458 13504 9463 13560
rect 5441 13502 9463 13504
rect 5441 13499 5507 13502
rect 9397 13499 9463 13502
rect 10777 13562 10843 13565
rect 18321 13562 18387 13565
rect 10777 13560 18387 13562
rect 10777 13504 10782 13560
rect 10838 13504 18326 13560
rect 18382 13504 18387 13560
rect 10777 13502 18387 13504
rect 10777 13499 10843 13502
rect 18321 13499 18387 13502
rect 1393 13426 1459 13429
rect 3693 13426 3759 13429
rect 1393 13424 3759 13426
rect 1393 13368 1398 13424
rect 1454 13368 3698 13424
rect 3754 13368 3759 13424
rect 1393 13366 3759 13368
rect 1393 13363 1459 13366
rect 3693 13363 3759 13366
rect 5165 13426 5231 13429
rect 14273 13426 14339 13429
rect 5165 13424 14339 13426
rect 5165 13368 5170 13424
rect 5226 13368 14278 13424
rect 14334 13368 14339 13424
rect 5165 13366 14339 13368
rect 5165 13363 5231 13366
rect 14273 13363 14339 13366
rect 15653 13426 15719 13429
rect 15837 13426 15903 13429
rect 15653 13424 15762 13426
rect 15653 13368 15658 13424
rect 15714 13368 15762 13424
rect 15653 13363 15762 13368
rect 15837 13424 16866 13426
rect 15837 13368 15842 13424
rect 15898 13368 16866 13424
rect 15837 13366 16866 13368
rect 15837 13363 15903 13366
rect 1669 13290 1735 13293
rect 3141 13290 3207 13293
rect 1669 13288 3207 13290
rect 1669 13232 1674 13288
rect 1730 13232 3146 13288
rect 3202 13232 3207 13288
rect 1669 13230 3207 13232
rect 1669 13227 1735 13230
rect 3141 13227 3207 13230
rect 5625 13290 5691 13293
rect 15702 13290 15762 13363
rect 16665 13290 16731 13293
rect 5625 13288 16731 13290
rect 5625 13232 5630 13288
rect 5686 13232 16670 13288
rect 16726 13232 16731 13288
rect 5625 13230 16731 13232
rect 16806 13290 16866 13366
rect 19149 13290 19215 13293
rect 26233 13290 26299 13293
rect 16806 13288 26299 13290
rect 16806 13232 19154 13288
rect 19210 13232 26238 13288
rect 26294 13232 26299 13288
rect 16806 13230 26299 13232
rect 5625 13227 5691 13230
rect 16665 13227 16731 13230
rect 19149 13227 19215 13230
rect 26233 13227 26299 13230
rect 0 13154 480 13184
rect 1577 13154 1643 13157
rect 0 13152 1643 13154
rect 0 13096 1582 13152
rect 1638 13096 1643 13152
rect 0 13094 1643 13096
rect 0 13064 480 13094
rect 1577 13091 1643 13094
rect 6177 13154 6243 13157
rect 8385 13154 8451 13157
rect 6177 13152 8451 13154
rect 6177 13096 6182 13152
rect 6238 13096 8390 13152
rect 8446 13096 8451 13152
rect 6177 13094 8451 13096
rect 6177 13091 6243 13094
rect 8385 13091 8451 13094
rect 8753 13154 8819 13157
rect 11973 13154 12039 13157
rect 8753 13152 12039 13154
rect 8753 13096 8758 13152
rect 8814 13096 11978 13152
rect 12034 13096 12039 13152
rect 8753 13094 12039 13096
rect 8753 13091 8819 13094
rect 11973 13091 12039 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 6361 13018 6427 13021
rect 8385 13018 8451 13021
rect 12341 13018 12407 13021
rect 6361 13016 12407 13018
rect 6361 12960 6366 13016
rect 6422 12960 8390 13016
rect 8446 12960 12346 13016
rect 12402 12960 12407 13016
rect 6361 12958 12407 12960
rect 6361 12955 6427 12958
rect 8385 12955 8451 12958
rect 12341 12955 12407 12958
rect 13 12882 79 12885
rect 3601 12882 3667 12885
rect 10777 12882 10843 12885
rect 13 12880 3480 12882
rect 13 12824 18 12880
rect 74 12824 3480 12880
rect 13 12822 3480 12824
rect 13 12819 79 12822
rect 3420 12746 3480 12822
rect 3601 12880 10843 12882
rect 3601 12824 3606 12880
rect 3662 12824 10782 12880
rect 10838 12824 10843 12880
rect 3601 12822 10843 12824
rect 3601 12819 3667 12822
rect 10777 12819 10843 12822
rect 11881 12882 11947 12885
rect 19333 12882 19399 12885
rect 11881 12880 19399 12882
rect 11881 12824 11886 12880
rect 11942 12824 19338 12880
rect 19394 12824 19399 12880
rect 11881 12822 19399 12824
rect 11881 12819 11947 12822
rect 19333 12819 19399 12822
rect 7189 12746 7255 12749
rect 9857 12746 9923 12749
rect 13629 12746 13695 12749
rect 3420 12686 6424 12746
rect 0 12610 480 12640
rect 1577 12610 1643 12613
rect 0 12608 1643 12610
rect 0 12552 1582 12608
rect 1638 12552 1643 12608
rect 0 12550 1643 12552
rect 0 12520 480 12550
rect 1577 12547 1643 12550
rect 2313 12610 2379 12613
rect 3233 12610 3299 12613
rect 2313 12608 3299 12610
rect 2313 12552 2318 12608
rect 2374 12552 3238 12608
rect 3294 12552 3299 12608
rect 2313 12550 3299 12552
rect 2313 12547 2379 12550
rect 3233 12547 3299 12550
rect 3877 12610 3943 12613
rect 5625 12610 5691 12613
rect 3877 12608 5691 12610
rect 3877 12552 3882 12608
rect 3938 12552 5630 12608
rect 5686 12552 5691 12608
rect 3877 12550 5691 12552
rect 6364 12610 6424 12686
rect 7189 12744 9923 12746
rect 7189 12688 7194 12744
rect 7250 12688 9862 12744
rect 9918 12688 9923 12744
rect 7189 12686 9923 12688
rect 7189 12683 7255 12686
rect 9857 12683 9923 12686
rect 10044 12744 13695 12746
rect 10044 12688 13634 12744
rect 13690 12688 13695 12744
rect 10044 12686 13695 12688
rect 10044 12613 10104 12686
rect 13629 12683 13695 12686
rect 15653 12746 15719 12749
rect 18505 12746 18571 12749
rect 15653 12744 18571 12746
rect 15653 12688 15658 12744
rect 15714 12688 18510 12744
rect 18566 12688 18571 12744
rect 15653 12686 18571 12688
rect 15653 12683 15719 12686
rect 18505 12683 18571 12686
rect 9397 12610 9463 12613
rect 10041 12610 10107 12613
rect 6364 12608 10107 12610
rect 6364 12552 9402 12608
rect 9458 12552 10046 12608
rect 10102 12552 10107 12608
rect 6364 12550 10107 12552
rect 3877 12547 3943 12550
rect 5625 12547 5691 12550
rect 9397 12547 9463 12550
rect 10041 12547 10107 12550
rect 11697 12610 11763 12613
rect 14641 12610 14707 12613
rect 11697 12608 14707 12610
rect 11697 12552 11702 12608
rect 11758 12552 14646 12608
rect 14702 12552 14707 12608
rect 11697 12550 14707 12552
rect 11697 12547 11763 12550
rect 14641 12547 14707 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 8569 12474 8635 12477
rect 11513 12474 11579 12477
rect 8569 12472 10196 12474
rect 8569 12416 8574 12472
rect 8630 12416 10196 12472
rect 8569 12414 10196 12416
rect 8569 12411 8635 12414
rect 10136 12338 10196 12414
rect 11513 12472 18338 12474
rect 11513 12416 11518 12472
rect 11574 12416 18338 12472
rect 11513 12414 18338 12416
rect 11513 12411 11579 12414
rect 12433 12338 12499 12341
rect 10136 12336 12499 12338
rect 10136 12280 12438 12336
rect 12494 12280 12499 12336
rect 10136 12278 12499 12280
rect 12433 12275 12499 12278
rect 13077 12338 13143 12341
rect 17769 12338 17835 12341
rect 13077 12336 17835 12338
rect 13077 12280 13082 12336
rect 13138 12280 17774 12336
rect 17830 12280 17835 12336
rect 13077 12278 17835 12280
rect 18278 12338 18338 12414
rect 20161 12338 20227 12341
rect 18278 12336 20227 12338
rect 18278 12280 20166 12336
rect 20222 12280 20227 12336
rect 18278 12278 20227 12280
rect 13077 12275 13143 12278
rect 17769 12275 17835 12278
rect 20161 12275 20227 12278
rect 8201 12202 8267 12205
rect 9949 12202 10015 12205
rect 8201 12200 10015 12202
rect 8201 12144 8206 12200
rect 8262 12144 9954 12200
rect 10010 12144 10015 12200
rect 8201 12142 10015 12144
rect 8201 12139 8267 12142
rect 9949 12139 10015 12142
rect 5993 12066 6059 12069
rect 12341 12066 12407 12069
rect 5993 12064 12407 12066
rect 5993 12008 5998 12064
rect 6054 12008 12346 12064
rect 12402 12008 12407 12064
rect 5993 12006 12407 12008
rect 5993 12003 6059 12006
rect 12341 12003 12407 12006
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 4245 11930 4311 11933
rect 0 11928 4311 11930
rect 0 11872 4250 11928
rect 4306 11872 4311 11928
rect 0 11870 4311 11872
rect 0 11840 480 11870
rect 4245 11867 4311 11870
rect 7097 11930 7163 11933
rect 8150 11930 8156 11932
rect 7097 11928 8156 11930
rect 7097 11872 7102 11928
rect 7158 11872 8156 11928
rect 7097 11870 8156 11872
rect 7097 11867 7163 11870
rect 8150 11868 8156 11870
rect 8220 11868 8226 11932
rect 9581 11930 9647 11933
rect 11605 11930 11671 11933
rect 9581 11928 11671 11930
rect 9581 11872 9586 11928
rect 9642 11872 11610 11928
rect 11666 11872 11671 11928
rect 9581 11870 11671 11872
rect 9581 11867 9647 11870
rect 11605 11867 11671 11870
rect 18270 11868 18276 11932
rect 18340 11930 18346 11932
rect 18413 11930 18479 11933
rect 18340 11928 18479 11930
rect 18340 11872 18418 11928
rect 18474 11872 18479 11928
rect 18340 11870 18479 11872
rect 18340 11868 18346 11870
rect 18413 11867 18479 11870
rect 4337 11658 4403 11661
rect 15009 11658 15075 11661
rect 4337 11656 15075 11658
rect 4337 11600 4342 11656
rect 4398 11600 15014 11656
rect 15070 11600 15075 11656
rect 4337 11598 15075 11600
rect 4337 11595 4403 11598
rect 15009 11595 15075 11598
rect 1761 11522 1827 11525
rect 4061 11522 4127 11525
rect 1761 11520 4127 11522
rect 1761 11464 1766 11520
rect 1822 11464 4066 11520
rect 4122 11464 4127 11520
rect 1761 11462 4127 11464
rect 1761 11459 1827 11462
rect 4061 11459 4127 11462
rect 14457 11522 14523 11525
rect 18045 11522 18111 11525
rect 14457 11520 18111 11522
rect 14457 11464 14462 11520
rect 14518 11464 18050 11520
rect 18106 11464 18111 11520
rect 14457 11462 18111 11464
rect 14457 11459 14523 11462
rect 18045 11459 18111 11462
rect 10277 11456 10597 11457
rect 0 11386 480 11416
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 3601 11386 3667 11389
rect 0 11384 3667 11386
rect 0 11328 3606 11384
rect 3662 11328 3667 11384
rect 0 11326 3667 11328
rect 0 11296 480 11326
rect 3601 11323 3667 11326
rect 7005 11386 7071 11389
rect 7833 11386 7899 11389
rect 8293 11386 8359 11389
rect 7005 11384 8359 11386
rect 7005 11328 7010 11384
rect 7066 11328 7838 11384
rect 7894 11328 8298 11384
rect 8354 11328 8359 11384
rect 7005 11326 8359 11328
rect 7005 11323 7071 11326
rect 7833 11323 7899 11326
rect 8293 11323 8359 11326
rect 13353 11386 13419 11389
rect 18045 11386 18111 11389
rect 13353 11384 18111 11386
rect 13353 11328 13358 11384
rect 13414 11328 18050 11384
rect 18106 11328 18111 11384
rect 13353 11326 18111 11328
rect 13353 11323 13419 11326
rect 18045 11323 18111 11326
rect 3877 11250 3943 11253
rect 14641 11250 14707 11253
rect 3877 11248 14707 11250
rect 3877 11192 3882 11248
rect 3938 11192 14646 11248
rect 14702 11192 14707 11248
rect 3877 11190 14707 11192
rect 3877 11187 3943 11190
rect 14641 11187 14707 11190
rect 17493 11250 17559 11253
rect 17718 11250 17724 11252
rect 17493 11248 17724 11250
rect 17493 11192 17498 11248
rect 17554 11192 17724 11248
rect 17493 11190 17724 11192
rect 17493 11187 17559 11190
rect 17718 11188 17724 11190
rect 17788 11188 17794 11252
rect 7925 11114 7991 11117
rect 8845 11114 8911 11117
rect 7925 11112 8911 11114
rect 7925 11056 7930 11112
rect 7986 11056 8850 11112
rect 8906 11056 8911 11112
rect 7925 11054 8911 11056
rect 7925 11051 7991 11054
rect 8845 11051 8911 11054
rect 9857 11114 9923 11117
rect 11237 11114 11303 11117
rect 15009 11114 15075 11117
rect 9857 11112 15075 11114
rect 9857 11056 9862 11112
rect 9918 11056 11242 11112
rect 11298 11056 15014 11112
rect 15070 11056 15075 11112
rect 9857 11054 15075 11056
rect 9857 11051 9923 11054
rect 11237 11051 11303 11054
rect 15009 11051 15075 11054
rect 1853 10978 1919 10981
rect 1853 10976 5458 10978
rect 1853 10920 1858 10976
rect 1914 10920 5458 10976
rect 1853 10918 5458 10920
rect 1853 10915 1919 10918
rect 0 10842 480 10872
rect 0 10782 2744 10842
rect 0 10752 480 10782
rect 2684 10706 2744 10782
rect 5398 10706 5458 10918
rect 9990 10916 9996 10980
rect 10060 10978 10066 10980
rect 14641 10978 14707 10981
rect 10060 10976 14707 10978
rect 10060 10920 14646 10976
rect 14702 10920 14707 10976
rect 10060 10918 14707 10920
rect 10060 10916 10066 10918
rect 14641 10915 14707 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 6361 10842 6427 10845
rect 10593 10842 10659 10845
rect 6361 10840 10659 10842
rect 6361 10784 6366 10840
rect 6422 10784 10598 10840
rect 10654 10784 10659 10840
rect 6361 10782 10659 10784
rect 6361 10779 6427 10782
rect 10593 10779 10659 10782
rect 12433 10842 12499 10845
rect 14641 10842 14707 10845
rect 12433 10840 14707 10842
rect 12433 10784 12438 10840
rect 12494 10784 14646 10840
rect 14702 10784 14707 10840
rect 12433 10782 14707 10784
rect 12433 10779 12499 10782
rect 14641 10779 14707 10782
rect 13905 10706 13971 10709
rect 2684 10646 2836 10706
rect 5398 10704 13971 10706
rect 5398 10648 13910 10704
rect 13966 10648 13971 10704
rect 5398 10646 13971 10648
rect 2776 10570 2836 10646
rect 13905 10643 13971 10646
rect 14365 10706 14431 10709
rect 16665 10706 16731 10709
rect 14365 10704 16731 10706
rect 14365 10648 14370 10704
rect 14426 10648 16670 10704
rect 16726 10648 16731 10704
rect 14365 10646 16731 10648
rect 14365 10643 14431 10646
rect 16665 10643 16731 10646
rect 6085 10570 6151 10573
rect 2776 10568 6151 10570
rect 2776 10512 6090 10568
rect 6146 10512 6151 10568
rect 2776 10510 6151 10512
rect 6085 10507 6151 10510
rect 8569 10570 8635 10573
rect 12157 10570 12223 10573
rect 8569 10568 12223 10570
rect 8569 10512 8574 10568
rect 8630 10512 12162 10568
rect 12218 10512 12223 10568
rect 8569 10510 12223 10512
rect 8569 10507 8635 10510
rect 12157 10507 12223 10510
rect 13077 10570 13143 10573
rect 17217 10570 17283 10573
rect 13077 10568 17283 10570
rect 13077 10512 13082 10568
rect 13138 10512 17222 10568
rect 17278 10512 17283 10568
rect 13077 10510 17283 10512
rect 13077 10507 13143 10510
rect 17217 10507 17283 10510
rect 3417 10434 3483 10437
rect 9990 10434 9996 10436
rect 3417 10432 9996 10434
rect 3417 10376 3422 10432
rect 3478 10376 9996 10432
rect 3417 10374 9996 10376
rect 3417 10371 3483 10374
rect 9990 10372 9996 10374
rect 10060 10372 10066 10436
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 9806 10236 9812 10300
rect 9876 10298 9882 10300
rect 10133 10298 10199 10301
rect 9876 10296 10199 10298
rect 9876 10240 10138 10296
rect 10194 10240 10199 10296
rect 9876 10238 10199 10240
rect 9876 10236 9882 10238
rect 10133 10235 10199 10238
rect 12893 10298 12959 10301
rect 18137 10298 18203 10301
rect 12893 10296 18203 10298
rect 12893 10240 12898 10296
rect 12954 10240 18142 10296
rect 18198 10240 18203 10296
rect 12893 10238 18203 10240
rect 12893 10235 12959 10238
rect 18137 10235 18203 10238
rect 0 10162 480 10192
rect 2865 10162 2931 10165
rect 14365 10162 14431 10165
rect 0 10102 1226 10162
rect 0 10072 480 10102
rect 1166 9890 1226 10102
rect 2865 10160 14431 10162
rect 2865 10104 2870 10160
rect 2926 10104 14370 10160
rect 14426 10104 14431 10160
rect 2865 10102 14431 10104
rect 2865 10099 2931 10102
rect 14365 10099 14431 10102
rect 14641 10162 14707 10165
rect 18597 10162 18663 10165
rect 14641 10160 18663 10162
rect 14641 10104 14646 10160
rect 14702 10104 18602 10160
rect 18658 10104 18663 10160
rect 14641 10102 18663 10104
rect 14641 10099 14707 10102
rect 18597 10099 18663 10102
rect 1393 10026 1459 10029
rect 14273 10026 14339 10029
rect 15469 10026 15535 10029
rect 1393 10024 14339 10026
rect 1393 9968 1398 10024
rect 1454 9968 14278 10024
rect 14334 9968 14339 10024
rect 1393 9966 14339 9968
rect 1393 9963 1459 9966
rect 14273 9963 14339 9966
rect 14782 10024 15535 10026
rect 14782 9968 15474 10024
rect 15530 9968 15535 10024
rect 14782 9966 15535 9968
rect 3969 9890 4035 9893
rect 1166 9888 4035 9890
rect 1166 9832 3974 9888
rect 4030 9832 4035 9888
rect 1166 9830 4035 9832
rect 3969 9827 4035 9830
rect 6085 9890 6151 9893
rect 14782 9890 14842 9966
rect 15469 9963 15535 9966
rect 6085 9888 14842 9890
rect 6085 9832 6090 9888
rect 6146 9832 14842 9888
rect 6085 9830 14842 9832
rect 16297 9890 16363 9893
rect 18781 9890 18847 9893
rect 16297 9888 18847 9890
rect 16297 9832 16302 9888
rect 16358 9832 18786 9888
rect 18842 9832 18847 9888
rect 16297 9830 18847 9832
rect 6085 9827 6151 9830
rect 16297 9827 16363 9830
rect 18781 9827 18847 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 8109 9754 8175 9757
rect 12525 9754 12591 9757
rect 8109 9752 12591 9754
rect 8109 9696 8114 9752
rect 8170 9696 12530 9752
rect 12586 9696 12591 9752
rect 8109 9694 12591 9696
rect 8109 9691 8175 9694
rect 12525 9691 12591 9694
rect 0 9618 480 9648
rect 1853 9618 1919 9621
rect 0 9616 1919 9618
rect 0 9560 1858 9616
rect 1914 9560 1919 9616
rect 0 9558 1919 9560
rect 0 9528 480 9558
rect 1853 9555 1919 9558
rect 3969 9618 4035 9621
rect 10593 9618 10659 9621
rect 3969 9616 10659 9618
rect 3969 9560 3974 9616
rect 4030 9560 10598 9616
rect 10654 9560 10659 9616
rect 3969 9558 10659 9560
rect 3969 9555 4035 9558
rect 10593 9555 10659 9558
rect 3785 9482 3851 9485
rect 4705 9482 4771 9485
rect 11053 9482 11119 9485
rect 3785 9480 11119 9482
rect 3785 9424 3790 9480
rect 3846 9424 4710 9480
rect 4766 9424 11058 9480
rect 11114 9424 11119 9480
rect 3785 9422 11119 9424
rect 3785 9419 3851 9422
rect 4705 9419 4771 9422
rect 11053 9419 11119 9422
rect 12433 9482 12499 9485
rect 13169 9482 13235 9485
rect 12433 9480 13235 9482
rect 12433 9424 12438 9480
rect 12494 9424 13174 9480
rect 13230 9424 13235 9480
rect 12433 9422 13235 9424
rect 12433 9419 12499 9422
rect 13169 9419 13235 9422
rect 7005 9346 7071 9349
rect 9029 9346 9095 9349
rect 7005 9344 9095 9346
rect 7005 9288 7010 9344
rect 7066 9288 9034 9344
rect 9090 9288 9095 9344
rect 7005 9286 9095 9288
rect 7005 9283 7071 9286
rect 9029 9283 9095 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 2497 9210 2563 9213
rect 2497 9208 4354 9210
rect 2497 9152 2502 9208
rect 2558 9152 4354 9208
rect 2497 9150 4354 9152
rect 2497 9147 2563 9150
rect 0 9074 480 9104
rect 4294 9074 4354 9150
rect 9806 9148 9812 9212
rect 9876 9210 9882 9212
rect 9949 9210 10015 9213
rect 9876 9208 10015 9210
rect 9876 9152 9954 9208
rect 10010 9152 10015 9208
rect 9876 9150 10015 9152
rect 9876 9148 9882 9150
rect 9949 9147 10015 9150
rect 4429 9074 4495 9077
rect 14917 9074 14983 9077
rect 0 9014 3986 9074
rect 4294 9072 14983 9074
rect 4294 9016 4434 9072
rect 4490 9016 14922 9072
rect 14978 9016 14983 9072
rect 4294 9014 14983 9016
rect 0 8984 480 9014
rect 0 8530 480 8560
rect 3785 8530 3851 8533
rect 0 8528 3851 8530
rect 0 8472 3790 8528
rect 3846 8472 3851 8528
rect 0 8470 3851 8472
rect 3926 8530 3986 9014
rect 4429 9011 4495 9014
rect 14917 9011 14983 9014
rect 4061 8938 4127 8941
rect 22369 8938 22435 8941
rect 4061 8936 22435 8938
rect 4061 8880 4066 8936
rect 4122 8880 22374 8936
rect 22430 8880 22435 8936
rect 4061 8878 22435 8880
rect 4061 8875 4127 8878
rect 22369 8875 22435 8878
rect 8017 8802 8083 8805
rect 9949 8802 10015 8805
rect 11053 8802 11119 8805
rect 14549 8802 14615 8805
rect 8017 8800 10196 8802
rect 8017 8744 8022 8800
rect 8078 8744 9954 8800
rect 10010 8744 10196 8800
rect 8017 8742 10196 8744
rect 8017 8739 8083 8742
rect 9949 8739 10015 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 10136 8666 10196 8742
rect 11053 8800 14615 8802
rect 11053 8744 11058 8800
rect 11114 8744 14554 8800
rect 14610 8744 14615 8800
rect 11053 8742 14615 8744
rect 11053 8739 11119 8742
rect 14549 8739 14615 8742
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 14181 8666 14247 8669
rect 10136 8664 14247 8666
rect 10136 8608 14186 8664
rect 14242 8608 14247 8664
rect 10136 8606 14247 8608
rect 14181 8603 14247 8606
rect 7189 8530 7255 8533
rect 20345 8530 20411 8533
rect 3926 8528 20411 8530
rect 3926 8472 7194 8528
rect 7250 8472 20350 8528
rect 20406 8472 20411 8528
rect 3926 8470 20411 8472
rect 0 8440 480 8470
rect 3785 8467 3851 8470
rect 7189 8467 7255 8470
rect 20345 8467 20411 8470
rect 1393 8394 1459 8397
rect 5533 8394 5599 8397
rect 12157 8394 12223 8397
rect 1393 8392 5599 8394
rect 1393 8336 1398 8392
rect 1454 8336 5538 8392
rect 5594 8336 5599 8392
rect 1393 8334 5599 8336
rect 1393 8331 1459 8334
rect 5533 8331 5599 8334
rect 9998 8392 12223 8394
rect 9998 8336 12162 8392
rect 12218 8336 12223 8392
rect 9998 8334 12223 8336
rect 3141 8258 3207 8261
rect 9998 8260 10058 8334
rect 12157 8331 12223 8334
rect 14273 8394 14339 8397
rect 17953 8394 18019 8397
rect 14273 8392 18019 8394
rect 14273 8336 14278 8392
rect 14334 8336 17958 8392
rect 18014 8336 18019 8392
rect 14273 8334 18019 8336
rect 14273 8331 14339 8334
rect 17953 8331 18019 8334
rect 9990 8258 9996 8260
rect 3141 8256 9996 8258
rect 3141 8200 3146 8256
rect 3202 8200 9996 8256
rect 3141 8198 9996 8200
rect 3141 8195 3207 8198
rect 9990 8196 9996 8198
rect 10060 8196 10066 8260
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 16389 8122 16455 8125
rect 18413 8122 18479 8125
rect 16389 8120 18479 8122
rect 16389 8064 16394 8120
rect 16450 8064 18418 8120
rect 18474 8064 18479 8120
rect 16389 8062 18479 8064
rect 16389 8059 16455 8062
rect 18413 8059 18479 8062
rect 17677 7986 17743 7989
rect 8526 7984 17743 7986
rect 8526 7928 17682 7984
rect 17738 7928 17743 7984
rect 8526 7926 17743 7928
rect 0 7850 480 7880
rect 8526 7853 8586 7926
rect 17677 7923 17743 7926
rect 8477 7850 8586 7853
rect 22737 7850 22803 7853
rect 0 7848 8586 7850
rect 0 7792 8482 7848
rect 8538 7792 8586 7848
rect 0 7790 8586 7792
rect 14460 7848 22803 7850
rect 14460 7792 22742 7848
rect 22798 7792 22803 7848
rect 14460 7790 22803 7792
rect 0 7760 480 7790
rect 8477 7787 8543 7790
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 8109 7578 8175 7581
rect 14460 7578 14520 7790
rect 22737 7787 22803 7790
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 8109 7576 14520 7578
rect 8109 7520 8114 7576
rect 8170 7520 14520 7576
rect 8109 7518 14520 7520
rect 8109 7515 8175 7518
rect 9305 7442 9371 7445
rect 15745 7442 15811 7445
rect 9305 7440 15811 7442
rect 9305 7384 9310 7440
rect 9366 7384 15750 7440
rect 15806 7384 15811 7440
rect 9305 7382 15811 7384
rect 9305 7379 9371 7382
rect 15745 7379 15811 7382
rect 0 7306 480 7336
rect 3417 7306 3483 7309
rect 0 7304 3483 7306
rect 0 7248 3422 7304
rect 3478 7248 3483 7304
rect 0 7246 3483 7248
rect 0 7216 480 7246
rect 3417 7243 3483 7246
rect 9305 7306 9371 7309
rect 15469 7306 15535 7309
rect 9305 7304 15535 7306
rect 9305 7248 9310 7304
rect 9366 7248 15474 7304
rect 15530 7248 15535 7304
rect 9305 7246 15535 7248
rect 9305 7243 9371 7246
rect 15469 7243 15535 7246
rect 18321 7306 18387 7309
rect 21357 7306 21423 7309
rect 18321 7304 21423 7306
rect 18321 7248 18326 7304
rect 18382 7248 21362 7304
rect 21418 7248 21423 7304
rect 18321 7246 21423 7248
rect 18321 7243 18387 7246
rect 21357 7243 21423 7246
rect 9213 7170 9279 7173
rect 9673 7170 9739 7173
rect 9213 7168 9739 7170
rect 9213 7112 9218 7168
rect 9274 7112 9678 7168
rect 9734 7112 9739 7168
rect 9213 7110 9739 7112
rect 9213 7107 9279 7110
rect 9673 7107 9739 7110
rect 10777 7170 10843 7173
rect 12157 7170 12223 7173
rect 10777 7168 12223 7170
rect 10777 7112 10782 7168
rect 10838 7112 12162 7168
rect 12218 7112 12223 7168
rect 10777 7110 12223 7112
rect 10777 7107 10843 7110
rect 12157 7107 12223 7110
rect 17718 7108 17724 7172
rect 17788 7170 17794 7172
rect 18781 7170 18847 7173
rect 17788 7168 18847 7170
rect 17788 7112 18786 7168
rect 18842 7112 18847 7168
rect 17788 7110 18847 7112
rect 17788 7108 17794 7110
rect 18781 7107 18847 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 4429 7034 4495 7037
rect 8569 7034 8635 7037
rect 4429 7032 8635 7034
rect 4429 6976 4434 7032
rect 4490 6976 8574 7032
rect 8630 6976 8635 7032
rect 4429 6974 8635 6976
rect 4429 6971 4495 6974
rect 8569 6971 8635 6974
rect 9581 7034 9647 7037
rect 14089 7034 14155 7037
rect 9581 7032 10196 7034
rect 9581 6976 9586 7032
rect 9642 6976 10196 7032
rect 9581 6974 10196 6976
rect 9581 6971 9647 6974
rect 4797 6898 4863 6901
rect 4294 6896 4863 6898
rect 4294 6840 4802 6896
rect 4858 6840 4863 6896
rect 4294 6838 4863 6840
rect 0 6762 480 6792
rect 4294 6762 4354 6838
rect 4797 6835 4863 6838
rect 6269 6898 6335 6901
rect 8477 6898 8543 6901
rect 6269 6896 8543 6898
rect 6269 6840 6274 6896
rect 6330 6840 8482 6896
rect 8538 6840 8543 6896
rect 6269 6838 8543 6840
rect 10136 6898 10196 6974
rect 10734 7032 14155 7034
rect 10734 6976 14094 7032
rect 14150 6976 14155 7032
rect 10734 6974 14155 6976
rect 10734 6898 10794 6974
rect 14089 6971 14155 6974
rect 14825 7034 14891 7037
rect 19333 7034 19399 7037
rect 14825 7032 19399 7034
rect 14825 6976 14830 7032
rect 14886 6976 19338 7032
rect 19394 6976 19399 7032
rect 14825 6974 19399 6976
rect 14825 6971 14891 6974
rect 19333 6971 19399 6974
rect 10136 6838 10794 6898
rect 12433 6898 12499 6901
rect 19977 6898 20043 6901
rect 12433 6896 20043 6898
rect 12433 6840 12438 6896
rect 12494 6840 19982 6896
rect 20038 6840 20043 6896
rect 12433 6838 20043 6840
rect 6269 6835 6335 6838
rect 8477 6835 8543 6838
rect 12433 6835 12499 6838
rect 19977 6835 20043 6838
rect 0 6702 4354 6762
rect 4521 6762 4587 6765
rect 8293 6762 8359 6765
rect 4521 6760 8359 6762
rect 4521 6704 4526 6760
rect 4582 6704 8298 6760
rect 8354 6704 8359 6760
rect 4521 6702 8359 6704
rect 0 6672 480 6702
rect 4521 6699 4587 6702
rect 8293 6699 8359 6702
rect 13077 6762 13143 6765
rect 18045 6762 18111 6765
rect 13077 6760 18111 6762
rect 13077 6704 13082 6760
rect 13138 6704 18050 6760
rect 18106 6704 18111 6760
rect 13077 6702 18111 6704
rect 13077 6699 13143 6702
rect 18045 6699 18111 6702
rect 10961 6626 11027 6629
rect 14641 6626 14707 6629
rect 10961 6624 14707 6626
rect 10961 6568 10966 6624
rect 11022 6568 14646 6624
rect 14702 6568 14707 6624
rect 10961 6566 14707 6568
rect 10961 6563 11027 6566
rect 14641 6563 14707 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 6678 6428 6684 6492
rect 6748 6490 6754 6492
rect 6821 6490 6887 6493
rect 6748 6488 6887 6490
rect 6748 6432 6826 6488
rect 6882 6432 6887 6488
rect 6748 6430 6887 6432
rect 6748 6428 6754 6430
rect 6821 6427 6887 6430
rect 16757 6490 16823 6493
rect 20253 6490 20319 6493
rect 16757 6488 20319 6490
rect 16757 6432 16762 6488
rect 16818 6432 20258 6488
rect 20314 6432 20319 6488
rect 16757 6430 20319 6432
rect 16757 6427 16823 6430
rect 20253 6427 20319 6430
rect 22134 6428 22140 6492
rect 22204 6490 22210 6492
rect 22277 6490 22343 6493
rect 22204 6488 22343 6490
rect 22204 6432 22282 6488
rect 22338 6432 22343 6488
rect 22204 6430 22343 6432
rect 22204 6428 22210 6430
rect 22277 6427 22343 6430
rect 3969 6354 4035 6357
rect 6913 6354 6979 6357
rect 3969 6352 6979 6354
rect 3969 6296 3974 6352
rect 4030 6296 6918 6352
rect 6974 6296 6979 6352
rect 3969 6294 6979 6296
rect 3969 6291 4035 6294
rect 6913 6291 6979 6294
rect 7281 6354 7347 6357
rect 10225 6354 10291 6357
rect 7281 6352 10291 6354
rect 7281 6296 7286 6352
rect 7342 6296 10230 6352
rect 10286 6296 10291 6352
rect 7281 6294 10291 6296
rect 7281 6291 7347 6294
rect 10225 6291 10291 6294
rect 4061 6218 4127 6221
rect 8293 6218 8359 6221
rect 4061 6216 8359 6218
rect 4061 6160 4066 6216
rect 4122 6160 8298 6216
rect 8354 6160 8359 6216
rect 4061 6158 8359 6160
rect 4061 6155 4127 6158
rect 8293 6155 8359 6158
rect 12525 6218 12591 6221
rect 18689 6218 18755 6221
rect 19333 6218 19399 6221
rect 12525 6216 19399 6218
rect 12525 6160 12530 6216
rect 12586 6160 18694 6216
rect 18750 6160 19338 6216
rect 19394 6160 19399 6216
rect 12525 6158 19399 6160
rect 12525 6155 12591 6158
rect 18689 6155 18755 6158
rect 19333 6155 19399 6158
rect 19517 6218 19583 6221
rect 22185 6218 22251 6221
rect 19517 6216 22251 6218
rect 19517 6160 19522 6216
rect 19578 6160 22190 6216
rect 22246 6160 22251 6216
rect 19517 6158 22251 6160
rect 19517 6155 19583 6158
rect 22185 6155 22251 6158
rect 0 6082 480 6112
rect 4889 6082 4955 6085
rect 9949 6082 10015 6085
rect 0 6080 4955 6082
rect 0 6024 4894 6080
rect 4950 6024 4955 6080
rect 0 6022 4955 6024
rect 0 5992 480 6022
rect 4889 6019 4955 6022
rect 7422 6080 10015 6082
rect 7422 6024 9954 6080
rect 10010 6024 10015 6080
rect 7422 6022 10015 6024
rect 3325 5946 3391 5949
rect 7422 5946 7482 6022
rect 9949 6019 10015 6022
rect 11513 6082 11579 6085
rect 14181 6082 14247 6085
rect 11513 6080 14247 6082
rect 11513 6024 11518 6080
rect 11574 6024 14186 6080
rect 14242 6024 14247 6080
rect 11513 6022 14247 6024
rect 11513 6019 11579 6022
rect 14181 6019 14247 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 3325 5944 7482 5946
rect 3325 5888 3330 5944
rect 3386 5888 7482 5944
rect 3325 5886 7482 5888
rect 7649 5946 7715 5949
rect 7925 5946 7991 5949
rect 9857 5946 9923 5949
rect 7649 5944 9923 5946
rect 7649 5888 7654 5944
rect 7710 5888 7930 5944
rect 7986 5888 9862 5944
rect 9918 5888 9923 5944
rect 7649 5886 9923 5888
rect 3325 5883 3391 5886
rect 7649 5883 7715 5886
rect 7925 5883 7991 5886
rect 9857 5883 9923 5886
rect 12433 5946 12499 5949
rect 12433 5944 17234 5946
rect 12433 5888 12438 5944
rect 12494 5888 17234 5944
rect 12433 5886 17234 5888
rect 12433 5883 12499 5886
rect 8569 5810 8635 5813
rect 13445 5810 13511 5813
rect 8569 5808 13511 5810
rect 8569 5752 8574 5808
rect 8630 5752 13450 5808
rect 13506 5752 13511 5808
rect 8569 5750 13511 5752
rect 8569 5747 8635 5750
rect 13445 5747 13511 5750
rect 13629 5810 13695 5813
rect 16665 5810 16731 5813
rect 13629 5808 16731 5810
rect 13629 5752 13634 5808
rect 13690 5752 16670 5808
rect 16726 5752 16731 5808
rect 13629 5750 16731 5752
rect 17174 5810 17234 5886
rect 22277 5810 22343 5813
rect 17174 5808 22343 5810
rect 17174 5752 22282 5808
rect 22338 5752 22343 5808
rect 17174 5750 22343 5752
rect 13629 5747 13695 5750
rect 16665 5747 16731 5750
rect 22277 5747 22343 5750
rect 4061 5674 4127 5677
rect 8937 5674 9003 5677
rect 4061 5672 9003 5674
rect 4061 5616 4066 5672
rect 4122 5616 8942 5672
rect 8998 5616 9003 5672
rect 4061 5614 9003 5616
rect 4061 5611 4127 5614
rect 8937 5611 9003 5614
rect 9397 5674 9463 5677
rect 11881 5674 11947 5677
rect 9397 5672 11947 5674
rect 9397 5616 9402 5672
rect 9458 5616 11886 5672
rect 11942 5616 11947 5672
rect 9397 5614 11947 5616
rect 9397 5611 9463 5614
rect 11881 5611 11947 5614
rect 12893 5674 12959 5677
rect 17953 5674 18019 5677
rect 12893 5672 18019 5674
rect 12893 5616 12898 5672
rect 12954 5616 17958 5672
rect 18014 5616 18019 5672
rect 12893 5614 18019 5616
rect 12893 5611 12959 5614
rect 17953 5611 18019 5614
rect 0 5538 480 5568
rect 2221 5538 2287 5541
rect 0 5536 2287 5538
rect 0 5480 2226 5536
rect 2282 5480 2287 5536
rect 0 5478 2287 5480
rect 0 5448 480 5478
rect 2221 5475 2287 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 8017 5402 8083 5405
rect 13721 5402 13787 5405
rect 20989 5402 21055 5405
rect 8017 5400 13787 5402
rect 8017 5344 8022 5400
rect 8078 5344 13726 5400
rect 13782 5344 13787 5400
rect 8017 5342 13787 5344
rect 8017 5339 8083 5342
rect 13721 5339 13787 5342
rect 16806 5400 21055 5402
rect 16806 5344 20994 5400
rect 21050 5344 21055 5400
rect 16806 5342 21055 5344
rect 1853 5266 1919 5269
rect 11237 5266 11303 5269
rect 1853 5264 11303 5266
rect 1853 5208 1858 5264
rect 1914 5208 11242 5264
rect 11298 5208 11303 5264
rect 1853 5206 11303 5208
rect 1853 5203 1919 5206
rect 11237 5203 11303 5206
rect 13629 5266 13695 5269
rect 16806 5266 16866 5342
rect 20989 5339 21055 5342
rect 13629 5264 16866 5266
rect 13629 5208 13634 5264
rect 13690 5208 16866 5264
rect 13629 5206 16866 5208
rect 16941 5266 17007 5269
rect 23565 5266 23631 5269
rect 16941 5264 23631 5266
rect 16941 5208 16946 5264
rect 17002 5208 23570 5264
rect 23626 5208 23631 5264
rect 16941 5206 23631 5208
rect 13629 5203 13695 5206
rect 16941 5203 17007 5206
rect 23565 5203 23631 5206
rect 3049 5130 3115 5133
rect 6269 5130 6335 5133
rect 3049 5128 6335 5130
rect 3049 5072 3054 5128
rect 3110 5072 6274 5128
rect 6330 5072 6335 5128
rect 3049 5070 6335 5072
rect 3049 5067 3115 5070
rect 6269 5067 6335 5070
rect 7557 5130 7623 5133
rect 11605 5130 11671 5133
rect 7557 5128 11671 5130
rect 7557 5072 7562 5128
rect 7618 5072 11610 5128
rect 11666 5072 11671 5128
rect 7557 5070 11671 5072
rect 7557 5067 7623 5070
rect 11605 5067 11671 5070
rect 13721 5130 13787 5133
rect 15285 5130 15351 5133
rect 15469 5132 15535 5133
rect 15469 5130 15516 5132
rect 13721 5128 15351 5130
rect 13721 5072 13726 5128
rect 13782 5072 15290 5128
rect 15346 5072 15351 5128
rect 13721 5070 15351 5072
rect 15424 5128 15516 5130
rect 15424 5072 15474 5128
rect 15424 5070 15516 5072
rect 13721 5067 13787 5070
rect 15285 5067 15351 5070
rect 15469 5068 15516 5070
rect 15580 5068 15586 5132
rect 15469 5067 15535 5068
rect 0 4994 480 5024
rect 1761 4994 1827 4997
rect 3969 4994 4035 4997
rect 0 4992 4035 4994
rect 0 4936 1766 4992
rect 1822 4936 3974 4992
rect 4030 4936 4035 4992
rect 0 4934 4035 4936
rect 0 4904 480 4934
rect 1761 4931 1827 4934
rect 3969 4931 4035 4934
rect 5165 4994 5231 4997
rect 8937 4994 9003 4997
rect 5165 4992 9003 4994
rect 5165 4936 5170 4992
rect 5226 4936 8942 4992
rect 8998 4936 9003 4992
rect 5165 4934 9003 4936
rect 5165 4931 5231 4934
rect 8937 4931 9003 4934
rect 11237 4994 11303 4997
rect 13077 4994 13143 4997
rect 19425 4994 19491 4997
rect 11237 4992 19491 4994
rect 11237 4936 11242 4992
rect 11298 4936 13082 4992
rect 13138 4936 19430 4992
rect 19486 4936 19491 4992
rect 11237 4934 19491 4936
rect 11237 4931 11303 4934
rect 13077 4931 13143 4934
rect 19425 4931 19491 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 3693 4858 3759 4861
rect 9806 4858 9812 4860
rect 3693 4856 9812 4858
rect 3693 4800 3698 4856
rect 3754 4800 9812 4856
rect 3693 4798 9812 4800
rect 3693 4795 3759 4798
rect 9806 4796 9812 4798
rect 9876 4796 9882 4860
rect 10685 4858 10751 4861
rect 19425 4858 19491 4861
rect 10685 4856 19491 4858
rect 10685 4800 10690 4856
rect 10746 4800 19430 4856
rect 19486 4800 19491 4856
rect 10685 4798 19491 4800
rect 10685 4795 10751 4798
rect 19425 4795 19491 4798
rect 2865 4722 2931 4725
rect 10777 4722 10843 4725
rect 2865 4720 10843 4722
rect 2865 4664 2870 4720
rect 2926 4664 10782 4720
rect 10838 4664 10843 4720
rect 2865 4662 10843 4664
rect 2865 4659 2931 4662
rect 10777 4659 10843 4662
rect 10961 4722 11027 4725
rect 14089 4722 14155 4725
rect 10961 4720 14155 4722
rect 10961 4664 10966 4720
rect 11022 4664 14094 4720
rect 14150 4664 14155 4720
rect 10961 4662 14155 4664
rect 10961 4659 11027 4662
rect 14089 4659 14155 4662
rect 18229 4722 18295 4725
rect 20897 4722 20963 4725
rect 27520 4722 28000 4752
rect 18229 4720 20963 4722
rect 18229 4664 18234 4720
rect 18290 4664 20902 4720
rect 20958 4664 20963 4720
rect 18229 4662 20963 4664
rect 18229 4659 18295 4662
rect 20897 4659 20963 4662
rect 21038 4662 28000 4722
rect 2681 4586 2747 4589
rect 5257 4586 5323 4589
rect 11237 4586 11303 4589
rect 2681 4584 5323 4586
rect 2681 4528 2686 4584
rect 2742 4528 5262 4584
rect 5318 4528 5323 4584
rect 2681 4526 5323 4528
rect 2681 4523 2747 4526
rect 5257 4523 5323 4526
rect 5398 4584 11303 4586
rect 5398 4528 11242 4584
rect 11298 4528 11303 4584
rect 5398 4526 11303 4528
rect 0 4450 480 4480
rect 3785 4450 3851 4453
rect 0 4448 3851 4450
rect 0 4392 3790 4448
rect 3846 4392 3851 4448
rect 0 4390 3851 4392
rect 0 4360 480 4390
rect 3785 4387 3851 4390
rect 289 4178 355 4181
rect 3417 4178 3483 4181
rect 5398 4178 5458 4526
rect 11237 4523 11303 4526
rect 11421 4586 11487 4589
rect 16757 4586 16823 4589
rect 11421 4584 16823 4586
rect 11421 4528 11426 4584
rect 11482 4528 16762 4584
rect 16818 4528 16823 4584
rect 11421 4526 16823 4528
rect 11421 4523 11487 4526
rect 16757 4523 16823 4526
rect 18413 4586 18479 4589
rect 21038 4586 21098 4662
rect 27520 4632 28000 4662
rect 18413 4584 21098 4586
rect 18413 4528 18418 4584
rect 18474 4528 21098 4584
rect 18413 4526 21098 4528
rect 18413 4523 18479 4526
rect 7925 4450 7991 4453
rect 12801 4450 12867 4453
rect 7925 4448 12867 4450
rect 7925 4392 7930 4448
rect 7986 4392 12806 4448
rect 12862 4392 12867 4448
rect 7925 4390 12867 4392
rect 7925 4387 7991 4390
rect 12801 4387 12867 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 289 4176 5458 4178
rect 289 4120 294 4176
rect 350 4120 3422 4176
rect 3478 4120 5458 4176
rect 289 4118 5458 4120
rect 5533 4178 5599 4181
rect 6177 4178 6243 4181
rect 10961 4178 11027 4181
rect 5533 4176 11027 4178
rect 5533 4120 5538 4176
rect 5594 4120 6182 4176
rect 6238 4120 10966 4176
rect 11022 4120 11027 4176
rect 5533 4118 11027 4120
rect 289 4115 355 4118
rect 3417 4115 3483 4118
rect 5533 4115 5599 4118
rect 6177 4115 6243 4118
rect 10961 4115 11027 4118
rect 14273 4178 14339 4181
rect 17953 4178 18019 4181
rect 20713 4178 20779 4181
rect 14273 4176 18019 4178
rect 14273 4120 14278 4176
rect 14334 4120 17958 4176
rect 18014 4120 18019 4176
rect 14273 4118 18019 4120
rect 14273 4115 14339 4118
rect 17953 4115 18019 4118
rect 19566 4176 20779 4178
rect 19566 4120 20718 4176
rect 20774 4120 20779 4176
rect 19566 4118 20779 4120
rect 7097 4042 7163 4045
rect 9489 4042 9555 4045
rect 7097 4040 9555 4042
rect 7097 3984 7102 4040
rect 7158 3984 9494 4040
rect 9550 3984 9555 4040
rect 7097 3982 9555 3984
rect 7097 3979 7163 3982
rect 9489 3979 9555 3982
rect 10133 4042 10199 4045
rect 15009 4042 15075 4045
rect 10133 4040 15075 4042
rect 10133 3984 10138 4040
rect 10194 3984 15014 4040
rect 15070 3984 15075 4040
rect 10133 3982 15075 3984
rect 10133 3979 10199 3982
rect 15009 3979 15075 3982
rect 16389 4042 16455 4045
rect 19566 4042 19626 4118
rect 20713 4115 20779 4118
rect 16389 4040 19626 4042
rect 16389 3984 16394 4040
rect 16450 3984 19626 4040
rect 16389 3982 19626 3984
rect 19793 4042 19859 4045
rect 21357 4042 21423 4045
rect 19793 4040 21423 4042
rect 19793 3984 19798 4040
rect 19854 3984 21362 4040
rect 21418 3984 21423 4040
rect 19793 3982 21423 3984
rect 16389 3979 16455 3982
rect 19793 3979 19859 3982
rect 21357 3979 21423 3982
rect 26366 3980 26372 4044
rect 26436 4042 26442 4044
rect 26509 4042 26575 4045
rect 26436 4040 26575 4042
rect 26436 3984 26514 4040
rect 26570 3984 26575 4040
rect 26436 3982 26575 3984
rect 26436 3980 26442 3982
rect 26509 3979 26575 3982
rect 3325 3906 3391 3909
rect 1350 3904 3391 3906
rect 1350 3848 3330 3904
rect 3386 3848 3391 3904
rect 1350 3846 3391 3848
rect 0 3770 480 3800
rect 1350 3770 1410 3846
rect 3325 3843 3391 3846
rect 3693 3906 3759 3909
rect 5993 3906 6059 3909
rect 7281 3906 7347 3909
rect 3693 3904 7347 3906
rect 3693 3848 3698 3904
rect 3754 3848 5998 3904
rect 6054 3848 7286 3904
rect 7342 3848 7347 3904
rect 3693 3846 7347 3848
rect 3693 3843 3759 3846
rect 5993 3843 6059 3846
rect 7281 3843 7347 3846
rect 11237 3906 11303 3909
rect 13813 3906 13879 3909
rect 17769 3906 17835 3909
rect 19241 3906 19307 3909
rect 11237 3904 13370 3906
rect 11237 3848 11242 3904
rect 11298 3848 13370 3904
rect 11237 3846 13370 3848
rect 11237 3843 11303 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 1669 3772 1735 3773
rect 1669 3770 1716 3772
rect 0 3710 1410 3770
rect 1624 3768 1716 3770
rect 1624 3712 1674 3768
rect 1624 3710 1716 3712
rect 0 3680 480 3710
rect 1669 3708 1716 3710
rect 1780 3708 1786 3772
rect 9213 3770 9279 3773
rect 5030 3768 9279 3770
rect 5030 3712 9218 3768
rect 9274 3712 9279 3768
rect 5030 3710 9279 3712
rect 1669 3707 1735 3708
rect 2497 3634 2563 3637
rect 4521 3634 4587 3637
rect 5030 3634 5090 3710
rect 9213 3707 9279 3710
rect 10685 3770 10751 3773
rect 12433 3770 12499 3773
rect 10685 3768 12499 3770
rect 10685 3712 10690 3768
rect 10746 3712 12438 3768
rect 12494 3712 12499 3768
rect 10685 3710 12499 3712
rect 13310 3770 13370 3846
rect 13813 3904 17835 3906
rect 13813 3848 13818 3904
rect 13874 3848 17774 3904
rect 17830 3848 17835 3904
rect 13813 3846 17835 3848
rect 13813 3843 13879 3846
rect 17769 3843 17835 3846
rect 18692 3904 19307 3906
rect 18692 3848 19246 3904
rect 19302 3848 19307 3904
rect 18692 3846 19307 3848
rect 14365 3770 14431 3773
rect 13310 3768 14431 3770
rect 13310 3712 14370 3768
rect 14426 3712 14431 3768
rect 13310 3710 14431 3712
rect 10685 3707 10751 3710
rect 12433 3707 12499 3710
rect 14365 3707 14431 3710
rect 14774 3708 14780 3772
rect 14844 3770 14850 3772
rect 18692 3770 18752 3846
rect 19241 3843 19307 3846
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 14844 3710 18752 3770
rect 14844 3708 14850 3710
rect 18822 3708 18828 3772
rect 18892 3770 18898 3772
rect 18965 3770 19031 3773
rect 18892 3768 19031 3770
rect 18892 3712 18970 3768
rect 19026 3712 19031 3768
rect 18892 3710 19031 3712
rect 18892 3708 18898 3710
rect 18965 3707 19031 3710
rect 20161 3770 20227 3773
rect 22277 3770 22343 3773
rect 20161 3768 22343 3770
rect 20161 3712 20166 3768
rect 20222 3712 22282 3768
rect 22338 3712 22343 3768
rect 20161 3710 22343 3712
rect 20161 3707 20227 3710
rect 22277 3707 22343 3710
rect 2497 3632 5090 3634
rect 2497 3576 2502 3632
rect 2558 3576 4526 3632
rect 4582 3576 5090 3632
rect 2497 3574 5090 3576
rect 5165 3634 5231 3637
rect 7649 3634 7715 3637
rect 5165 3632 7715 3634
rect 5165 3576 5170 3632
rect 5226 3576 7654 3632
rect 7710 3576 7715 3632
rect 5165 3574 7715 3576
rect 2497 3571 2563 3574
rect 4521 3571 4587 3574
rect 5165 3571 5231 3574
rect 7649 3571 7715 3574
rect 7925 3634 7991 3637
rect 12341 3634 12407 3637
rect 14641 3634 14707 3637
rect 7925 3632 11898 3634
rect 7925 3576 7930 3632
rect 7986 3576 11898 3632
rect 7925 3574 11898 3576
rect 7925 3571 7991 3574
rect 2865 3498 2931 3501
rect 9397 3498 9463 3501
rect 9857 3498 9923 3501
rect 11605 3498 11671 3501
rect 2865 3496 6194 3498
rect 2865 3440 2870 3496
rect 2926 3440 6194 3496
rect 2865 3438 6194 3440
rect 2865 3435 2931 3438
rect 841 3362 907 3365
rect 4429 3362 4495 3365
rect 841 3360 5458 3362
rect 841 3304 846 3360
rect 902 3304 4434 3360
rect 4490 3304 5458 3360
rect 841 3302 5458 3304
rect 841 3299 907 3302
rect 4429 3299 4495 3302
rect 0 3226 480 3256
rect 2681 3226 2747 3229
rect 5165 3226 5231 3229
rect 0 3166 2514 3226
rect 0 3136 480 3166
rect 2454 3090 2514 3166
rect 2681 3224 5231 3226
rect 2681 3168 2686 3224
rect 2742 3168 5170 3224
rect 5226 3168 5231 3224
rect 2681 3166 5231 3168
rect 2681 3163 2747 3166
rect 5165 3163 5231 3166
rect 3417 3090 3483 3093
rect 2454 3088 3483 3090
rect 2454 3032 3422 3088
rect 3478 3032 3483 3088
rect 2454 3030 3483 3032
rect 5398 3090 5458 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 6134 3226 6194 3438
rect 9397 3496 11671 3498
rect 9397 3440 9402 3496
rect 9458 3440 9862 3496
rect 9918 3440 11610 3496
rect 11666 3440 11671 3496
rect 9397 3438 11671 3440
rect 11838 3498 11898 3574
rect 12341 3632 14707 3634
rect 12341 3576 12346 3632
rect 12402 3576 14646 3632
rect 14702 3576 14707 3632
rect 12341 3574 14707 3576
rect 12341 3571 12407 3574
rect 14641 3571 14707 3574
rect 16481 3634 16547 3637
rect 21633 3634 21699 3637
rect 16481 3632 21699 3634
rect 16481 3576 16486 3632
rect 16542 3576 21638 3632
rect 21694 3576 21699 3632
rect 16481 3574 21699 3576
rect 16481 3571 16547 3574
rect 21633 3571 21699 3574
rect 19057 3498 19123 3501
rect 27613 3498 27679 3501
rect 11838 3496 19123 3498
rect 11838 3440 19062 3496
rect 19118 3440 19123 3496
rect 11838 3438 19123 3440
rect 9397 3435 9463 3438
rect 9857 3435 9923 3438
rect 11605 3435 11671 3438
rect 19057 3435 19123 3438
rect 23982 3496 27679 3498
rect 23982 3440 27618 3496
rect 27674 3440 27679 3496
rect 23982 3438 27679 3440
rect 11053 3362 11119 3365
rect 12157 3362 12223 3365
rect 11053 3360 12223 3362
rect 11053 3304 11058 3360
rect 11114 3304 12162 3360
rect 12218 3304 12223 3360
rect 11053 3302 12223 3304
rect 11053 3299 11119 3302
rect 12157 3299 12223 3302
rect 18045 3362 18111 3365
rect 22185 3362 22251 3365
rect 18045 3360 22251 3362
rect 18045 3304 18050 3360
rect 18106 3304 22190 3360
rect 22246 3304 22251 3360
rect 18045 3302 22251 3304
rect 18045 3299 18111 3302
rect 22185 3299 22251 3302
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 13905 3226 13971 3229
rect 14774 3226 14780 3228
rect 6134 3224 13971 3226
rect 6134 3168 13910 3224
rect 13966 3168 13971 3224
rect 6134 3166 13971 3168
rect 13905 3163 13971 3166
rect 14414 3166 14780 3226
rect 7741 3090 7807 3093
rect 5398 3088 7807 3090
rect 5398 3032 7746 3088
rect 7802 3032 7807 3088
rect 5398 3030 7807 3032
rect 3417 3027 3483 3030
rect 7741 3027 7807 3030
rect 8017 3090 8083 3093
rect 9673 3090 9739 3093
rect 8017 3088 9739 3090
rect 8017 3032 8022 3088
rect 8078 3032 9678 3088
rect 9734 3032 9739 3088
rect 8017 3030 9739 3032
rect 8017 3027 8083 3030
rect 9673 3027 9739 3030
rect 10133 3090 10199 3093
rect 14414 3090 14474 3166
rect 14774 3164 14780 3166
rect 14844 3164 14850 3228
rect 18505 3226 18571 3229
rect 23841 3226 23907 3229
rect 18505 3224 23907 3226
rect 18505 3168 18510 3224
rect 18566 3168 23846 3224
rect 23902 3168 23907 3224
rect 18505 3166 23907 3168
rect 18505 3163 18571 3166
rect 23841 3163 23907 3166
rect 10133 3088 14474 3090
rect 10133 3032 10138 3088
rect 10194 3032 14474 3088
rect 10133 3030 14474 3032
rect 15193 3090 15259 3093
rect 19425 3090 19491 3093
rect 23982 3090 24042 3438
rect 27613 3435 27679 3438
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 15193 3088 19491 3090
rect 15193 3032 15198 3088
rect 15254 3032 19430 3088
rect 19486 3032 19491 3088
rect 15193 3030 19491 3032
rect 10133 3027 10199 3030
rect 15193 3027 15259 3030
rect 19425 3027 19491 3030
rect 19566 3030 24042 3090
rect 2865 2954 2931 2957
rect 7373 2954 7439 2957
rect 17401 2954 17467 2957
rect 2865 2952 17467 2954
rect 2865 2896 2870 2952
rect 2926 2896 7378 2952
rect 7434 2896 17406 2952
rect 17462 2896 17467 2952
rect 2865 2894 17467 2896
rect 2865 2891 2931 2894
rect 7373 2891 7439 2894
rect 17401 2891 17467 2894
rect 17677 2954 17743 2957
rect 19566 2954 19626 3030
rect 17677 2952 19626 2954
rect 17677 2896 17682 2952
rect 17738 2896 19626 2952
rect 17677 2894 19626 2896
rect 21817 2954 21883 2957
rect 23657 2954 23723 2957
rect 21817 2952 23723 2954
rect 21817 2896 21822 2952
rect 21878 2896 23662 2952
rect 23718 2896 23723 2952
rect 21817 2894 23723 2896
rect 17677 2891 17743 2894
rect 21817 2891 21883 2894
rect 23657 2891 23723 2894
rect 9121 2818 9187 2821
rect 4846 2816 9187 2818
rect 4846 2760 9126 2816
rect 9182 2760 9187 2816
rect 4846 2758 9187 2760
rect 0 2682 480 2712
rect 4846 2682 4906 2758
rect 9121 2755 9187 2758
rect 10961 2818 11027 2821
rect 11237 2818 11303 2821
rect 10961 2816 11303 2818
rect 10961 2760 10966 2816
rect 11022 2760 11242 2816
rect 11298 2760 11303 2816
rect 10961 2758 11303 2760
rect 10961 2755 11027 2758
rect 11237 2755 11303 2758
rect 11421 2818 11487 2821
rect 17401 2818 17467 2821
rect 11421 2816 17467 2818
rect 11421 2760 11426 2816
rect 11482 2760 17406 2816
rect 17462 2760 17467 2816
rect 11421 2758 17467 2760
rect 11421 2755 11487 2758
rect 17401 2755 17467 2758
rect 21265 2818 21331 2821
rect 23105 2818 23171 2821
rect 21265 2816 23171 2818
rect 21265 2760 21270 2816
rect 21326 2760 23110 2816
rect 23166 2760 23171 2816
rect 21265 2758 23171 2760
rect 21265 2755 21331 2758
rect 23105 2755 23171 2758
rect 23473 2818 23539 2821
rect 25313 2818 25379 2821
rect 23473 2816 25379 2818
rect 23473 2760 23478 2816
rect 23534 2760 25318 2816
rect 25374 2760 25379 2816
rect 23473 2758 25379 2760
rect 23473 2755 23539 2758
rect 25313 2755 25379 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 0 2622 4906 2682
rect 5257 2682 5323 2685
rect 6913 2682 6979 2685
rect 5257 2680 6979 2682
rect 5257 2624 5262 2680
rect 5318 2624 6918 2680
rect 6974 2624 6979 2680
rect 5257 2622 6979 2624
rect 0 2592 480 2622
rect 5257 2619 5323 2622
rect 6913 2619 6979 2622
rect 11145 2682 11211 2685
rect 18689 2682 18755 2685
rect 11145 2680 18890 2682
rect 11145 2624 11150 2680
rect 11206 2624 18694 2680
rect 18750 2624 18890 2680
rect 11145 2622 18890 2624
rect 11145 2619 11211 2622
rect 18689 2619 18755 2622
rect 2957 2546 3023 2549
rect 8385 2546 8451 2549
rect 2957 2544 8451 2546
rect 2957 2488 2962 2544
rect 3018 2488 8390 2544
rect 8446 2488 8451 2544
rect 2957 2486 8451 2488
rect 2957 2483 3023 2486
rect 8385 2483 8451 2486
rect 8569 2546 8635 2549
rect 14733 2546 14799 2549
rect 17125 2546 17191 2549
rect 8569 2544 14799 2546
rect 8569 2488 8574 2544
rect 8630 2488 14738 2544
rect 14794 2488 14799 2544
rect 8569 2486 14799 2488
rect 8569 2483 8635 2486
rect 14733 2483 14799 2486
rect 14966 2544 17191 2546
rect 14966 2488 17130 2544
rect 17186 2488 17191 2544
rect 14966 2486 17191 2488
rect 18830 2546 18890 2622
rect 23473 2546 23539 2549
rect 18830 2544 23539 2546
rect 18830 2488 23478 2544
rect 23534 2488 23539 2544
rect 18830 2486 23539 2488
rect 4981 2412 5047 2413
rect 4981 2410 5028 2412
rect 4936 2408 5028 2410
rect 4936 2352 4986 2408
rect 4936 2350 5028 2352
rect 4981 2348 5028 2350
rect 5092 2348 5098 2412
rect 6269 2410 6335 2413
rect 11973 2410 12039 2413
rect 6269 2408 12039 2410
rect 6269 2352 6274 2408
rect 6330 2352 11978 2408
rect 12034 2352 12039 2408
rect 6269 2350 12039 2352
rect 4981 2347 5047 2348
rect 6269 2347 6335 2350
rect 11973 2347 12039 2350
rect 12157 2410 12223 2413
rect 13169 2410 13235 2413
rect 12157 2408 13235 2410
rect 12157 2352 12162 2408
rect 12218 2352 13174 2408
rect 13230 2352 13235 2408
rect 12157 2350 13235 2352
rect 12157 2347 12223 2350
rect 13169 2347 13235 2350
rect 13537 2410 13603 2413
rect 14966 2410 15026 2486
rect 17125 2483 17191 2486
rect 23473 2483 23539 2486
rect 13537 2408 15026 2410
rect 13537 2352 13542 2408
rect 13598 2352 15026 2408
rect 13537 2350 15026 2352
rect 19149 2410 19215 2413
rect 21541 2410 21607 2413
rect 24025 2412 24091 2413
rect 19149 2408 21607 2410
rect 19149 2352 19154 2408
rect 19210 2352 21546 2408
rect 21602 2352 21607 2408
rect 19149 2350 21607 2352
rect 13537 2347 13603 2350
rect 19149 2347 19215 2350
rect 21541 2347 21607 2350
rect 23974 2348 23980 2412
rect 24044 2410 24091 2412
rect 24044 2408 24136 2410
rect 24086 2352 24136 2408
rect 24044 2350 24136 2352
rect 24044 2348 24091 2350
rect 24025 2347 24091 2348
rect 9990 2212 9996 2276
rect 10060 2274 10066 2276
rect 10501 2274 10567 2277
rect 10060 2272 10567 2274
rect 10060 2216 10506 2272
rect 10562 2216 10567 2272
rect 10060 2214 10567 2216
rect 10060 2212 10066 2214
rect 10501 2211 10567 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 6453 2138 6519 2141
rect 8477 2138 8543 2141
rect 13813 2138 13879 2141
rect 6453 2136 8402 2138
rect 6453 2080 6458 2136
rect 6514 2080 8402 2136
rect 6453 2078 8402 2080
rect 6453 2075 6519 2078
rect 0 2002 480 2032
rect 8109 2002 8175 2005
rect 0 2000 8175 2002
rect 0 1944 8114 2000
rect 8170 1944 8175 2000
rect 0 1942 8175 1944
rect 8342 2002 8402 2078
rect 8477 2136 13879 2138
rect 8477 2080 8482 2136
rect 8538 2080 13818 2136
rect 13874 2080 13879 2136
rect 8477 2078 13879 2080
rect 8477 2075 8543 2078
rect 13813 2075 13879 2078
rect 16849 2138 16915 2141
rect 19517 2138 19583 2141
rect 16849 2136 19583 2138
rect 16849 2080 16854 2136
rect 16910 2080 19522 2136
rect 19578 2080 19583 2136
rect 16849 2078 19583 2080
rect 16849 2075 16915 2078
rect 19517 2075 19583 2078
rect 12157 2002 12223 2005
rect 8342 2000 12223 2002
rect 8342 1944 12162 2000
rect 12218 1944 12223 2000
rect 8342 1942 12223 1944
rect 0 1912 480 1942
rect 8109 1939 8175 1942
rect 12157 1939 12223 1942
rect 13721 2002 13787 2005
rect 16941 2002 17007 2005
rect 13721 2000 17007 2002
rect 13721 1944 13726 2000
rect 13782 1944 16946 2000
rect 17002 1944 17007 2000
rect 13721 1942 17007 1944
rect 13721 1939 13787 1942
rect 16941 1939 17007 1942
rect 18873 2002 18939 2005
rect 21633 2002 21699 2005
rect 18873 2000 21699 2002
rect 18873 1944 18878 2000
rect 18934 1944 21638 2000
rect 21694 1944 21699 2000
rect 18873 1942 21699 1944
rect 18873 1939 18939 1942
rect 21633 1939 21699 1942
rect 1393 1866 1459 1869
rect 16849 1866 16915 1869
rect 1393 1864 16915 1866
rect 1393 1808 1398 1864
rect 1454 1808 16854 1864
rect 16910 1808 16915 1864
rect 1393 1806 16915 1808
rect 1393 1803 1459 1806
rect 16849 1803 16915 1806
rect 17125 1866 17191 1869
rect 20897 1866 20963 1869
rect 17125 1864 20963 1866
rect 17125 1808 17130 1864
rect 17186 1808 20902 1864
rect 20958 1808 20963 1864
rect 17125 1806 20963 1808
rect 17125 1803 17191 1806
rect 20897 1803 20963 1806
rect 10685 1730 10751 1733
rect 21173 1730 21239 1733
rect 10685 1728 21239 1730
rect 10685 1672 10690 1728
rect 10746 1672 21178 1728
rect 21234 1672 21239 1728
rect 10685 1670 21239 1672
rect 10685 1667 10751 1670
rect 21173 1667 21239 1670
rect 2313 1594 2379 1597
rect 18873 1594 18939 1597
rect 2313 1592 18939 1594
rect 2313 1536 2318 1592
rect 2374 1536 18878 1592
rect 18934 1536 18939 1592
rect 2313 1534 18939 1536
rect 2313 1531 2379 1534
rect 18873 1531 18939 1534
rect 19057 1594 19123 1597
rect 24209 1594 24275 1597
rect 19057 1592 24275 1594
rect 19057 1536 19062 1592
rect 19118 1536 24214 1592
rect 24270 1536 24275 1592
rect 19057 1534 24275 1536
rect 19057 1531 19123 1534
rect 24209 1531 24275 1534
rect 0 1458 480 1488
rect 1577 1458 1643 1461
rect 0 1456 1643 1458
rect 0 1400 1582 1456
rect 1638 1400 1643 1456
rect 0 1398 1643 1400
rect 0 1368 480 1398
rect 1577 1395 1643 1398
rect 5441 1458 5507 1461
rect 17125 1458 17191 1461
rect 5441 1456 17191 1458
rect 5441 1400 5446 1456
rect 5502 1400 17130 1456
rect 17186 1400 17191 1456
rect 5441 1398 17191 1400
rect 5441 1395 5507 1398
rect 17125 1395 17191 1398
rect 17309 1458 17375 1461
rect 19609 1458 19675 1461
rect 17309 1456 19675 1458
rect 17309 1400 17314 1456
rect 17370 1400 19614 1456
rect 19670 1400 19675 1456
rect 17309 1398 19675 1400
rect 17309 1395 17375 1398
rect 19609 1395 19675 1398
rect 20069 1458 20135 1461
rect 25957 1458 26023 1461
rect 20069 1456 26023 1458
rect 20069 1400 20074 1456
rect 20130 1400 25962 1456
rect 26018 1400 26023 1456
rect 20069 1398 26023 1400
rect 20069 1395 20135 1398
rect 25957 1395 26023 1398
rect 10869 1322 10935 1325
rect 15285 1322 15351 1325
rect 10869 1320 15351 1322
rect 10869 1264 10874 1320
rect 10930 1264 15290 1320
rect 15346 1264 15351 1320
rect 10869 1262 15351 1264
rect 10869 1259 10935 1262
rect 15285 1259 15351 1262
rect 15469 1322 15535 1325
rect 21081 1322 21147 1325
rect 15469 1320 21147 1322
rect 15469 1264 15474 1320
rect 15530 1264 21086 1320
rect 21142 1264 21147 1320
rect 15469 1262 21147 1264
rect 15469 1259 15535 1262
rect 21081 1259 21147 1262
rect 9806 1124 9812 1188
rect 9876 1186 9882 1188
rect 21449 1186 21515 1189
rect 9876 1184 21515 1186
rect 9876 1128 21454 1184
rect 21510 1128 21515 1184
rect 9876 1126 21515 1128
rect 9876 1124 9882 1126
rect 21449 1123 21515 1126
rect 3417 1050 3483 1053
rect 18781 1050 18847 1053
rect 3417 1048 18847 1050
rect 3417 992 3422 1048
rect 3478 992 18786 1048
rect 18842 992 18847 1048
rect 3417 990 18847 992
rect 3417 987 3483 990
rect 18781 987 18847 990
rect 0 914 480 944
rect 1669 914 1735 917
rect 0 912 1735 914
rect 0 856 1674 912
rect 1730 856 1735 912
rect 0 854 1735 856
rect 0 824 480 854
rect 1669 851 1735 854
rect 14457 914 14523 917
rect 27061 914 27127 917
rect 14457 912 27127 914
rect 14457 856 14462 912
rect 14518 856 27066 912
rect 27122 856 27127 912
rect 14457 854 27127 856
rect 14457 851 14523 854
rect 27061 851 27127 854
rect 0 370 480 400
rect 6361 370 6427 373
rect 0 368 6427 370
rect 0 312 6366 368
rect 6422 312 6427 368
rect 0 310 6427 312
rect 0 280 480 310
rect 6361 307 6427 310
rect 11605 98 11671 101
rect 24669 98 24735 101
rect 11605 96 24735 98
rect 11605 40 11610 96
rect 11666 40 24674 96
rect 24730 40 24735 96
rect 11605 38 24735 40
rect 11605 35 11671 38
rect 24669 35 24735 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 9812 18668 9876 18732
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 8156 11868 8220 11932
rect 18276 11868 18340 11932
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 17724 11188 17788 11252
rect 9996 10916 10060 10980
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 9996 10372 10060 10436
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 9812 10236 9876 10300
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 9812 9148 9876 9212
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 9996 8196 10060 8260
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 17724 7108 17788 7172
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 6684 6428 6748 6492
rect 22140 6428 22204 6492
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 15516 5128 15580 5132
rect 15516 5072 15530 5128
rect 15530 5072 15580 5128
rect 15516 5068 15580 5072
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 9812 4796 9876 4860
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 26372 3980 26436 4044
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 1716 3768 1780 3772
rect 1716 3712 1730 3768
rect 1730 3712 1780 3768
rect 1716 3708 1780 3712
rect 14780 3708 14844 3772
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 18828 3708 18892 3772
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 14780 3164 14844 3228
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5028 2408 5092 2412
rect 5028 2352 5042 2408
rect 5042 2352 5092 2408
rect 5028 2348 5092 2352
rect 23980 2408 24044 2412
rect 23980 2352 24030 2408
rect 24030 2352 24044 2408
rect 23980 2348 24044 2352
rect 9996 2212 10060 2276
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 9812 1124 9876 1188
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 9811 18732 9877 18733
rect 9811 18668 9812 18732
rect 9876 18668 9877 18732
rect 9811 18667 9877 18668
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 9814 10301 9874 18667
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 9995 10980 10061 10981
rect 9995 10916 9996 10980
rect 10060 10916 10061 10980
rect 9995 10915 10061 10916
rect 9998 10437 10058 10915
rect 9995 10436 10061 10437
rect 9995 10372 9996 10436
rect 10060 10372 10061 10436
rect 9995 10371 10061 10372
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 9811 10300 9877 10301
rect 9811 10236 9812 10300
rect 9876 10236 9877 10300
rect 9811 10235 9877 10236
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 9811 9212 9877 9213
rect 9811 9148 9812 9212
rect 9876 9148 9877 9212
rect 9811 9147 9877 9148
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 9814 4861 9874 9147
rect 9995 8260 10061 8261
rect 9995 8196 9996 8260
rect 10060 8196 10061 8260
rect 9995 8195 10061 8196
rect 9811 4860 9877 4861
rect 9811 4796 9812 4860
rect 9876 4796 9877 4860
rect 9811 4795 9877 4796
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 9814 1189 9874 4795
rect 9998 2277 10058 8195
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 17723 11252 17789 11253
rect 17723 11188 17724 11252
rect 17788 11188 17789 11252
rect 17723 11187 17789 11188
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 17726 7173 17786 11187
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 17723 7172 17789 7173
rect 17723 7108 17724 7172
rect 17788 7108 17789 7172
rect 17723 7107 17789 7108
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14779 3772 14845 3773
rect 14779 3708 14780 3772
rect 14844 3708 14845 3772
rect 14779 3707 14845 3708
rect 14782 3229 14842 3707
rect 14944 3296 15264 4320
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14779 3228 14845 3229
rect 14779 3164 14780 3228
rect 14844 3164 14845 3228
rect 14779 3163 14845 3164
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 9995 2276 10061 2277
rect 9995 2212 9996 2276
rect 10060 2212 10061 2276
rect 9995 2211 10061 2212
rect 10277 2128 10597 2688
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 26374 4045 26434 4982
rect 26371 4044 26437 4045
rect 26371 3980 26372 4044
rect 26436 3980 26437 4044
rect 26371 3979 26437 3980
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 9811 1188 9877 1189
rect 9811 1124 9812 1188
rect 9876 1124 9877 1188
rect 9811 1123 9877 1124
<< via4 >>
rect 8070 11932 8306 12018
rect 8070 11868 8156 11932
rect 8156 11868 8220 11932
rect 8220 11868 8306 11932
rect 8070 11782 8306 11868
rect 6598 6492 6834 6578
rect 6598 6428 6684 6492
rect 6684 6428 6748 6492
rect 6748 6428 6834 6492
rect 6598 6342 6834 6428
rect 1630 3772 1866 3858
rect 1630 3708 1716 3772
rect 1716 3708 1780 3772
rect 1780 3708 1866 3772
rect 1630 3622 1866 3708
rect 4942 2412 5178 2498
rect 4942 2348 5028 2412
rect 5028 2348 5092 2412
rect 5092 2348 5178 2412
rect 4942 2262 5178 2348
rect 18190 11932 18426 12018
rect 18190 11868 18276 11932
rect 18276 11868 18340 11932
rect 18340 11868 18426 11932
rect 18190 11782 18426 11868
rect 22054 6492 22290 6578
rect 22054 6428 22140 6492
rect 22140 6428 22204 6492
rect 22204 6428 22290 6492
rect 22054 6342 22290 6428
rect 15430 5132 15666 5218
rect 15430 5068 15516 5132
rect 15516 5068 15580 5132
rect 15580 5068 15666 5132
rect 15430 4982 15666 5068
rect 18742 3772 18978 3858
rect 18742 3708 18828 3772
rect 18828 3708 18892 3772
rect 18892 3708 18978 3772
rect 18742 3622 18978 3708
rect 26286 4982 26522 5218
rect 23894 2412 24130 2498
rect 23894 2348 23980 2412
rect 23980 2348 24044 2412
rect 24044 2348 24130 2412
rect 23894 2262 24130 2348
<< metal5 >>
rect 8028 12018 18468 12060
rect 8028 11782 8070 12018
rect 8306 11782 18190 12018
rect 18426 11782 18468 12018
rect 8028 11740 18468 11782
rect 6556 6578 22332 6620
rect 6556 6342 6598 6578
rect 6834 6342 22054 6578
rect 22290 6342 22332 6578
rect 6556 6300 22332 6342
rect 15388 5218 26564 5260
rect 15388 4982 15430 5218
rect 15666 4982 26286 5218
rect 26522 4982 26564 5218
rect 15388 4940 26564 4982
rect 1588 3858 19020 3900
rect 1588 3622 1630 3858
rect 1866 3622 18742 3858
rect 18978 3622 19020 3858
rect 1588 3580 19020 3622
rect 4900 2498 24172 2540
rect 4900 2262 4942 2498
rect 5178 2262 23894 2498
rect 24130 2262 24172 2498
rect 4900 2220 24172 2262
use sky130_fd_sc_hd__fill_2  FILLER_1_8 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1840 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6
timestamp 1604666999
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604666999
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604666999
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10
timestamp 1604666999
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 2024 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_29
timestamp 1604666999
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1604666999
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604666999
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_37
timestamp 1604666999
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_33
timestamp 1604666999
transform 1 0 4140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 4048 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604666999
transform 1 0 4876 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 5888 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51
timestamp 1604666999
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_50
timestamp 1604666999
transform 1 0 5704 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_54 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 6072 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 6348 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55
timestamp 1604666999
transform 1 0 6164 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59
timestamp 1604666999
transform 1 0 6532 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_58 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 6440 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_62
timestamp 1604666999
transform 1 0 6808 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67
timestamp 1604666999
transform 1 0 7268 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63
timestamp 1604666999
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 7084 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604666999
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604666999
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_4_
timestamp 1604666999
transform 1 0 6900 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_1_77
timestamp 1604666999
transform 1 0 8188 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_72
timestamp 1604666999
transform 1 0 7728 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1604666999
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__A1
timestamp 1604666999
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_5_
timestamp 1604666999
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 8464 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604666999
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604666999
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__A0
timestamp 1604666999
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_5__S
timestamp 1604666999
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604666999
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604666999
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_99
timestamp 1604666999
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_103
timestamp 1604666999
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1604666999
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_107
timestamp 1604666999
transform 1 0 10948 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_107
timestamp 1604666999
transform 1 0 10948 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 10764 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604666999
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604666999
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604666999
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604666999
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604666999
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_123
timestamp 1604666999
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604666999
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604666999
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604666999
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1604666999
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_0_138
timestamp 1604666999
transform 1 0 13800 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1604666999
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 12604 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_148
timestamp 1604666999
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_144
timestamp 1604666999
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1604666999
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604666999
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604666999
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604666999
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604666999
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1604666999
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 15088 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1604666999
transform 1 0 16284 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 16560 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_171
timestamp 1604666999
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_170
timestamp 1604666999
transform 1 0 16744 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_175
timestamp 1604666999
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1604666999
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604666999
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_179
timestamp 1604666999
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1604666999
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604666999
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604666999
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604666999
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604666999
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604666999
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1604666999
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_193
timestamp 1604666999
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_196
timestamp 1604666999
transform 1 0 19136 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_208
timestamp 1604666999
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_203
timestamp 1604666999
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_200
timestamp 1604666999
transform 1 0 19504 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1604666999
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604666999
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604666999
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_212
timestamp 1604666999
transform 1 0 20608 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_210
timestamp 1604666999
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604666999
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_214
timestamp 1604666999
transform 1 0 20792 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_218
timestamp 1604666999
transform 1 0 21160 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1604666999
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_227
timestamp 1604666999
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_222
timestamp 1604666999
transform 1 0 21528 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_227
timestamp 1604666999
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604666999
transform 1 0 21344 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604666999
transform 1 0 21620 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_235 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 22724 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_231
timestamp 1604666999
transform 1 0 22356 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_231
timestamp 1604666999
transform 1 0 22356 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 22540 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604666999
transform 1 0 22540 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604666999
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604666999
transform 1 0 22724 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1604666999
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_247
timestamp 1604666999
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_243
timestamp 1604666999
transform 1 0 23460 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_239
timestamp 1604666999
transform 1 0 23092 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 23644 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604666999
transform 1 0 23276 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604666999
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604666999
transform 1 0 23644 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_249
timestamp 1604666999
transform 1 0 24012 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1604666999
transform 1 0 24380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604666999
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604666999
transform 1 0 24564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604666999
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604666999
transform 1 0 24012 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_253 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 24380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_257
timestamp 1604666999
transform 1 0 24748 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604666999
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604666999
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_269
timestamp 1604666999
transform 1 0 25852 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_265
timestamp 1604666999
transform 1 0 25484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1604666999
transform 1 0 1656 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604666999
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 2668 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1604666999
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_15
timestamp 1604666999
transform 1 0 2484 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_19
timestamp 1604666999
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604666999
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 4416 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 3036 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1604666999
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1604666999
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1604666999
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_38
timestamp 1604666999
transform 1 0 4600 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 5520 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 4784 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_42
timestamp 1604666999
transform 1 0 4968 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_46
timestamp 1604666999
transform 1 0 5336 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1604666999
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_67
timestamp 1604666999
transform 1 0 7268 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_72
timestamp 1604666999
transform 1 0 7728 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604666999
transform 1 0 10120 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604666999
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9844 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1604666999
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_88
timestamp 1604666999
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1604666999
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_97
timestamp 1604666999
transform 1 0 10028 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 11684 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 11500 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604666999
transform 1 0 11132 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_107
timestamp 1604666999
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_111
timestamp 1604666999
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_134
timestamp 1604666999
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1604666999
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604666999
transform 1 0 14168 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604666999
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604666999
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604666999
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604666999
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_145
timestamp 1604666999
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1604666999
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_158
timestamp 1604666999
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 16652 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_162
timestamp 1604666999
transform 1 0 16008 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_166
timestamp 1604666999
transform 1 0 16376 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1604666999
transform 1 0 19136 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1604666999
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_192
timestamp 1604666999
transform 1 0 18768 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604666999
transform 1 0 21068 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604666999
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 20516 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_205
timestamp 1604666999
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_209
timestamp 1604666999
transform 1 0 20332 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1604666999
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_215
timestamp 1604666999
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604666999
transform 1 0 22172 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 21620 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1604666999
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_225
timestamp 1604666999
transform 1 0 21804 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1604666999
transform 1 0 22540 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_245
timestamp 1604666999
transform 1 0 23644 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_257
timestamp 1604666999
transform 1 0 24748 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604666999
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604666999
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_269 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 25852 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604666999
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604666999
transform 1 0 2300 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604666999
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 1656 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1604666999
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_8
timestamp 1604666999
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_12
timestamp 1604666999
transform 1 0 2208 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 3864 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 3312 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_22
timestamp 1604666999
transform 1 0 3128 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_26
timestamp 1604666999
transform 1 0 3496 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_49
timestamp 1604666999
transform 1 0 5612 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_55
timestamp 1604666999
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604666999
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1604666999
transform 1 0 7820 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604666999
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1604666999
transform 1 0 6808 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_68
timestamp 1604666999
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_72
timestamp 1604666999
transform 1 0 7728 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1604666999
transform 1 0 9384 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 8832 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_82
timestamp 1604666999
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_86
timestamp 1604666999
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_99
timestamp 1604666999
transform 1 0 10212 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604666999
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__A1
timestamp 1604666999
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__A0
timestamp 1604666999
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__S
timestamp 1604666999
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_105
timestamp 1604666999
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_109
timestamp 1604666999
transform 1 0 11132 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1604666999
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604666999
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604666999
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604666999
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1604666999
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_136
timestamp 1604666999
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1604666999
transform 1 0 13984 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604666999
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_149
timestamp 1604666999
transform 1 0 14812 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_153
timestamp 1604666999
transform 1 0 15180 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_156
timestamp 1604666999
transform 1 0 15456 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1604666999
transform 1 0 16100 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 15916 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_160
timestamp 1604666999
transform 1 0 15824 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_172
timestamp 1604666999
transform 1 0 16928 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_176
timestamp 1604666999
transform 1 0 17296 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604666999
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604666999
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1604666999
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1604666999
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_197
timestamp 1604666999
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604666999
transform 1 0 21160 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604666999
transform 1 0 19596 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604666999
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_210
timestamp 1604666999
transform 1 0 20424 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_214
timestamp 1604666999
transform 1 0 20792 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_217
timestamp 1604666999
transform 1 0 21068 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 22264 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604666999
transform 1 0 21712 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 22080 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1604666999
transform 1 0 21528 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_226
timestamp 1604666999
transform 1 0 21896 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_233
timestamp 1604666999
transform 1 0 22540 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_237
timestamp 1604666999
transform 1 0 22908 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604666999
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_243
timestamp 1604666999
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604666999
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604666999
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604666999
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_269
timestamp 1604666999
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604666999
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 1564 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1604666999
transform 1 0 1380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_7
timestamp 1604666999
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_11
timestamp 1604666999
transform 1 0 2116 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604666999
transform 1 0 4416 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604666999
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1604666999
transform 1 0 3220 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1604666999
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1604666999
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1604666999
transform 1 0 5980 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_45
timestamp 1604666999
transform 1 0 5244 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_49
timestamp 1604666999
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1604666999
transform 1 0 7544 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_62
timestamp 1604666999
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp 1604666999
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_79
timestamp 1604666999
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_83
timestamp 1604666999
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_87
timestamp 1604666999
transform 1 0 9108 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 8924 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9292 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_93
timestamp 1604666999
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1604666999
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604666999
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 9936 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_99
timestamp 1604666999
transform 1 0 10212 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_6_
timestamp 1604666999
transform 1 0 10948 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 11960 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 10396 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_103
timestamp 1604666999
transform 1 0 10580 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_116
timestamp 1604666999
transform 1 0 11776 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1604666999
transform 1 0 12512 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 13524 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_120
timestamp 1604666999
transform 1 0 12144 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_133
timestamp 1604666999
transform 1 0 13340 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_137
timestamp 1604666999
transform 1 0 13708 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604666999
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604666999
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604666999
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13892 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_145
timestamp 1604666999
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_149
timestamp 1604666999
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_158
timestamp 1604666999
transform 1 0 15640 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604666999
transform 1 0 16468 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 17480 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_162
timestamp 1604666999
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_165
timestamp 1604666999
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_176
timestamp 1604666999
transform 1 0 17296 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604666999
transform 1 0 18032 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_180
timestamp 1604666999
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_193
timestamp 1604666999
transform 1 0 18860 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1604666999
transform 1 0 19228 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604666999
transform 1 0 19596 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604666999
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604666999
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 20516 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 20148 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 19412 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_205
timestamp 1604666999
transform 1 0 19964 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_209
timestamp 1604666999
transform 1 0 20332 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1604666999
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 21436 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 21804 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_219
timestamp 1604666999
transform 1 0 21252 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_223
timestamp 1604666999
transform 1 0 21620 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1604666999
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1604666999
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1604666999
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604666999
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604666999
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1604666999
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604666999
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1604666999
transform 1 0 1380 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604666999
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_12
timestamp 1604666999
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_16
timestamp 1604666999
transform 1 0 2576 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 3588 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 3404 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_20
timestamp 1604666999
transform 1 0 2944 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_23
timestamp 1604666999
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_36
timestamp 1604666999
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_40
timestamp 1604666999
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1604666999
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1604666999
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 6808 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604666999
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9292 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_81
timestamp 1604666999
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_85
timestamp 1604666999
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_108
timestamp 1604666999
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_112
timestamp 1604666999
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_116
timestamp 1604666999
transform 1 0 11776 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 13524 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 12512 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604666999
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12972 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_123
timestamp 1604666999
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_127
timestamp 1604666999
transform 1 0 12788 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_131
timestamp 1604666999
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_154
timestamp 1604666999
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_158
timestamp 1604666999
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_162
timestamp 1604666999
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1604666999
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 18032 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604666999
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1604666999
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1604666999
transform 1 0 20516 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 20332 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604666999
transform 1 0 19964 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_203
timestamp 1604666999
transform 1 0 19780 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_207
timestamp 1604666999
transform 1 0 20148 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 22080 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 21528 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 21896 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 22540 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_220
timestamp 1604666999
transform 1 0 21344 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_224
timestamp 1604666999
transform 1 0 21712 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_231
timestamp 1604666999
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_235
timestamp 1604666999
transform 1 0 22724 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604666999
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604666999
transform 1 0 23276 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_243
timestamp 1604666999
transform 1 0 23460 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604666999
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604666999
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604666999
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_269
timestamp 1604666999
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 1380 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 2208 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604666999
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604666999
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1604666999
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_7
timestamp 1604666999
transform 1 0 1748 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1604666999
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_26
timestamp 1604666999
transform 1 0 3496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_22
timestamp 1604666999
transform 1 0 3128 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_35
timestamp 1604666999
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_31
timestamp 1604666999
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604666999
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604666999
transform 1 0 4692 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 4048 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_7_48
timestamp 1604666999
transform 1 0 5520 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 5980 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_51
timestamp 1604666999
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_52
timestamp 1604666999
transform 1 0 5888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 6348 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_55
timestamp 1604666999
transform 1 0 6164 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_55
timestamp 1604666999
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604666999
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1604666999
transform 1 0 6532 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_68
timestamp 1604666999
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604666999
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1604666999
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 7544 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_72
timestamp 1604666999
transform 1 0 7728 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1604666999
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 7912 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_75
timestamp 1604666999
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_76
timestamp 1604666999
transform 1 0 8096 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 8280 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_79
timestamp 1604666999
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604666999
transform 1 0 8556 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_80
timestamp 1604666999
transform 1 0 8464 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_84
timestamp 1604666999
transform 1 0 8832 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_83
timestamp 1604666999
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9292 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_88
timestamp 1604666999
transform 1 0 9200 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_87
timestamp 1604666999
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1604666999
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604666999
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9476 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 9660 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 11592 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11960 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_112
timestamp 1604666999
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_116
timestamp 1604666999
transform 1 0 11776 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1604666999
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_114
timestamp 1604666999
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1604666999
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12144 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604666999
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_132
timestamp 1604666999
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_136
timestamp 1604666999
transform 1 0 13616 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_140
timestamp 1604666999
transform 1 0 13984 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_145
timestamp 1604666999
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_139
timestamp 1604666999
transform 1 0 13892 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 14076 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_149
timestamp 1604666999
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604666999
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1604666999
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 14260 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_168
timestamp 1604666999
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_162
timestamp 1604666999
transform 1 0 16008 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_167
timestamp 1604666999
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_163
timestamp 1604666999
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_173
timestamp 1604666999
transform 1 0 17020 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 16652 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 16744 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 16836 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604666999
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604666999
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1604666999
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_197
timestamp 1604666999
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1604666999
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_195
timestamp 1604666999
transform 1 0 19044 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_190
timestamp 1604666999
transform 1 0 18584 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604666999
transform 1 0 19320 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_206
timestamp 1604666999
transform 1 0 20056 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_202
timestamp 1604666999
transform 1 0 19688 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 19872 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_3_
timestamp 1604666999
transform 1 0 19596 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 20608 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 20516 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_210
timestamp 1604666999
transform 1 0 20424 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1604666999
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_210
timestamp 1604666999
transform 1 0 20424 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604666999
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 20976 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_214
timestamp 1604666999
transform 1 0 20792 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604666999
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1604666999
transform 1 0 21160 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 22264 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_224
timestamp 1604666999
transform 1 0 21712 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_236
timestamp 1604666999
transform 1 0 22816 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_227
timestamp 1604666999
transform 1 0 21988 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1604666999
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604666999
transform 1 0 23276 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604666999
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_240
timestamp 1604666999
transform 1 0 23184 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_245
timestamp 1604666999
transform 1 0 23644 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_257
timestamp 1604666999
transform 1 0 24748 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604666999
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604666999
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604666999
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604666999
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604666999
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_269
timestamp 1604666999
transform 1 0 25852 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604666999
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1604666999
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604666999
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604666999
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_6
timestamp 1604666999
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_10
timestamp 1604666999
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604666999
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604666999
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1604666999
transform 1 0 3220 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1604666999
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 5980 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp 1604666999
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_46
timestamp 1604666999
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_50
timestamp 1604666999
transform 1 0 5704 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_72
timestamp 1604666999
transform 1 0 7728 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_77
timestamp 1604666999
transform 1 0 8188 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_83
timestamp 1604666999
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604666999
transform 1 0 8464 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_87
timestamp 1604666999
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9292 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1604666999
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1604666999
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604666999
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_97
timestamp 1604666999
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 10212 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1604666999
transform 1 0 11040 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 10764 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 12052 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_101
timestamp 1604666999
transform 1 0 10396 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_107
timestamp 1604666999
transform 1 0 10948 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_117
timestamp 1604666999
transform 1 0 11868 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1604666999
transform 1 0 12604 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_121
timestamp 1604666999
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_134
timestamp 1604666999
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1604666999
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 14168 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1604666999
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_149
timestamp 1604666999
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604666999
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_158
timestamp 1604666999
transform 1 0 15640 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_154
timestamp 1604666999
transform 1 0 15272 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604666999
transform 1 0 15364 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 16376 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_162
timestamp 1604666999
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_165
timestamp 1604666999
transform 1 0 16284 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1604666999
transform 1 0 18860 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 18308 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_185
timestamp 1604666999
transform 1 0 18124 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_189
timestamp 1604666999
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604666999
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 19872 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 21160 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_202
timestamp 1604666999
transform 1 0 19688 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_206
timestamp 1604666999
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_210
timestamp 1604666999
transform 1 0 20424 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_215
timestamp 1604666999
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 22264 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 21528 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_220
timestamp 1604666999
transform 1 0 21344 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_224
timestamp 1604666999
transform 1 0 21712 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1604666999
transform 1 0 22540 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_245
timestamp 1604666999
transform 1 0 23644 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_257
timestamp 1604666999
transform 1 0 24748 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604666999
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604666999
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_269
timestamp 1604666999
transform 1 0 25852 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604666999
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1604666999
transform 1 0 1380 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604666999
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_12
timestamp 1604666999
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_16
timestamp 1604666999
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604666999
transform 1 0 3588 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_20
timestamp 1604666999
transform 1 0 2944 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_24
timestamp 1604666999
transform 1 0 3312 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1604666999
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1604666999
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1604666999
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_53
timestamp 1604666999
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1604666999
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 6808 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604666999
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604666999
transform 1 0 9292 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_81
timestamp 1604666999
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_85
timestamp 1604666999
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_92
timestamp 1604666999
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_96
timestamp 1604666999
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1604666999
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_100
timestamp 1604666999
transform 1 0 10304 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604666999
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604666999
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604666999
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604666999
transform 1 0 13616 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604666999
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_126
timestamp 1604666999
transform 1 0 12696 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1604666999
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_145
timestamp 1604666999
transform 1 0 14444 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_151
timestamp 1604666999
transform 1 0 14996 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_155
timestamp 1604666999
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1604666999
transform 1 0 15732 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_168
timestamp 1604666999
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_172
timestamp 1604666999
transform 1 0 16928 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_178
timestamp 1604666999
transform 1 0 17480 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604666999
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604666999
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 17664 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1604666999
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_193
timestamp 1604666999
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_197
timestamp 1604666999
transform 1 0 19228 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1604666999
transform 1 0 19596 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_210
timestamp 1604666999
transform 1 0 20424 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_222
timestamp 1604666999
transform 1 0 21528 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_234
timestamp 1604666999
transform 1 0 22632 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604666999
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_242
timestamp 1604666999
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604666999
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604666999
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604666999
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_269
timestamp 1604666999
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1604666999
transform 1 0 1380 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604666999
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 2668 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_12
timestamp 1604666999
transform 1 0 2208 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_16
timestamp 1604666999
transform 1 0 2576 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_19
timestamp 1604666999
transform 1 0 2852 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604666999
transform 1 0 4324 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604666999
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 3036 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1604666999
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1604666999
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_32
timestamp 1604666999
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1604666999
transform 1 0 5888 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 5336 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_44
timestamp 1604666999
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_48
timestamp 1604666999
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1604666999
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 6900 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_61
timestamp 1604666999
transform 1 0 6716 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_65
timestamp 1604666999
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_69
timestamp 1604666999
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_73
timestamp 1604666999
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1604666999
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604666999
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1604666999
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_88
timestamp 1604666999
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1604666999
transform 1 0 11684 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 11500 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_102
timestamp 1604666999
transform 1 0 10488 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_107
timestamp 1604666999
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_111
timestamp 1604666999
transform 1 0 11316 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13248 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_124
timestamp 1604666999
transform 1 0 12512 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_128
timestamp 1604666999
transform 1 0 12880 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_131
timestamp 1604666999
transform 1 0 13156 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604666999
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1604666999
transform 1 0 14076 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_145
timestamp 1604666999
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_149
timestamp 1604666999
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1604666999
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_158
timestamp 1604666999
transform 1 0 15640 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1604666999
transform 1 0 16100 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 17480 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 17112 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_161
timestamp 1604666999
transform 1 0 15916 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_172
timestamp 1604666999
transform 1 0 16928 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_176
timestamp 1604666999
transform 1 0 17296 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1604666999
transform 1 0 17664 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_189
timestamp 1604666999
transform 1 0 18492 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604666999
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_203
timestamp 1604666999
transform 1 0 19780 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_207
timestamp 1604666999
transform 1 0 20148 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1604666999
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604666999
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604666999
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1604666999
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1604666999
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604666999
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604666999
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1604666999
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604666999
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604666999
transform 1 0 1656 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1604666999
transform 1 0 2668 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604666999
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1604666999
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_9
timestamp 1604666999
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_13
timestamp 1604666999
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4232 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_26
timestamp 1604666999
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_30
timestamp 1604666999
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1604666999
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604666999
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1604666999
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604666999
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_71
timestamp 1604666999
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_75
timestamp 1604666999
transform 1 0 8004 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_79
timestamp 1604666999
transform 1 0 8372 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 8648 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604666999
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1604666999
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_105
timestamp 1604666999
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_109
timestamp 1604666999
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_114
timestamp 1604666999
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1604666999
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 12972 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604666999
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 12788 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_123
timestamp 1604666999
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 15180 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_148
timestamp 1604666999
transform 1 0 14720 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_152
timestamp 1604666999
transform 1 0 15088 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_155
timestamp 1604666999
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1604666999
transform 1 0 15732 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 17480 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_168
timestamp 1604666999
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1604666999
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_176
timestamp 1604666999
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604666999
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_180
timestamp 1604666999
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604666999
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1604666999
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1604666999
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1604666999
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1604666999
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604666999
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1604666999
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1604666999
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604666999
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1604666999
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 1472 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604666999
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1604666999
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1604666999
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604666999
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1604666999
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1604666999
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 6348 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 5796 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1604666999
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_45
timestamp 1604666999
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_49
timestamp 1604666999
transform 1 0 5612 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_53
timestamp 1604666999
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 8280 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_76
timestamp 1604666999
transform 1 0 8096 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1604666999
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604666999
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_80
timestamp 1604666999
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1604666999
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_88
timestamp 1604666999
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 11776 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 11592 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_102
timestamp 1604666999
transform 1 0 10488 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_107
timestamp 1604666999
transform 1 0 10948 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_112
timestamp 1604666999
transform 1 0 11408 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_135
timestamp 1604666999
transform 1 0 13524 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_140
timestamp 1604666999
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_144
timestamp 1604666999
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_148
timestamp 1604666999
transform 1 0 14720 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 14904 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_154
timestamp 1604666999
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1604666999
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604666999
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604666999
transform 1 0 15548 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 16560 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 16008 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_160
timestamp 1604666999
transform 1 0 15824 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_164
timestamp 1604666999
transform 1 0 16192 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_187
timestamp 1604666999
transform 1 0 18308 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604666999
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_199
timestamp 1604666999
transform 1 0 19412 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_211
timestamp 1604666999
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604666999
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604666999
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1604666999
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1604666999
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604666999
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604666999
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1604666999
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604666999
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604666999
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604666999
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_3_
timestamp 1604666999
transform 1 0 1380 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1604666999
transform 1 0 1380 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_16
timestamp 1604666999
transform 1 0 2576 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_12
timestamp 1604666999
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_16
timestamp 1604666999
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_12
timestamp 1604666999
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1604666999
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1604666999
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_20
timestamp 1604666999
transform 1 0 2944 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_20
timestamp 1604666999
transform 1 0 2944 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_36
timestamp 1604666999
transform 1 0 4416 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1604666999
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604666999
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 3036 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 4784 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_40
timestamp 1604666999
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_44
timestamp 1604666999
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_42
timestamp 1604666999
transform 1 0 4968 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604666999
transform 1 0 5520 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_46
timestamp 1604666999
transform 1 0 5336 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1604666999
transform 1 0 5428 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_56
timestamp 1604666999
transform 1 0 6256 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_55
timestamp 1604666999
transform 1 0 6164 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_51
timestamp 1604666999
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 6440 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_68
timestamp 1604666999
transform 1 0 7360 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_64
timestamp 1604666999
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_60
timestamp 1604666999
transform 1 0 6624 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604666999
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1604666999
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_72
timestamp 1604666999
transform 1 0 7728 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_77
timestamp 1604666999
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_71
timestamp 1604666999
transform 1 0 7636 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604666999
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1604666999
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_84
timestamp 1604666999
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_81
timestamp 1604666999
transform 1 0 8556 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604666999
transform 1 0 8648 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_95
timestamp 1604666999
transform 1 0 9844 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_91
timestamp 1604666999
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604666999
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 9660 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1604666999
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_3_
timestamp 1604666999
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_116
timestamp 1604666999
transform 1 0 11776 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_112
timestamp 1604666999
transform 1 0 11408 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1604666999
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_114
timestamp 1604666999
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 11960 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11592 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_125
timestamp 1604666999
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_120
timestamp 1604666999
transform 1 0 12144 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_123
timestamp 1604666999
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 12788 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604666999
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1604666999
transform 1 0 12788 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1604666999
transform 1 0 13616 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_134
timestamp 1604666999
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_129
timestamp 1604666999
transform 1 0 12972 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13800 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_14_142
timestamp 1604666999
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_146
timestamp 1604666999
transform 1 0 14536 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 14720 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_150
timestamp 1604666999
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604666999
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_154
timestamp 1604666999
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_157
timestamp 1604666999
transform 1 0 15548 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 15548 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 16008 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1604666999
transform 1 0 16284 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_161
timestamp 1604666999
transform 1 0 15916 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_164
timestamp 1604666999
transform 1 0 16192 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_174
timestamp 1604666999
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_178
timestamp 1604666999
transform 1 0 17480 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_159
timestamp 1604666999
transform 1 0 15732 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_186
timestamp 1604666999
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_181
timestamp 1604666999
transform 1 0 17756 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1604666999
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1604666999
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 18216 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 17664 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__S
timestamp 1604666999
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__A0
timestamp 1604666999
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604666999
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_190
timestamp 1604666999
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 18768 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_194
timestamp 1604666999
transform 1 0 18952 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_188
timestamp 1604666999
transform 1 0 18400 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604666999
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_200
timestamp 1604666999
transform 1 0 19504 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_212
timestamp 1604666999
transform 1 0 20608 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_206
timestamp 1604666999
transform 1 0 20056 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604666999
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_224
timestamp 1604666999
transform 1 0 21712 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_236
timestamp 1604666999
transform 1 0 22816 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1604666999
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604666999
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1604666999
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1604666999
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1604666999
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1604666999
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604666999
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604666999
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604666999
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1604666999
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1604666999
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604666999
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1604666999
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604666999
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 2668 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_12
timestamp 1604666999
transform 1 0 2208 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_16
timestamp 1604666999
transform 1 0 2576 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_19
timestamp 1604666999
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1604666999
transform 1 0 3220 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_32
timestamp 1604666999
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_36
timestamp 1604666999
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1604666999
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_40
timestamp 1604666999
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1604666999
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1604666999
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 7820 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604666999
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1604666999
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_66
timestamp 1604666999
transform 1 0 7176 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_69
timestamp 1604666999
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_92
timestamp 1604666999
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_96
timestamp 1604666999
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604666999
transform 1 0 10304 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_109
timestamp 1604666999
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1604666999
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_117
timestamp 1604666999
transform 1 0 11868 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604666999
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1604666999
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_136
timestamp 1604666999
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1604666999
transform 1 0 13984 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604666999
transform 1 0 15548 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_149
timestamp 1604666999
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_153
timestamp 1604666999
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 16560 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1604666999
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_170
timestamp 1604666999
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_174
timestamp 1604666999
transform 1 0 17112 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1604666999
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604666999
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_6__A1
timestamp 1604666999
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1604666999
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_193
timestamp 1604666999
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_197
timestamp 1604666999
transform 1 0 19228 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_209
timestamp 1604666999
transform 1 0 20332 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_221
timestamp 1604666999
transform 1 0 21436 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_233
timestamp 1604666999
transform 1 0 22540 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604666999
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_241
timestamp 1604666999
transform 1 0 23276 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1604666999
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1604666999
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604666999
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_269
timestamp 1604666999
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604666999
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604666999
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_6
timestamp 1604666999
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_10
timestamp 1604666999
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604666999
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 4508 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1604666999
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1604666999
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_35
timestamp 1604666999
transform 1 0 4324 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_39
timestamp 1604666999
transform 1 0 4692 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 5428 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_43
timestamp 1604666999
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604666999
transform 1 0 7912 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 7728 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_66
timestamp 1604666999
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_70
timestamp 1604666999
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_83
timestamp 1604666999
transform 1 0 8740 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 8924 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_87
timestamp 1604666999
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 9292 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1604666999
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1604666999
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604666999
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_97
timestamp 1604666999
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 10396 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1604666999
transform 1 0 12880 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_120
timestamp 1604666999
transform 1 0 12144 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_125
timestamp 1604666999
transform 1 0 12604 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_137
timestamp 1604666999
transform 1 0 13708 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_145
timestamp 1604666999
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1604666999
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1604666999
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_149
timestamp 1604666999
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604666999
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 15548 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 17480 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_176
timestamp 1604666999
transform 1 0 17296 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_6_
timestamp 1604666999
transform 1 0 18032 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_180
timestamp 1604666999
transform 1 0 17664 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_193
timestamp 1604666999
transform 1 0 18860 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604666999
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_205
timestamp 1604666999
transform 1 0 19964 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1604666999
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604666999
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1604666999
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1604666999
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1604666999
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604666999
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604666999
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1604666999
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604666999
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604666999
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 2852 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604666999
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 2668 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1604666999
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_11
timestamp 1604666999
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_15
timestamp 1604666999
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_38
timestamp 1604666999
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_42
timestamp 1604666999
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604666999
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 5336 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_49
timestamp 1604666999
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_53
timestamp 1604666999
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1604666999
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 6808 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604666999
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1604666999
transform 1 0 9292 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_81
timestamp 1604666999
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_85
timestamp 1604666999
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_98
timestamp 1604666999
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604666999
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_102
timestamp 1604666999
transform 1 0 10488 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_107
timestamp 1604666999
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1604666999
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604666999
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12512 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604666999
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_123
timestamp 1604666999
transform 1 0 12420 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604666999
transform 1 0 14996 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_143
timestamp 1604666999
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_147
timestamp 1604666999
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A0
timestamp 1604666999
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__S
timestamp 1604666999
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_160
timestamp 1604666999
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_164
timestamp 1604666999
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_168
timestamp 1604666999
transform 1 0 16560 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_172
timestamp 1604666999
transform 1 0 16928 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1604666999
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_4_
timestamp 1604666999
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604666999
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A1
timestamp 1604666999
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1604666999
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1604666999
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_197
timestamp 1604666999
transform 1 0 19228 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_209
timestamp 1604666999
transform 1 0 20332 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_221
timestamp 1604666999
transform 1 0 21436 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_233
timestamp 1604666999
transform 1 0 22540 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604666999
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_241
timestamp 1604666999
transform 1 0 23276 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1604666999
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1604666999
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604666999
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1604666999
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 1380 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604666999
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604666999
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604666999
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604666999
transform 1 0 3312 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 3680 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_22
timestamp 1604666999
transform 1 0 3128 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1604666999
transform 1 0 3496 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1604666999
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_36
timestamp 1604666999
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 5336 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_40
timestamp 1604666999
transform 1 0 4784 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 7820 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 7268 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_65
timestamp 1604666999
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_69
timestamp 1604666999
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604666999
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604666999
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_82
timestamp 1604666999
transform 1 0 8648 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_88
timestamp 1604666999
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604666999
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1604666999
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_106
timestamp 1604666999
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_119
timestamp 1604666999
transform 1 0 12052 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604666999
transform 1 0 12788 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 13800 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_123
timestamp 1604666999
transform 1 0 12420 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_126
timestamp 1604666999
transform 1 0 12696 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_136
timestamp 1604666999
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_140
timestamp 1604666999
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 14168 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_144
timestamp 1604666999
transform 1 0 14352 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_149
timestamp 1604666999
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1604666999
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604666999
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_158
timestamp 1604666999
transform 1 0 15640 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 15456 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_5_
timestamp 1604666999
transform 1 0 17388 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604666999
transform 1 0 15824 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_169
timestamp 1604666999
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_173
timestamp 1604666999
transform 1 0 17020 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_186
timestamp 1604666999
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_190
timestamp 1604666999
transform 1 0 18584 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_194
timestamp 1604666999
transform 1 0 18952 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604666999
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_206
timestamp 1604666999
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_215
timestamp 1604666999
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_227
timestamp 1604666999
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1604666999
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_251
timestamp 1604666999
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604666999
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604666999
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_263
timestamp 1604666999
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604666999
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_6
timestamp 1604666999
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1604666999
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1604666999
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604666999
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604666999
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_10
timestamp 1604666999
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 2024 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1604666999
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1604666999
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_29
timestamp 1604666999
transform 1 0 3772 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_38
timestamp 1604666999
transform 1 0 4600 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_34
timestamp 1604666999
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604666999
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604666999
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_46
timestamp 1604666999
transform 1 0 5336 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_41
timestamp 1604666999
transform 1 0 4876 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1604666999
transform 1 0 5612 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1604666999
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_58
timestamp 1604666999
transform 1 0 6440 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604666999
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604666999
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_62
timestamp 1604666999
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604666999
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604666999
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604666999
transform 1 0 7176 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_75
timestamp 1604666999
transform 1 0 8004 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_79
timestamp 1604666999
transform 1 0 8372 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_75
timestamp 1604666999
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_71
timestamp 1604666999
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_88
timestamp 1604666999
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1604666999
transform 1 0 8924 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_81
timestamp 1604666999
transform 1 0 8556 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_83
timestamp 1604666999
transform 1 0 8740 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604666999
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9016 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_20_106
timestamp 1604666999
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1604666999
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_109
timestamp 1604666999
transform 1 0 11132 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_105
timestamp 1604666999
transform 1 0 10764 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_116
timestamp 1604666999
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_112
timestamp 1604666999
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1604666999
transform 1 0 11224 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_119
timestamp 1604666999
transform 1 0 12052 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_128
timestamp 1604666999
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_124
timestamp 1604666999
transform 1 0 12512 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1604666999
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 12328 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 12696 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604666999
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1604666999
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_132
timestamp 1604666999
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_138
timestamp 1604666999
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_132
timestamp 1604666999
transform 1 0 13248 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_145
timestamp 1604666999
transform 1 0 14444 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_146
timestamp 1604666999
transform 1 0 14536 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_142
timestamp 1604666999
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1604666999
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_152
timestamp 1604666999
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604666999
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 15456 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 16652 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1604666999
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1604666999
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_167
timestamp 1604666999
transform 1 0 16468 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_171
timestamp 1604666999
transform 1 0 16836 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 17940 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604666999
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 18216 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 18584 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_179
timestamp 1604666999
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1604666999
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_188
timestamp 1604666999
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_192
timestamp 1604666999
transform 1 0 18768 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604666999
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_204
timestamp 1604666999
transform 1 0 19872 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_216
timestamp 1604666999
transform 1 0 20976 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1604666999
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1604666999
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_228
timestamp 1604666999
transform 1 0 22080 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_227
timestamp 1604666999
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604666999
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_240
timestamp 1604666999
transform 1 0 23184 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_245
timestamp 1604666999
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_257
timestamp 1604666999
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_239
timestamp 1604666999
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_251
timestamp 1604666999
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604666999
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604666999
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604666999
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1604666999
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_263
timestamp 1604666999
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604666999
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604666999
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1604666999
transform 1 0 2852 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604666999
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 2024 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_7
timestamp 1604666999
transform 1 0 1748 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_12
timestamp 1604666999
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_16
timestamp 1604666999
transform 1 0 2576 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_28
timestamp 1604666999
transform 1 0 3680 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_34
timestamp 1604666999
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_38
timestamp 1604666999
transform 1 0 4600 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604666999
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1604666999
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604666999
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604666999
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604666999
transform 1 0 8372 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604666999
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1604666999
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_75
timestamp 1604666999
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_1_
timestamp 1604666999
transform 1 0 9936 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_88
timestamp 1604666999
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_92
timestamp 1604666999
transform 1 0 9568 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 10948 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 11316 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_105
timestamp 1604666999
transform 1 0 10764 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_109
timestamp 1604666999
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1604666999
transform 1 0 11500 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp 1604666999
transform 1 0 12052 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1604666999
transform 1 0 13248 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604666999
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 12696 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_123
timestamp 1604666999
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_128
timestamp 1604666999
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 14812 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 14260 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_141
timestamp 1604666999
transform 1 0 14076 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_145
timestamp 1604666999
transform 1 0 14444 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_168
timestamp 1604666999
transform 1 0 16560 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_173
timestamp 1604666999
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_177
timestamp 1604666999
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604666999
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1604666999
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604666999
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1604666999
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1604666999
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_220
timestamp 1604666999
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_232
timestamp 1604666999
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604666999
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1604666999
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1604666999
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604666999
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_269
timestamp 1604666999
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1604666999
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604666999
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604666999
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_6
timestamp 1604666999
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_10
timestamp 1604666999
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4048 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604666999
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_23
timestamp 1604666999
transform 1 0 3220 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1604666999
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 6532 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 5980 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 6348 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_51
timestamp 1604666999
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_55
timestamp 1604666999
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_78
timestamp 1604666999
transform 1 0 8280 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l3_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604666999
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1604666999
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1604666999
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_102
timestamp 1604666999
transform 1 0 10488 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_114
timestamp 1604666999
transform 1 0 11592 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 12696 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_122
timestamp 1604666999
transform 1 0 12328 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_125
timestamp 1604666999
transform 1 0 12604 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604666999
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604666999
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1604666999
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1604666999
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604666999
transform 1 0 16836 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 16376 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_163
timestamp 1604666999
transform 1 0 16100 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_168
timestamp 1604666999
transform 1 0 16560 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_180
timestamp 1604666999
transform 1 0 17664 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_192
timestamp 1604666999
transform 1 0 18768 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604666999
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_204
timestamp 1604666999
transform 1 0 19872 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1604666999
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604666999
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1604666999
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1604666999
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_251
timestamp 1604666999
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604666999
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604666999
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_263
timestamp 1604666999
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604666999
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604666999
transform 1 0 2484 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604666999
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604666999
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604666999
transform 1 0 2300 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1604666999
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_11
timestamp 1604666999
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_19
timestamp 1604666999
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 3588 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_23
timestamp 1604666999
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_30
timestamp 1604666999
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_34
timestamp 1604666999
transform 1 0 4232 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1604666999
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_40
timestamp 1604666999
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604666999
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604666999
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1604666999
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604666999
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1604666999
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_75
timestamp 1604666999
transform 1 0 8004 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_79
timestamp 1604666999
transform 1 0 8372 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 8648 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 10764 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_101
timestamp 1604666999
transform 1 0 10396 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_107
timestamp 1604666999
transform 1 0 10948 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_111
timestamp 1604666999
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_115
timestamp 1604666999
transform 1 0 11684 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_119
timestamp 1604666999
transform 1 0 12052 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1604666999
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604666999
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_127
timestamp 1604666999
transform 1 0 12788 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 12972 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_131
timestamp 1604666999
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_135
timestamp 1604666999
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 13892 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_23_158
timestamp 1604666999
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_162
timestamp 1604666999
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_175
timestamp 1604666999
transform 1 0 17204 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604666999
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604666999
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1604666999
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1604666999
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_220
timestamp 1604666999
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_232
timestamp 1604666999
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604666999
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1604666999
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1604666999
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604666999
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_269
timestamp 1604666999
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604666999
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1604666999
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_6
timestamp 1604666999
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_10
timestamp 1604666999
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604666999
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 4508 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604666999
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_23
timestamp 1604666999
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1604666999
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_35
timestamp 1604666999
transform 1 0 4324 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_39
timestamp 1604666999
transform 1 0 4692 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 5704 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 5520 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_43
timestamp 1604666999
transform 1 0 5060 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_46
timestamp 1604666999
transform 1 0 5336 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 8004 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_69
timestamp 1604666999
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_73
timestamp 1604666999
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_77
timestamp 1604666999
transform 1 0 8188 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604666999
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1604666999
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_88
timestamp 1604666999
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1604666999
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604666999
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_97
timestamp 1604666999
transform 1 0 10028 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 10212 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l3_in_0_
timestamp 1604666999
transform 1 0 10764 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_101
timestamp 1604666999
transform 1 0 10396 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_114
timestamp 1604666999
transform 1 0 11592 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12328 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 13708 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_131
timestamp 1604666999
transform 1 0 13156 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 14168 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604666999
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_139
timestamp 1604666999
transform 1 0 13892 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_145
timestamp 1604666999
transform 1 0 14444 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_149
timestamp 1604666999
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_163
timestamp 1604666999
transform 1 0 16100 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_168
timestamp 1604666999
transform 1 0 16560 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_180
timestamp 1604666999
transform 1 0 17664 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_192
timestamp 1604666999
transform 1 0 18768 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604666999
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_204
timestamp 1604666999
transform 1 0 19872 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1604666999
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604666999
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1604666999
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1604666999
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_251
timestamp 1604666999
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604666999
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604666999
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1604666999
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604666999
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604666999
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 2852 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604666999
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604666999
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1604666999
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1604666999
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_15
timestamp 1604666999
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_38
timestamp 1604666999
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_42
timestamp 1604666999
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_46
timestamp 1604666999
transform 1 0 5336 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 5152 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604666999
transform 1 0 5704 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1604666999
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1604666999
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 7084 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604666999
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_62
timestamp 1604666999
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 9752 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_84
timestamp 1604666999
transform 1 0 8832 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_90
timestamp 1604666999
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12052 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1604666999
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_117
timestamp 1604666999
transform 1 0 11868 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604666999
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 13708 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604666999
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1604666999
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_126
timestamp 1604666999
transform 1 0 12696 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_134
timestamp 1604666999
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_156
timestamp 1604666999
transform 1 0 15456 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_168
timestamp 1604666999
transform 1 0 16560 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604666999
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1604666999
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1604666999
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1604666999
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1604666999
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1604666999
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_232
timestamp 1604666999
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604666999
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1604666999
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1604666999
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604666999
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_269
timestamp 1604666999
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604666999
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604666999
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604666999
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604666999
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_7
timestamp 1604666999
transform 1 0 1748 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1604666999
transform 1 0 1748 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_12
timestamp 1604666999
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_11
timestamp 1604666999
transform 1 0 2116 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 2300 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 2024 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_16
timestamp 1604666999
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_19
timestamp 1604666999
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1604666999
transform 1 0 2484 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 2944 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1604666999
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604666999
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1604666999
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1604666999
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1604666999
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_39
timestamp 1604666999
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_43
timestamp 1604666999
transform 1 0 5060 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_45
timestamp 1604666999
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_41
timestamp 1604666999
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 5428 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 5244 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 4876 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1604666999
transform 1 0 5612 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 5428 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1604666999
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_54
timestamp 1604666999
transform 1 0 6072 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_50
timestamp 1604666999
transform 1 0 5704 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_58
timestamp 1604666999
transform 1 0 6440 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_62
timestamp 1604666999
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604666999
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1604666999
transform 1 0 7176 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l3_in_0_
timestamp 1604666999
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_75
timestamp 1604666999
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_71
timestamp 1604666999
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_79
timestamp 1604666999
transform 1 0 8372 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_75
timestamp 1604666999
transform 1 0 8004 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 8188 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 8372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_86
timestamp 1604666999
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_82
timestamp 1604666999
transform 1 0 8648 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_89
timestamp 1604666999
transform 1 0 9292 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_83
timestamp 1604666999
transform 1 0 8740 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 8556 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 8832 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604666999
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9384 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_109
timestamp 1604666999
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_106
timestamp 1604666999
transform 1 0 10856 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_102
timestamp 1604666999
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_117
timestamp 1604666999
transform 1 0 11868 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1604666999
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_114
timestamp 1604666999
transform 1 0 11592 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 11316 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 11684 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_128
timestamp 1604666999
transform 1 0 12880 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_123
timestamp 1604666999
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1604666999
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12696 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604666999
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1604666999
transform 1 0 13800 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_134
timestamp 1604666999
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 13616 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 13064 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 13248 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604666999
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_142
timestamp 1604666999
transform 1 0 14168 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_150
timestamp 1604666999
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1604666999
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_151
timestamp 1604666999
transform 1 0 14996 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1604666999
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1604666999
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_163
timestamp 1604666999
transform 1 0 16100 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_175
timestamp 1604666999
transform 1 0 17204 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604666999
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1604666999
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604666999
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604666999
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604666999
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1604666999
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604666999
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604666999
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1604666999
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1604666999
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1604666999
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604666999
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1604666999
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1604666999
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1604666999
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1604666999
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604666999
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604666999
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604666999
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1604666999
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604666999
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1604666999
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1604666999
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1604666999
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604666999
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1604666999
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1604666999
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_6
timestamp 1604666999
transform 1 0 1656 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_10
timestamp 1604666999
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_3_
timestamp 1604666999
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604666999
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1604666999
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1604666999
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604666999
transform 1 0 5612 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 6440 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 6072 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 5428 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_41
timestamp 1604666999
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_45
timestamp 1604666999
transform 1 0 5244 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_52
timestamp 1604666999
transform 1 0 5888 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_56
timestamp 1604666999
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 6624 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_28_79
timestamp 1604666999
transform 1 0 8372 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 9936 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604666999
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_83
timestamp 1604666999
transform 1 0 8740 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1604666999
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_93
timestamp 1604666999
transform 1 0 9660 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_99
timestamp 1604666999
transform 1 0 10212 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 10948 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10396 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_103
timestamp 1604666999
transform 1 0 10580 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13432 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12880 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_126
timestamp 1604666999
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_130
timestamp 1604666999
transform 1 0 13064 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604666999
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_143
timestamp 1604666999
transform 1 0 14260 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_147
timestamp 1604666999
transform 1 0 14628 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604666999
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1604666999
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1604666999
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1604666999
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604666999
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1604666999
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604666999
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604666999
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604666999
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1604666999
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604666999
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604666999
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1604666999
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604666999
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1604666999
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_2_
timestamp 1604666999
transform 1 0 2668 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604666999
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1604666999
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_7
timestamp 1604666999
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_13
timestamp 1604666999
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4232 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 3680 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_26
timestamp 1604666999
transform 1 0 3496 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_30
timestamp 1604666999
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1604666999
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1604666999
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 7084 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604666999
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_62
timestamp 1604666999
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1604666999
transform 1 0 9936 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 9292 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_84
timestamp 1604666999
transform 1 0 8832 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_88
timestamp 1604666999
transform 1 0 9200 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_91
timestamp 1604666999
transform 1 0 9476 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_95
timestamp 1604666999
transform 1 0 9844 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 10948 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 11316 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_105
timestamp 1604666999
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_109
timestamp 1604666999
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1604666999
transform 1 0 11500 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604666999
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_1_
timestamp 1604666999
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604666999
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13432 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_132
timestamp 1604666999
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_136
timestamp 1604666999
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_1_
timestamp 1604666999
transform 1 0 13984 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 14996 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_149
timestamp 1604666999
transform 1 0 14812 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_153
timestamp 1604666999
transform 1 0 15180 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_165
timestamp 1604666999
transform 1 0 16284 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_177
timestamp 1604666999
transform 1 0 17388 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604666999
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604666999
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604666999
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604666999
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1604666999
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1604666999
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604666999
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1604666999
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1604666999
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604666999
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp 1604666999
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1604666999
transform 1 0 2484 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1604666999
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604666999
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1604666999
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 2300 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1604666999
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1604666999
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_19
timestamp 1604666999
transform 1 0 2852 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1604666999
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_23
timestamp 1604666999
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 3036 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_36
timestamp 1604666999
transform 1 0 4416 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_32
timestamp 1604666999
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 4232 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604666999
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604666999
transform 1 0 4508 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604666999
transform 1 0 6072 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_46
timestamp 1604666999
transform 1 0 5336 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_1_
timestamp 1604666999
transform 1 0 7636 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_63
timestamp 1604666999
transform 1 0 6900 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_67
timestamp 1604666999
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604666999
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_80
timestamp 1604666999
transform 1 0 8464 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1604666999
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _027_
timestamp 1604666999
transform 1 0 11224 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11040 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 11684 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12052 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_102
timestamp 1604666999
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_106
timestamp 1604666999
transform 1 0 10856 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_113
timestamp 1604666999
transform 1 0 11500 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_117
timestamp 1604666999
transform 1 0 11868 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 12696 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_121
timestamp 1604666999
transform 1 0 12236 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_125
timestamp 1604666999
transform 1 0 12604 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1604666999
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604666999
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_145
timestamp 1604666999
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1604666999
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_157
timestamp 1604666999
transform 1 0 15548 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_169
timestamp 1604666999
transform 1 0 16652 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_181
timestamp 1604666999
transform 1 0 17756 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_193
timestamp 1604666999
transform 1 0 18860 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604666999
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_205
timestamp 1604666999
transform 1 0 19964 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_213
timestamp 1604666999
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604666999
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1604666999
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1604666999
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1604666999
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604666999
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604666999
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1604666999
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604666999
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1604666999
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 2484 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604666999
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1604666999
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2300 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_7
timestamp 1604666999
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1604666999
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_18
timestamp 1604666999
transform 1 0 2760 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604666999
transform 1 0 3772 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_22
timestamp 1604666999
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_25
timestamp 1604666999
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_38
timestamp 1604666999
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1604666999
transform 1 0 5336 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 5152 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_42
timestamp 1604666999
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_49
timestamp 1604666999
transform 1 0 5612 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604666999
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604666999
transform 1 0 7636 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604666999
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 7452 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 6992 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1604666999
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_66
timestamp 1604666999
transform 1 0 7176 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9200 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 9016 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_80
timestamp 1604666999
transform 1 0 8464 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_84
timestamp 1604666999
transform 1 0 8832 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_97
timestamp 1604666999
transform 1 0 10028 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1604666999
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 10488 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_101
timestamp 1604666999
transform 1 0 10396 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_104
timestamp 1604666999
transform 1 0 10672 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_114
timestamp 1604666999
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604666999
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1604666999
transform 1 0 12604 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604666999
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_123
timestamp 1604666999
transform 1 0 12420 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_134
timestamp 1604666999
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_138
timestamp 1604666999
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 14168 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 13984 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_161
timestamp 1604666999
transform 1 0 15916 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_173
timestamp 1604666999
transform 1 0 17020 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604666999
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1604666999
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604666999
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604666999
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1604666999
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1604666999
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1604666999
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604666999
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1604666999
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1604666999
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604666999
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_269
timestamp 1604666999
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1604666999
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604666999
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1604666999
transform 1 0 1932 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_7
timestamp 1604666999
transform 1 0 1748 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_11
timestamp 1604666999
transform 1 0 2116 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_19
timestamp 1604666999
transform 1 0 2852 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604666999
transform 1 0 2944 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 4048 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604666999
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_23
timestamp 1604666999
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1604666999
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604666999
transform 1 0 6532 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_51
timestamp 1604666999
transform 1 0 5796 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 7636 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 8004 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 8372 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_68
timestamp 1604666999
transform 1 0 7360 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_73
timestamp 1604666999
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_77
timestamp 1604666999
transform 1 0 8188 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604666999
transform 1 0 8556 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604666999
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9844 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 10212 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_84
timestamp 1604666999
transform 1 0 8832 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_90
timestamp 1604666999
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1604666999
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_97
timestamp 1604666999
transform 1 0 10028 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 10488 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_32_101
timestamp 1604666999
transform 1 0 10396 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13340 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 12604 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12972 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_121
timestamp 1604666999
transform 1 0 12236 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_127
timestamp 1604666999
transform 1 0 12788 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_131
timestamp 1604666999
transform 1 0 13156 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604666999
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14720 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_142
timestamp 1604666999
transform 1 0 14168 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_146
timestamp 1604666999
transform 1 0 14536 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_150
timestamp 1604666999
transform 1 0 14904 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1604666999
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1604666999
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1604666999
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1604666999
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604666999
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1604666999
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604666999
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604666999
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1604666999
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1604666999
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604666999
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604666999
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1604666999
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604666999
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1604666999
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_3
timestamp 1604666999
transform 1 0 1380 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 1564 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604666999
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604666999
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1472 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_11
timestamp 1604666999
transform 1 0 2116 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_7
timestamp 1604666999
transform 1 0 1748 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_11
timestamp 1604666999
transform 1 0 2116 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1604666999
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 2208 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_18
timestamp 1604666999
transform 1 0 2760 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_14
timestamp 1604666999
transform 1 0 2392 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_15
timestamp 1604666999
transform 1 0 2484 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 2852 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 2576 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1604666999
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_24
timestamp 1604666999
transform 1 0 3312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_21
timestamp 1604666999
transform 1 0 3036 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_32
timestamp 1604666999
transform 1 0 4048 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604666999
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604666999
transform 1 0 4324 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 3404 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_34_48
timestamp 1604666999
transform 1 0 5520 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_44
timestamp 1604666999
transform 1 0 5152 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_44
timestamp 1604666999
transform 1 0 5152 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 5520 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 5336 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_58
timestamp 1604666999
transform 1 0 6440 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1604666999
transform 1 0 6072 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_50
timestamp 1604666999
transform 1 0 5704 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 5704 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 6256 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604666999
transform 1 0 5888 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_65
timestamp 1604666999
transform 1 0 7084 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_61
timestamp 1604666999
transform 1 0 6716 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_62
timestamp 1604666999
transform 1 0 6808 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 6900 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 7268 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 7176 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604666999
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1604666999
transform 1 0 7452 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_78
timestamp 1604666999
transform 1 0 8280 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 7360 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_34_87
timestamp 1604666999
transform 1 0 9108 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_82
timestamp 1604666999
transform 1 0 8648 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_87
timestamp 1604666999
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 8464 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 8924 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1604666999
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_91
timestamp 1604666999
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604666999
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9660 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_19.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9844 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 11592 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_114
timestamp 1604666999
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_118
timestamp 1604666999
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_112
timestamp 1604666999
transform 1 0 11408 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_116
timestamp 1604666999
transform 1 0 11776 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_127
timestamp 1604666999
transform 1 0 12788 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_123
timestamp 1604666999
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604666999
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 12144 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_135
timestamp 1604666999
transform 1 0 13524 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_131
timestamp 1604666999
transform 1 0 13156 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 12972 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13340 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_21.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12420 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_34_145
timestamp 1604666999
transform 1 0 14444 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_146
timestamp 1604666999
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_142
timestamp 1604666999
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_154
timestamp 1604666999
transform 1 0 15272 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_150
timestamp 1604666999
transform 1 0 14904 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 15456 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 15088 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604666999
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_158
timestamp 1604666999
transform 1 0 15640 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_154
timestamp 1604666999
transform 1 0 15272 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_166
timestamp 1604666999
transform 1 0 16376 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_178
timestamp 1604666999
transform 1 0 17480 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_170
timestamp 1604666999
transform 1 0 16744 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604666999
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_182
timestamp 1604666999
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604666999
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604666999
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_182
timestamp 1604666999
transform 1 0 17848 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_194
timestamp 1604666999
transform 1 0 18952 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604666999
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1604666999
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_206
timestamp 1604666999
transform 1 0 20056 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604666999
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1604666999
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1604666999
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604666999
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604666999
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1604666999
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1604666999
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1604666999
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1604666999
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604666999
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604666999
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604666999
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1604666999
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1604666999
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604666999
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 2208 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604666999
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 2024 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 1564 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1604666999
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_7
timestamp 1604666999
transform 1 0 1748 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 4692 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 4324 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_31
timestamp 1604666999
transform 1 0 3956 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_37
timestamp 1604666999
transform 1 0 4508 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1604666999
transform 1 0 4876 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 6440 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 6072 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_50
timestamp 1604666999
transform 1 0 5704 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_56
timestamp 1604666999
transform 1 0 6256 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604666999
transform 1 0 6992 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604666999
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 8372 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_60
timestamp 1604666999
transform 1 0 6624 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_62
timestamp 1604666999
transform 1 0 6808 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_73
timestamp 1604666999
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_77
timestamp 1604666999
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_1_
timestamp 1604666999
transform 1 0 8924 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10120 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 8740 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_81
timestamp 1604666999
transform 1 0 8556 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_94
timestamp 1604666999
transform 1 0 9752 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_1_
timestamp 1604666999
transform 1 0 10764 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10488 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_100
timestamp 1604666999
transform 1 0 10304 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_104
timestamp 1604666999
transform 1 0 10672 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_114
timestamp 1604666999
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1604666999
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604666999
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_132
timestamp 1604666999
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_136
timestamp 1604666999
transform 1 0 13616 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 14168 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13984 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 16100 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_161
timestamp 1604666999
transform 1 0 15916 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_165
timestamp 1604666999
transform 1 0 16284 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_177
timestamp 1604666999
transform 1 0 17388 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604666999
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1604666999
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1604666999
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1604666999
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1604666999
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1604666999
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604666999
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_245
timestamp 1604666999
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_257
timestamp 1604666999
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604666999
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1604666999
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 1380 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604666999
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604666999
transform 1 0 4048 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604666999
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_22
timestamp 1604666999
transform 1 0 3128 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1604666999
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604666999
transform 1 0 6440 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6256 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 5152 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 5888 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 5520 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_41
timestamp 1604666999
transform 1 0 4876 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_46
timestamp 1604666999
transform 1 0 5336 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_50
timestamp 1604666999
transform 1 0 5704 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_54
timestamp 1604666999
transform 1 0 6072 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604666999
transform 1 0 8004 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 7452 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_67
timestamp 1604666999
transform 1 0 7268 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_71
timestamp 1604666999
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_78
timestamp 1604666999
transform 1 0 8280 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604666999
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 8924 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_84
timestamp 1604666999
transform 1 0 8832 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_87
timestamp 1604666999
transform 1 0 9108 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_91
timestamp 1604666999
transform 1 0 9476 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_93
timestamp 1604666999
transform 1 0 9660 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_99
timestamp 1604666999
transform 1 0 10212 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10488 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 11500 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 10304 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_111
timestamp 1604666999
transform 1 0 11316 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_115
timestamp 1604666999
transform 1 0 11684 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1604666999
transform 1 0 12328 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13340 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 13156 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_121
timestamp 1604666999
transform 1 0 12236 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_125
timestamp 1604666999
transform 1 0 12604 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 15272 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604666999
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 14352 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_142
timestamp 1604666999
transform 1 0 14168 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_146
timestamp 1604666999
transform 1 0 14536 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_152
timestamp 1604666999
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_173
timestamp 1604666999
transform 1 0 17020 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_185
timestamp 1604666999
transform 1 0 18124 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1604666999
transform 1 0 19228 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604666999
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_209
timestamp 1604666999
transform 1 0 20332 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp 1604666999
transform 1 0 20700 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1604666999
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1604666999
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1604666999
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_251
timestamp 1604666999
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604666999
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604666999
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_263
timestamp 1604666999
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604666999
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1604666999
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 2668 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604666999
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__A
timestamp 1604666999
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 2484 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_7
timestamp 1604666999
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_11
timestamp 1604666999
transform 1 0 2116 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 4692 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_36
timestamp 1604666999
transform 1 0 4416 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604666999
transform 1 0 5152 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_41
timestamp 1604666999
transform 1 0 4876 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_53
timestamp 1604666999
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1604666999
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1604666999
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1604666999
transform 1 0 8372 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604666999
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_71
timestamp 1604666999
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_75
timestamp 1604666999
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 9660 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_88
timestamp 1604666999
transform 1 0 9200 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_92
timestamp 1604666999
transform 1 0 9568 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_95
timestamp 1604666999
transform 1 0 9844 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 10764 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_103
timestamp 1604666999
transform 1 0 10580 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_107
timestamp 1604666999
transform 1 0 10948 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_119
timestamp 1604666999
transform 1 0 12052 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604666999
transform 1 0 13524 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604666999
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604666999
transform 1 0 12696 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 13340 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_123
timestamp 1604666999
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_128
timestamp 1604666999
transform 1 0 12880 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_132
timestamp 1604666999
transform 1 0 13248 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604666999
transform 1 0 15456 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604666999
transform 1 0 15272 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 14536 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_144
timestamp 1604666999
transform 1 0 14352 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_148
timestamp 1604666999
transform 1 0 14720 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 16560 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604666999
transform 1 0 17020 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604666999
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_160
timestamp 1604666999
transform 1 0 15824 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1604666999
transform 1 0 16192 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_171
timestamp 1604666999
transform 1 0 16836 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_175
timestamp 1604666999
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604666999
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 18216 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_179
timestamp 1604666999
transform 1 0 17572 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_184
timestamp 1604666999
transform 1 0 18032 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_188
timestamp 1604666999
transform 1 0 18400 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 20884 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_200
timestamp 1604666999
transform 1 0 19504 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_212
timestamp 1604666999
transform 1 0 20608 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_217
timestamp 1604666999
transform 1 0 21068 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 22356 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_229
timestamp 1604666999
transform 1 0 22172 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_233
timestamp 1604666999
transform 1 0 22540 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604666999
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_241
timestamp 1604666999
transform 1 0 23276 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1604666999
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1604666999
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604666999
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1604666999
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604666999
transform 1 0 1748 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604666999
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 1564 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 2760 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1604666999
transform 1 0 1380 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_16
timestamp 1604666999
transform 1 0 2576 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_28
timestamp 1604666999
transform 1 0 3680 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1604666999
transform 1 0 3312 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_20
timestamp 1604666999
transform 1 0 2944 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 3128 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_36
timestamp 1604666999
transform 1 0 4416 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_32
timestamp 1604666999
transform 1 0 4048 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 4232 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604666999
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604666999
transform 1 0 4692 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 6256 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 5888 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_48
timestamp 1604666999
transform 1 0 5520 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_54
timestamp 1604666999
transform 1 0 6072 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 8372 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_75
timestamp 1604666999
transform 1 0 8004 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 9660 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604666999
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_81
timestamp 1604666999
transform 1 0 8556 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_89
timestamp 1604666999
transform 1 0 9292 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_96
timestamp 1604666999
transform 1 0 9936 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_108
timestamp 1604666999
transform 1 0 11040 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604666999
transform 1 0 12696 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 13800 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 13524 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_120
timestamp 1604666999
transform 1 0 12144 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_130
timestamp 1604666999
transform 1 0 13064 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_134
timestamp 1604666999
transform 1 0 13432 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_137
timestamp 1604666999
transform 1 0 13708 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604666999
transform 1 0 15272 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604666999
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 14260 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1604666999
transform 1 0 14076 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_145
timestamp 1604666999
transform 1 0 14444 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_158
timestamp 1604666999
transform 1 0 15640 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604666999
transform 1 0 17020 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_170
timestamp 1604666999
transform 1 0 16744 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_177
timestamp 1604666999
transform 1 0 17388 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 18124 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_188
timestamp 1604666999
transform 1 0 18400 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 20884 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604666999
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_200
timestamp 1604666999
transform 1 0 19504 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_212
timestamp 1604666999
transform 1 0 20608 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_218
timestamp 1604666999
transform 1 0 21160 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 22356 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_230
timestamp 1604666999
transform 1 0 22264 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_234
timestamp 1604666999
transform 1 0 22632 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_246
timestamp 1604666999
transform 1 0 23736 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604666999
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604666999
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_258
timestamp 1604666999
transform 1 0 24840 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_270
timestamp 1604666999
transform 1 0 25944 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_274
timestamp 1604666999
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604666999
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_6
timestamp 1604666999
transform 1 0 1656 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_7
timestamp 1604666999
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1604666999
transform 1 0 1380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 1564 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__055__A
timestamp 1604666999
transform 1 0 1840 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604666999
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604666999
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1604666999
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_10
timestamp 1604666999
transform 1 0 2024 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 2208 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604666999
transform 1 0 2116 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1604666999
transform 1 0 2392 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_27
timestamp 1604666999
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_23
timestamp 1604666999
transform 1 0 3220 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_24
timestamp 1604666999
transform 1 0 3312 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_20
timestamp 1604666999
transform 1 0 2944 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 3128 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 3404 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 3680 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_32
timestamp 1604666999
transform 1 0 4048 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_30
timestamp 1604666999
transform 1 0 3864 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 4048 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604666999
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604666999
transform 1 0 4140 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4232 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 5888 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_53
timestamp 1604666999
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1604666999
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_42
timestamp 1604666999
transform 1 0 4968 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_46
timestamp 1604666999
transform 1 0 5336 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 7084 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 7452 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604666999
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 7084 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_62
timestamp 1604666999
transform 1 0 6808 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_61
timestamp 1604666999
transform 1 0 6716 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_67
timestamp 1604666999
transform 1 0 7268 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_78
timestamp 1604666999
transform 1 0 8280 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604666999
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 9016 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_84
timestamp 1604666999
transform 1 0 8832 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_88
timestamp 1604666999
transform 1 0 9200 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_90
timestamp 1604666999
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_93
timestamp 1604666999
transform 1 0 9660 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_101
timestamp 1604666999
transform 1 0 10396 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_109
timestamp 1604666999
transform 1 0 11132 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_105
timestamp 1604666999
transform 1 0 10764 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_100
timestamp 1604666999
transform 1 0 10304 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604666999
transform 1 0 10580 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604666999
transform 1 0 10580 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1604666999
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_114
timestamp 1604666999
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604666999
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604666999
transform 1 0 11224 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604666999
transform 1 0 12052 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_107
timestamp 1604666999
transform 1 0 10948 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_127
timestamp 1604666999
transform 1 0 12788 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604666999
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604666999
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1604666999
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_135
timestamp 1604666999
transform 1 0 13524 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_135
timestamp 1604666999
transform 1 0 13524 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_131
timestamp 1604666999
transform 1 0 13156 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1604666999
transform 1 0 13616 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__058__A
timestamp 1604666999
transform 1 0 12972 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1604666999
transform 1 0 13800 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_123
timestamp 1604666999
transform 1 0 12420 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_145
timestamp 1604666999
transform 1 0 14444 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_146
timestamp 1604666999
transform 1 0 14536 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_142
timestamp 1604666999
transform 1 0 14168 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A
timestamp 1604666999
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604666999
transform 1 0 14076 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_155
timestamp 1604666999
transform 1 0 15364 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604666999
transform 1 0 14812 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604666999
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604666999
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604666999
transform 1 0 14996 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_158
timestamp 1604666999
transform 1 0 15640 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604666999
transform 1 0 15548 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_166
timestamp 1604666999
transform 1 0 16376 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_159
timestamp 1604666999
transform 1 0 15732 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604666999
transform 1 0 16468 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604666999
transform 1 0 16468 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_171
timestamp 1604666999
transform 1 0 16836 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_174
timestamp 1604666999
transform 1 0 17112 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_169
timestamp 1604666999
transform 1 0 16652 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604666999
transform 1 0 17296 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604666999
transform 1 0 16744 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_178
timestamp 1604666999
transform 1 0 17480 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_183
timestamp 1604666999
transform 1 0 17940 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_184
timestamp 1604666999
transform 1 0 18032 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_182
timestamp 1604666999
transform 1 0 17848 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604666999
transform 1 0 17664 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604666999
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604666999
transform 1 0 17572 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604666999
transform 1 0 18124 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_191
timestamp 1604666999
transform 1 0 18676 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_197
timestamp 1604666999
transform 1 0 19228 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_193
timestamp 1604666999
transform 1 0 18860 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_189
timestamp 1604666999
transform 1 0 18492 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604666999
transform 1 0 19044 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604666999
transform 1 0 18676 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604666999
transform 1 0 18768 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604666999
transform 1 0 19320 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_196
timestamp 1604666999
transform 1 0 19136 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604666999
transform 1 0 21068 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604666999
transform 1 0 20884 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604666999
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604666999
transform 1 0 20884 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604666999
transform 1 0 19872 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_202
timestamp 1604666999
transform 1 0 19688 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_206
timestamp 1604666999
transform 1 0 20056 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_214
timestamp 1604666999
transform 1 0 20792 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_208
timestamp 1604666999
transform 1 0 20240 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604666999
transform 1 0 21620 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_221
timestamp 1604666999
transform 1 0 21436 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1604666999
transform 1 0 21804 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_237
timestamp 1604666999
transform 1 0 22908 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_219
timestamp 1604666999
transform 1 0 21252 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_231
timestamp 1604666999
transform 1 0 22356 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604666999
transform 1 0 23644 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604666999
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604666999
transform 1 0 24196 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_243
timestamp 1604666999
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_249
timestamp 1604666999
transform 1 0 24012 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_253
timestamp 1604666999
transform 1 0 24380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_243
timestamp 1604666999
transform 1 0 23460 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_255
timestamp 1604666999
transform 1 0 24564 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604666999
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604666999
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604666999
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_265
timestamp 1604666999
transform 1 0 25484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_267
timestamp 1604666999
transform 1 0 25668 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604666999
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1604666999
transform 1 0 1380 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1604666999
transform 1 0 2576 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604666999
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__057__A
timestamp 1604666999
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__054__A
timestamp 1604666999
transform 1 0 2392 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_7
timestamp 1604666999
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_11
timestamp 1604666999
transform 1 0 2116 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604666999
transform 1 0 4140 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 3956 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 3588 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_25
timestamp 1604666999
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_29
timestamp 1604666999
transform 1 0 3772 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_42
timestamp 1604666999
transform 1 0 4968 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_54
timestamp 1604666999
transform 1 0 6072 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604666999
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 7084 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 7452 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 7820 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_60
timestamp 1604666999
transform 1 0 6624 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_62
timestamp 1604666999
transform 1 0 6808 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_67
timestamp 1604666999
transform 1 0 7268 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_71
timestamp 1604666999
transform 1 0 7636 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_75
timestamp 1604666999
transform 1 0 8004 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_87
timestamp 1604666999
transform 1 0 9108 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_99
timestamp 1604666999
transform 1 0 10212 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_111
timestamp 1604666999
transform 1 0 11316 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_119
timestamp 1604666999
transform 1 0 12052 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604666999
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1604666999
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_135
timestamp 1604666999
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_147
timestamp 1604666999
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604666999
transform 1 0 16008 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604666999
transform 1 0 16560 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_159
timestamp 1604666999
transform 1 0 15732 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1604666999
transform 1 0 16376 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_170
timestamp 1604666999
transform 1 0 16744 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604666999
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_182
timestamp 1604666999
transform 1 0 17848 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1604666999
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1604666999
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1604666999
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1604666999
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1604666999
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604666999
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1604666999
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1604666999
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604666999
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1604666999
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _054_
timestamp 1604666999
transform 1 0 2484 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _055_
timestamp 1604666999
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604666999
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 2116 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_7
timestamp 1604666999
transform 1 0 1748 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_13
timestamp 1604666999
transform 1 0 2300 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_19
timestamp 1604666999
transform 1 0 2852 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604666999
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 3036 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 3404 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 4232 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_23
timestamp 1604666999
transform 1 0 3220 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604666999
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_32
timestamp 1604666999
transform 1 0 4048 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_36
timestamp 1604666999
transform 1 0 4416 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_48
timestamp 1604666999
transform 1 0 5520 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604666999
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_60
timestamp 1604666999
transform 1 0 6624 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_63
timestamp 1604666999
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604666999
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604666999
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_87
timestamp 1604666999
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_94
timestamp 1604666999
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1604666999
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_118
timestamp 1604666999
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604666999
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_125
timestamp 1604666999
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_137
timestamp 1604666999
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604666999
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_149
timestamp 1604666999
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1604666999
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604666999
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604666999
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_180
timestamp 1604666999
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604666999
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604666999
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604666999
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604666999
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604666999
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1604666999
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604666999
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1604666999
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604666999
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604666999
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604666999
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604666999
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_34_
port 0 nsew default input
rlabel metal2 s 846 0 902 480 6 bottom_left_grid_pin_35_
port 1 nsew default input
rlabel metal2 s 1398 0 1454 480 6 bottom_left_grid_pin_36_
port 2 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_left_grid_pin_37_
port 3 nsew default input
rlabel metal2 s 2502 0 2558 480 6 bottom_left_grid_pin_38_
port 4 nsew default input
rlabel metal2 s 3146 0 3202 480 6 bottom_left_grid_pin_39_
port 5 nsew default input
rlabel metal2 s 3698 0 3754 480 6 bottom_left_grid_pin_40_
port 6 nsew default input
rlabel metal2 s 4250 0 4306 480 6 bottom_left_grid_pin_41_
port 7 nsew default input
rlabel metal2 s 27618 0 27674 480 6 bottom_right_grid_pin_1_
port 8 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 ccff_head
port 9 nsew default input
rlabel metal3 s 27520 23264 28000 23384 6 ccff_tail
port 10 nsew default tristate
rlabel metal3 s 0 280 480 400 6 chanx_left_in[0]
port 11 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[10]
port 12 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[11]
port 13 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[12]
port 14 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[13]
port 15 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[14]
port 16 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[15]
port 17 nsew default input
rlabel metal3 s 0 9528 480 9648 6 chanx_left_in[16]
port 18 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[17]
port 19 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[18]
port 20 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[19]
port 21 nsew default input
rlabel metal3 s 0 824 480 944 6 chanx_left_in[1]
port 22 nsew default input
rlabel metal3 s 0 1368 480 1488 6 chanx_left_in[2]
port 23 nsew default input
rlabel metal3 s 0 1912 480 2032 6 chanx_left_in[3]
port 24 nsew default input
rlabel metal3 s 0 2592 480 2712 6 chanx_left_in[4]
port 25 nsew default input
rlabel metal3 s 0 3136 480 3256 6 chanx_left_in[5]
port 26 nsew default input
rlabel metal3 s 0 3680 480 3800 6 chanx_left_in[6]
port 27 nsew default input
rlabel metal3 s 0 4360 480 4480 6 chanx_left_in[7]
port 28 nsew default input
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[8]
port 29 nsew default input
rlabel metal3 s 0 5448 480 5568 6 chanx_left_in[9]
port 30 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_out[0]
port 31 nsew default tristate
rlabel metal3 s 0 17688 480 17808 6 chanx_left_out[10]
port 32 nsew default tristate
rlabel metal3 s 0 18368 480 18488 6 chanx_left_out[11]
port 33 nsew default tristate
rlabel metal3 s 0 18912 480 19032 6 chanx_left_out[12]
port 34 nsew default tristate
rlabel metal3 s 0 19456 480 19576 6 chanx_left_out[13]
port 35 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 chanx_left_out[14]
port 36 nsew default tristate
rlabel metal3 s 0 20680 480 20800 6 chanx_left_out[15]
port 37 nsew default tristate
rlabel metal3 s 0 21224 480 21344 6 chanx_left_out[16]
port 38 nsew default tristate
rlabel metal3 s 0 21768 480 21888 6 chanx_left_out[17]
port 39 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[18]
port 40 nsew default tristate
rlabel metal3 s 0 22992 480 23112 6 chanx_left_out[19]
port 41 nsew default tristate
rlabel metal3 s 0 12520 480 12640 6 chanx_left_out[1]
port 42 nsew default tristate
rlabel metal3 s 0 13064 480 13184 6 chanx_left_out[2]
port 43 nsew default tristate
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[3]
port 44 nsew default tristate
rlabel metal3 s 0 14288 480 14408 6 chanx_left_out[4]
port 45 nsew default tristate
rlabel metal3 s 0 14832 480 14952 6 chanx_left_out[5]
port 46 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chanx_left_out[6]
port 47 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[7]
port 48 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[8]
port 49 nsew default tristate
rlabel metal3 s 0 17144 480 17264 6 chanx_left_out[9]
port 50 nsew default tristate
rlabel metal2 s 4802 0 4858 480 6 chany_bottom_in[0]
port 51 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[10]
port 52 nsew default input
rlabel metal2 s 11058 0 11114 480 6 chany_bottom_in[11]
port 53 nsew default input
rlabel metal2 s 11702 0 11758 480 6 chany_bottom_in[12]
port 54 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[13]
port 55 nsew default input
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_in[14]
port 56 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[15]
port 57 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[16]
port 58 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_in[17]
port 59 nsew default input
rlabel metal2 s 15106 0 15162 480 6 chany_bottom_in[18]
port 60 nsew default input
rlabel metal2 s 15658 0 15714 480 6 chany_bottom_in[19]
port 61 nsew default input
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_in[1]
port 62 nsew default input
rlabel metal2 s 5998 0 6054 480 6 chany_bottom_in[2]
port 63 nsew default input
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_in[3]
port 64 nsew default input
rlabel metal2 s 7102 0 7158 480 6 chany_bottom_in[4]
port 65 nsew default input
rlabel metal2 s 7654 0 7710 480 6 chany_bottom_in[5]
port 66 nsew default input
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[6]
port 67 nsew default input
rlabel metal2 s 8850 0 8906 480 6 chany_bottom_in[7]
port 68 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[8]
port 69 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[9]
port 70 nsew default input
rlabel metal2 s 16210 0 16266 480 6 chany_bottom_out[0]
port 71 nsew default tristate
rlabel metal2 s 21914 0 21970 480 6 chany_bottom_out[10]
port 72 nsew default tristate
rlabel metal2 s 22466 0 22522 480 6 chany_bottom_out[11]
port 73 nsew default tristate
rlabel metal2 s 23110 0 23166 480 6 chany_bottom_out[12]
port 74 nsew default tristate
rlabel metal2 s 23662 0 23718 480 6 chany_bottom_out[13]
port 75 nsew default tristate
rlabel metal2 s 24214 0 24270 480 6 chany_bottom_out[14]
port 76 nsew default tristate
rlabel metal2 s 24766 0 24822 480 6 chany_bottom_out[15]
port 77 nsew default tristate
rlabel metal2 s 25318 0 25374 480 6 chany_bottom_out[16]
port 78 nsew default tristate
rlabel metal2 s 25962 0 26018 480 6 chany_bottom_out[17]
port 79 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[18]
port 80 nsew default tristate
rlabel metal2 s 27066 0 27122 480 6 chany_bottom_out[19]
port 81 nsew default tristate
rlabel metal2 s 16762 0 16818 480 6 chany_bottom_out[1]
port 82 nsew default tristate
rlabel metal2 s 17406 0 17462 480 6 chany_bottom_out[2]
port 83 nsew default tristate
rlabel metal2 s 17958 0 18014 480 6 chany_bottom_out[3]
port 84 nsew default tristate
rlabel metal2 s 18510 0 18566 480 6 chany_bottom_out[4]
port 85 nsew default tristate
rlabel metal2 s 19062 0 19118 480 6 chany_bottom_out[5]
port 86 nsew default tristate
rlabel metal2 s 19614 0 19670 480 6 chany_bottom_out[6]
port 87 nsew default tristate
rlabel metal2 s 20258 0 20314 480 6 chany_bottom_out[7]
port 88 nsew default tristate
rlabel metal2 s 20810 0 20866 480 6 chany_bottom_out[8]
port 89 nsew default tristate
rlabel metal2 s 21362 0 21418 480 6 chany_bottom_out[9]
port 90 nsew default tristate
rlabel metal2 s 4802 27520 4858 28000 6 chany_top_in[0]
port 91 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 chany_top_in[10]
port 92 nsew default input
rlabel metal2 s 11058 27520 11114 28000 6 chany_top_in[11]
port 93 nsew default input
rlabel metal2 s 11702 27520 11758 28000 6 chany_top_in[12]
port 94 nsew default input
rlabel metal2 s 12254 27520 12310 28000 6 chany_top_in[13]
port 95 nsew default input
rlabel metal2 s 12806 27520 12862 28000 6 chany_top_in[14]
port 96 nsew default input
rlabel metal2 s 13358 27520 13414 28000 6 chany_top_in[15]
port 97 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[16]
port 98 nsew default input
rlabel metal2 s 14554 27520 14610 28000 6 chany_top_in[17]
port 99 nsew default input
rlabel metal2 s 15106 27520 15162 28000 6 chany_top_in[18]
port 100 nsew default input
rlabel metal2 s 15658 27520 15714 28000 6 chany_top_in[19]
port 101 nsew default input
rlabel metal2 s 5354 27520 5410 28000 6 chany_top_in[1]
port 102 nsew default input
rlabel metal2 s 5998 27520 6054 28000 6 chany_top_in[2]
port 103 nsew default input
rlabel metal2 s 6550 27520 6606 28000 6 chany_top_in[3]
port 104 nsew default input
rlabel metal2 s 7102 27520 7158 28000 6 chany_top_in[4]
port 105 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chany_top_in[5]
port 106 nsew default input
rlabel metal2 s 8206 27520 8262 28000 6 chany_top_in[6]
port 107 nsew default input
rlabel metal2 s 8850 27520 8906 28000 6 chany_top_in[7]
port 108 nsew default input
rlabel metal2 s 9402 27520 9458 28000 6 chany_top_in[8]
port 109 nsew default input
rlabel metal2 s 9954 27520 10010 28000 6 chany_top_in[9]
port 110 nsew default input
rlabel metal2 s 16210 27520 16266 28000 6 chany_top_out[0]
port 111 nsew default tristate
rlabel metal2 s 21914 27520 21970 28000 6 chany_top_out[10]
port 112 nsew default tristate
rlabel metal2 s 22466 27520 22522 28000 6 chany_top_out[11]
port 113 nsew default tristate
rlabel metal2 s 23110 27520 23166 28000 6 chany_top_out[12]
port 114 nsew default tristate
rlabel metal2 s 23662 27520 23718 28000 6 chany_top_out[13]
port 115 nsew default tristate
rlabel metal2 s 24214 27520 24270 28000 6 chany_top_out[14]
port 116 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[15]
port 117 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[16]
port 118 nsew default tristate
rlabel metal2 s 25962 27520 26018 28000 6 chany_top_out[17]
port 119 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[18]
port 120 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 chany_top_out[19]
port 121 nsew default tristate
rlabel metal2 s 16762 27520 16818 28000 6 chany_top_out[1]
port 122 nsew default tristate
rlabel metal2 s 17406 27520 17462 28000 6 chany_top_out[2]
port 123 nsew default tristate
rlabel metal2 s 17958 27520 18014 28000 6 chany_top_out[3]
port 124 nsew default tristate
rlabel metal2 s 18510 27520 18566 28000 6 chany_top_out[4]
port 125 nsew default tristate
rlabel metal2 s 19062 27520 19118 28000 6 chany_top_out[5]
port 126 nsew default tristate
rlabel metal2 s 19614 27520 19670 28000 6 chany_top_out[6]
port 127 nsew default tristate
rlabel metal2 s 20258 27520 20314 28000 6 chany_top_out[7]
port 128 nsew default tristate
rlabel metal2 s 20810 27520 20866 28000 6 chany_top_out[8]
port 129 nsew default tristate
rlabel metal2 s 21362 27520 21418 28000 6 chany_top_out[9]
port 130 nsew default tristate
rlabel metal3 s 0 23536 480 23656 6 left_top_grid_pin_42_
port 131 nsew default input
rlabel metal3 s 0 24080 480 24200 6 left_top_grid_pin_43_
port 132 nsew default input
rlabel metal3 s 0 24760 480 24880 6 left_top_grid_pin_44_
port 133 nsew default input
rlabel metal3 s 0 25304 480 25424 6 left_top_grid_pin_45_
port 134 nsew default input
rlabel metal3 s 0 25848 480 25968 6 left_top_grid_pin_46_
port 135 nsew default input
rlabel metal3 s 0 26528 480 26648 6 left_top_grid_pin_47_
port 136 nsew default input
rlabel metal3 s 0 27072 480 27192 6 left_top_grid_pin_48_
port 137 nsew default input
rlabel metal3 s 0 27616 480 27736 6 left_top_grid_pin_49_
port 138 nsew default input
rlabel metal3 s 27520 4632 28000 4752 6 prog_clk
port 139 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_34_
port 140 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_35_
port 141 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_36_
port 142 nsew default input
rlabel metal2 s 1950 27520 2006 28000 6 top_left_grid_pin_37_
port 143 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 top_left_grid_pin_38_
port 144 nsew default input
rlabel metal2 s 3146 27520 3202 28000 6 top_left_grid_pin_39_
port 145 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 top_left_grid_pin_40_
port 146 nsew default input
rlabel metal2 s 4250 27520 4306 28000 6 top_left_grid_pin_41_
port 147 nsew default input
rlabel metal2 s 27618 27520 27674 28000 6 top_right_grid_pin_1_
port 148 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 149 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 150 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
