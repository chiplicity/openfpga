magic
tech sky130A
magscale 1 2
timestamp 1608761905
<< checkpaint >>
rect -1260 -1260 24060 24060
<< locali >>
rect 18705 19907 18739 20009
rect 18647 19873 18739 19907
rect 14381 19703 14415 19873
rect 19809 19703 19843 19873
rect 9413 18683 9447 18921
rect 12173 18207 12207 18377
rect 21741 18003 21775 19125
rect 11253 17527 11287 17697
rect 17785 17663 17819 17765
rect 9413 15895 9447 16065
rect 18337 15011 18371 15113
rect 18429 14875 18463 15113
rect 20085 14807 20119 15045
rect 12449 10523 12483 10761
rect 16129 10523 16163 10625
rect 18981 8347 19015 8449
rect 16681 5083 16715 5321
rect 10425 3451 10459 3621
rect 12909 2839 12943 3145
rect 17877 2839 17911 2941
<< viali >>
rect 12817 20009 12851 20043
rect 14197 20009 14231 20043
rect 14749 20009 14783 20043
rect 15669 20009 15703 20043
rect 16865 20009 16899 20043
rect 17417 20009 17451 20043
rect 18521 20009 18555 20043
rect 18705 20009 18739 20043
rect 19073 20009 19107 20043
rect 19625 20009 19659 20043
rect 12633 19873 12667 19907
rect 13461 19873 13495 19907
rect 14013 19873 14047 19907
rect 14381 19873 14415 19907
rect 14565 19873 14599 19907
rect 15485 19873 15519 19907
rect 16129 19873 16163 19907
rect 16681 19873 16715 19907
rect 17233 19873 17267 19907
rect 18337 19873 18371 19907
rect 18613 19873 18647 19907
rect 18889 19873 18923 19907
rect 19441 19873 19475 19907
rect 19809 19873 19843 19907
rect 19993 19873 20027 19907
rect 20545 19873 20579 19907
rect 13645 19737 13679 19771
rect 16313 19737 16347 19771
rect 14381 19669 14415 19703
rect 19809 19669 19843 19703
rect 20177 19669 20211 19703
rect 20729 19669 20763 19703
rect 19165 19465 19199 19499
rect 8677 19261 8711 19295
rect 10977 19261 11011 19295
rect 11805 19261 11839 19295
rect 12449 19261 12483 19295
rect 14105 19261 14139 19295
rect 14657 19261 14691 19295
rect 14933 19261 14967 19295
rect 15577 19261 15611 19295
rect 16497 19261 16531 19295
rect 17049 19261 17083 19295
rect 18061 19261 18095 19295
rect 18981 19261 19015 19295
rect 19533 19261 19567 19295
rect 20821 19261 20855 19295
rect 8944 19193 8978 19227
rect 12716 19193 12750 19227
rect 20361 19193 20395 19227
rect 10057 19125 10091 19159
rect 11161 19125 11195 19159
rect 11989 19125 12023 19159
rect 13829 19125 13863 19159
rect 14289 19125 14323 19159
rect 15761 19125 15795 19159
rect 16681 19125 16715 19159
rect 17233 19125 17267 19159
rect 18245 19125 18279 19159
rect 21005 19125 21039 19159
rect 21741 19125 21775 19159
rect 8953 18921 8987 18955
rect 9413 18921 9447 18955
rect 13369 18921 13403 18955
rect 14657 18921 14691 18955
rect 18061 18921 18095 18955
rect 9045 18717 9079 18751
rect 9137 18717 9171 18751
rect 13461 18853 13495 18887
rect 17233 18853 17267 18887
rect 18705 18853 18739 18887
rect 19901 18853 19935 18887
rect 9956 18785 9990 18819
rect 11601 18785 11635 18819
rect 14473 18785 14507 18819
rect 15301 18785 15335 18819
rect 15568 18785 15602 18819
rect 16957 18785 16991 18819
rect 17877 18785 17911 18819
rect 18429 18785 18463 18819
rect 19625 18785 19659 18819
rect 9689 18717 9723 18751
rect 11345 18717 11379 18751
rect 13645 18717 13679 18751
rect 14013 18717 14047 18751
rect 19165 18717 19199 18751
rect 9413 18649 9447 18683
rect 12725 18649 12759 18683
rect 8585 18581 8619 18615
rect 11069 18581 11103 18615
rect 13001 18581 13035 18615
rect 16681 18581 16715 18615
rect 9229 18377 9263 18411
rect 12173 18377 12207 18411
rect 15853 18377 15887 18411
rect 17601 18377 17635 18411
rect 9597 18309 9631 18343
rect 10057 18241 10091 18275
rect 10241 18241 10275 18275
rect 11161 18241 11195 18275
rect 12817 18241 12851 18275
rect 16681 18241 16715 18275
rect 18613 18241 18647 18275
rect 7113 18173 7147 18207
rect 7849 18173 7883 18207
rect 11069 18173 11103 18207
rect 11621 18173 11655 18207
rect 11897 18173 11931 18207
rect 12173 18173 12207 18207
rect 13084 18173 13118 18207
rect 14473 18173 14507 18207
rect 16589 18173 16623 18207
rect 17417 18173 17451 18207
rect 18429 18173 18463 18207
rect 19441 18173 19475 18207
rect 19993 18173 20027 18207
rect 20545 18173 20579 18207
rect 7389 18105 7423 18139
rect 8116 18105 8150 18139
rect 14718 18105 14752 18139
rect 9965 18037 9999 18071
rect 10609 18037 10643 18071
rect 10977 18037 11011 18071
rect 14197 18037 14231 18071
rect 16129 18037 16163 18071
rect 16497 18037 16531 18071
rect 18061 18037 18095 18071
rect 18521 18037 18555 18071
rect 19625 18037 19659 18071
rect 20177 18037 20211 18071
rect 20729 18037 20763 18071
rect 21741 17969 21775 18003
rect 7389 17833 7423 17867
rect 7481 17833 7515 17867
rect 9873 17833 9907 17867
rect 10701 17833 10735 17867
rect 10793 17833 10827 17867
rect 13093 17833 13127 17867
rect 13185 17833 13219 17867
rect 14105 17833 14139 17867
rect 14197 17833 14231 17867
rect 14749 17833 14783 17867
rect 8677 17765 8711 17799
rect 16580 17765 16614 17799
rect 17785 17765 17819 17799
rect 18236 17765 18270 17799
rect 19993 17765 20027 17799
rect 8585 17697 8619 17731
rect 11253 17697 11287 17731
rect 11345 17697 11379 17731
rect 11621 17697 11655 17731
rect 15669 17697 15703 17731
rect 15761 17697 15795 17731
rect 7665 17629 7699 17663
rect 8769 17629 8803 17663
rect 10977 17629 11011 17663
rect 7021 17561 7055 17595
rect 19717 17697 19751 17731
rect 13277 17629 13311 17663
rect 14289 17629 14323 17663
rect 15853 17629 15887 17663
rect 16313 17629 16347 17663
rect 17785 17629 17819 17663
rect 17969 17629 18003 17663
rect 17693 17561 17727 17595
rect 8217 17493 8251 17527
rect 10333 17493 10367 17527
rect 11253 17493 11287 17527
rect 12725 17493 12759 17527
rect 13737 17493 13771 17527
rect 15301 17493 15335 17527
rect 19349 17493 19383 17527
rect 8861 17289 8895 17323
rect 16957 17289 16991 17323
rect 13093 17221 13127 17255
rect 15761 17221 15795 17255
rect 7481 17153 7515 17187
rect 9689 17153 9723 17187
rect 10885 17153 10919 17187
rect 11897 17153 11931 17187
rect 13553 17153 13587 17187
rect 13737 17153 13771 17187
rect 16221 17153 16255 17187
rect 16405 17153 16439 17187
rect 17601 17153 17635 17187
rect 18705 17153 18739 17187
rect 19993 17153 20027 17187
rect 20821 17153 20855 17187
rect 9505 17085 9539 17119
rect 14105 17085 14139 17119
rect 15209 17085 15243 17119
rect 16129 17085 16163 17119
rect 17325 17085 17359 17119
rect 18429 17085 18463 17119
rect 19257 17085 19291 17119
rect 19809 17085 19843 17119
rect 20545 17085 20579 17119
rect 7748 17017 7782 17051
rect 10701 17017 10735 17051
rect 11713 17017 11747 17051
rect 12541 17017 12575 17051
rect 13461 17017 13495 17051
rect 14381 17017 14415 17051
rect 9137 16949 9171 16983
rect 9597 16949 9631 16983
rect 10241 16949 10275 16983
rect 10609 16949 10643 16983
rect 11345 16949 11379 16983
rect 11805 16949 11839 16983
rect 15393 16949 15427 16983
rect 17417 16949 17451 16983
rect 18061 16949 18095 16983
rect 18521 16949 18555 16983
rect 19441 16949 19475 16983
rect 14105 16745 14139 16779
rect 15761 16745 15795 16779
rect 17141 16745 17175 16779
rect 8953 16677 8987 16711
rect 10692 16677 10726 16711
rect 7021 16609 7055 16643
rect 7288 16609 7322 16643
rect 8677 16609 8711 16643
rect 9689 16609 9723 16643
rect 10425 16609 10459 16643
rect 12173 16609 12207 16643
rect 12440 16609 12474 16643
rect 14473 16609 14507 16643
rect 15669 16609 15703 16643
rect 16405 16609 16439 16643
rect 16957 16609 16991 16643
rect 17776 16609 17810 16643
rect 19533 16609 19567 16643
rect 20269 16609 20303 16643
rect 9965 16541 9999 16575
rect 14565 16541 14599 16575
rect 14749 16541 14783 16575
rect 15853 16541 15887 16575
rect 17509 16541 17543 16575
rect 19625 16541 19659 16575
rect 19717 16541 19751 16575
rect 8401 16405 8435 16439
rect 11805 16405 11839 16439
rect 13553 16405 13587 16439
rect 15301 16405 15335 16439
rect 16589 16405 16623 16439
rect 18889 16405 18923 16439
rect 19165 16405 19199 16439
rect 20453 16405 20487 16439
rect 8493 16201 8527 16235
rect 15577 16201 15611 16235
rect 19625 16201 19659 16235
rect 6837 16065 6871 16099
rect 9045 16065 9079 16099
rect 9413 16065 9447 16099
rect 11621 16065 11655 16099
rect 11805 16065 11839 16099
rect 13553 16065 13587 16099
rect 16221 16065 16255 16099
rect 17233 16065 17267 16099
rect 19165 16065 19199 16099
rect 20177 16065 20211 16099
rect 20821 16065 20855 16099
rect 8953 15997 8987 16031
rect 7104 15929 7138 15963
rect 9505 15997 9539 16031
rect 13277 15997 13311 16031
rect 13369 15997 13403 16031
rect 13921 15997 13955 16031
rect 16037 15997 16071 16031
rect 17785 15997 17819 16031
rect 18061 15997 18095 16031
rect 19073 15997 19107 16031
rect 19993 15997 20027 16031
rect 20637 15997 20671 16031
rect 9772 15929 9806 15963
rect 11529 15929 11563 15963
rect 14188 15929 14222 15963
rect 15945 15929 15979 15963
rect 17049 15929 17083 15963
rect 20085 15929 20119 15963
rect 8217 15861 8251 15895
rect 8861 15861 8895 15895
rect 9413 15861 9447 15895
rect 10885 15861 10919 15895
rect 11161 15861 11195 15895
rect 12909 15861 12943 15895
rect 15301 15861 15335 15895
rect 16589 15861 16623 15895
rect 16957 15861 16991 15895
rect 17601 15861 17635 15895
rect 18245 15861 18279 15895
rect 18613 15861 18647 15895
rect 18981 15861 19015 15895
rect 7757 15657 7791 15691
rect 8125 15657 8159 15691
rect 10057 15657 10091 15691
rect 10701 15657 10735 15691
rect 11805 15657 11839 15691
rect 15761 15657 15795 15691
rect 17785 15657 17819 15691
rect 19441 15657 19475 15691
rect 19717 15657 19751 15691
rect 10793 15589 10827 15623
rect 11713 15589 11747 15623
rect 13820 15589 13854 15623
rect 15853 15589 15887 15623
rect 18328 15589 18362 15623
rect 6377 15521 6411 15555
rect 6644 15521 6678 15555
rect 8953 15521 8987 15555
rect 9045 15521 9079 15555
rect 10241 15521 10275 15555
rect 12725 15521 12759 15555
rect 16672 15521 16706 15555
rect 20085 15521 20119 15555
rect 9137 15453 9171 15487
rect 10977 15453 11011 15487
rect 11989 15453 12023 15487
rect 12817 15453 12851 15487
rect 13001 15453 13035 15487
rect 13553 15453 13587 15487
rect 16037 15453 16071 15487
rect 16405 15453 16439 15487
rect 18061 15453 18095 15487
rect 20177 15453 20211 15487
rect 20269 15453 20303 15487
rect 8585 15317 8619 15351
rect 10333 15317 10367 15351
rect 11345 15317 11379 15351
rect 12357 15317 12391 15351
rect 14933 15317 14967 15351
rect 15393 15317 15427 15351
rect 9321 15113 9355 15147
rect 10057 15113 10091 15147
rect 12909 15113 12943 15147
rect 18337 15113 18371 15147
rect 7297 14977 7331 15011
rect 7481 14977 7515 15011
rect 10517 14977 10551 15011
rect 10609 14977 10643 15011
rect 11621 14977 11655 15011
rect 13461 14977 13495 15011
rect 16129 14977 16163 15011
rect 18061 14977 18095 15011
rect 18337 14977 18371 15011
rect 18429 15113 18463 15147
rect 20177 15113 20211 15147
rect 7205 14909 7239 14943
rect 7941 14909 7975 14943
rect 10425 14909 10459 14943
rect 13921 14909 13955 14943
rect 15945 14909 15979 14943
rect 16037 14909 16071 14943
rect 17233 14909 17267 14943
rect 17417 14909 17451 14943
rect 19901 15045 19935 15079
rect 20085 15045 20119 15079
rect 18521 14909 18555 14943
rect 8208 14841 8242 14875
rect 9597 14841 9631 14875
rect 11529 14841 11563 14875
rect 14188 14841 14222 14875
rect 18429 14841 18463 14875
rect 18788 14841 18822 14875
rect 20729 14977 20763 15011
rect 20545 14909 20579 14943
rect 6837 14773 6871 14807
rect 11069 14773 11103 14807
rect 11437 14773 11471 14807
rect 13277 14773 13311 14807
rect 13369 14773 13403 14807
rect 15301 14773 15335 14807
rect 15577 14773 15611 14807
rect 16589 14773 16623 14807
rect 17049 14773 17083 14807
rect 17601 14773 17635 14807
rect 20085 14773 20119 14807
rect 20637 14773 20671 14807
rect 9689 14569 9723 14603
rect 10057 14569 10091 14603
rect 12541 14569 12575 14603
rect 14197 14569 14231 14603
rect 15669 14569 15703 14603
rect 7288 14501 7322 14535
rect 9137 14501 9171 14535
rect 10149 14501 10183 14535
rect 11428 14501 11462 14535
rect 13084 14501 13118 14535
rect 15761 14501 15795 14535
rect 17509 14501 17543 14535
rect 19248 14501 19282 14535
rect 7021 14433 7055 14467
rect 8861 14433 8895 14467
rect 11069 14433 11103 14467
rect 12817 14433 12851 14467
rect 14473 14433 14507 14467
rect 16313 14433 16347 14467
rect 16589 14433 16623 14467
rect 17601 14433 17635 14467
rect 18429 14433 18463 14467
rect 18981 14433 19015 14467
rect 10241 14365 10275 14399
rect 11161 14365 11195 14399
rect 14749 14365 14783 14399
rect 15853 14365 15887 14399
rect 17785 14365 17819 14399
rect 20913 14365 20947 14399
rect 8401 14297 8435 14331
rect 15301 14297 15335 14331
rect 18613 14297 18647 14331
rect 10885 14229 10919 14263
rect 17141 14229 17175 14263
rect 20361 14229 20395 14263
rect 8217 14025 8251 14059
rect 11345 14025 11379 14059
rect 14105 14025 14139 14059
rect 19809 14025 19843 14059
rect 21005 13957 21039 13991
rect 8861 13889 8895 13923
rect 9229 13889 9263 13923
rect 11805 13889 11839 13923
rect 11989 13889 12023 13923
rect 13093 13889 13127 13923
rect 14749 13889 14783 13923
rect 15669 13889 15703 13923
rect 18613 13889 18647 13923
rect 20361 13889 20395 13923
rect 8585 13821 8619 13855
rect 9496 13821 9530 13855
rect 14565 13821 14599 13855
rect 15577 13821 15611 13855
rect 16129 13821 16163 13855
rect 16396 13821 16430 13855
rect 19073 13821 19107 13855
rect 19349 13821 19383 13855
rect 20821 13821 20855 13855
rect 15485 13753 15519 13787
rect 20177 13753 20211 13787
rect 8677 13685 8711 13719
rect 10609 13685 10643 13719
rect 11713 13685 11747 13719
rect 12449 13685 12483 13719
rect 12817 13685 12851 13719
rect 12909 13685 12943 13719
rect 13645 13685 13679 13719
rect 14473 13685 14507 13719
rect 15117 13685 15151 13719
rect 17509 13685 17543 13719
rect 18061 13685 18095 13719
rect 18429 13685 18463 13719
rect 18521 13685 18555 13719
rect 20269 13685 20303 13719
rect 9321 13481 9355 13515
rect 9781 13481 9815 13515
rect 12449 13481 12483 13515
rect 13461 13481 13495 13515
rect 13829 13481 13863 13515
rect 15669 13481 15703 13515
rect 17877 13481 17911 13515
rect 18153 13481 18187 13515
rect 19625 13481 19659 13515
rect 20453 13481 20487 13515
rect 11989 13413 12023 13447
rect 12909 13413 12943 13447
rect 14749 13413 14783 13447
rect 9505 13345 9539 13379
rect 10149 13345 10183 13379
rect 11713 13345 11747 13379
rect 12817 13345 12851 13379
rect 13921 13345 13955 13379
rect 14473 13345 14507 13379
rect 15761 13345 15795 13379
rect 16497 13345 16531 13379
rect 16764 13345 16798 13379
rect 18521 13345 18555 13379
rect 19533 13345 19567 13379
rect 20269 13345 20303 13379
rect 10241 13277 10275 13311
rect 10333 13277 10367 13311
rect 13093 13277 13127 13311
rect 14105 13277 14139 13311
rect 15853 13277 15887 13311
rect 18613 13277 18647 13311
rect 18705 13277 18739 13311
rect 19717 13277 19751 13311
rect 15301 13141 15335 13175
rect 19165 13141 19199 13175
rect 12081 12937 12115 12971
rect 12449 12937 12483 12971
rect 16497 12937 16531 12971
rect 18061 12937 18095 12971
rect 20453 12937 20487 12971
rect 20913 12937 20947 12971
rect 16773 12869 16807 12903
rect 9321 12801 9355 12835
rect 11529 12801 11563 12835
rect 13093 12801 13127 12835
rect 13461 12801 13495 12835
rect 15117 12801 15151 12835
rect 17233 12801 17267 12835
rect 17417 12801 17451 12835
rect 18705 12801 18739 12835
rect 9588 12733 9622 12767
rect 12265 12733 12299 12767
rect 12909 12733 12943 12767
rect 15384 12733 15418 12767
rect 17141 12733 17175 12767
rect 19073 12733 19107 12767
rect 20729 12733 20763 12767
rect 11345 12665 11379 12699
rect 13728 12665 13762 12699
rect 18521 12665 18555 12699
rect 19340 12665 19374 12699
rect 10701 12597 10735 12631
rect 10977 12597 11011 12631
rect 11437 12597 11471 12631
rect 12817 12597 12851 12631
rect 14841 12597 14875 12631
rect 18429 12597 18463 12631
rect 10057 12393 10091 12427
rect 10517 12393 10551 12427
rect 14749 12393 14783 12427
rect 15485 12393 15519 12427
rect 16129 12393 16163 12427
rect 17233 12393 17267 12427
rect 20453 12393 20487 12427
rect 10425 12257 10459 12291
rect 11704 12257 11738 12291
rect 13360 12257 13394 12291
rect 15669 12257 15703 12291
rect 17141 12257 17175 12291
rect 17785 12257 17819 12291
rect 18613 12257 18647 12291
rect 18880 12257 18914 12291
rect 20269 12257 20303 12291
rect 10609 12189 10643 12223
rect 11437 12189 11471 12223
rect 13093 12189 13127 12223
rect 16221 12189 16255 12223
rect 16405 12189 16439 12223
rect 17417 12189 17451 12223
rect 18061 12189 18095 12223
rect 12817 12121 12851 12155
rect 14473 12121 14507 12155
rect 15761 12053 15795 12087
rect 16773 12053 16807 12087
rect 19993 12053 20027 12087
rect 10425 11849 10459 11883
rect 14381 11849 14415 11883
rect 18613 11849 18647 11883
rect 8769 11713 8803 11747
rect 10977 11713 11011 11747
rect 13185 11713 13219 11747
rect 14105 11713 14139 11747
rect 14933 11713 14967 11747
rect 15761 11713 15795 11747
rect 17417 11713 17451 11747
rect 19257 11713 19291 11747
rect 20177 11713 20211 11747
rect 20821 11713 20855 11747
rect 9036 11645 9070 11679
rect 14841 11645 14875 11679
rect 16028 11645 16062 11679
rect 20637 11645 20671 11679
rect 10793 11577 10827 11611
rect 11437 11577 11471 11611
rect 14749 11577 14783 11611
rect 18153 11577 18187 11611
rect 19993 11577 20027 11611
rect 10149 11509 10183 11543
rect 10885 11509 10919 11543
rect 12541 11509 12575 11543
rect 12909 11509 12943 11543
rect 13001 11509 13035 11543
rect 13553 11509 13587 11543
rect 13921 11509 13955 11543
rect 14013 11509 14047 11543
rect 17141 11509 17175 11543
rect 18981 11509 19015 11543
rect 19073 11509 19107 11543
rect 19625 11509 19659 11543
rect 20085 11509 20119 11543
rect 12265 11305 12299 11339
rect 15301 11305 15335 11339
rect 15669 11305 15703 11339
rect 20545 11305 20579 11339
rect 8208 11237 8242 11271
rect 9965 11237 9999 11271
rect 16856 11237 16890 11271
rect 18705 11237 18739 11271
rect 7941 11169 7975 11203
rect 9689 11169 9723 11203
rect 10885 11169 10919 11203
rect 11152 11169 11186 11203
rect 13001 11169 13035 11203
rect 18429 11169 18463 11203
rect 19432 11169 19466 11203
rect 15761 11101 15795 11135
rect 15853 11101 15887 11135
rect 16589 11101 16623 11135
rect 19165 11101 19199 11135
rect 14289 11033 14323 11067
rect 9321 10965 9355 10999
rect 17969 10965 18003 10999
rect 12449 10761 12483 10795
rect 13369 10761 13403 10795
rect 14473 10761 14507 10795
rect 15301 10761 15335 10795
rect 18061 10761 18095 10795
rect 10425 10625 10459 10659
rect 11437 10625 11471 10659
rect 8217 10557 8251 10591
rect 8484 10557 8518 10591
rect 10333 10557 10367 10591
rect 12081 10557 12115 10591
rect 12541 10693 12575 10727
rect 13093 10625 13127 10659
rect 13921 10625 13955 10659
rect 15025 10625 15059 10659
rect 15945 10625 15979 10659
rect 16129 10625 16163 10659
rect 18613 10625 18647 10659
rect 13737 10557 13771 10591
rect 14841 10557 14875 10591
rect 15669 10557 15703 10591
rect 10241 10489 10275 10523
rect 11253 10489 11287 10523
rect 12449 10489 12483 10523
rect 16313 10557 16347 10591
rect 16580 10557 16614 10591
rect 19717 10557 19751 10591
rect 16129 10489 16163 10523
rect 18429 10489 18463 10523
rect 19073 10489 19107 10523
rect 19984 10489 20018 10523
rect 9597 10421 9631 10455
rect 9873 10421 9907 10455
rect 10885 10421 10919 10455
rect 11345 10421 11379 10455
rect 12909 10421 12943 10455
rect 13001 10421 13035 10455
rect 13829 10421 13863 10455
rect 14933 10421 14967 10455
rect 15761 10421 15795 10455
rect 17693 10421 17727 10455
rect 18521 10421 18555 10455
rect 21097 10421 21131 10455
rect 9045 10217 9079 10251
rect 11989 10217 12023 10251
rect 13185 10217 13219 10251
rect 14565 10217 14599 10251
rect 15301 10217 15335 10251
rect 16865 10217 16899 10251
rect 18245 10217 18279 10251
rect 10876 10149 10910 10183
rect 13645 10149 13679 10183
rect 19625 10149 19659 10183
rect 8953 10081 8987 10115
rect 9689 10081 9723 10115
rect 13553 10081 13587 10115
rect 14657 10081 14691 10115
rect 15669 10081 15703 10115
rect 17233 10081 17267 10115
rect 9229 10013 9263 10047
rect 10609 10013 10643 10047
rect 13737 10013 13771 10047
rect 14749 10013 14783 10047
rect 15761 10013 15795 10047
rect 15945 10013 15979 10047
rect 17325 10013 17359 10047
rect 17509 10013 17543 10047
rect 18337 10013 18371 10047
rect 18521 10013 18555 10047
rect 19717 10013 19751 10047
rect 19901 10013 19935 10047
rect 8585 9945 8619 9979
rect 17877 9945 17911 9979
rect 14197 9877 14231 9911
rect 19257 9877 19291 9911
rect 11345 9673 11379 9707
rect 18061 9673 18095 9707
rect 16037 9605 16071 9639
rect 9965 9537 9999 9571
rect 11897 9537 11931 9571
rect 12541 9537 12575 9571
rect 14657 9537 14691 9571
rect 16865 9537 16899 9571
rect 18613 9537 18647 9571
rect 20821 9537 20855 9571
rect 7757 9469 7791 9503
rect 8024 9469 8058 9503
rect 9873 9469 9907 9503
rect 11621 9469 11655 9503
rect 12808 9469 12842 9503
rect 19165 9469 19199 9503
rect 10232 9401 10266 9435
rect 14924 9401 14958 9435
rect 16681 9401 16715 9435
rect 16773 9401 16807 9435
rect 18429 9401 18463 9435
rect 19432 9401 19466 9435
rect 9137 9333 9171 9367
rect 9689 9333 9723 9367
rect 13921 9333 13955 9367
rect 14197 9333 14231 9367
rect 16313 9333 16347 9367
rect 18521 9333 18555 9367
rect 20545 9333 20579 9367
rect 9873 9129 9907 9163
rect 11345 9129 11379 9163
rect 11897 9129 11931 9163
rect 12265 9129 12299 9163
rect 14013 9129 14047 9163
rect 15301 9129 15335 9163
rect 18889 9129 18923 9163
rect 20545 9129 20579 9163
rect 9045 9061 9079 9095
rect 10241 9061 10275 9095
rect 12909 9061 12943 9095
rect 13921 9061 13955 9095
rect 17754 9061 17788 9095
rect 19410 9061 19444 9095
rect 8953 8993 8987 9027
rect 11253 8993 11287 9027
rect 12357 8993 12391 9027
rect 14749 8993 14783 9027
rect 15669 8993 15703 9027
rect 16773 8993 16807 9027
rect 19165 8993 19199 9027
rect 9137 8925 9171 8959
rect 10333 8925 10367 8959
rect 10425 8925 10459 8959
rect 11437 8925 11471 8959
rect 12449 8925 12483 8959
rect 14105 8925 14139 8959
rect 15761 8925 15795 8959
rect 15945 8925 15979 8959
rect 17509 8925 17543 8959
rect 10885 8857 10919 8891
rect 14565 8857 14599 8891
rect 8585 8789 8619 8823
rect 13553 8789 13587 8823
rect 16589 8789 16623 8823
rect 11253 8585 11287 8619
rect 15117 8585 15151 8619
rect 17325 8585 17359 8619
rect 18061 8585 18095 8619
rect 19073 8585 19107 8619
rect 12633 8517 12667 8551
rect 11713 8449 11747 8483
rect 13093 8449 13127 8483
rect 15945 8449 15979 8483
rect 18521 8449 18555 8483
rect 18705 8449 18739 8483
rect 18981 8449 19015 8483
rect 19625 8449 19659 8483
rect 20545 8449 20579 8483
rect 20637 8449 20671 8483
rect 8033 8381 8067 8415
rect 8300 8381 8334 8415
rect 9873 8381 9907 8415
rect 11529 8381 11563 8415
rect 12817 8381 12851 8415
rect 13360 8381 13394 8415
rect 15301 8381 15335 8415
rect 18429 8381 18463 8415
rect 19441 8381 19475 8415
rect 10140 8313 10174 8347
rect 16212 8313 16246 8347
rect 18981 8313 19015 8347
rect 19533 8313 19567 8347
rect 9413 8245 9447 8279
rect 14473 8245 14507 8279
rect 20085 8245 20119 8279
rect 20453 8245 20487 8279
rect 9045 8041 9079 8075
rect 10149 8041 10183 8075
rect 14289 8041 14323 8075
rect 18061 8041 18095 8075
rect 20913 8041 20947 8075
rect 10609 7973 10643 8007
rect 13185 7973 13219 8007
rect 8953 7905 8987 7939
rect 9689 7905 9723 7939
rect 10517 7905 10551 7939
rect 11428 7905 11462 7939
rect 14197 7905 14231 7939
rect 15577 7905 15611 7939
rect 15844 7905 15878 7939
rect 17233 7905 17267 7939
rect 18153 7905 18187 7939
rect 19993 7905 20027 7939
rect 9229 7837 9263 7871
rect 10793 7837 10827 7871
rect 11161 7837 11195 7871
rect 13277 7837 13311 7871
rect 13461 7837 13495 7871
rect 14473 7837 14507 7871
rect 18245 7837 18279 7871
rect 20085 7837 20119 7871
rect 20269 7837 20303 7871
rect 8585 7769 8619 7803
rect 12541 7701 12575 7735
rect 12817 7701 12851 7735
rect 13829 7701 13863 7735
rect 16957 7701 16991 7735
rect 17693 7701 17727 7735
rect 19625 7701 19659 7735
rect 8217 7497 8251 7531
rect 15025 7497 15059 7531
rect 10609 7429 10643 7463
rect 8861 7361 8895 7395
rect 11989 7361 12023 7395
rect 13093 7361 13127 7395
rect 13185 7361 13219 7395
rect 15945 7361 15979 7395
rect 9229 7293 9263 7327
rect 9485 7293 9519 7327
rect 13001 7293 13035 7327
rect 13645 7293 13679 7327
rect 13912 7293 13946 7327
rect 15669 7293 15703 7327
rect 16313 7293 16347 7327
rect 18797 7293 18831 7327
rect 20453 7293 20487 7327
rect 11713 7225 11747 7259
rect 16580 7225 16614 7259
rect 19064 7225 19098 7259
rect 8585 7157 8619 7191
rect 8677 7157 8711 7191
rect 11345 7157 11379 7191
rect 11805 7157 11839 7191
rect 12633 7157 12667 7191
rect 15301 7157 15335 7191
rect 15761 7157 15795 7191
rect 17693 7157 17727 7191
rect 20177 7157 20211 7191
rect 20637 7157 20671 7191
rect 9321 6953 9355 6987
rect 9689 6953 9723 6987
rect 16221 6953 16255 6987
rect 16681 6953 16715 6987
rect 17601 6953 17635 6987
rect 19165 6953 19199 6987
rect 10057 6885 10091 6919
rect 11520 6885 11554 6919
rect 14197 6885 14231 6919
rect 16589 6885 16623 6919
rect 20177 6885 20211 6919
rect 8208 6817 8242 6851
rect 10885 6817 10919 6851
rect 18245 6817 18279 6851
rect 19257 6817 19291 6851
rect 20269 6817 20303 6851
rect 7941 6749 7975 6783
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 11253 6749 11287 6783
rect 13369 6749 13403 6783
rect 14289 6749 14323 6783
rect 14473 6749 14507 6783
rect 16865 6749 16899 6783
rect 17693 6749 17727 6783
rect 17877 6749 17911 6783
rect 19441 6749 19475 6783
rect 20361 6749 20395 6783
rect 18429 6681 18463 6715
rect 10701 6613 10735 6647
rect 12633 6613 12667 6647
rect 13829 6613 13863 6647
rect 17233 6613 17267 6647
rect 18797 6613 18831 6647
rect 19809 6613 19843 6647
rect 9137 6409 9171 6443
rect 10149 6409 10183 6443
rect 11161 6409 11195 6443
rect 13277 6409 13311 6443
rect 15853 6409 15887 6443
rect 18153 6409 18187 6443
rect 20545 6409 20579 6443
rect 8861 6341 8895 6375
rect 14841 6341 14875 6375
rect 7481 6273 7515 6307
rect 9689 6273 9723 6307
rect 10793 6273 10827 6307
rect 11713 6273 11747 6307
rect 13829 6273 13863 6307
rect 15301 6273 15335 6307
rect 15393 6273 15427 6307
rect 16497 6273 16531 6307
rect 17325 6273 17359 6307
rect 17509 6273 17543 6307
rect 18797 6273 18831 6307
rect 7748 6205 7782 6239
rect 10609 6205 10643 6239
rect 11529 6205 11563 6239
rect 16221 6205 16255 6239
rect 17233 6205 17267 6239
rect 19165 6205 19199 6239
rect 20821 6205 20855 6239
rect 10517 6137 10551 6171
rect 13645 6137 13679 6171
rect 13737 6137 13771 6171
rect 15209 6137 15243 6171
rect 18521 6137 18555 6171
rect 19410 6137 19444 6171
rect 9505 6069 9539 6103
rect 9597 6069 9631 6103
rect 11621 6069 11655 6103
rect 12449 6069 12483 6103
rect 16313 6069 16347 6103
rect 16865 6069 16899 6103
rect 18613 6069 18647 6103
rect 21005 6069 21039 6103
rect 7665 5865 7699 5899
rect 9137 5865 9171 5899
rect 9689 5865 9723 5899
rect 10057 5865 10091 5899
rect 13921 5865 13955 5899
rect 15669 5865 15703 5899
rect 15761 5865 15795 5899
rect 16773 5865 16807 5899
rect 18521 5865 18555 5899
rect 6530 5797 6564 5831
rect 13001 5797 13035 5831
rect 14749 5797 14783 5831
rect 19248 5797 19282 5831
rect 6285 5729 6319 5763
rect 11152 5729 11186 5763
rect 12909 5729 12943 5763
rect 16497 5729 16531 5763
rect 16589 5729 16623 5763
rect 17408 5729 17442 5763
rect 10149 5661 10183 5695
rect 10333 5661 10367 5695
rect 10885 5661 10919 5695
rect 13093 5661 13127 5695
rect 14013 5661 14047 5695
rect 14105 5661 14139 5695
rect 15945 5661 15979 5695
rect 17141 5661 17175 5695
rect 18981 5661 19015 5695
rect 12265 5525 12299 5559
rect 12541 5525 12575 5559
rect 13553 5525 13587 5559
rect 15301 5525 15335 5559
rect 16313 5525 16347 5559
rect 20361 5525 20395 5559
rect 16681 5321 16715 5355
rect 19625 5321 19659 5355
rect 11989 5185 12023 5219
rect 12909 5185 12943 5219
rect 13093 5185 13127 5219
rect 13461 5185 13495 5219
rect 11805 5117 11839 5151
rect 12817 5117 12851 5151
rect 15117 5117 15151 5151
rect 15384 5117 15418 5151
rect 17325 5185 17359 5219
rect 18245 5185 18279 5219
rect 20453 5185 20487 5219
rect 20913 5185 20947 5219
rect 17141 5117 17175 5151
rect 20269 5117 20303 5151
rect 11713 5049 11747 5083
rect 13728 5049 13762 5083
rect 16681 5049 16715 5083
rect 18512 5049 18546 5083
rect 20361 5049 20395 5083
rect 11345 4981 11379 5015
rect 12449 4981 12483 5015
rect 14841 4981 14875 5015
rect 16497 4981 16531 5015
rect 16773 4981 16807 5015
rect 17233 4981 17267 5015
rect 19901 4981 19935 5015
rect 14105 4777 14139 4811
rect 18705 4777 18739 4811
rect 15936 4709 15970 4743
rect 17570 4709 17604 4743
rect 20177 4709 20211 4743
rect 11989 4641 12023 4675
rect 12256 4641 12290 4675
rect 14013 4641 14047 4675
rect 14657 4641 14691 4675
rect 15669 4641 15703 4675
rect 17325 4641 17359 4675
rect 18981 4641 19015 4675
rect 14197 4573 14231 4607
rect 20269 4573 20303 4607
rect 20453 4573 20487 4607
rect 20913 4573 20947 4607
rect 13369 4505 13403 4539
rect 17049 4505 17083 4539
rect 19165 4505 19199 4539
rect 13645 4437 13679 4471
rect 14841 4437 14875 4471
rect 19809 4437 19843 4471
rect 12909 4097 12943 4131
rect 13001 4097 13035 4131
rect 15669 4097 15703 4131
rect 15853 4097 15887 4131
rect 16681 4097 16715 4131
rect 16773 4097 16807 4131
rect 19257 4097 19291 4131
rect 20085 4097 20119 4131
rect 20177 4097 20211 4131
rect 9045 4029 9079 4063
rect 11621 4029 11655 4063
rect 12817 4029 12851 4063
rect 13461 4029 13495 4063
rect 14197 4029 14231 4063
rect 14749 4029 14783 4063
rect 15577 4029 15611 4063
rect 17233 4029 17267 4063
rect 18061 4029 18095 4063
rect 18981 4029 19015 4063
rect 19993 4029 20027 4063
rect 20637 4029 20671 4063
rect 9290 3961 9324 3995
rect 11897 3961 11931 3995
rect 13737 3961 13771 3995
rect 10425 3893 10459 3927
rect 12449 3893 12483 3927
rect 14381 3893 14415 3927
rect 15209 3893 15243 3927
rect 16221 3893 16255 3927
rect 16589 3893 16623 3927
rect 17417 3893 17451 3927
rect 18245 3893 18279 3927
rect 18613 3893 18647 3927
rect 19073 3893 19107 3927
rect 19625 3893 19659 3927
rect 20821 3893 20855 3927
rect 15853 3689 15887 3723
rect 15945 3689 15979 3723
rect 18153 3689 18187 3723
rect 19809 3689 19843 3723
rect 10425 3621 10459 3655
rect 13829 3621 13863 3655
rect 13921 3621 13955 3655
rect 18674 3621 18708 3655
rect 20913 3621 20947 3655
rect 10609 3553 10643 3587
rect 11336 3553 11370 3587
rect 12725 3553 12759 3587
rect 14473 3553 14507 3587
rect 16773 3553 16807 3587
rect 17040 3553 17074 3587
rect 18429 3553 18463 3587
rect 20085 3553 20119 3587
rect 11069 3485 11103 3519
rect 12909 3485 12943 3519
rect 14013 3485 14047 3519
rect 16037 3485 16071 3519
rect 10425 3417 10459 3451
rect 20269 3417 20303 3451
rect 12449 3349 12483 3383
rect 13461 3349 13495 3383
rect 14657 3349 14691 3383
rect 15485 3349 15519 3383
rect 12909 3145 12943 3179
rect 16037 3145 16071 3179
rect 17693 3145 17727 3179
rect 12633 3077 12667 3111
rect 10057 3009 10091 3043
rect 10324 2941 10358 2975
rect 11805 2941 11839 2975
rect 12449 2941 12483 2975
rect 14381 3077 14415 3111
rect 13001 3009 13035 3043
rect 18613 3009 18647 3043
rect 18889 3009 18923 3043
rect 19349 3009 19383 3043
rect 13257 2941 13291 2975
rect 14657 2941 14691 2975
rect 16313 2941 16347 2975
rect 16569 2941 16603 2975
rect 17877 2941 17911 2975
rect 18429 2941 18463 2975
rect 19073 2941 19107 2975
rect 19809 2941 19843 2975
rect 20545 2941 20579 2975
rect 14902 2873 14936 2907
rect 11437 2805 11471 2839
rect 11989 2805 12023 2839
rect 12909 2805 12943 2839
rect 20085 2873 20119 2907
rect 17877 2805 17911 2839
rect 18061 2805 18095 2839
rect 18521 2805 18555 2839
rect 20729 2805 20763 2839
rect 10701 2601 10735 2635
rect 10793 2601 10827 2635
rect 11713 2601 11747 2635
rect 14013 2601 14047 2635
rect 14381 2601 14415 2635
rect 14473 2601 14507 2635
rect 16497 2601 16531 2635
rect 16957 2601 16991 2635
rect 18337 2601 18371 2635
rect 19533 2601 19567 2635
rect 13185 2533 13219 2567
rect 9781 2465 9815 2499
rect 12909 2465 12943 2499
rect 15761 2465 15795 2499
rect 16865 2465 16899 2499
rect 17509 2465 17543 2499
rect 18705 2465 18739 2499
rect 19349 2465 19383 2499
rect 19901 2465 19935 2499
rect 20453 2465 20487 2499
rect 10885 2397 10919 2431
rect 11805 2397 11839 2431
rect 11897 2397 11931 2431
rect 14565 2397 14599 2431
rect 16037 2397 16071 2431
rect 17141 2397 17175 2431
rect 18797 2397 18831 2431
rect 18981 2397 19015 2431
rect 9965 2329 9999 2363
rect 11345 2329 11379 2363
rect 17693 2329 17727 2363
rect 20637 2329 20671 2363
rect 10333 2261 10367 2295
rect 20085 2261 20119 2295
<< metal1 >>
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 12805 20043 12863 20049
rect 12805 20009 12817 20043
rect 12851 20040 12863 20043
rect 13078 20040 13084 20052
rect 12851 20012 13084 20040
rect 12851 20009 12863 20012
rect 12805 20003 12863 20009
rect 13078 20000 13084 20012
rect 13136 20000 13142 20052
rect 14182 20040 14188 20052
rect 14143 20012 14188 20040
rect 14182 20000 14188 20012
rect 14240 20000 14246 20052
rect 14550 20000 14556 20052
rect 14608 20040 14614 20052
rect 14737 20043 14795 20049
rect 14737 20040 14749 20043
rect 14608 20012 14749 20040
rect 14608 20000 14614 20012
rect 14737 20009 14749 20012
rect 14783 20009 14795 20043
rect 14737 20003 14795 20009
rect 15657 20043 15715 20049
rect 15657 20009 15669 20043
rect 15703 20040 15715 20043
rect 15838 20040 15844 20052
rect 15703 20012 15844 20040
rect 15703 20009 15715 20012
rect 15657 20003 15715 20009
rect 15838 20000 15844 20012
rect 15896 20000 15902 20052
rect 16853 20043 16911 20049
rect 16853 20009 16865 20043
rect 16899 20009 16911 20043
rect 16853 20003 16911 20009
rect 17405 20043 17463 20049
rect 17405 20009 17417 20043
rect 17451 20040 17463 20043
rect 17494 20040 17500 20052
rect 17451 20012 17500 20040
rect 17451 20009 17463 20012
rect 17405 20003 17463 20009
rect 16868 19972 16896 20003
rect 17494 20000 17500 20012
rect 17552 20000 17558 20052
rect 18046 20000 18052 20052
rect 18104 20040 18110 20052
rect 18509 20043 18567 20049
rect 18509 20040 18521 20043
rect 18104 20012 18521 20040
rect 18104 20000 18110 20012
rect 18509 20009 18521 20012
rect 18555 20009 18567 20043
rect 18509 20003 18567 20009
rect 18693 20043 18751 20049
rect 18693 20009 18705 20043
rect 18739 20040 18751 20043
rect 18874 20040 18880 20052
rect 18739 20012 18880 20040
rect 18739 20009 18751 20012
rect 18693 20003 18751 20009
rect 18874 20000 18880 20012
rect 18932 20000 18938 20052
rect 19058 20040 19064 20052
rect 19019 20012 19064 20040
rect 19058 20000 19064 20012
rect 19116 20000 19122 20052
rect 19610 20040 19616 20052
rect 19571 20012 19616 20040
rect 19610 20000 19616 20012
rect 19668 20000 19674 20052
rect 19150 19972 19156 19984
rect 16868 19944 19156 19972
rect 19150 19932 19156 19944
rect 19208 19932 19214 19984
rect 12618 19904 12624 19916
rect 12579 19876 12624 19904
rect 12618 19864 12624 19876
rect 12676 19864 12682 19916
rect 13354 19864 13360 19916
rect 13412 19904 13418 19916
rect 13449 19907 13507 19913
rect 13449 19904 13461 19907
rect 13412 19876 13461 19904
rect 13412 19864 13418 19876
rect 13449 19873 13461 19876
rect 13495 19873 13507 19907
rect 13449 19867 13507 19873
rect 14001 19907 14059 19913
rect 14001 19873 14013 19907
rect 14047 19904 14059 19907
rect 14369 19907 14427 19913
rect 14369 19904 14381 19907
rect 14047 19876 14381 19904
rect 14047 19873 14059 19876
rect 14001 19867 14059 19873
rect 14369 19873 14381 19876
rect 14415 19873 14427 19907
rect 14369 19867 14427 19873
rect 14458 19864 14464 19916
rect 14516 19904 14522 19916
rect 14553 19907 14611 19913
rect 14553 19904 14565 19907
rect 14516 19876 14565 19904
rect 14516 19864 14522 19876
rect 14553 19873 14565 19876
rect 14599 19873 14611 19907
rect 15470 19904 15476 19916
rect 15431 19876 15476 19904
rect 14553 19867 14611 19873
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 16022 19864 16028 19916
rect 16080 19904 16086 19916
rect 16117 19907 16175 19913
rect 16117 19904 16129 19907
rect 16080 19876 16129 19904
rect 16080 19864 16086 19876
rect 16117 19873 16129 19876
rect 16163 19873 16175 19907
rect 16117 19867 16175 19873
rect 16574 19864 16580 19916
rect 16632 19904 16638 19916
rect 16669 19907 16727 19913
rect 16669 19904 16681 19907
rect 16632 19876 16681 19904
rect 16632 19864 16638 19876
rect 16669 19873 16681 19876
rect 16715 19873 16727 19907
rect 16669 19867 16727 19873
rect 16850 19864 16856 19916
rect 16908 19904 16914 19916
rect 17221 19907 17279 19913
rect 17221 19904 17233 19907
rect 16908 19876 17233 19904
rect 16908 19864 16914 19876
rect 17221 19873 17233 19876
rect 17267 19873 17279 19907
rect 17221 19867 17279 19873
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19904 18383 19907
rect 18601 19907 18659 19913
rect 18601 19904 18613 19907
rect 18371 19876 18613 19904
rect 18371 19873 18383 19876
rect 18325 19867 18383 19873
rect 18601 19873 18613 19876
rect 18647 19873 18659 19907
rect 18601 19867 18659 19873
rect 18690 19864 18696 19916
rect 18748 19904 18754 19916
rect 18877 19907 18935 19913
rect 18877 19904 18889 19907
rect 18748 19876 18889 19904
rect 18748 19864 18754 19876
rect 18877 19873 18889 19876
rect 18923 19873 18935 19907
rect 19426 19904 19432 19916
rect 19387 19876 19432 19904
rect 18877 19867 18935 19873
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 19797 19907 19855 19913
rect 19797 19873 19809 19907
rect 19843 19904 19855 19907
rect 19981 19907 20039 19913
rect 19981 19904 19993 19907
rect 19843 19876 19993 19904
rect 19843 19873 19855 19876
rect 19797 19867 19855 19873
rect 19981 19873 19993 19876
rect 20027 19873 20039 19907
rect 20530 19904 20536 19916
rect 20491 19876 20536 19904
rect 19981 19867 20039 19873
rect 20530 19864 20536 19876
rect 20588 19864 20594 19916
rect 20806 19836 20812 19848
rect 13648 19808 20812 19836
rect 13648 19777 13676 19808
rect 20806 19796 20812 19808
rect 20864 19796 20870 19848
rect 13633 19771 13691 19777
rect 13633 19737 13645 19771
rect 13679 19737 13691 19771
rect 13633 19731 13691 19737
rect 16301 19771 16359 19777
rect 16301 19737 16313 19771
rect 16347 19768 16359 19771
rect 19702 19768 19708 19780
rect 16347 19740 19708 19768
rect 16347 19737 16359 19740
rect 16301 19731 16359 19737
rect 19702 19728 19708 19740
rect 19760 19728 19766 19780
rect 14369 19703 14427 19709
rect 14369 19669 14381 19703
rect 14415 19700 14427 19703
rect 17126 19700 17132 19712
rect 14415 19672 17132 19700
rect 14415 19669 14427 19672
rect 14369 19663 14427 19669
rect 17126 19660 17132 19672
rect 17184 19660 17190 19712
rect 17954 19660 17960 19712
rect 18012 19700 18018 19712
rect 19797 19703 19855 19709
rect 19797 19700 19809 19703
rect 18012 19672 19809 19700
rect 18012 19660 18018 19672
rect 19797 19669 19809 19672
rect 19843 19669 19855 19703
rect 20162 19700 20168 19712
rect 20123 19672 20168 19700
rect 19797 19663 19855 19669
rect 20162 19660 20168 19672
rect 20220 19660 20226 19712
rect 20622 19660 20628 19712
rect 20680 19700 20686 19712
rect 20717 19703 20775 19709
rect 20717 19700 20729 19703
rect 20680 19672 20729 19700
rect 20680 19660 20686 19672
rect 20717 19669 20729 19672
rect 20763 19669 20775 19703
rect 20717 19663 20775 19669
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 9582 19496 9588 19508
rect 8680 19468 9588 19496
rect 7742 19252 7748 19304
rect 7800 19292 7806 19304
rect 8680 19301 8708 19468
rect 9582 19456 9588 19468
rect 9640 19456 9646 19508
rect 19150 19496 19156 19508
rect 12452 19468 13492 19496
rect 19111 19468 19156 19496
rect 12452 19428 12480 19468
rect 12360 19400 12480 19428
rect 8665 19295 8723 19301
rect 8665 19292 8677 19295
rect 7800 19264 8677 19292
rect 7800 19252 7806 19264
rect 8665 19261 8677 19264
rect 8711 19261 8723 19295
rect 10042 19292 10048 19304
rect 8665 19255 8723 19261
rect 8864 19264 10048 19292
rect 1394 19184 1400 19236
rect 1452 19224 1458 19236
rect 2682 19224 2688 19236
rect 1452 19196 2688 19224
rect 1452 19184 1458 19196
rect 2682 19184 2688 19196
rect 2740 19184 2746 19236
rect 8202 19184 8208 19236
rect 8260 19224 8266 19236
rect 8864 19224 8892 19264
rect 10042 19252 10048 19264
rect 10100 19252 10106 19304
rect 10965 19295 11023 19301
rect 10965 19261 10977 19295
rect 11011 19292 11023 19295
rect 11422 19292 11428 19304
rect 11011 19264 11428 19292
rect 11011 19261 11023 19264
rect 10965 19255 11023 19261
rect 11422 19252 11428 19264
rect 11480 19252 11486 19304
rect 11790 19292 11796 19304
rect 11751 19264 11796 19292
rect 11790 19252 11796 19264
rect 11848 19252 11854 19304
rect 8938 19233 8944 19236
rect 8260 19196 8892 19224
rect 8260 19184 8266 19196
rect 8932 19187 8944 19233
rect 8996 19224 9002 19236
rect 8996 19196 9032 19224
rect 8938 19184 8944 19187
rect 8996 19184 9002 19196
rect 9674 19184 9680 19236
rect 9732 19224 9738 19236
rect 9732 19196 10272 19224
rect 9732 19184 9738 19196
rect 2498 19116 2504 19168
rect 2556 19156 2562 19168
rect 9766 19156 9772 19168
rect 2556 19128 9772 19156
rect 2556 19116 2562 19128
rect 9766 19116 9772 19128
rect 9824 19116 9830 19168
rect 10045 19159 10103 19165
rect 10045 19125 10057 19159
rect 10091 19156 10103 19159
rect 10134 19156 10140 19168
rect 10091 19128 10140 19156
rect 10091 19125 10103 19128
rect 10045 19119 10103 19125
rect 10134 19116 10140 19128
rect 10192 19116 10198 19168
rect 10244 19156 10272 19196
rect 10318 19184 10324 19236
rect 10376 19224 10382 19236
rect 12360 19224 12388 19400
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19292 12495 19295
rect 13464 19292 13492 19468
rect 19150 19456 19156 19468
rect 19208 19456 19214 19508
rect 14016 19332 15700 19360
rect 14016 19292 14044 19332
rect 12483 19264 12848 19292
rect 13464 19264 14044 19292
rect 14093 19295 14151 19301
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 12820 19236 12848 19264
rect 14093 19261 14105 19295
rect 14139 19292 14151 19295
rect 14274 19292 14280 19304
rect 14139 19264 14280 19292
rect 14139 19261 14151 19264
rect 14093 19255 14151 19261
rect 14274 19252 14280 19264
rect 14332 19252 14338 19304
rect 14366 19252 14372 19304
rect 14424 19292 14430 19304
rect 14645 19295 14703 19301
rect 14645 19292 14657 19295
rect 14424 19264 14657 19292
rect 14424 19252 14430 19264
rect 14645 19261 14657 19264
rect 14691 19261 14703 19295
rect 14645 19255 14703 19261
rect 14921 19295 14979 19301
rect 14921 19261 14933 19295
rect 14967 19292 14979 19295
rect 15565 19295 15623 19301
rect 15565 19292 15577 19295
rect 14967 19264 15577 19292
rect 14967 19261 14979 19264
rect 14921 19255 14979 19261
rect 15565 19261 15577 19264
rect 15611 19261 15623 19295
rect 15672 19292 15700 19332
rect 16298 19292 16304 19304
rect 15672 19264 16304 19292
rect 15565 19255 15623 19261
rect 16298 19252 16304 19264
rect 16356 19252 16362 19304
rect 16482 19292 16488 19304
rect 16443 19264 16488 19292
rect 16482 19252 16488 19264
rect 16540 19252 16546 19304
rect 16758 19252 16764 19304
rect 16816 19292 16822 19304
rect 17037 19295 17095 19301
rect 17037 19292 17049 19295
rect 16816 19264 17049 19292
rect 16816 19252 16822 19264
rect 17037 19261 17049 19264
rect 17083 19261 17095 19295
rect 17037 19255 17095 19261
rect 17218 19252 17224 19304
rect 17276 19292 17282 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17276 19264 18061 19292
rect 17276 19252 17282 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18966 19292 18972 19304
rect 18927 19264 18972 19292
rect 18049 19255 18107 19261
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 19242 19252 19248 19304
rect 19300 19292 19306 19304
rect 19521 19295 19579 19301
rect 19521 19292 19533 19295
rect 19300 19264 19533 19292
rect 19300 19252 19306 19264
rect 19521 19261 19533 19264
rect 19567 19261 19579 19295
rect 20806 19292 20812 19304
rect 20767 19264 20812 19292
rect 19521 19255 19579 19261
rect 20806 19252 20812 19264
rect 20864 19252 20870 19304
rect 12710 19233 12716 19236
rect 12704 19224 12716 19233
rect 10376 19196 12388 19224
rect 12671 19196 12716 19224
rect 10376 19184 10382 19196
rect 12704 19187 12716 19196
rect 12710 19184 12716 19187
rect 12768 19184 12774 19236
rect 12802 19184 12808 19236
rect 12860 19184 12866 19236
rect 13630 19184 13636 19236
rect 13688 19224 13694 19236
rect 17862 19224 17868 19236
rect 13688 19196 14320 19224
rect 13688 19184 13694 19196
rect 10870 19156 10876 19168
rect 10244 19128 10876 19156
rect 10870 19116 10876 19128
rect 10928 19116 10934 19168
rect 11149 19159 11207 19165
rect 11149 19125 11161 19159
rect 11195 19156 11207 19159
rect 11882 19156 11888 19168
rect 11195 19128 11888 19156
rect 11195 19125 11207 19128
rect 11149 19119 11207 19125
rect 11882 19116 11888 19128
rect 11940 19116 11946 19168
rect 11977 19159 12035 19165
rect 11977 19125 11989 19159
rect 12023 19156 12035 19159
rect 12526 19156 12532 19168
rect 12023 19128 12532 19156
rect 12023 19125 12035 19128
rect 11977 19119 12035 19125
rect 12526 19116 12532 19128
rect 12584 19116 12590 19168
rect 13078 19116 13084 19168
rect 13136 19156 13142 19168
rect 14292 19165 14320 19196
rect 15764 19196 17868 19224
rect 15764 19165 15792 19196
rect 17862 19184 17868 19196
rect 17920 19184 17926 19236
rect 19702 19184 19708 19236
rect 19760 19224 19766 19236
rect 20349 19227 20407 19233
rect 20349 19224 20361 19227
rect 19760 19196 20361 19224
rect 19760 19184 19766 19196
rect 20349 19193 20361 19196
rect 20395 19193 20407 19227
rect 20349 19187 20407 19193
rect 13817 19159 13875 19165
rect 13817 19156 13829 19159
rect 13136 19128 13829 19156
rect 13136 19116 13142 19128
rect 13817 19125 13829 19128
rect 13863 19125 13875 19159
rect 13817 19119 13875 19125
rect 14277 19159 14335 19165
rect 14277 19125 14289 19159
rect 14323 19125 14335 19159
rect 14277 19119 14335 19125
rect 15749 19159 15807 19165
rect 15749 19125 15761 19159
rect 15795 19125 15807 19159
rect 15749 19119 15807 19125
rect 16390 19116 16396 19168
rect 16448 19156 16454 19168
rect 16669 19159 16727 19165
rect 16669 19156 16681 19159
rect 16448 19128 16681 19156
rect 16448 19116 16454 19128
rect 16669 19125 16681 19128
rect 16715 19125 16727 19159
rect 16669 19119 16727 19125
rect 16942 19116 16948 19168
rect 17000 19156 17006 19168
rect 17221 19159 17279 19165
rect 17221 19156 17233 19159
rect 17000 19128 17233 19156
rect 17000 19116 17006 19128
rect 17221 19125 17233 19128
rect 17267 19125 17279 19159
rect 17221 19119 17279 19125
rect 18233 19159 18291 19165
rect 18233 19125 18245 19159
rect 18279 19156 18291 19159
rect 18506 19156 18512 19168
rect 18279 19128 18512 19156
rect 18279 19125 18291 19128
rect 18233 19119 18291 19125
rect 18506 19116 18512 19128
rect 18564 19116 18570 19168
rect 20993 19159 21051 19165
rect 20993 19125 21005 19159
rect 21039 19156 21051 19159
rect 21729 19159 21787 19165
rect 21729 19156 21741 19159
rect 21039 19128 21741 19156
rect 21039 19125 21051 19128
rect 20993 19119 21051 19125
rect 21729 19125 21741 19128
rect 21775 19125 21787 19159
rect 21729 19119 21787 19125
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 2682 18912 2688 18964
rect 2740 18952 2746 18964
rect 8754 18952 8760 18964
rect 2740 18924 8760 18952
rect 2740 18912 2746 18924
rect 8754 18912 8760 18924
rect 8812 18912 8818 18964
rect 8941 18955 8999 18961
rect 8941 18921 8953 18955
rect 8987 18952 8999 18955
rect 9122 18952 9128 18964
rect 8987 18924 9128 18952
rect 8987 18921 8999 18924
rect 8941 18915 8999 18921
rect 9122 18912 9128 18924
rect 9180 18912 9186 18964
rect 9401 18955 9459 18961
rect 9401 18921 9413 18955
rect 9447 18952 9459 18955
rect 11514 18952 11520 18964
rect 9447 18924 11520 18952
rect 9447 18921 9459 18924
rect 9401 18915 9459 18921
rect 11514 18912 11520 18924
rect 11572 18912 11578 18964
rect 11606 18912 11612 18964
rect 11664 18952 11670 18964
rect 13357 18955 13415 18961
rect 13357 18952 13369 18955
rect 11664 18924 13369 18952
rect 11664 18912 11670 18924
rect 13357 18921 13369 18924
rect 13403 18921 13415 18955
rect 13357 18915 13415 18921
rect 14645 18955 14703 18961
rect 14645 18921 14657 18955
rect 14691 18952 14703 18955
rect 15286 18952 15292 18964
rect 14691 18924 15292 18952
rect 14691 18921 14703 18924
rect 14645 18915 14703 18921
rect 15286 18912 15292 18924
rect 15344 18912 15350 18964
rect 18049 18955 18107 18961
rect 18049 18921 18061 18955
rect 18095 18952 18107 18955
rect 18782 18952 18788 18964
rect 18095 18924 18788 18952
rect 18095 18921 18107 18924
rect 18049 18915 18107 18921
rect 18782 18912 18788 18924
rect 18840 18912 18846 18964
rect 8570 18844 8576 18896
rect 8628 18884 8634 18896
rect 11974 18884 11980 18896
rect 8628 18856 11980 18884
rect 8628 18844 8634 18856
rect 11974 18844 11980 18856
rect 12032 18844 12038 18896
rect 13449 18887 13507 18893
rect 13449 18853 13461 18887
rect 13495 18884 13507 18887
rect 15378 18884 15384 18896
rect 13495 18856 15384 18884
rect 13495 18853 13507 18856
rect 13449 18847 13507 18853
rect 4154 18776 4160 18828
rect 4212 18816 4218 18828
rect 8846 18816 8852 18828
rect 4212 18788 8852 18816
rect 4212 18776 4218 18788
rect 8846 18776 8852 18788
rect 8904 18776 8910 18828
rect 8938 18776 8944 18828
rect 8996 18816 9002 18828
rect 9944 18819 10002 18825
rect 8996 18788 9168 18816
rect 8996 18776 9002 18788
rect 6362 18708 6368 18760
rect 6420 18748 6426 18760
rect 9140 18757 9168 18788
rect 9944 18785 9956 18819
rect 9990 18816 10002 18819
rect 10226 18816 10232 18828
rect 9990 18788 10232 18816
rect 9990 18785 10002 18788
rect 9944 18779 10002 18785
rect 10226 18776 10232 18788
rect 10284 18776 10290 18828
rect 11054 18776 11060 18828
rect 11112 18816 11118 18828
rect 11589 18819 11647 18825
rect 11589 18816 11601 18819
rect 11112 18788 11601 18816
rect 11112 18776 11118 18788
rect 11589 18785 11601 18788
rect 11635 18785 11647 18819
rect 11589 18779 11647 18785
rect 11882 18776 11888 18828
rect 11940 18816 11946 18828
rect 13464 18816 13492 18847
rect 15378 18844 15384 18856
rect 15436 18844 15442 18896
rect 17218 18884 17224 18896
rect 17179 18856 17224 18884
rect 17218 18844 17224 18856
rect 17276 18844 17282 18896
rect 18690 18884 18696 18896
rect 18651 18856 18696 18884
rect 18690 18844 18696 18856
rect 18748 18844 18754 18896
rect 19426 18844 19432 18896
rect 19484 18884 19490 18896
rect 19889 18887 19947 18893
rect 19889 18884 19901 18887
rect 19484 18856 19901 18884
rect 19484 18844 19490 18856
rect 19889 18853 19901 18856
rect 19935 18853 19947 18887
rect 19889 18847 19947 18853
rect 11940 18788 13492 18816
rect 11940 18776 11946 18788
rect 14090 18776 14096 18828
rect 14148 18816 14154 18828
rect 14461 18819 14519 18825
rect 14461 18816 14473 18819
rect 14148 18788 14473 18816
rect 14148 18776 14154 18788
rect 14461 18785 14473 18788
rect 14507 18785 14519 18819
rect 15286 18816 15292 18828
rect 15247 18788 15292 18816
rect 14461 18779 14519 18785
rect 15286 18776 15292 18788
rect 15344 18776 15350 18828
rect 15556 18819 15614 18825
rect 15556 18785 15568 18819
rect 15602 18816 15614 18819
rect 15838 18816 15844 18828
rect 15602 18788 15844 18816
rect 15602 18785 15614 18788
rect 15556 18779 15614 18785
rect 15838 18776 15844 18788
rect 15896 18776 15902 18828
rect 16945 18819 17003 18825
rect 16945 18785 16957 18819
rect 16991 18816 17003 18819
rect 17678 18816 17684 18828
rect 16991 18788 17684 18816
rect 16991 18785 17003 18788
rect 16945 18779 17003 18785
rect 17678 18776 17684 18788
rect 17736 18776 17742 18828
rect 17865 18819 17923 18825
rect 17865 18785 17877 18819
rect 17911 18785 17923 18819
rect 17865 18779 17923 18785
rect 18417 18819 18475 18825
rect 18417 18785 18429 18819
rect 18463 18816 18475 18819
rect 18782 18816 18788 18828
rect 18463 18788 18788 18816
rect 18463 18785 18475 18788
rect 18417 18779 18475 18785
rect 9033 18751 9091 18757
rect 9033 18748 9045 18751
rect 6420 18720 9045 18748
rect 6420 18708 6426 18720
rect 9033 18717 9045 18720
rect 9079 18717 9091 18751
rect 9033 18711 9091 18717
rect 9125 18751 9183 18757
rect 9125 18717 9137 18751
rect 9171 18717 9183 18751
rect 9674 18748 9680 18760
rect 9635 18720 9680 18748
rect 9125 18711 9183 18717
rect 3050 18640 3056 18692
rect 3108 18680 3114 18692
rect 8754 18680 8760 18692
rect 3108 18652 8760 18680
rect 3108 18640 3114 18652
rect 8754 18640 8760 18652
rect 8812 18640 8818 18692
rect 9048 18680 9076 18711
rect 9674 18708 9680 18720
rect 9732 18708 9738 18760
rect 10962 18708 10968 18760
rect 11020 18748 11026 18760
rect 11333 18751 11391 18757
rect 11333 18748 11345 18751
rect 11020 18720 11345 18748
rect 11020 18708 11026 18720
rect 11333 18717 11345 18720
rect 11379 18717 11391 18751
rect 11333 18711 11391 18717
rect 13633 18751 13691 18757
rect 13633 18717 13645 18751
rect 13679 18717 13691 18751
rect 13998 18748 14004 18760
rect 13959 18720 14004 18748
rect 13633 18711 13691 18717
rect 9401 18683 9459 18689
rect 9401 18680 9413 18683
rect 9048 18652 9413 18680
rect 9401 18649 9413 18652
rect 9447 18649 9459 18683
rect 9401 18643 9459 18649
rect 10778 18640 10784 18692
rect 10836 18680 10842 18692
rect 12710 18680 12716 18692
rect 10836 18652 11183 18680
rect 12623 18652 12716 18680
rect 10836 18640 10842 18652
rect 3602 18572 3608 18624
rect 3660 18612 3666 18624
rect 8478 18612 8484 18624
rect 3660 18584 8484 18612
rect 3660 18572 3666 18584
rect 8478 18572 8484 18584
rect 8536 18572 8542 18624
rect 8573 18615 8631 18621
rect 8573 18581 8585 18615
rect 8619 18612 8631 18615
rect 10042 18612 10048 18624
rect 8619 18584 10048 18612
rect 8619 18581 8631 18584
rect 8573 18575 8631 18581
rect 10042 18572 10048 18584
rect 10100 18572 10106 18624
rect 11054 18612 11060 18624
rect 11015 18584 11060 18612
rect 11054 18572 11060 18584
rect 11112 18572 11118 18624
rect 11155 18612 11183 18652
rect 12710 18640 12716 18652
rect 12768 18680 12774 18692
rect 13648 18680 13676 18711
rect 13998 18708 14004 18720
rect 14056 18708 14062 18760
rect 17310 18708 17316 18760
rect 17368 18748 17374 18760
rect 17880 18748 17908 18779
rect 18782 18776 18788 18788
rect 18840 18776 18846 18828
rect 19613 18819 19671 18825
rect 19613 18785 19625 18819
rect 19659 18816 19671 18819
rect 19794 18816 19800 18828
rect 19659 18788 19800 18816
rect 19659 18785 19671 18788
rect 19613 18779 19671 18785
rect 19794 18776 19800 18788
rect 19852 18776 19858 18828
rect 19150 18748 19156 18760
rect 17368 18720 17908 18748
rect 19111 18720 19156 18748
rect 17368 18708 17374 18720
rect 19150 18708 19156 18720
rect 19208 18708 19214 18760
rect 17954 18680 17960 18692
rect 12768 18652 13676 18680
rect 16224 18652 17960 18680
rect 12768 18640 12774 18652
rect 12066 18612 12072 18624
rect 11155 18584 12072 18612
rect 12066 18572 12072 18584
rect 12124 18572 12130 18624
rect 12342 18572 12348 18624
rect 12400 18612 12406 18624
rect 12802 18612 12808 18624
rect 12400 18584 12808 18612
rect 12400 18572 12406 18584
rect 12802 18572 12808 18584
rect 12860 18572 12866 18624
rect 12989 18615 13047 18621
rect 12989 18581 13001 18615
rect 13035 18612 13047 18615
rect 13262 18612 13268 18624
rect 13035 18584 13268 18612
rect 13035 18581 13047 18584
rect 12989 18575 13047 18581
rect 13262 18572 13268 18584
rect 13320 18572 13326 18624
rect 13906 18572 13912 18624
rect 13964 18612 13970 18624
rect 16224 18612 16252 18652
rect 17954 18640 17960 18652
rect 18012 18640 18018 18692
rect 18506 18640 18512 18692
rect 18564 18680 18570 18692
rect 20254 18680 20260 18692
rect 18564 18652 20260 18680
rect 18564 18640 18570 18652
rect 20254 18640 20260 18652
rect 20312 18640 20318 18692
rect 16666 18612 16672 18624
rect 13964 18584 16252 18612
rect 16627 18584 16672 18612
rect 13964 18572 13970 18584
rect 16666 18572 16672 18584
rect 16724 18572 16730 18624
rect 16850 18572 16856 18624
rect 16908 18612 16914 18624
rect 19518 18612 19524 18624
rect 16908 18584 19524 18612
rect 16908 18572 16914 18584
rect 19518 18572 19524 18584
rect 19576 18572 19582 18624
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 7466 18368 7472 18420
rect 7524 18408 7530 18420
rect 7524 18380 8892 18408
rect 7524 18368 7530 18380
rect 8864 18340 8892 18380
rect 8938 18368 8944 18420
rect 8996 18408 9002 18420
rect 9217 18411 9275 18417
rect 9217 18408 9229 18411
rect 8996 18380 9229 18408
rect 8996 18368 9002 18380
rect 9217 18377 9229 18380
rect 9263 18377 9275 18411
rect 11882 18408 11888 18420
rect 9217 18371 9275 18377
rect 9508 18380 11888 18408
rect 9508 18340 9536 18380
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 12161 18411 12219 18417
rect 12161 18377 12173 18411
rect 12207 18408 12219 18411
rect 13906 18408 13912 18420
rect 12207 18380 13912 18408
rect 12207 18377 12219 18380
rect 12161 18371 12219 18377
rect 13906 18368 13912 18380
rect 13964 18368 13970 18420
rect 15838 18408 15844 18420
rect 15799 18380 15844 18408
rect 15838 18368 15844 18380
rect 15896 18368 15902 18420
rect 17589 18411 17647 18417
rect 17589 18377 17601 18411
rect 17635 18408 17647 18411
rect 18598 18408 18604 18420
rect 17635 18380 18604 18408
rect 17635 18377 17647 18380
rect 17589 18371 17647 18377
rect 18598 18368 18604 18380
rect 18656 18368 18662 18420
rect 8864 18312 9536 18340
rect 9585 18343 9643 18349
rect 9585 18309 9597 18343
rect 9631 18340 9643 18343
rect 10778 18340 10784 18352
rect 9631 18312 10784 18340
rect 9631 18309 9643 18312
rect 9585 18303 9643 18309
rect 10778 18300 10784 18312
rect 10836 18300 10842 18352
rect 5810 18232 5816 18284
rect 5868 18272 5874 18284
rect 7466 18272 7472 18284
rect 5868 18244 7472 18272
rect 5868 18232 5874 18244
rect 7466 18232 7472 18244
rect 7524 18232 7530 18284
rect 8846 18232 8852 18284
rect 8904 18272 8910 18284
rect 9858 18272 9864 18284
rect 8904 18244 9864 18272
rect 8904 18232 8910 18244
rect 9858 18232 9864 18244
rect 9916 18232 9922 18284
rect 10042 18272 10048 18284
rect 10003 18244 10048 18272
rect 10042 18232 10048 18244
rect 10100 18232 10106 18284
rect 10226 18272 10232 18284
rect 10139 18244 10232 18272
rect 10226 18232 10232 18244
rect 10284 18272 10290 18284
rect 11149 18275 11207 18281
rect 11149 18272 11161 18275
rect 10284 18244 11161 18272
rect 10284 18232 10290 18244
rect 11149 18241 11161 18244
rect 11195 18241 11207 18275
rect 12802 18272 12808 18284
rect 12763 18244 12808 18272
rect 11149 18235 11207 18241
rect 12802 18232 12808 18244
rect 12860 18232 12866 18284
rect 15838 18232 15844 18284
rect 15896 18272 15902 18284
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 15896 18244 16681 18272
rect 15896 18232 15902 18244
rect 16669 18241 16681 18244
rect 16715 18241 16727 18275
rect 18598 18272 18604 18284
rect 18559 18244 18604 18272
rect 16669 18235 16727 18241
rect 18598 18232 18604 18244
rect 18656 18232 18662 18284
rect 7101 18207 7159 18213
rect 7101 18173 7113 18207
rect 7147 18204 7159 18207
rect 7147 18176 7328 18204
rect 7147 18173 7159 18176
rect 7101 18167 7159 18173
rect 4706 18096 4712 18148
rect 4764 18136 4770 18148
rect 6822 18136 6828 18148
rect 4764 18108 6828 18136
rect 4764 18096 4770 18108
rect 6822 18096 6828 18108
rect 6880 18096 6886 18148
rect 5258 18028 5264 18080
rect 5316 18068 5322 18080
rect 7190 18068 7196 18080
rect 5316 18040 7196 18068
rect 5316 18028 5322 18040
rect 7190 18028 7196 18040
rect 7248 18028 7254 18080
rect 7300 18068 7328 18176
rect 7742 18164 7748 18216
rect 7800 18204 7806 18216
rect 7837 18207 7895 18213
rect 7837 18204 7849 18207
rect 7800 18176 7849 18204
rect 7800 18164 7806 18176
rect 7837 18173 7849 18176
rect 7883 18173 7895 18207
rect 10318 18204 10324 18216
rect 7837 18167 7895 18173
rect 8036 18176 10324 18204
rect 7377 18139 7435 18145
rect 7377 18105 7389 18139
rect 7423 18136 7435 18139
rect 8036 18136 8064 18176
rect 10318 18164 10324 18176
rect 10376 18164 10382 18216
rect 10962 18164 10968 18216
rect 11020 18204 11026 18216
rect 13078 18213 13084 18216
rect 11057 18207 11115 18213
rect 11057 18204 11069 18207
rect 11020 18176 11069 18204
rect 11020 18164 11026 18176
rect 11057 18173 11069 18176
rect 11103 18173 11115 18207
rect 11057 18167 11115 18173
rect 11609 18207 11667 18213
rect 11609 18173 11621 18207
rect 11655 18173 11667 18207
rect 11609 18167 11667 18173
rect 11885 18207 11943 18213
rect 11885 18173 11897 18207
rect 11931 18204 11943 18207
rect 12161 18207 12219 18213
rect 12161 18204 12173 18207
rect 11931 18176 12173 18204
rect 11931 18173 11943 18176
rect 11885 18167 11943 18173
rect 12161 18173 12173 18176
rect 12207 18173 12219 18207
rect 13072 18204 13084 18213
rect 13039 18176 13084 18204
rect 12161 18167 12219 18173
rect 13072 18167 13084 18176
rect 7423 18108 8064 18136
rect 8104 18139 8162 18145
rect 7423 18105 7435 18108
rect 7377 18099 7435 18105
rect 8104 18105 8116 18139
rect 8150 18136 8162 18139
rect 8846 18136 8852 18148
rect 8150 18108 8852 18136
rect 8150 18105 8162 18108
rect 8104 18099 8162 18105
rect 8846 18096 8852 18108
rect 8904 18096 8910 18148
rect 9858 18096 9864 18148
rect 9916 18136 9922 18148
rect 9916 18108 10916 18136
rect 9916 18096 9922 18108
rect 8662 18068 8668 18080
rect 7300 18040 8668 18068
rect 8662 18028 8668 18040
rect 8720 18028 8726 18080
rect 9953 18071 10011 18077
rect 9953 18037 9965 18071
rect 9999 18068 10011 18071
rect 10042 18068 10048 18080
rect 9999 18040 10048 18068
rect 9999 18037 10011 18040
rect 9953 18031 10011 18037
rect 10042 18028 10048 18040
rect 10100 18028 10106 18080
rect 10594 18068 10600 18080
rect 10555 18040 10600 18068
rect 10594 18028 10600 18040
rect 10652 18028 10658 18080
rect 10888 18068 10916 18108
rect 11146 18096 11152 18148
rect 11204 18136 11210 18148
rect 11624 18136 11652 18167
rect 13078 18164 13084 18167
rect 13136 18164 13142 18216
rect 14461 18207 14519 18213
rect 14461 18173 14473 18207
rect 14507 18204 14519 18207
rect 14507 18176 15148 18204
rect 14507 18173 14519 18176
rect 14461 18167 14519 18173
rect 14706 18139 14764 18145
rect 14706 18136 14718 18139
rect 11204 18108 11652 18136
rect 14200 18108 14718 18136
rect 11204 18096 11210 18108
rect 14200 18080 14228 18108
rect 14706 18105 14718 18108
rect 14752 18105 14764 18139
rect 15120 18136 15148 18176
rect 15194 18164 15200 18216
rect 15252 18204 15258 18216
rect 16022 18204 16028 18216
rect 15252 18176 16028 18204
rect 15252 18164 15258 18176
rect 16022 18164 16028 18176
rect 16080 18204 16086 18216
rect 16577 18207 16635 18213
rect 16577 18204 16589 18207
rect 16080 18176 16589 18204
rect 16080 18164 16086 18176
rect 16577 18173 16589 18176
rect 16623 18173 16635 18207
rect 16577 18167 16635 18173
rect 17405 18207 17463 18213
rect 17405 18173 17417 18207
rect 17451 18173 17463 18207
rect 17405 18167 17463 18173
rect 18417 18207 18475 18213
rect 18417 18173 18429 18207
rect 18463 18204 18475 18207
rect 19150 18204 19156 18216
rect 18463 18176 19156 18204
rect 18463 18173 18475 18176
rect 18417 18167 18475 18173
rect 17420 18136 17448 18167
rect 19150 18164 19156 18176
rect 19208 18164 19214 18216
rect 19426 18204 19432 18216
rect 19387 18176 19432 18204
rect 19426 18164 19432 18176
rect 19484 18164 19490 18216
rect 19978 18204 19984 18216
rect 19939 18176 19984 18204
rect 19978 18164 19984 18176
rect 20036 18164 20042 18216
rect 20070 18164 20076 18216
rect 20128 18204 20134 18216
rect 20533 18207 20591 18213
rect 20533 18204 20545 18207
rect 20128 18176 20545 18204
rect 20128 18164 20134 18176
rect 20533 18173 20545 18176
rect 20579 18173 20591 18207
rect 20533 18167 20591 18173
rect 18874 18136 18880 18148
rect 15120 18108 15332 18136
rect 17420 18108 18880 18136
rect 14706 18099 14764 18105
rect 15304 18080 15332 18108
rect 18874 18096 18880 18108
rect 18932 18096 18938 18148
rect 10965 18071 11023 18077
rect 10965 18068 10977 18071
rect 10888 18040 10977 18068
rect 10965 18037 10977 18040
rect 11011 18037 11023 18071
rect 10965 18031 11023 18037
rect 11238 18028 11244 18080
rect 11296 18068 11302 18080
rect 12710 18068 12716 18080
rect 11296 18040 12716 18068
rect 11296 18028 11302 18040
rect 12710 18028 12716 18040
rect 12768 18028 12774 18080
rect 14182 18068 14188 18080
rect 14143 18040 14188 18068
rect 14182 18028 14188 18040
rect 14240 18028 14246 18080
rect 15286 18028 15292 18080
rect 15344 18068 15350 18080
rect 15930 18068 15936 18080
rect 15344 18040 15936 18068
rect 15344 18028 15350 18040
rect 15930 18028 15936 18040
rect 15988 18028 15994 18080
rect 16114 18068 16120 18080
rect 16075 18040 16120 18068
rect 16114 18028 16120 18040
rect 16172 18028 16178 18080
rect 16206 18028 16212 18080
rect 16264 18068 16270 18080
rect 16485 18071 16543 18077
rect 16485 18068 16497 18071
rect 16264 18040 16497 18068
rect 16264 18028 16270 18040
rect 16485 18037 16497 18040
rect 16531 18037 16543 18071
rect 16485 18031 16543 18037
rect 17954 18028 17960 18080
rect 18012 18068 18018 18080
rect 18049 18071 18107 18077
rect 18049 18068 18061 18071
rect 18012 18040 18061 18068
rect 18012 18028 18018 18040
rect 18049 18037 18061 18040
rect 18095 18037 18107 18071
rect 18049 18031 18107 18037
rect 18138 18028 18144 18080
rect 18196 18068 18202 18080
rect 18509 18071 18567 18077
rect 18509 18068 18521 18071
rect 18196 18040 18521 18068
rect 18196 18028 18202 18040
rect 18509 18037 18521 18040
rect 18555 18037 18567 18071
rect 18509 18031 18567 18037
rect 19242 18028 19248 18080
rect 19300 18068 19306 18080
rect 19613 18071 19671 18077
rect 19613 18068 19625 18071
rect 19300 18040 19625 18068
rect 19300 18028 19306 18040
rect 19613 18037 19625 18040
rect 19659 18037 19671 18071
rect 20162 18068 20168 18080
rect 20123 18040 20168 18068
rect 19613 18031 19671 18037
rect 20162 18028 20168 18040
rect 20220 18028 20226 18080
rect 20714 18068 20720 18080
rect 20675 18040 20720 18068
rect 20714 18028 20720 18040
rect 20772 18028 20778 18080
rect 21726 18000 21732 18012
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 21687 17972 21732 18000
rect 21726 17960 21732 17972
rect 21784 17960 21790 18012
rect 1104 17904 21620 17926
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 7377 17867 7435 17873
rect 7377 17864 7389 17867
rect 6972 17836 7389 17864
rect 6972 17824 6978 17836
rect 7377 17833 7389 17836
rect 7423 17833 7435 17867
rect 7377 17827 7435 17833
rect 7466 17824 7472 17876
rect 7524 17864 7530 17876
rect 9858 17864 9864 17876
rect 7524 17836 7569 17864
rect 9819 17836 9864 17864
rect 7524 17824 7530 17836
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 10594 17824 10600 17876
rect 10652 17864 10658 17876
rect 10689 17867 10747 17873
rect 10689 17864 10701 17867
rect 10652 17836 10701 17864
rect 10652 17824 10658 17836
rect 10689 17833 10701 17836
rect 10735 17833 10747 17867
rect 10689 17827 10747 17833
rect 10778 17824 10784 17876
rect 10836 17864 10842 17876
rect 10836 17836 10881 17864
rect 10836 17824 10842 17836
rect 12342 17824 12348 17876
rect 12400 17864 12406 17876
rect 13081 17867 13139 17873
rect 13081 17864 13093 17867
rect 12400 17836 13093 17864
rect 12400 17824 12406 17836
rect 13081 17833 13093 17836
rect 13127 17833 13139 17867
rect 13081 17827 13139 17833
rect 13173 17867 13231 17873
rect 13173 17833 13185 17867
rect 13219 17864 13231 17867
rect 13262 17864 13268 17876
rect 13219 17836 13268 17864
rect 13219 17833 13231 17836
rect 13173 17827 13231 17833
rect 13262 17824 13268 17836
rect 13320 17824 13326 17876
rect 13998 17824 14004 17876
rect 14056 17864 14062 17876
rect 14093 17867 14151 17873
rect 14093 17864 14105 17867
rect 14056 17836 14105 17864
rect 14056 17824 14062 17836
rect 14093 17833 14105 17836
rect 14139 17833 14151 17867
rect 14093 17827 14151 17833
rect 14185 17867 14243 17873
rect 14185 17833 14197 17867
rect 14231 17864 14243 17867
rect 14550 17864 14556 17876
rect 14231 17836 14556 17864
rect 14231 17833 14243 17836
rect 14185 17827 14243 17833
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 14737 17867 14795 17873
rect 14737 17833 14749 17867
rect 14783 17864 14795 17867
rect 16206 17864 16212 17876
rect 14783 17836 16212 17864
rect 14783 17833 14795 17836
rect 14737 17827 14795 17833
rect 16206 17824 16212 17836
rect 16264 17824 16270 17876
rect 20070 17864 20076 17876
rect 16316 17836 20076 17864
rect 8665 17799 8723 17805
rect 8665 17765 8677 17799
rect 8711 17796 8723 17799
rect 9398 17796 9404 17808
rect 8711 17768 9404 17796
rect 8711 17765 8723 17768
rect 8665 17759 8723 17765
rect 9398 17756 9404 17768
rect 9456 17796 9462 17808
rect 10502 17796 10508 17808
rect 9456 17768 10508 17796
rect 9456 17756 9462 17768
rect 10502 17756 10508 17768
rect 10560 17756 10566 17808
rect 16316 17796 16344 17836
rect 20070 17824 20076 17836
rect 20128 17824 20134 17876
rect 13004 17768 16344 17796
rect 16568 17799 16626 17805
rect 8570 17728 8576 17740
rect 8531 17700 8576 17728
rect 8570 17688 8576 17700
rect 8628 17688 8634 17740
rect 11241 17731 11299 17737
rect 11241 17697 11253 17731
rect 11287 17728 11299 17731
rect 11333 17731 11391 17737
rect 11333 17728 11345 17731
rect 11287 17700 11345 17728
rect 11287 17697 11299 17700
rect 11241 17691 11299 17697
rect 11333 17697 11345 17700
rect 11379 17697 11391 17731
rect 11333 17691 11391 17697
rect 11609 17731 11667 17737
rect 11609 17697 11621 17731
rect 11655 17728 11667 17731
rect 13004 17728 13032 17768
rect 16568 17765 16580 17799
rect 16614 17796 16626 17799
rect 16666 17796 16672 17808
rect 16614 17768 16672 17796
rect 16614 17765 16626 17768
rect 16568 17759 16626 17765
rect 16666 17756 16672 17768
rect 16724 17756 16730 17808
rect 17773 17799 17831 17805
rect 17773 17765 17785 17799
rect 17819 17796 17831 17799
rect 18224 17799 18282 17805
rect 18224 17796 18236 17799
rect 17819 17768 18236 17796
rect 17819 17765 17831 17768
rect 17773 17759 17831 17765
rect 18224 17765 18236 17768
rect 18270 17796 18282 17799
rect 18598 17796 18604 17808
rect 18270 17768 18604 17796
rect 18270 17765 18282 17768
rect 18224 17759 18282 17765
rect 18598 17756 18604 17768
rect 18656 17756 18662 17808
rect 19426 17756 19432 17808
rect 19484 17796 19490 17808
rect 19981 17799 20039 17805
rect 19981 17796 19993 17799
rect 19484 17768 19993 17796
rect 19484 17756 19490 17768
rect 19981 17765 19993 17768
rect 20027 17765 20039 17799
rect 19981 17759 20039 17765
rect 15654 17728 15660 17740
rect 11655 17700 13032 17728
rect 15615 17700 15660 17728
rect 11655 17697 11667 17700
rect 11609 17691 11667 17697
rect 15654 17688 15660 17700
rect 15712 17688 15718 17740
rect 15746 17688 15752 17740
rect 15804 17728 15810 17740
rect 15804 17700 15849 17728
rect 15804 17688 15810 17700
rect 16390 17688 16396 17740
rect 16448 17728 16454 17740
rect 16448 17700 19012 17728
rect 16448 17688 16454 17700
rect 7653 17663 7711 17669
rect 7653 17629 7665 17663
rect 7699 17660 7711 17663
rect 7742 17660 7748 17672
rect 7699 17632 7748 17660
rect 7699 17629 7711 17632
rect 7653 17623 7711 17629
rect 7742 17620 7748 17632
rect 7800 17620 7806 17672
rect 8757 17663 8815 17669
rect 8757 17629 8769 17663
rect 8803 17629 8815 17663
rect 8757 17623 8815 17629
rect 10965 17663 11023 17669
rect 10965 17629 10977 17663
rect 11011 17660 11023 17663
rect 11054 17660 11060 17672
rect 11011 17632 11060 17660
rect 11011 17629 11023 17632
rect 10965 17623 11023 17629
rect 7009 17595 7067 17601
rect 7009 17561 7021 17595
rect 7055 17592 7067 17595
rect 8294 17592 8300 17604
rect 7055 17564 8300 17592
rect 7055 17561 7067 17564
rect 7009 17555 7067 17561
rect 8294 17552 8300 17564
rect 8352 17552 8358 17604
rect 8386 17552 8392 17604
rect 8444 17592 8450 17604
rect 8772 17592 8800 17623
rect 11054 17620 11060 17632
rect 11112 17620 11118 17672
rect 13170 17620 13176 17672
rect 13228 17660 13234 17672
rect 13265 17663 13323 17669
rect 13265 17660 13277 17663
rect 13228 17632 13277 17660
rect 13228 17620 13234 17632
rect 13265 17629 13277 17632
rect 13311 17629 13323 17663
rect 13265 17623 13323 17629
rect 14277 17663 14335 17669
rect 14277 17629 14289 17663
rect 14323 17629 14335 17663
rect 15838 17660 15844 17672
rect 15799 17632 15844 17660
rect 14277 17623 14335 17629
rect 8444 17564 8800 17592
rect 13280 17592 13308 17623
rect 14292 17592 14320 17623
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 16022 17620 16028 17672
rect 16080 17660 16086 17672
rect 16301 17663 16359 17669
rect 16301 17660 16313 17663
rect 16080 17632 16313 17660
rect 16080 17620 16086 17632
rect 16301 17629 16313 17632
rect 16347 17629 16359 17663
rect 17773 17663 17831 17669
rect 17773 17660 17785 17663
rect 16301 17623 16359 17629
rect 17696 17632 17785 17660
rect 13280 17564 14320 17592
rect 8444 17552 8450 17564
rect 8205 17527 8263 17533
rect 8205 17493 8217 17527
rect 8251 17524 8263 17527
rect 9490 17524 9496 17536
rect 8251 17496 9496 17524
rect 8251 17493 8263 17496
rect 8205 17487 8263 17493
rect 9490 17484 9496 17496
rect 9548 17484 9554 17536
rect 10321 17527 10379 17533
rect 10321 17493 10333 17527
rect 10367 17524 10379 17527
rect 11241 17527 11299 17533
rect 11241 17524 11253 17527
rect 10367 17496 11253 17524
rect 10367 17493 10379 17496
rect 10321 17487 10379 17493
rect 11241 17493 11253 17496
rect 11287 17493 11299 17527
rect 11241 17487 11299 17493
rect 12713 17527 12771 17533
rect 12713 17493 12725 17527
rect 12759 17524 12771 17527
rect 13262 17524 13268 17536
rect 12759 17496 13268 17524
rect 12759 17493 12771 17496
rect 12713 17487 12771 17493
rect 13262 17484 13268 17496
rect 13320 17484 13326 17536
rect 13446 17484 13452 17536
rect 13504 17524 13510 17536
rect 13725 17527 13783 17533
rect 13725 17524 13737 17527
rect 13504 17496 13737 17524
rect 13504 17484 13510 17496
rect 13725 17493 13737 17496
rect 13771 17493 13783 17527
rect 13725 17487 13783 17493
rect 15289 17527 15347 17533
rect 15289 17493 15301 17527
rect 15335 17524 15347 17527
rect 16206 17524 16212 17536
rect 15335 17496 16212 17524
rect 15335 17493 15347 17496
rect 15289 17487 15347 17493
rect 16206 17484 16212 17496
rect 16264 17484 16270 17536
rect 16316 17524 16344 17623
rect 17494 17592 17500 17604
rect 17236 17564 17500 17592
rect 17236 17524 17264 17564
rect 17494 17552 17500 17564
rect 17552 17552 17558 17604
rect 17696 17601 17724 17632
rect 17773 17629 17785 17632
rect 17819 17629 17831 17663
rect 17773 17623 17831 17629
rect 17862 17620 17868 17672
rect 17920 17660 17926 17672
rect 17957 17663 18015 17669
rect 17957 17660 17969 17663
rect 17920 17632 17969 17660
rect 17920 17620 17926 17632
rect 17957 17629 17969 17632
rect 18003 17629 18015 17663
rect 18984 17660 19012 17700
rect 19150 17688 19156 17740
rect 19208 17728 19214 17740
rect 19705 17731 19763 17737
rect 19705 17728 19717 17731
rect 19208 17700 19717 17728
rect 19208 17688 19214 17700
rect 19705 17697 19717 17700
rect 19751 17697 19763 17731
rect 19705 17691 19763 17697
rect 21910 17660 21916 17672
rect 18984 17632 21916 17660
rect 17957 17623 18015 17629
rect 21910 17620 21916 17632
rect 21968 17620 21974 17672
rect 17681 17595 17739 17601
rect 17681 17561 17693 17595
rect 17727 17561 17739 17595
rect 17681 17555 17739 17561
rect 16316 17496 17264 17524
rect 17770 17484 17776 17536
rect 17828 17524 17834 17536
rect 19337 17527 19395 17533
rect 19337 17524 19349 17527
rect 17828 17496 19349 17524
rect 17828 17484 17834 17496
rect 19337 17493 19349 17496
rect 19383 17493 19395 17527
rect 19337 17487 19395 17493
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 7834 17320 7840 17332
rect 7484 17292 7840 17320
rect 7006 17144 7012 17196
rect 7064 17184 7070 17196
rect 7484 17193 7512 17292
rect 7834 17280 7840 17292
rect 7892 17280 7898 17332
rect 8846 17320 8852 17332
rect 8807 17292 8852 17320
rect 8846 17280 8852 17292
rect 8904 17280 8910 17332
rect 12250 17280 12256 17332
rect 12308 17320 12314 17332
rect 15470 17320 15476 17332
rect 12308 17292 15476 17320
rect 12308 17280 12314 17292
rect 15470 17280 15476 17292
rect 15528 17280 15534 17332
rect 16574 17320 16580 17332
rect 15672 17292 16580 17320
rect 13081 17255 13139 17261
rect 8496 17224 13032 17252
rect 7469 17187 7527 17193
rect 7469 17184 7481 17187
rect 7064 17156 7481 17184
rect 7064 17144 7070 17156
rect 7469 17153 7481 17156
rect 7515 17153 7527 17187
rect 7469 17147 7527 17153
rect 842 17076 848 17128
rect 900 17116 906 17128
rect 8496 17116 8524 17224
rect 8846 17144 8852 17196
rect 8904 17184 8910 17196
rect 9677 17187 9735 17193
rect 9677 17184 9689 17187
rect 8904 17156 9689 17184
rect 8904 17144 8910 17156
rect 9677 17153 9689 17156
rect 9723 17153 9735 17187
rect 10870 17184 10876 17196
rect 10783 17156 10876 17184
rect 9677 17147 9735 17153
rect 10870 17144 10876 17156
rect 10928 17184 10934 17196
rect 11882 17184 11888 17196
rect 10928 17156 11888 17184
rect 10928 17144 10934 17156
rect 11882 17144 11888 17156
rect 11940 17144 11946 17196
rect 9490 17116 9496 17128
rect 900 17088 8524 17116
rect 9451 17088 9496 17116
rect 900 17076 906 17088
rect 9490 17076 9496 17088
rect 9548 17076 9554 17128
rect 9950 17076 9956 17128
rect 10008 17116 10014 17128
rect 10008 17088 10824 17116
rect 10008 17076 10014 17088
rect 7736 17051 7794 17057
rect 7736 17017 7748 17051
rect 7782 17048 7794 17051
rect 8386 17048 8392 17060
rect 7782 17020 8392 17048
rect 7782 17017 7794 17020
rect 7736 17011 7794 17017
rect 8386 17008 8392 17020
rect 8444 17008 8450 17060
rect 9766 17008 9772 17060
rect 9824 17048 9830 17060
rect 10689 17051 10747 17057
rect 10689 17048 10701 17051
rect 9824 17020 10701 17048
rect 9824 17008 9830 17020
rect 10689 17017 10701 17020
rect 10735 17017 10747 17051
rect 10689 17011 10747 17017
rect 9122 16980 9128 16992
rect 9083 16952 9128 16980
rect 9122 16940 9128 16952
rect 9180 16940 9186 16992
rect 9214 16940 9220 16992
rect 9272 16980 9278 16992
rect 9585 16983 9643 16989
rect 9585 16980 9597 16983
rect 9272 16952 9597 16980
rect 9272 16940 9278 16952
rect 9585 16949 9597 16952
rect 9631 16949 9643 16983
rect 9585 16943 9643 16949
rect 10229 16983 10287 16989
rect 10229 16949 10241 16983
rect 10275 16980 10287 16983
rect 10502 16980 10508 16992
rect 10275 16952 10508 16980
rect 10275 16949 10287 16952
rect 10229 16943 10287 16949
rect 10502 16940 10508 16952
rect 10560 16940 10566 16992
rect 10597 16983 10655 16989
rect 10597 16949 10609 16983
rect 10643 16980 10655 16983
rect 10796 16980 10824 17088
rect 11701 17051 11759 17057
rect 11701 17017 11713 17051
rect 11747 17048 11759 17051
rect 12529 17051 12587 17057
rect 12529 17048 12541 17051
rect 11747 17020 12541 17048
rect 11747 17017 11759 17020
rect 11701 17011 11759 17017
rect 12529 17017 12541 17020
rect 12575 17017 12587 17051
rect 12529 17011 12587 17017
rect 10962 16980 10968 16992
rect 10643 16952 10968 16980
rect 10643 16949 10655 16952
rect 10597 16943 10655 16949
rect 10962 16940 10968 16952
rect 11020 16940 11026 16992
rect 11333 16983 11391 16989
rect 11333 16949 11345 16983
rect 11379 16980 11391 16983
rect 11606 16980 11612 16992
rect 11379 16952 11612 16980
rect 11379 16949 11391 16952
rect 11333 16943 11391 16949
rect 11606 16940 11612 16952
rect 11664 16940 11670 16992
rect 11793 16983 11851 16989
rect 11793 16949 11805 16983
rect 11839 16980 11851 16983
rect 12250 16980 12256 16992
rect 11839 16952 12256 16980
rect 11839 16949 11851 16952
rect 11793 16943 11851 16949
rect 12250 16940 12256 16952
rect 12308 16940 12314 16992
rect 13004 16980 13032 17224
rect 13081 17221 13093 17255
rect 13127 17221 13139 17255
rect 13081 17215 13139 17221
rect 13096 17116 13124 17215
rect 14550 17212 14556 17264
rect 14608 17252 14614 17264
rect 15672 17252 15700 17292
rect 16574 17280 16580 17292
rect 16632 17280 16638 17332
rect 16945 17323 17003 17329
rect 16945 17289 16957 17323
rect 16991 17320 17003 17323
rect 19150 17320 19156 17332
rect 16991 17292 19156 17320
rect 16991 17289 17003 17292
rect 16945 17283 17003 17289
rect 19150 17280 19156 17292
rect 19208 17280 19214 17332
rect 14608 17224 15700 17252
rect 15749 17255 15807 17261
rect 14608 17212 14614 17224
rect 15749 17221 15761 17255
rect 15795 17252 15807 17255
rect 15795 17224 19840 17252
rect 15795 17221 15807 17224
rect 15749 17215 15807 17221
rect 13262 17144 13268 17196
rect 13320 17184 13326 17196
rect 13541 17187 13599 17193
rect 13541 17184 13553 17187
rect 13320 17156 13553 17184
rect 13320 17144 13326 17156
rect 13541 17153 13553 17156
rect 13587 17153 13599 17187
rect 13541 17147 13599 17153
rect 13725 17187 13783 17193
rect 13725 17153 13737 17187
rect 13771 17184 13783 17187
rect 14182 17184 14188 17196
rect 13771 17156 14188 17184
rect 13771 17153 13783 17156
rect 13725 17147 13783 17153
rect 14182 17144 14188 17156
rect 14240 17144 14246 17196
rect 16206 17184 16212 17196
rect 16167 17156 16212 17184
rect 16206 17144 16212 17156
rect 16264 17144 16270 17196
rect 16393 17187 16451 17193
rect 16393 17153 16405 17187
rect 16439 17184 16451 17187
rect 16666 17184 16672 17196
rect 16439 17156 16672 17184
rect 16439 17153 16451 17156
rect 16393 17147 16451 17153
rect 16666 17144 16672 17156
rect 16724 17144 16730 17196
rect 17589 17187 17647 17193
rect 17589 17153 17601 17187
rect 17635 17184 17647 17187
rect 17770 17184 17776 17196
rect 17635 17156 17776 17184
rect 17635 17153 17647 17156
rect 17589 17147 17647 17153
rect 17770 17144 17776 17156
rect 17828 17144 17834 17196
rect 17862 17144 17868 17196
rect 17920 17184 17926 17196
rect 18690 17184 18696 17196
rect 17920 17156 18460 17184
rect 18651 17156 18696 17184
rect 17920 17144 17926 17156
rect 14093 17119 14151 17125
rect 14093 17116 14105 17119
rect 13096 17088 14105 17116
rect 14093 17085 14105 17088
rect 14139 17085 14151 17119
rect 14093 17079 14151 17085
rect 15197 17119 15255 17125
rect 15197 17085 15209 17119
rect 15243 17116 15255 17119
rect 16022 17116 16028 17128
rect 15243 17088 16028 17116
rect 15243 17085 15255 17088
rect 15197 17079 15255 17085
rect 16022 17076 16028 17088
rect 16080 17076 16086 17128
rect 16114 17076 16120 17128
rect 16172 17116 16178 17128
rect 17313 17119 17371 17125
rect 16172 17088 16217 17116
rect 16172 17076 16178 17088
rect 17313 17085 17325 17119
rect 17359 17116 17371 17119
rect 17954 17116 17960 17128
rect 17359 17088 17960 17116
rect 17359 17085 17371 17088
rect 17313 17079 17371 17085
rect 17954 17076 17960 17088
rect 18012 17076 18018 17128
rect 18432 17125 18460 17156
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 19812 17125 19840 17224
rect 19978 17184 19984 17196
rect 19939 17156 19984 17184
rect 19978 17144 19984 17156
rect 20036 17144 20042 17196
rect 20806 17184 20812 17196
rect 20767 17156 20812 17184
rect 20806 17144 20812 17156
rect 20864 17144 20870 17196
rect 18417 17119 18475 17125
rect 18417 17085 18429 17119
rect 18463 17085 18475 17119
rect 18417 17079 18475 17085
rect 19245 17119 19303 17125
rect 19245 17085 19257 17119
rect 19291 17085 19303 17119
rect 19245 17079 19303 17085
rect 19797 17119 19855 17125
rect 19797 17085 19809 17119
rect 19843 17085 19855 17119
rect 19797 17079 19855 17085
rect 13446 17048 13452 17060
rect 13407 17020 13452 17048
rect 13446 17008 13452 17020
rect 13504 17008 13510 17060
rect 14369 17051 14427 17057
rect 14369 17017 14381 17051
rect 14415 17048 14427 17051
rect 19260 17048 19288 17079
rect 20070 17076 20076 17128
rect 20128 17116 20134 17128
rect 20533 17119 20591 17125
rect 20533 17116 20545 17119
rect 20128 17088 20545 17116
rect 20128 17076 20134 17088
rect 20533 17085 20545 17088
rect 20579 17085 20591 17119
rect 20533 17079 20591 17085
rect 14415 17020 19288 17048
rect 14415 17017 14427 17020
rect 14369 17011 14427 17017
rect 14274 16980 14280 16992
rect 13004 16952 14280 16980
rect 14274 16940 14280 16952
rect 14332 16940 14338 16992
rect 15381 16983 15439 16989
rect 15381 16949 15393 16983
rect 15427 16980 15439 16983
rect 16390 16980 16396 16992
rect 15427 16952 16396 16980
rect 15427 16949 15439 16952
rect 15381 16943 15439 16949
rect 16390 16940 16396 16952
rect 16448 16940 16454 16992
rect 17405 16983 17463 16989
rect 17405 16949 17417 16983
rect 17451 16980 17463 16983
rect 18049 16983 18107 16989
rect 18049 16980 18061 16983
rect 17451 16952 18061 16980
rect 17451 16949 17463 16952
rect 17405 16943 17463 16949
rect 18049 16949 18061 16952
rect 18095 16949 18107 16983
rect 18049 16943 18107 16949
rect 18414 16940 18420 16992
rect 18472 16980 18478 16992
rect 18509 16983 18567 16989
rect 18509 16980 18521 16983
rect 18472 16952 18521 16980
rect 18472 16940 18478 16952
rect 18509 16949 18521 16952
rect 18555 16949 18567 16983
rect 19426 16980 19432 16992
rect 19387 16952 19432 16980
rect 18509 16943 18567 16949
rect 19426 16940 19432 16952
rect 19484 16940 19490 16992
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 10318 16776 10324 16788
rect 8956 16748 10324 16776
rect 8956 16717 8984 16748
rect 10318 16736 10324 16748
rect 10376 16736 10382 16788
rect 14093 16779 14151 16785
rect 14093 16745 14105 16779
rect 14139 16776 14151 16779
rect 15749 16779 15807 16785
rect 15749 16776 15761 16779
rect 14139 16748 15761 16776
rect 14139 16745 14151 16748
rect 14093 16739 14151 16745
rect 15749 16745 15761 16748
rect 15795 16745 15807 16779
rect 15749 16739 15807 16745
rect 17129 16779 17187 16785
rect 17129 16745 17141 16779
rect 17175 16776 17187 16779
rect 18506 16776 18512 16788
rect 17175 16748 18512 16776
rect 17175 16745 17187 16748
rect 17129 16739 17187 16745
rect 18506 16736 18512 16748
rect 18564 16736 18570 16788
rect 18598 16736 18604 16788
rect 18656 16776 18662 16788
rect 21358 16776 21364 16788
rect 18656 16748 21364 16776
rect 18656 16736 18662 16748
rect 21358 16736 21364 16748
rect 21416 16736 21422 16788
rect 8941 16711 8999 16717
rect 8941 16677 8953 16711
rect 8987 16677 8999 16711
rect 8941 16671 8999 16677
rect 10680 16711 10738 16717
rect 10680 16677 10692 16711
rect 10726 16708 10738 16711
rect 10870 16708 10876 16720
rect 10726 16680 10876 16708
rect 10726 16677 10738 16680
rect 10680 16671 10738 16677
rect 10870 16668 10876 16680
rect 10928 16668 10934 16720
rect 12360 16680 20300 16708
rect 7006 16640 7012 16652
rect 6967 16612 7012 16640
rect 7006 16600 7012 16612
rect 7064 16600 7070 16652
rect 7276 16643 7334 16649
rect 7276 16609 7288 16643
rect 7322 16640 7334 16643
rect 7742 16640 7748 16652
rect 7322 16612 7748 16640
rect 7322 16609 7334 16612
rect 7276 16603 7334 16609
rect 7742 16600 7748 16612
rect 7800 16600 7806 16652
rect 8665 16643 8723 16649
rect 8665 16609 8677 16643
rect 8711 16640 8723 16643
rect 9122 16640 9128 16652
rect 8711 16612 9128 16640
rect 8711 16609 8723 16612
rect 8665 16603 8723 16609
rect 9122 16600 9128 16612
rect 9180 16600 9186 16652
rect 9674 16640 9680 16652
rect 9635 16612 9680 16640
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 10410 16640 10416 16652
rect 10371 16612 10416 16640
rect 10410 16600 10416 16612
rect 10468 16640 10474 16652
rect 12161 16643 12219 16649
rect 12161 16640 12173 16643
rect 10468 16612 12173 16640
rect 10468 16600 10474 16612
rect 12161 16609 12173 16612
rect 12207 16609 12219 16643
rect 12360 16640 12388 16680
rect 12161 16603 12219 16609
rect 12268 16612 12388 16640
rect 12428 16643 12486 16649
rect 9953 16575 10011 16581
rect 9953 16541 9965 16575
rect 9999 16541 10011 16575
rect 12268 16572 12296 16612
rect 12428 16609 12440 16643
rect 12474 16640 12486 16643
rect 14182 16640 14188 16652
rect 12474 16612 14188 16640
rect 12474 16609 12486 16612
rect 12428 16603 12486 16609
rect 14182 16600 14188 16612
rect 14240 16600 14246 16652
rect 14461 16643 14519 16649
rect 14461 16609 14473 16643
rect 14507 16609 14519 16643
rect 15654 16640 15660 16652
rect 15615 16612 15660 16640
rect 14461 16603 14519 16609
rect 9953 16535 10011 16541
rect 11431 16544 12296 16572
rect 8386 16436 8392 16448
rect 8347 16408 8392 16436
rect 8386 16396 8392 16408
rect 8444 16396 8450 16448
rect 9968 16436 9996 16535
rect 11431 16436 11459 16544
rect 13906 16532 13912 16584
rect 13964 16572 13970 16584
rect 14476 16572 14504 16603
rect 15654 16600 15660 16612
rect 15712 16600 15718 16652
rect 16390 16640 16396 16652
rect 16351 16612 16396 16640
rect 16390 16600 16396 16612
rect 16448 16600 16454 16652
rect 16945 16643 17003 16649
rect 16945 16609 16957 16643
rect 16991 16640 17003 16643
rect 17034 16640 17040 16652
rect 16991 16612 17040 16640
rect 16991 16609 17003 16612
rect 16945 16603 17003 16609
rect 13964 16544 14504 16572
rect 14553 16575 14611 16581
rect 13964 16532 13970 16544
rect 14553 16541 14565 16575
rect 14599 16541 14611 16575
rect 14553 16535 14611 16541
rect 14737 16575 14795 16581
rect 14737 16541 14749 16575
rect 14783 16572 14795 16575
rect 14918 16572 14924 16584
rect 14783 16544 14924 16572
rect 14783 16541 14795 16544
rect 14737 16535 14795 16541
rect 14274 16464 14280 16516
rect 14332 16504 14338 16516
rect 14568 16504 14596 16535
rect 14918 16532 14924 16544
rect 14976 16532 14982 16584
rect 15470 16532 15476 16584
rect 15528 16572 15534 16584
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 15528 16544 15853 16572
rect 15528 16532 15534 16544
rect 15841 16541 15853 16544
rect 15887 16541 15899 16575
rect 15841 16535 15899 16541
rect 16960 16504 16988 16603
rect 17034 16600 17040 16612
rect 17092 16600 17098 16652
rect 17770 16649 17776 16652
rect 17764 16640 17776 16649
rect 17731 16612 17776 16640
rect 17764 16603 17776 16612
rect 17770 16600 17776 16603
rect 17828 16600 17834 16652
rect 18690 16600 18696 16652
rect 18748 16640 18754 16652
rect 20272 16649 20300 16680
rect 19521 16643 19579 16649
rect 19521 16640 19533 16643
rect 18748 16612 19533 16640
rect 18748 16600 18754 16612
rect 19521 16609 19533 16612
rect 19567 16609 19579 16643
rect 19521 16603 19579 16609
rect 20257 16643 20315 16649
rect 20257 16609 20269 16643
rect 20303 16609 20315 16643
rect 20257 16603 20315 16609
rect 17494 16572 17500 16584
rect 17455 16544 17500 16572
rect 17494 16532 17500 16544
rect 17552 16532 17558 16584
rect 18506 16532 18512 16584
rect 18564 16572 18570 16584
rect 19613 16575 19671 16581
rect 19613 16572 19625 16575
rect 18564 16544 19625 16572
rect 18564 16532 18570 16544
rect 19613 16541 19625 16544
rect 19659 16541 19671 16575
rect 19613 16535 19671 16541
rect 19705 16575 19763 16581
rect 19705 16541 19717 16575
rect 19751 16541 19763 16575
rect 19705 16535 19763 16541
rect 19720 16504 19748 16535
rect 14332 16476 14596 16504
rect 14660 16476 16988 16504
rect 19076 16476 19748 16504
rect 14332 16464 14338 16476
rect 9968 16408 11459 16436
rect 11793 16439 11851 16445
rect 11793 16405 11805 16439
rect 11839 16436 11851 16439
rect 11974 16436 11980 16448
rect 11839 16408 11980 16436
rect 11839 16405 11851 16408
rect 11793 16399 11851 16405
rect 11974 16396 11980 16408
rect 12032 16396 12038 16448
rect 13538 16436 13544 16448
rect 13499 16408 13544 16436
rect 13538 16396 13544 16408
rect 13596 16396 13602 16448
rect 13630 16396 13636 16448
rect 13688 16436 13694 16448
rect 14660 16436 14688 16476
rect 19076 16448 19104 16476
rect 15286 16436 15292 16448
rect 13688 16408 14688 16436
rect 15247 16408 15292 16436
rect 13688 16396 13694 16408
rect 15286 16396 15292 16408
rect 15344 16396 15350 16448
rect 16577 16439 16635 16445
rect 16577 16405 16589 16439
rect 16623 16436 16635 16439
rect 18598 16436 18604 16448
rect 16623 16408 18604 16436
rect 16623 16405 16635 16408
rect 16577 16399 16635 16405
rect 18598 16396 18604 16408
rect 18656 16396 18662 16448
rect 18877 16439 18935 16445
rect 18877 16405 18889 16439
rect 18923 16436 18935 16439
rect 19058 16436 19064 16448
rect 18923 16408 19064 16436
rect 18923 16405 18935 16408
rect 18877 16399 18935 16405
rect 19058 16396 19064 16408
rect 19116 16396 19122 16448
rect 19153 16439 19211 16445
rect 19153 16405 19165 16439
rect 19199 16436 19211 16439
rect 19242 16436 19248 16448
rect 19199 16408 19248 16436
rect 19199 16405 19211 16408
rect 19153 16399 19211 16405
rect 19242 16396 19248 16408
rect 19300 16396 19306 16448
rect 20438 16436 20444 16448
rect 20399 16408 20444 16436
rect 20438 16396 20444 16408
rect 20496 16396 20502 16448
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 7006 16232 7012 16244
rect 6840 16204 7012 16232
rect 6840 16105 6868 16204
rect 7006 16192 7012 16204
rect 7064 16192 7070 16244
rect 8481 16235 8539 16241
rect 8481 16201 8493 16235
rect 8527 16232 8539 16235
rect 9214 16232 9220 16244
rect 8527 16204 9220 16232
rect 8527 16201 8539 16204
rect 8481 16195 8539 16201
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 10410 16232 10416 16244
rect 9324 16204 10416 16232
rect 6825 16099 6883 16105
rect 6825 16065 6837 16099
rect 6871 16065 6883 16099
rect 6825 16059 6883 16065
rect 8386 16056 8392 16108
rect 8444 16096 8450 16108
rect 9033 16099 9091 16105
rect 9033 16096 9045 16099
rect 8444 16068 9045 16096
rect 8444 16056 8450 16068
rect 9033 16065 9045 16068
rect 9079 16065 9091 16099
rect 9033 16059 9091 16065
rect 8294 15988 8300 16040
rect 8352 16028 8358 16040
rect 8941 16031 8999 16037
rect 8941 16028 8953 16031
rect 8352 16000 8953 16028
rect 8352 15988 8358 16000
rect 8941 15997 8953 16000
rect 8987 15997 8999 16031
rect 9324 16028 9352 16204
rect 10410 16192 10416 16204
rect 10468 16192 10474 16244
rect 12710 16192 12716 16244
rect 12768 16232 12774 16244
rect 13722 16232 13728 16244
rect 12768 16204 13728 16232
rect 12768 16192 12774 16204
rect 13722 16192 13728 16204
rect 13780 16192 13786 16244
rect 15565 16235 15623 16241
rect 15565 16201 15577 16235
rect 15611 16232 15623 16235
rect 15654 16232 15660 16244
rect 15611 16204 15660 16232
rect 15611 16201 15623 16204
rect 15565 16195 15623 16201
rect 15654 16192 15660 16204
rect 15712 16192 15718 16244
rect 15838 16192 15844 16244
rect 15896 16232 15902 16244
rect 19613 16235 19671 16241
rect 15896 16204 18184 16232
rect 15896 16192 15902 16204
rect 11624 16136 13676 16164
rect 11624 16105 11652 16136
rect 9401 16099 9459 16105
rect 9401 16065 9413 16099
rect 9447 16096 9459 16099
rect 11609 16099 11667 16105
rect 9447 16068 9628 16096
rect 9447 16065 9459 16068
rect 9401 16059 9459 16065
rect 9493 16031 9551 16037
rect 9493 16028 9505 16031
rect 9324 16000 9505 16028
rect 8941 15991 8999 15997
rect 9493 15997 9505 16000
rect 9539 15997 9551 16031
rect 9600 16028 9628 16068
rect 11609 16065 11621 16099
rect 11655 16065 11667 16099
rect 11609 16059 11667 16065
rect 11793 16099 11851 16105
rect 11793 16065 11805 16099
rect 11839 16096 11851 16099
rect 11882 16096 11888 16108
rect 11839 16068 11888 16096
rect 11839 16065 11851 16068
rect 11793 16059 11851 16065
rect 10318 16028 10324 16040
rect 9600 16000 10324 16028
rect 9493 15991 9551 15997
rect 10318 15988 10324 16000
rect 10376 16028 10382 16040
rect 11624 16028 11652 16059
rect 11882 16056 11888 16068
rect 11940 16096 11946 16108
rect 13538 16096 13544 16108
rect 11940 16068 13544 16096
rect 11940 16056 11946 16068
rect 13538 16056 13544 16068
rect 13596 16056 13602 16108
rect 13648 16096 13676 16136
rect 15102 16124 15108 16176
rect 15160 16164 15166 16176
rect 15160 16136 18092 16164
rect 15160 16124 15166 16136
rect 13648 16068 14044 16096
rect 13262 16028 13268 16040
rect 10376 16000 11652 16028
rect 13223 16000 13268 16028
rect 10376 15988 10382 16000
rect 13262 15988 13268 16000
rect 13320 15988 13326 16040
rect 13357 16031 13415 16037
rect 13357 15997 13369 16031
rect 13403 16028 13415 16031
rect 13446 16028 13452 16040
rect 13403 16000 13452 16028
rect 13403 15997 13415 16000
rect 13357 15991 13415 15997
rect 13446 15988 13452 16000
rect 13504 15988 13510 16040
rect 13909 16031 13967 16037
rect 13909 15997 13921 16031
rect 13955 15997 13967 16031
rect 14016 16028 14044 16068
rect 14918 16056 14924 16108
rect 14976 16096 14982 16108
rect 16206 16096 16212 16108
rect 14976 16068 16212 16096
rect 14976 16056 14982 16068
rect 16206 16056 16212 16068
rect 16264 16096 16270 16108
rect 17218 16096 17224 16108
rect 16264 16068 17224 16096
rect 16264 16056 16270 16068
rect 17218 16056 17224 16068
rect 17276 16056 17282 16108
rect 16025 16031 16083 16037
rect 16025 16028 16037 16031
rect 14016 16000 16037 16028
rect 13909 15991 13967 15997
rect 16025 15997 16037 16000
rect 16071 15997 16083 16031
rect 17770 16028 17776 16040
rect 17731 16000 17776 16028
rect 16025 15991 16083 15997
rect 7092 15963 7150 15969
rect 7092 15929 7104 15963
rect 7138 15960 7150 15963
rect 9760 15963 9818 15969
rect 7138 15932 9536 15960
rect 7138 15929 7150 15932
rect 7092 15923 7150 15929
rect 7466 15852 7472 15904
rect 7524 15892 7530 15904
rect 8205 15895 8263 15901
rect 8205 15892 8217 15895
rect 7524 15864 8217 15892
rect 7524 15852 7530 15864
rect 8205 15861 8217 15864
rect 8251 15861 8263 15895
rect 8205 15855 8263 15861
rect 8849 15895 8907 15901
rect 8849 15861 8861 15895
rect 8895 15892 8907 15895
rect 9401 15895 9459 15901
rect 9401 15892 9413 15895
rect 8895 15864 9413 15892
rect 8895 15861 8907 15864
rect 8849 15855 8907 15861
rect 9401 15861 9413 15864
rect 9447 15861 9459 15895
rect 9508 15892 9536 15932
rect 9760 15929 9772 15963
rect 9806 15960 9818 15963
rect 11054 15960 11060 15972
rect 9806 15932 11060 15960
rect 9806 15929 9818 15932
rect 9760 15923 9818 15929
rect 11054 15920 11060 15932
rect 11112 15920 11118 15972
rect 11517 15963 11575 15969
rect 11517 15929 11529 15963
rect 11563 15960 11575 15963
rect 12342 15960 12348 15972
rect 11563 15932 12348 15960
rect 11563 15929 11575 15932
rect 11517 15923 11575 15929
rect 12342 15920 12348 15932
rect 12400 15960 12406 15972
rect 12400 15932 13391 15960
rect 12400 15920 12406 15932
rect 10594 15892 10600 15904
rect 9508 15864 10600 15892
rect 9401 15855 9459 15861
rect 10594 15852 10600 15864
rect 10652 15892 10658 15904
rect 10873 15895 10931 15901
rect 10873 15892 10885 15895
rect 10652 15864 10885 15892
rect 10652 15852 10658 15864
rect 10873 15861 10885 15864
rect 10919 15861 10931 15895
rect 11146 15892 11152 15904
rect 11107 15864 11152 15892
rect 10873 15855 10931 15861
rect 11146 15852 11152 15864
rect 11204 15852 11210 15904
rect 11790 15852 11796 15904
rect 11848 15892 11854 15904
rect 12897 15895 12955 15901
rect 12897 15892 12909 15895
rect 11848 15864 12909 15892
rect 11848 15852 11854 15864
rect 12897 15861 12909 15864
rect 12943 15861 12955 15895
rect 13363 15892 13391 15932
rect 13538 15920 13544 15972
rect 13596 15960 13602 15972
rect 13924 15960 13952 15991
rect 17770 15988 17776 16000
rect 17828 15988 17834 16040
rect 18064 16037 18092 16136
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 15997 18107 16031
rect 18156 16028 18184 16204
rect 19613 16201 19625 16235
rect 19659 16232 19671 16235
rect 20070 16232 20076 16244
rect 19659 16204 20076 16232
rect 19659 16201 19671 16204
rect 19613 16195 19671 16201
rect 20070 16192 20076 16204
rect 20128 16192 20134 16244
rect 19150 16096 19156 16108
rect 19111 16068 19156 16096
rect 19150 16056 19156 16068
rect 19208 16056 19214 16108
rect 19426 16056 19432 16108
rect 19484 16096 19490 16108
rect 20165 16099 20223 16105
rect 20165 16096 20177 16099
rect 19484 16068 20177 16096
rect 19484 16056 19490 16068
rect 20165 16065 20177 16068
rect 20211 16065 20223 16099
rect 20165 16059 20223 16065
rect 20530 16056 20536 16108
rect 20588 16096 20594 16108
rect 20809 16099 20867 16105
rect 20809 16096 20821 16099
rect 20588 16068 20821 16096
rect 20588 16056 20594 16068
rect 20809 16065 20821 16068
rect 20855 16065 20867 16099
rect 20809 16059 20867 16065
rect 19061 16031 19119 16037
rect 19061 16028 19073 16031
rect 18156 16000 19073 16028
rect 18049 15991 18107 15997
rect 19061 15997 19073 16000
rect 19107 15997 19119 16031
rect 19061 15991 19119 15997
rect 19242 15988 19248 16040
rect 19300 16028 19306 16040
rect 19981 16031 20039 16037
rect 19981 16028 19993 16031
rect 19300 16000 19993 16028
rect 19300 15988 19306 16000
rect 19981 15997 19993 16000
rect 20027 15997 20039 16031
rect 20622 16028 20628 16040
rect 20583 16000 20628 16028
rect 19981 15991 20039 15997
rect 20622 15988 20628 16000
rect 20680 15988 20686 16040
rect 13998 15960 14004 15972
rect 13596 15932 14004 15960
rect 13596 15920 13602 15932
rect 13998 15920 14004 15932
rect 14056 15920 14062 15972
rect 14176 15963 14234 15969
rect 14176 15929 14188 15963
rect 14222 15960 14234 15963
rect 14918 15960 14924 15972
rect 14222 15932 14924 15960
rect 14222 15929 14234 15932
rect 14176 15923 14234 15929
rect 14918 15920 14924 15932
rect 14976 15920 14982 15972
rect 15933 15963 15991 15969
rect 15933 15960 15945 15963
rect 15028 15932 15945 15960
rect 15028 15892 15056 15932
rect 15933 15929 15945 15932
rect 15979 15929 15991 15963
rect 15933 15923 15991 15929
rect 16850 15920 16856 15972
rect 16908 15960 16914 15972
rect 17037 15963 17095 15969
rect 17037 15960 17049 15963
rect 16908 15932 17049 15960
rect 16908 15920 16914 15932
rect 17037 15929 17049 15932
rect 17083 15960 17095 15963
rect 17862 15960 17868 15972
rect 17083 15932 17868 15960
rect 17083 15929 17095 15932
rect 17037 15923 17095 15929
rect 17862 15920 17868 15932
rect 17920 15920 17926 15972
rect 20073 15963 20131 15969
rect 20073 15960 20085 15963
rect 18616 15932 20085 15960
rect 13363 15864 15056 15892
rect 15289 15895 15347 15901
rect 12897 15855 12955 15861
rect 15289 15861 15301 15895
rect 15335 15892 15347 15895
rect 15470 15892 15476 15904
rect 15335 15864 15476 15892
rect 15335 15861 15347 15864
rect 15289 15855 15347 15861
rect 15470 15852 15476 15864
rect 15528 15852 15534 15904
rect 16574 15892 16580 15904
rect 16535 15864 16580 15892
rect 16574 15852 16580 15864
rect 16632 15852 16638 15904
rect 16945 15895 17003 15901
rect 16945 15861 16957 15895
rect 16991 15892 17003 15895
rect 17310 15892 17316 15904
rect 16991 15864 17316 15892
rect 16991 15861 17003 15864
rect 16945 15855 17003 15861
rect 17310 15852 17316 15864
rect 17368 15852 17374 15904
rect 17494 15852 17500 15904
rect 17552 15892 17558 15904
rect 17589 15895 17647 15901
rect 17589 15892 17601 15895
rect 17552 15864 17601 15892
rect 17552 15852 17558 15864
rect 17589 15861 17601 15864
rect 17635 15892 17647 15895
rect 17954 15892 17960 15904
rect 17635 15864 17960 15892
rect 17635 15861 17647 15864
rect 17589 15855 17647 15861
rect 17954 15852 17960 15864
rect 18012 15852 18018 15904
rect 18230 15892 18236 15904
rect 18191 15864 18236 15892
rect 18230 15852 18236 15864
rect 18288 15852 18294 15904
rect 18616 15901 18644 15932
rect 20073 15929 20085 15932
rect 20119 15929 20131 15963
rect 20073 15923 20131 15929
rect 18601 15895 18659 15901
rect 18601 15861 18613 15895
rect 18647 15861 18659 15895
rect 18966 15892 18972 15904
rect 18927 15864 18972 15892
rect 18601 15855 18659 15861
rect 18966 15852 18972 15864
rect 19024 15852 19030 15904
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 7742 15688 7748 15700
rect 7703 15660 7748 15688
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 8113 15691 8171 15697
rect 8113 15657 8125 15691
rect 8159 15688 8171 15691
rect 8570 15688 8576 15700
rect 8159 15660 8576 15688
rect 8159 15657 8171 15660
rect 8113 15651 8171 15657
rect 8570 15648 8576 15660
rect 8628 15648 8634 15700
rect 10045 15691 10103 15697
rect 10045 15657 10057 15691
rect 10091 15688 10103 15691
rect 10410 15688 10416 15700
rect 10091 15660 10416 15688
rect 10091 15657 10103 15660
rect 10045 15651 10103 15657
rect 10410 15648 10416 15660
rect 10468 15648 10474 15700
rect 10689 15691 10747 15697
rect 10689 15657 10701 15691
rect 10735 15688 10747 15691
rect 11146 15688 11152 15700
rect 10735 15660 11152 15688
rect 10735 15657 10747 15660
rect 10689 15651 10747 15657
rect 11146 15648 11152 15660
rect 11204 15648 11210 15700
rect 11790 15688 11796 15700
rect 11751 15660 11796 15688
rect 11790 15648 11796 15660
rect 11848 15648 11854 15700
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 12710 15688 12716 15700
rect 12492 15660 12716 15688
rect 12492 15648 12498 15660
rect 12710 15648 12716 15660
rect 12768 15648 12774 15700
rect 13906 15648 13912 15700
rect 13964 15688 13970 15700
rect 14458 15688 14464 15700
rect 13964 15660 14464 15688
rect 13964 15648 13970 15660
rect 14458 15648 14464 15660
rect 14516 15688 14522 15700
rect 15749 15691 15807 15697
rect 14516 15660 15608 15688
rect 14516 15648 14522 15660
rect 7006 15620 7012 15632
rect 6380 15592 7012 15620
rect 6380 15561 6408 15592
rect 7006 15580 7012 15592
rect 7064 15580 7070 15632
rect 10502 15580 10508 15632
rect 10560 15620 10566 15632
rect 10781 15623 10839 15629
rect 10781 15620 10793 15623
rect 10560 15592 10793 15620
rect 10560 15580 10566 15592
rect 10781 15589 10793 15592
rect 10827 15589 10839 15623
rect 10781 15583 10839 15589
rect 11606 15580 11612 15632
rect 11664 15620 11670 15632
rect 11701 15623 11759 15629
rect 11701 15620 11713 15623
rect 11664 15592 11713 15620
rect 11664 15580 11670 15592
rect 11701 15589 11713 15592
rect 11747 15589 11759 15623
rect 11701 15583 11759 15589
rect 13808 15623 13866 15629
rect 13808 15589 13820 15623
rect 13854 15620 13866 15623
rect 15470 15620 15476 15632
rect 13854 15592 15476 15620
rect 13854 15589 13866 15592
rect 13808 15583 13866 15589
rect 15470 15580 15476 15592
rect 15528 15580 15534 15632
rect 15580 15620 15608 15660
rect 15749 15657 15761 15691
rect 15795 15688 15807 15691
rect 16666 15688 16672 15700
rect 15795 15660 16672 15688
rect 15795 15657 15807 15660
rect 15749 15651 15807 15657
rect 16666 15648 16672 15660
rect 16724 15648 16730 15700
rect 17218 15648 17224 15700
rect 17276 15688 17282 15700
rect 17773 15691 17831 15697
rect 17773 15688 17785 15691
rect 17276 15660 17785 15688
rect 17276 15648 17282 15660
rect 17773 15657 17785 15660
rect 17819 15657 17831 15691
rect 19426 15688 19432 15700
rect 19387 15660 19432 15688
rect 17773 15651 17831 15657
rect 19426 15648 19432 15660
rect 19484 15648 19490 15700
rect 19705 15691 19763 15697
rect 19705 15657 19717 15691
rect 19751 15688 19763 15691
rect 20622 15688 20628 15700
rect 19751 15660 20628 15688
rect 19751 15657 19763 15660
rect 19705 15651 19763 15657
rect 20622 15648 20628 15660
rect 20680 15648 20686 15700
rect 15841 15623 15899 15629
rect 15841 15620 15853 15623
rect 15580 15592 15853 15620
rect 15841 15589 15853 15592
rect 15887 15589 15899 15623
rect 15841 15583 15899 15589
rect 16942 15580 16948 15632
rect 17000 15620 17006 15632
rect 17862 15620 17868 15632
rect 17000 15592 17868 15620
rect 17000 15580 17006 15592
rect 17862 15580 17868 15592
rect 17920 15580 17926 15632
rect 18316 15623 18374 15629
rect 18316 15589 18328 15623
rect 18362 15620 18374 15623
rect 19150 15620 19156 15632
rect 18362 15592 19156 15620
rect 18362 15589 18374 15592
rect 18316 15583 18374 15589
rect 19150 15580 19156 15592
rect 19208 15580 19214 15632
rect 6365 15555 6423 15561
rect 6365 15521 6377 15555
rect 6411 15521 6423 15555
rect 6365 15515 6423 15521
rect 6632 15555 6690 15561
rect 6632 15521 6644 15555
rect 6678 15552 6690 15555
rect 8938 15552 8944 15564
rect 6678 15524 8432 15552
rect 8899 15524 8944 15552
rect 6678 15521 6690 15524
rect 6632 15515 6690 15521
rect 8404 15484 8432 15524
rect 8938 15512 8944 15524
rect 8996 15512 9002 15564
rect 9033 15555 9091 15561
rect 9033 15521 9045 15555
rect 9079 15552 9091 15555
rect 9766 15552 9772 15564
rect 9079 15524 9772 15552
rect 9079 15521 9091 15524
rect 9033 15515 9091 15521
rect 9766 15512 9772 15524
rect 9824 15512 9830 15564
rect 9950 15512 9956 15564
rect 10008 15552 10014 15564
rect 10229 15555 10287 15561
rect 10229 15552 10241 15555
rect 10008 15524 10241 15552
rect 10008 15512 10014 15524
rect 10229 15521 10241 15524
rect 10275 15521 10287 15555
rect 12710 15552 12716 15564
rect 12671 15524 12716 15552
rect 10229 15515 10287 15521
rect 12710 15512 12716 15524
rect 12768 15512 12774 15564
rect 14274 15552 14280 15564
rect 12912 15524 14280 15552
rect 9125 15487 9183 15493
rect 9125 15484 9137 15487
rect 8404 15456 9137 15484
rect 9125 15453 9137 15456
rect 9171 15484 9183 15487
rect 9306 15484 9312 15496
rect 9171 15456 9312 15484
rect 9171 15453 9183 15456
rect 9125 15447 9183 15453
rect 9306 15444 9312 15456
rect 9364 15444 9370 15496
rect 10965 15487 11023 15493
rect 10965 15453 10977 15487
rect 11011 15484 11023 15487
rect 11054 15484 11060 15496
rect 11011 15456 11060 15484
rect 11011 15453 11023 15456
rect 10965 15447 11023 15453
rect 11054 15444 11060 15456
rect 11112 15484 11118 15496
rect 11974 15484 11980 15496
rect 11112 15456 11980 15484
rect 11112 15444 11118 15456
rect 11974 15444 11980 15456
rect 12032 15444 12038 15496
rect 12802 15484 12808 15496
rect 12763 15456 12808 15484
rect 12802 15444 12808 15456
rect 12860 15444 12866 15496
rect 8573 15351 8631 15357
rect 8573 15317 8585 15351
rect 8619 15348 8631 15351
rect 8846 15348 8852 15360
rect 8619 15320 8852 15348
rect 8619 15317 8631 15320
rect 8573 15311 8631 15317
rect 8846 15308 8852 15320
rect 8904 15308 8910 15360
rect 10318 15348 10324 15360
rect 10279 15320 10324 15348
rect 10318 15308 10324 15320
rect 10376 15308 10382 15360
rect 11054 15308 11060 15360
rect 11112 15348 11118 15360
rect 11333 15351 11391 15357
rect 11333 15348 11345 15351
rect 11112 15320 11345 15348
rect 11112 15308 11118 15320
rect 11333 15317 11345 15320
rect 11379 15317 11391 15351
rect 11333 15311 11391 15317
rect 12345 15351 12403 15357
rect 12345 15317 12357 15351
rect 12391 15348 12403 15351
rect 12912 15348 12940 15524
rect 14274 15512 14280 15524
rect 14332 15512 14338 15564
rect 16660 15555 16718 15561
rect 16660 15521 16672 15555
rect 16706 15552 16718 15555
rect 17494 15552 17500 15564
rect 16706 15524 17500 15552
rect 16706 15521 16718 15524
rect 16660 15515 16718 15521
rect 17494 15512 17500 15524
rect 17552 15512 17558 15564
rect 18138 15512 18144 15564
rect 18196 15552 18202 15564
rect 19334 15552 19340 15564
rect 18196 15524 19340 15552
rect 18196 15512 18202 15524
rect 19334 15512 19340 15524
rect 19392 15512 19398 15564
rect 20070 15552 20076 15564
rect 20031 15524 20076 15552
rect 20070 15512 20076 15524
rect 20128 15512 20134 15564
rect 12989 15487 13047 15493
rect 12989 15453 13001 15487
rect 13035 15453 13047 15487
rect 13538 15484 13544 15496
rect 13499 15456 13544 15484
rect 12989 15447 13047 15453
rect 12391 15320 12940 15348
rect 13004 15348 13032 15447
rect 13538 15444 13544 15456
rect 13596 15444 13602 15496
rect 16025 15487 16083 15493
rect 16025 15453 16037 15487
rect 16071 15484 16083 15487
rect 16206 15484 16212 15496
rect 16071 15456 16212 15484
rect 16071 15453 16083 15456
rect 16025 15447 16083 15453
rect 16206 15444 16212 15456
rect 16264 15444 16270 15496
rect 16393 15487 16451 15493
rect 16393 15453 16405 15487
rect 16439 15453 16451 15487
rect 16393 15447 16451 15453
rect 14642 15376 14648 15428
rect 14700 15416 14706 15428
rect 16408 15416 16436 15447
rect 17954 15444 17960 15496
rect 18012 15484 18018 15496
rect 18049 15487 18107 15493
rect 18049 15484 18061 15487
rect 18012 15456 18061 15484
rect 18012 15444 18018 15456
rect 18049 15453 18061 15456
rect 18095 15453 18107 15487
rect 20162 15484 20168 15496
rect 20123 15456 20168 15484
rect 18049 15447 18107 15453
rect 20162 15444 20168 15456
rect 20220 15444 20226 15496
rect 20254 15444 20260 15496
rect 20312 15484 20318 15496
rect 20312 15456 20357 15484
rect 20312 15444 20318 15456
rect 14700 15388 16436 15416
rect 14700 15376 14706 15388
rect 14182 15348 14188 15360
rect 13004 15320 14188 15348
rect 12391 15317 12403 15320
rect 12345 15311 12403 15317
rect 14182 15308 14188 15320
rect 14240 15308 14246 15360
rect 14921 15351 14979 15357
rect 14921 15317 14933 15351
rect 14967 15348 14979 15351
rect 15010 15348 15016 15360
rect 14967 15320 15016 15348
rect 14967 15317 14979 15320
rect 14921 15311 14979 15317
rect 15010 15308 15016 15320
rect 15068 15308 15074 15360
rect 15378 15348 15384 15360
rect 15339 15320 15384 15348
rect 15378 15308 15384 15320
rect 15436 15308 15442 15360
rect 16408 15348 16436 15388
rect 17954 15348 17960 15360
rect 16408 15320 17960 15348
rect 17954 15308 17960 15320
rect 18012 15308 18018 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 9306 15144 9312 15156
rect 9267 15116 9312 15144
rect 9306 15104 9312 15116
rect 9364 15104 9370 15156
rect 9674 15104 9680 15156
rect 9732 15144 9738 15156
rect 10045 15147 10103 15153
rect 10045 15144 10057 15147
rect 9732 15116 10057 15144
rect 9732 15104 9738 15116
rect 10045 15113 10057 15116
rect 10091 15113 10103 15147
rect 10045 15107 10103 15113
rect 12710 15104 12716 15156
rect 12768 15144 12774 15156
rect 12897 15147 12955 15153
rect 12897 15144 12909 15147
rect 12768 15116 12909 15144
rect 12768 15104 12774 15116
rect 12897 15113 12909 15116
rect 12943 15113 12955 15147
rect 18325 15147 18383 15153
rect 18325 15144 18337 15147
rect 12897 15107 12955 15113
rect 13924 15116 18337 15144
rect 9122 15036 9128 15088
rect 9180 15076 9186 15088
rect 13924 15076 13952 15116
rect 18325 15113 18337 15116
rect 18371 15113 18383 15147
rect 18325 15107 18383 15113
rect 18417 15147 18475 15153
rect 18417 15113 18429 15147
rect 18463 15144 18475 15147
rect 20162 15144 20168 15156
rect 18463 15116 20024 15144
rect 20123 15116 20168 15144
rect 18463 15113 18475 15116
rect 18417 15107 18475 15113
rect 18506 15076 18512 15088
rect 9180 15048 13952 15076
rect 18064 15048 18512 15076
rect 9180 15036 9186 15048
rect 6822 14968 6828 15020
rect 6880 15008 6886 15020
rect 7285 15011 7343 15017
rect 7285 15008 7297 15011
rect 6880 14980 7297 15008
rect 6880 14968 6886 14980
rect 7285 14977 7297 14980
rect 7331 14977 7343 15011
rect 7466 15008 7472 15020
rect 7427 14980 7472 15008
rect 7285 14971 7343 14977
rect 7466 14968 7472 14980
rect 7524 14968 7530 15020
rect 10318 14968 10324 15020
rect 10376 15008 10382 15020
rect 10505 15011 10563 15017
rect 10505 15008 10517 15011
rect 10376 14980 10517 15008
rect 10376 14968 10382 14980
rect 10505 14977 10517 14980
rect 10551 14977 10563 15011
rect 10505 14971 10563 14977
rect 10594 14968 10600 15020
rect 10652 15008 10658 15020
rect 11609 15011 11667 15017
rect 10652 14980 10697 15008
rect 10652 14968 10658 14980
rect 11609 14977 11621 15011
rect 11655 14977 11667 15011
rect 11609 14971 11667 14977
rect 7190 14940 7196 14952
rect 7151 14912 7196 14940
rect 7190 14900 7196 14912
rect 7248 14900 7254 14952
rect 7742 14900 7748 14952
rect 7800 14940 7806 14952
rect 7929 14943 7987 14949
rect 7929 14940 7941 14943
rect 7800 14912 7941 14940
rect 7800 14900 7806 14912
rect 7929 14909 7941 14912
rect 7975 14909 7987 14943
rect 7929 14903 7987 14909
rect 10413 14943 10471 14949
rect 10413 14909 10425 14943
rect 10459 14940 10471 14943
rect 11054 14940 11060 14952
rect 10459 14912 11060 14940
rect 10459 14909 10471 14912
rect 10413 14903 10471 14909
rect 11054 14900 11060 14912
rect 11112 14900 11118 14952
rect 11624 14940 11652 14971
rect 12342 14968 12348 15020
rect 12400 15008 12406 15020
rect 12710 15008 12716 15020
rect 12400 14980 12716 15008
rect 12400 14968 12406 14980
rect 12710 14968 12716 14980
rect 12768 14968 12774 15020
rect 13446 15008 13452 15020
rect 13407 14980 13452 15008
rect 13446 14968 13452 14980
rect 13504 14968 13510 15020
rect 15470 14968 15476 15020
rect 15528 15008 15534 15020
rect 18064 15017 18092 15048
rect 18506 15036 18512 15048
rect 18564 15036 18570 15088
rect 19889 15079 19947 15085
rect 19889 15045 19901 15079
rect 19935 15045 19947 15079
rect 19996 15076 20024 15116
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 20073 15079 20131 15085
rect 20073 15076 20085 15079
rect 19996 15048 20085 15076
rect 19889 15039 19947 15045
rect 20073 15045 20085 15048
rect 20119 15045 20131 15079
rect 20073 15039 20131 15045
rect 16117 15011 16175 15017
rect 16117 15008 16129 15011
rect 15528 14980 16129 15008
rect 15528 14968 15534 14980
rect 16117 14977 16129 14980
rect 16163 14977 16175 15011
rect 16117 14971 16175 14977
rect 18049 15011 18107 15017
rect 18049 14977 18061 15011
rect 18095 14977 18107 15011
rect 18049 14971 18107 14977
rect 18325 15011 18383 15017
rect 18325 14977 18337 15011
rect 18371 15008 18383 15011
rect 18414 15008 18420 15020
rect 18371 14980 18420 15008
rect 18371 14977 18383 14980
rect 18325 14971 18383 14977
rect 18414 14968 18420 14980
rect 18472 14968 18478 15020
rect 19904 15008 19932 15039
rect 20346 15008 20352 15020
rect 19904 14980 20352 15008
rect 20346 14968 20352 14980
rect 20404 15008 20410 15020
rect 20717 15011 20775 15017
rect 20717 15008 20729 15011
rect 20404 14980 20729 15008
rect 20404 14968 20410 14980
rect 20717 14977 20729 14980
rect 20763 14977 20775 15011
rect 20717 14971 20775 14977
rect 11698 14940 11704 14952
rect 11624 14912 11704 14940
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 13909 14943 13967 14949
rect 13909 14909 13921 14943
rect 13955 14940 13967 14943
rect 13998 14940 14004 14952
rect 13955 14912 14004 14940
rect 13955 14909 13967 14912
rect 13909 14903 13967 14909
rect 13998 14900 14004 14912
rect 14056 14940 14062 14952
rect 14642 14940 14648 14952
rect 14056 14912 14648 14940
rect 14056 14900 14062 14912
rect 14642 14900 14648 14912
rect 14700 14900 14706 14952
rect 15378 14900 15384 14952
rect 15436 14940 15442 14952
rect 15933 14943 15991 14949
rect 15933 14940 15945 14943
rect 15436 14912 15945 14940
rect 15436 14900 15442 14912
rect 15933 14909 15945 14912
rect 15979 14909 15991 14943
rect 15933 14903 15991 14909
rect 16025 14943 16083 14949
rect 16025 14909 16037 14943
rect 16071 14940 16083 14943
rect 16574 14940 16580 14952
rect 16071 14912 16580 14940
rect 16071 14909 16083 14912
rect 16025 14903 16083 14909
rect 16574 14900 16580 14912
rect 16632 14900 16638 14952
rect 16850 14900 16856 14952
rect 16908 14940 16914 14952
rect 17221 14943 17279 14949
rect 17221 14940 17233 14943
rect 16908 14912 17233 14940
rect 16908 14900 16914 14912
rect 17221 14909 17233 14912
rect 17267 14909 17279 14943
rect 17402 14940 17408 14952
rect 17363 14912 17408 14940
rect 17221 14903 17279 14909
rect 17402 14900 17408 14912
rect 17460 14900 17466 14952
rect 17954 14900 17960 14952
rect 18012 14940 18018 14952
rect 18506 14940 18512 14952
rect 18012 14912 18512 14940
rect 18012 14900 18018 14912
rect 18506 14900 18512 14912
rect 18564 14900 18570 14952
rect 20530 14940 20536 14952
rect 20491 14912 20536 14940
rect 20530 14900 20536 14912
rect 20588 14900 20594 14952
rect 8196 14875 8254 14881
rect 8196 14841 8208 14875
rect 8242 14872 8254 14875
rect 8386 14872 8392 14884
rect 8242 14844 8392 14872
rect 8242 14841 8254 14844
rect 8196 14835 8254 14841
rect 8386 14832 8392 14844
rect 8444 14832 8450 14884
rect 8570 14832 8576 14884
rect 8628 14872 8634 14884
rect 9585 14875 9643 14881
rect 9585 14872 9597 14875
rect 8628 14844 9597 14872
rect 8628 14832 8634 14844
rect 9585 14841 9597 14844
rect 9631 14841 9643 14875
rect 11517 14875 11575 14881
rect 9585 14835 9643 14841
rect 10888 14844 11468 14872
rect 6822 14804 6828 14816
rect 6783 14776 6828 14804
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 8478 14764 8484 14816
rect 8536 14804 8542 14816
rect 10888 14804 10916 14844
rect 11054 14804 11060 14816
rect 8536 14776 10916 14804
rect 11015 14776 11060 14804
rect 8536 14764 8542 14776
rect 11054 14764 11060 14776
rect 11112 14764 11118 14816
rect 11440 14813 11468 14844
rect 11517 14841 11529 14875
rect 11563 14872 11575 14875
rect 12158 14872 12164 14884
rect 11563 14844 12164 14872
rect 11563 14841 11575 14844
rect 11517 14835 11575 14841
rect 12158 14832 12164 14844
rect 12216 14832 12222 14884
rect 14176 14875 14234 14881
rect 14176 14841 14188 14875
rect 14222 14872 14234 14875
rect 15010 14872 15016 14884
rect 14222 14844 15016 14872
rect 14222 14841 14234 14844
rect 14176 14835 14234 14841
rect 15010 14832 15016 14844
rect 15068 14832 15074 14884
rect 16298 14832 16304 14884
rect 16356 14872 16362 14884
rect 18417 14875 18475 14881
rect 18417 14872 18429 14875
rect 16356 14844 18429 14872
rect 16356 14832 16362 14844
rect 18417 14841 18429 14844
rect 18463 14841 18475 14875
rect 18417 14835 18475 14841
rect 18776 14875 18834 14881
rect 18776 14841 18788 14875
rect 18822 14872 18834 14875
rect 19426 14872 19432 14884
rect 18822 14844 19432 14872
rect 18822 14841 18834 14844
rect 18776 14835 18834 14841
rect 19426 14832 19432 14844
rect 19484 14832 19490 14884
rect 22462 14872 22468 14884
rect 19996 14844 22468 14872
rect 11425 14807 11483 14813
rect 11425 14773 11437 14807
rect 11471 14804 11483 14807
rect 11790 14804 11796 14816
rect 11471 14776 11796 14804
rect 11471 14773 11483 14776
rect 11425 14767 11483 14773
rect 11790 14764 11796 14776
rect 11848 14764 11854 14816
rect 13262 14804 13268 14816
rect 13223 14776 13268 14804
rect 13262 14764 13268 14776
rect 13320 14764 13326 14816
rect 13354 14764 13360 14816
rect 13412 14804 13418 14816
rect 13412 14776 13457 14804
rect 13412 14764 13418 14776
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 13998 14804 14004 14816
rect 13872 14776 14004 14804
rect 13872 14764 13878 14776
rect 13998 14764 14004 14776
rect 14056 14764 14062 14816
rect 15102 14764 15108 14816
rect 15160 14804 15166 14816
rect 15289 14807 15347 14813
rect 15289 14804 15301 14807
rect 15160 14776 15301 14804
rect 15160 14764 15166 14776
rect 15289 14773 15301 14776
rect 15335 14773 15347 14807
rect 15289 14767 15347 14773
rect 15565 14807 15623 14813
rect 15565 14773 15577 14807
rect 15611 14804 15623 14807
rect 15654 14804 15660 14816
rect 15611 14776 15660 14804
rect 15611 14773 15623 14776
rect 15565 14767 15623 14773
rect 15654 14764 15660 14776
rect 15712 14764 15718 14816
rect 16577 14807 16635 14813
rect 16577 14773 16589 14807
rect 16623 14804 16635 14807
rect 16666 14804 16672 14816
rect 16623 14776 16672 14804
rect 16623 14773 16635 14776
rect 16577 14767 16635 14773
rect 16666 14764 16672 14776
rect 16724 14764 16730 14816
rect 16942 14764 16948 14816
rect 17000 14804 17006 14816
rect 17037 14807 17095 14813
rect 17037 14804 17049 14807
rect 17000 14776 17049 14804
rect 17000 14764 17006 14776
rect 17037 14773 17049 14776
rect 17083 14773 17095 14807
rect 17037 14767 17095 14773
rect 17589 14807 17647 14813
rect 17589 14773 17601 14807
rect 17635 14804 17647 14807
rect 19996 14804 20024 14844
rect 22462 14832 22468 14844
rect 22520 14832 22526 14884
rect 17635 14776 20024 14804
rect 20073 14807 20131 14813
rect 17635 14773 17647 14776
rect 17589 14767 17647 14773
rect 20073 14773 20085 14807
rect 20119 14804 20131 14807
rect 20625 14807 20683 14813
rect 20625 14804 20637 14807
rect 20119 14776 20637 14804
rect 20119 14773 20131 14776
rect 20073 14767 20131 14773
rect 20625 14773 20637 14776
rect 20671 14773 20683 14807
rect 20625 14767 20683 14773
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 6822 14560 6828 14612
rect 6880 14600 6886 14612
rect 9677 14603 9735 14609
rect 6880 14572 9352 14600
rect 6880 14560 6886 14572
rect 7276 14535 7334 14541
rect 7276 14501 7288 14535
rect 7322 14532 7334 14535
rect 7466 14532 7472 14544
rect 7322 14504 7472 14532
rect 7322 14501 7334 14504
rect 7276 14495 7334 14501
rect 7466 14492 7472 14504
rect 7524 14492 7530 14544
rect 9122 14532 9128 14544
rect 9083 14504 9128 14532
rect 9122 14492 9128 14504
rect 9180 14492 9186 14544
rect 9324 14532 9352 14572
rect 9677 14569 9689 14603
rect 9723 14600 9735 14603
rect 9766 14600 9772 14612
rect 9723 14572 9772 14600
rect 9723 14569 9735 14572
rect 9677 14563 9735 14569
rect 9766 14560 9772 14572
rect 9824 14560 9830 14612
rect 10045 14603 10103 14609
rect 10045 14569 10057 14603
rect 10091 14600 10103 14603
rect 10502 14600 10508 14612
rect 10091 14572 10508 14600
rect 10091 14569 10103 14572
rect 10045 14563 10103 14569
rect 10502 14560 10508 14572
rect 10560 14560 10566 14612
rect 12529 14603 12587 14609
rect 12529 14569 12541 14603
rect 12575 14569 12587 14603
rect 14182 14600 14188 14612
rect 14143 14572 14188 14600
rect 12529 14563 12587 14569
rect 10137 14535 10195 14541
rect 10137 14532 10149 14535
rect 9324 14504 10149 14532
rect 10137 14501 10149 14504
rect 10183 14501 10195 14535
rect 10137 14495 10195 14501
rect 11416 14535 11474 14541
rect 11416 14501 11428 14535
rect 11462 14532 11474 14535
rect 11698 14532 11704 14544
rect 11462 14504 11704 14532
rect 11462 14501 11474 14504
rect 11416 14495 11474 14501
rect 11698 14492 11704 14504
rect 11756 14492 11762 14544
rect 11974 14492 11980 14544
rect 12032 14532 12038 14544
rect 12544 14532 12572 14563
rect 14182 14560 14188 14572
rect 14240 14560 14246 14612
rect 15654 14600 15660 14612
rect 15615 14572 15660 14600
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 16022 14560 16028 14612
rect 16080 14600 16086 14612
rect 18690 14600 18696 14612
rect 16080 14572 18696 14600
rect 16080 14560 16086 14572
rect 18690 14560 18696 14572
rect 18748 14600 18754 14612
rect 19978 14600 19984 14612
rect 18748 14572 19984 14600
rect 18748 14560 18754 14572
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 13072 14535 13130 14541
rect 13072 14532 13084 14535
rect 12032 14504 13084 14532
rect 12032 14492 12038 14504
rect 13072 14501 13084 14504
rect 13118 14532 13130 14535
rect 13446 14532 13452 14544
rect 13118 14504 13452 14532
rect 13118 14501 13130 14504
rect 13072 14495 13130 14501
rect 13446 14492 13452 14504
rect 13504 14492 13510 14544
rect 14292 14504 14596 14532
rect 7009 14467 7067 14473
rect 7009 14433 7021 14467
rect 7055 14464 7067 14467
rect 7742 14464 7748 14476
rect 7055 14436 7748 14464
rect 7055 14433 7067 14436
rect 7009 14427 7067 14433
rect 7742 14424 7748 14436
rect 7800 14424 7806 14476
rect 8846 14464 8852 14476
rect 8807 14436 8852 14464
rect 8846 14424 8852 14436
rect 8904 14424 8910 14476
rect 9306 14424 9312 14476
rect 9364 14464 9370 14476
rect 11057 14467 11115 14473
rect 9364 14436 10364 14464
rect 9364 14424 9370 14436
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14365 10287 14399
rect 10336 14396 10364 14436
rect 11057 14433 11069 14467
rect 11103 14464 11115 14467
rect 12158 14464 12164 14476
rect 11103 14436 12164 14464
rect 11103 14433 11115 14436
rect 11057 14427 11115 14433
rect 12158 14424 12164 14436
rect 12216 14464 12222 14476
rect 12805 14467 12863 14473
rect 12216 14436 12756 14464
rect 12216 14424 12222 14436
rect 11149 14399 11207 14405
rect 11149 14396 11161 14399
rect 10336 14368 11161 14396
rect 10229 14359 10287 14365
rect 11149 14365 11161 14368
rect 11195 14365 11207 14399
rect 11149 14359 11207 14365
rect 8386 14328 8392 14340
rect 8299 14300 8392 14328
rect 8386 14288 8392 14300
rect 8444 14328 8450 14340
rect 8846 14328 8852 14340
rect 8444 14300 8852 14328
rect 8444 14288 8450 14300
rect 8846 14288 8852 14300
rect 8904 14328 8910 14340
rect 10244 14328 10272 14359
rect 8904 14300 10272 14328
rect 8904 14288 8910 14300
rect 9950 14220 9956 14272
rect 10008 14260 10014 14272
rect 10873 14263 10931 14269
rect 10873 14260 10885 14263
rect 10008 14232 10885 14260
rect 10008 14220 10014 14232
rect 10873 14229 10885 14232
rect 10919 14229 10931 14263
rect 12728 14260 12756 14436
rect 12805 14433 12817 14467
rect 12851 14464 12863 14467
rect 12894 14464 12900 14476
rect 12851 14436 12900 14464
rect 12851 14433 12863 14436
rect 12805 14427 12863 14433
rect 12894 14424 12900 14436
rect 12952 14424 12958 14476
rect 13814 14288 13820 14340
rect 13872 14328 13878 14340
rect 14292 14328 14320 14504
rect 14461 14467 14519 14473
rect 14461 14433 14473 14467
rect 14507 14433 14519 14467
rect 14568 14464 14596 14504
rect 15286 14492 15292 14544
rect 15344 14532 15350 14544
rect 15749 14535 15807 14541
rect 15749 14532 15761 14535
rect 15344 14504 15761 14532
rect 15344 14492 15350 14504
rect 15749 14501 15761 14504
rect 15795 14501 15807 14535
rect 15749 14495 15807 14501
rect 17497 14535 17555 14541
rect 17497 14501 17509 14535
rect 17543 14532 17555 14535
rect 17543 14504 18276 14532
rect 17543 14501 17555 14504
rect 17497 14495 17555 14501
rect 16301 14467 16359 14473
rect 16301 14464 16313 14467
rect 14568 14436 16313 14464
rect 14461 14427 14519 14433
rect 16301 14433 16313 14436
rect 16347 14433 16359 14467
rect 16301 14427 16359 14433
rect 16577 14467 16635 14473
rect 16577 14433 16589 14467
rect 16623 14464 16635 14467
rect 17126 14464 17132 14476
rect 16623 14436 17132 14464
rect 16623 14433 16635 14436
rect 16577 14427 16635 14433
rect 13872 14300 14320 14328
rect 14476 14328 14504 14427
rect 17126 14424 17132 14436
rect 17184 14424 17190 14476
rect 17589 14467 17647 14473
rect 17589 14433 17601 14467
rect 17635 14464 17647 14467
rect 17954 14464 17960 14476
rect 17635 14436 17960 14464
rect 17635 14433 17647 14436
rect 17589 14427 17647 14433
rect 17954 14424 17960 14436
rect 18012 14424 18018 14476
rect 14734 14396 14740 14408
rect 14695 14368 14740 14396
rect 14734 14356 14740 14368
rect 14792 14356 14798 14408
rect 15010 14356 15016 14408
rect 15068 14396 15074 14408
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 15068 14368 15853 14396
rect 15068 14356 15074 14368
rect 15841 14365 15853 14368
rect 15887 14365 15899 14399
rect 16206 14396 16212 14408
rect 15841 14359 15899 14365
rect 15948 14368 16212 14396
rect 15289 14331 15347 14337
rect 15289 14328 15301 14331
rect 14476 14300 15301 14328
rect 13872 14288 13878 14300
rect 15289 14297 15301 14300
rect 15335 14297 15347 14331
rect 15289 14291 15347 14297
rect 15654 14288 15660 14340
rect 15712 14328 15718 14340
rect 15948 14328 15976 14368
rect 16206 14356 16212 14368
rect 16264 14356 16270 14408
rect 17773 14399 17831 14405
rect 17773 14365 17785 14399
rect 17819 14396 17831 14399
rect 17862 14396 17868 14408
rect 17819 14368 17868 14396
rect 17819 14365 17831 14368
rect 17773 14359 17831 14365
rect 17862 14356 17868 14368
rect 17920 14356 17926 14408
rect 18248 14396 18276 14504
rect 18506 14492 18512 14544
rect 18564 14532 18570 14544
rect 19236 14535 19294 14541
rect 18564 14504 19012 14532
rect 18564 14492 18570 14504
rect 18414 14464 18420 14476
rect 18375 14436 18420 14464
rect 18414 14424 18420 14436
rect 18472 14424 18478 14476
rect 18984 14473 19012 14504
rect 19236 14501 19248 14535
rect 19282 14532 19294 14535
rect 20346 14532 20352 14544
rect 19282 14504 20352 14532
rect 19282 14501 19294 14504
rect 19236 14495 19294 14501
rect 20346 14492 20352 14504
rect 20404 14492 20410 14544
rect 18969 14467 19027 14473
rect 18969 14433 18981 14467
rect 19015 14433 19027 14467
rect 18969 14427 19027 14433
rect 18506 14396 18512 14408
rect 18248 14368 18512 14396
rect 18506 14356 18512 14368
rect 18564 14356 18570 14408
rect 20162 14356 20168 14408
rect 20220 14396 20226 14408
rect 20901 14399 20959 14405
rect 20901 14396 20913 14399
rect 20220 14368 20913 14396
rect 20220 14356 20226 14368
rect 20901 14365 20913 14368
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 15712 14300 15976 14328
rect 15712 14288 15718 14300
rect 16114 14288 16120 14340
rect 16172 14328 16178 14340
rect 18598 14328 18604 14340
rect 16172 14300 17724 14328
rect 18559 14300 18604 14328
rect 16172 14288 16178 14300
rect 16850 14260 16856 14272
rect 12728 14232 16856 14260
rect 10873 14223 10931 14229
rect 16850 14220 16856 14232
rect 16908 14220 16914 14272
rect 17034 14220 17040 14272
rect 17092 14260 17098 14272
rect 17129 14263 17187 14269
rect 17129 14260 17141 14263
rect 17092 14232 17141 14260
rect 17092 14220 17098 14232
rect 17129 14229 17141 14232
rect 17175 14229 17187 14263
rect 17696 14260 17724 14300
rect 18598 14288 18604 14300
rect 18656 14288 18662 14340
rect 20254 14260 20260 14272
rect 17696 14232 20260 14260
rect 17129 14223 17187 14229
rect 20254 14220 20260 14232
rect 20312 14260 20318 14272
rect 20349 14263 20407 14269
rect 20349 14260 20361 14263
rect 20312 14232 20361 14260
rect 20312 14220 20318 14232
rect 20349 14229 20361 14232
rect 20395 14229 20407 14263
rect 20349 14223 20407 14229
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 8205 14059 8263 14065
rect 8205 14025 8217 14059
rect 8251 14056 8263 14059
rect 8938 14056 8944 14068
rect 8251 14028 8944 14056
rect 8251 14025 8263 14028
rect 8205 14019 8263 14025
rect 8938 14016 8944 14028
rect 8996 14016 9002 14068
rect 11333 14059 11391 14065
rect 11333 14025 11345 14059
rect 11379 14056 11391 14059
rect 12802 14056 12808 14068
rect 11379 14028 12808 14056
rect 11379 14025 11391 14028
rect 11333 14019 11391 14025
rect 12802 14016 12808 14028
rect 12860 14016 12866 14068
rect 13354 14016 13360 14068
rect 13412 14056 13418 14068
rect 14093 14059 14151 14065
rect 14093 14056 14105 14059
rect 13412 14028 14105 14056
rect 13412 14016 13418 14028
rect 14093 14025 14105 14028
rect 14139 14025 14151 14059
rect 14093 14019 14151 14025
rect 14734 14016 14740 14068
rect 14792 14056 14798 14068
rect 19797 14059 19855 14065
rect 14792 14028 19748 14056
rect 14792 14016 14798 14028
rect 7742 13948 7748 14000
rect 7800 13988 7806 14000
rect 16114 13988 16120 14000
rect 7800 13960 9260 13988
rect 7800 13948 7806 13960
rect 9232 13932 9260 13960
rect 10980 13960 16120 13988
rect 8846 13920 8852 13932
rect 8807 13892 8852 13920
rect 8846 13880 8852 13892
rect 8904 13880 8910 13932
rect 9214 13920 9220 13932
rect 9127 13892 9220 13920
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 8570 13852 8576 13864
rect 8531 13824 8576 13852
rect 8570 13812 8576 13824
rect 8628 13812 8634 13864
rect 9484 13855 9542 13861
rect 9484 13821 9496 13855
rect 9530 13852 9542 13855
rect 10980 13852 11008 13960
rect 16114 13948 16120 13960
rect 16172 13948 16178 14000
rect 19720 13988 19748 14028
rect 19797 14025 19809 14059
rect 19843 14056 19855 14059
rect 20070 14056 20076 14068
rect 19843 14028 20076 14056
rect 19843 14025 19855 14028
rect 19797 14019 19855 14025
rect 20070 14016 20076 14028
rect 20128 14016 20134 14068
rect 18156 13960 19104 13988
rect 19720 13960 20576 13988
rect 11054 13880 11060 13932
rect 11112 13920 11118 13932
rect 11793 13923 11851 13929
rect 11793 13920 11805 13923
rect 11112 13892 11805 13920
rect 11112 13880 11118 13892
rect 11793 13889 11805 13892
rect 11839 13889 11851 13923
rect 11974 13920 11980 13932
rect 11935 13892 11980 13920
rect 11793 13883 11851 13889
rect 11974 13880 11980 13892
rect 12032 13880 12038 13932
rect 13081 13923 13139 13929
rect 13081 13889 13093 13923
rect 13127 13920 13139 13923
rect 14182 13920 14188 13932
rect 13127 13892 14188 13920
rect 13127 13889 13139 13892
rect 13081 13883 13139 13889
rect 9530 13824 11008 13852
rect 9530 13821 9542 13824
rect 9484 13815 9542 13821
rect 11698 13812 11704 13864
rect 11756 13852 11762 13864
rect 13096 13852 13124 13883
rect 14182 13880 14188 13892
rect 14240 13920 14246 13932
rect 14737 13923 14795 13929
rect 14737 13920 14749 13923
rect 14240 13892 14749 13920
rect 14240 13880 14246 13892
rect 14737 13889 14749 13892
rect 14783 13920 14795 13923
rect 15102 13920 15108 13932
rect 14783 13892 15108 13920
rect 14783 13889 14795 13892
rect 14737 13883 14795 13889
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 15470 13920 15476 13932
rect 15396 13892 15476 13920
rect 11756 13824 13124 13852
rect 14553 13855 14611 13861
rect 11756 13812 11762 13824
rect 14553 13821 14565 13855
rect 14599 13852 14611 13855
rect 15396 13852 15424 13892
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 15654 13920 15660 13932
rect 15615 13892 15660 13920
rect 15654 13880 15660 13892
rect 15712 13880 15718 13932
rect 17586 13880 17592 13932
rect 17644 13920 17650 13932
rect 18156 13920 18184 13960
rect 17644 13892 18184 13920
rect 18601 13923 18659 13929
rect 17644 13880 17650 13892
rect 18601 13889 18613 13923
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 15562 13852 15568 13864
rect 14599 13824 15424 13852
rect 15523 13824 15568 13852
rect 14599 13821 14611 13824
rect 14553 13815 14611 13821
rect 15562 13812 15568 13824
rect 15620 13812 15626 13864
rect 15838 13812 15844 13864
rect 15896 13852 15902 13864
rect 16117 13855 16175 13861
rect 16117 13852 16129 13855
rect 15896 13824 16129 13852
rect 15896 13812 15902 13824
rect 16117 13821 16129 13824
rect 16163 13852 16175 13855
rect 16384 13855 16442 13861
rect 16163 13824 16344 13852
rect 16163 13821 16175 13824
rect 16117 13815 16175 13821
rect 16316 13796 16344 13824
rect 16384 13821 16396 13855
rect 16430 13852 16442 13855
rect 17862 13852 17868 13864
rect 16430 13824 17868 13852
rect 16430 13821 16442 13824
rect 16384 13815 16442 13821
rect 17862 13812 17868 13824
rect 17920 13852 17926 13864
rect 18616 13852 18644 13883
rect 19076 13861 19104 13960
rect 20346 13920 20352 13932
rect 20307 13892 20352 13920
rect 20346 13880 20352 13892
rect 20404 13880 20410 13932
rect 20548 13920 20576 13960
rect 20622 13948 20628 14000
rect 20680 13988 20686 14000
rect 20993 13991 21051 13997
rect 20993 13988 21005 13991
rect 20680 13960 21005 13988
rect 20680 13948 20686 13960
rect 20993 13957 21005 13960
rect 21039 13957 21051 13991
rect 20993 13951 21051 13957
rect 20548 13892 20852 13920
rect 17920 13824 18644 13852
rect 19061 13855 19119 13861
rect 17920 13812 17926 13824
rect 19061 13821 19073 13855
rect 19107 13821 19119 13855
rect 19061 13815 19119 13821
rect 19337 13855 19395 13861
rect 19337 13821 19349 13855
rect 19383 13852 19395 13855
rect 20714 13852 20720 13864
rect 19383 13824 20720 13852
rect 19383 13821 19395 13824
rect 19337 13815 19395 13821
rect 20714 13812 20720 13824
rect 20772 13812 20778 13864
rect 20824 13861 20852 13892
rect 20809 13855 20867 13861
rect 20809 13821 20821 13855
rect 20855 13821 20867 13855
rect 20809 13815 20867 13821
rect 12986 13744 12992 13796
rect 13044 13784 13050 13796
rect 13722 13784 13728 13796
rect 13044 13756 13728 13784
rect 13044 13744 13050 13756
rect 13722 13744 13728 13756
rect 13780 13744 13786 13796
rect 15010 13744 15016 13796
rect 15068 13784 15074 13796
rect 15473 13787 15531 13793
rect 15473 13784 15485 13787
rect 15068 13756 15485 13784
rect 15068 13744 15074 13756
rect 15473 13753 15485 13756
rect 15519 13753 15531 13787
rect 15473 13747 15531 13753
rect 16298 13744 16304 13796
rect 16356 13744 16362 13796
rect 16666 13744 16672 13796
rect 16724 13784 16730 13796
rect 20162 13784 20168 13796
rect 16724 13756 18092 13784
rect 20123 13756 20168 13784
rect 16724 13744 16730 13756
rect 8665 13719 8723 13725
rect 8665 13685 8677 13719
rect 8711 13716 8723 13719
rect 8846 13716 8852 13728
rect 8711 13688 8852 13716
rect 8711 13685 8723 13688
rect 8665 13679 8723 13685
rect 8846 13676 8852 13688
rect 8904 13676 8910 13728
rect 10594 13716 10600 13728
rect 10555 13688 10600 13716
rect 10594 13676 10600 13688
rect 10652 13676 10658 13728
rect 11701 13719 11759 13725
rect 11701 13685 11713 13719
rect 11747 13716 11759 13719
rect 12437 13719 12495 13725
rect 12437 13716 12449 13719
rect 11747 13688 12449 13716
rect 11747 13685 11759 13688
rect 11701 13679 11759 13685
rect 12437 13685 12449 13688
rect 12483 13685 12495 13719
rect 12802 13716 12808 13728
rect 12763 13688 12808 13716
rect 12437 13679 12495 13685
rect 12802 13676 12808 13688
rect 12860 13676 12866 13728
rect 12897 13719 12955 13725
rect 12897 13685 12909 13719
rect 12943 13716 12955 13719
rect 13078 13716 13084 13728
rect 12943 13688 13084 13716
rect 12943 13685 12955 13688
rect 12897 13679 12955 13685
rect 13078 13676 13084 13688
rect 13136 13676 13142 13728
rect 13633 13719 13691 13725
rect 13633 13685 13645 13719
rect 13679 13716 13691 13719
rect 13814 13716 13820 13728
rect 13679 13688 13820 13716
rect 13679 13685 13691 13688
rect 13633 13679 13691 13685
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 14458 13716 14464 13728
rect 14419 13688 14464 13716
rect 14458 13676 14464 13688
rect 14516 13676 14522 13728
rect 15102 13716 15108 13728
rect 15063 13688 15108 13716
rect 15102 13676 15108 13688
rect 15160 13676 15166 13728
rect 15746 13676 15752 13728
rect 15804 13716 15810 13728
rect 16206 13716 16212 13728
rect 15804 13688 16212 13716
rect 15804 13676 15810 13688
rect 16206 13676 16212 13688
rect 16264 13716 16270 13728
rect 17310 13716 17316 13728
rect 16264 13688 17316 13716
rect 16264 13676 16270 13688
rect 17310 13676 17316 13688
rect 17368 13676 17374 13728
rect 17494 13716 17500 13728
rect 17455 13688 17500 13716
rect 17494 13676 17500 13688
rect 17552 13676 17558 13728
rect 18064 13725 18092 13756
rect 20162 13744 20168 13756
rect 20220 13744 20226 13796
rect 18049 13719 18107 13725
rect 18049 13685 18061 13719
rect 18095 13685 18107 13719
rect 18049 13679 18107 13685
rect 18138 13676 18144 13728
rect 18196 13716 18202 13728
rect 18417 13719 18475 13725
rect 18417 13716 18429 13719
rect 18196 13688 18429 13716
rect 18196 13676 18202 13688
rect 18417 13685 18429 13688
rect 18463 13685 18475 13719
rect 18417 13679 18475 13685
rect 18509 13719 18567 13725
rect 18509 13685 18521 13719
rect 18555 13716 18567 13719
rect 18598 13716 18604 13728
rect 18555 13688 18604 13716
rect 18555 13685 18567 13688
rect 18509 13679 18567 13685
rect 18598 13676 18604 13688
rect 18656 13676 18662 13728
rect 19978 13676 19984 13728
rect 20036 13716 20042 13728
rect 20257 13719 20315 13725
rect 20257 13716 20269 13719
rect 20036 13688 20269 13716
rect 20036 13676 20042 13688
rect 20257 13685 20269 13688
rect 20303 13685 20315 13719
rect 20257 13679 20315 13685
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 9214 13472 9220 13524
rect 9272 13512 9278 13524
rect 9309 13515 9367 13521
rect 9309 13512 9321 13515
rect 9272 13484 9321 13512
rect 9272 13472 9278 13484
rect 9309 13481 9321 13484
rect 9355 13481 9367 13515
rect 9309 13475 9367 13481
rect 9769 13515 9827 13521
rect 9769 13481 9781 13515
rect 9815 13512 9827 13515
rect 11146 13512 11152 13524
rect 9815 13484 11152 13512
rect 9815 13481 9827 13484
rect 9769 13475 9827 13481
rect 11146 13472 11152 13484
rect 11204 13472 11210 13524
rect 12437 13515 12495 13521
rect 12437 13481 12449 13515
rect 12483 13512 12495 13515
rect 12986 13512 12992 13524
rect 12483 13484 12992 13512
rect 12483 13481 12495 13484
rect 12437 13475 12495 13481
rect 12986 13472 12992 13484
rect 13044 13472 13050 13524
rect 13262 13472 13268 13524
rect 13320 13512 13326 13524
rect 13449 13515 13507 13521
rect 13449 13512 13461 13515
rect 13320 13484 13461 13512
rect 13320 13472 13326 13484
rect 13449 13481 13461 13484
rect 13495 13481 13507 13515
rect 13814 13512 13820 13524
rect 13775 13484 13820 13512
rect 13449 13475 13507 13481
rect 13814 13472 13820 13484
rect 13872 13472 13878 13524
rect 15102 13512 15108 13524
rect 14016 13484 15108 13512
rect 11977 13447 12035 13453
rect 11977 13413 11989 13447
rect 12023 13444 12035 13447
rect 12618 13444 12624 13456
rect 12023 13416 12624 13444
rect 12023 13413 12035 13416
rect 11977 13407 12035 13413
rect 12618 13404 12624 13416
rect 12676 13404 12682 13456
rect 12897 13447 12955 13453
rect 12897 13413 12909 13447
rect 12943 13444 12955 13447
rect 14016 13444 14044 13484
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 15657 13515 15715 13521
rect 15657 13481 15669 13515
rect 15703 13512 15715 13515
rect 16114 13512 16120 13524
rect 15703 13484 16120 13512
rect 15703 13481 15715 13484
rect 15657 13475 15715 13481
rect 16114 13472 16120 13484
rect 16172 13512 16178 13524
rect 16390 13512 16396 13524
rect 16172 13484 16396 13512
rect 16172 13472 16178 13484
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 17862 13512 17868 13524
rect 17823 13484 17868 13512
rect 17862 13472 17868 13484
rect 17920 13472 17926 13524
rect 17954 13472 17960 13524
rect 18012 13512 18018 13524
rect 18141 13515 18199 13521
rect 18141 13512 18153 13515
rect 18012 13484 18153 13512
rect 18012 13472 18018 13484
rect 18141 13481 18153 13484
rect 18187 13481 18199 13515
rect 18141 13475 18199 13481
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19613 13515 19671 13521
rect 19613 13512 19625 13515
rect 19392 13484 19625 13512
rect 19392 13472 19398 13484
rect 19613 13481 19625 13484
rect 19659 13481 19671 13515
rect 20438 13512 20444 13524
rect 20399 13484 20444 13512
rect 19613 13475 19671 13481
rect 20438 13472 20444 13484
rect 20496 13472 20502 13524
rect 12943 13416 14044 13444
rect 12943 13413 12955 13416
rect 12897 13407 12955 13413
rect 14090 13404 14096 13456
rect 14148 13404 14154 13456
rect 14737 13447 14795 13453
rect 14737 13413 14749 13447
rect 14783 13444 14795 13447
rect 14783 13416 16252 13444
rect 14783 13413 14795 13416
rect 14737 13407 14795 13413
rect 9493 13379 9551 13385
rect 9493 13345 9505 13379
rect 9539 13376 9551 13379
rect 9950 13376 9956 13388
rect 9539 13348 9956 13376
rect 9539 13345 9551 13348
rect 9493 13339 9551 13345
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 10134 13376 10140 13388
rect 10095 13348 10140 13376
rect 10134 13336 10140 13348
rect 10192 13336 10198 13388
rect 11701 13379 11759 13385
rect 11701 13345 11713 13379
rect 11747 13345 11759 13379
rect 11701 13339 11759 13345
rect 10226 13308 10232 13320
rect 10187 13280 10232 13308
rect 10226 13268 10232 13280
rect 10284 13268 10290 13320
rect 10318 13268 10324 13320
rect 10376 13308 10382 13320
rect 10376 13280 10421 13308
rect 10376 13268 10382 13280
rect 11716 13240 11744 13339
rect 12434 13336 12440 13388
rect 12492 13376 12498 13388
rect 12805 13379 12863 13385
rect 12805 13376 12817 13379
rect 12492 13348 12817 13376
rect 12492 13336 12498 13348
rect 12805 13345 12817 13348
rect 12851 13345 12863 13379
rect 12805 13339 12863 13345
rect 13538 13336 13544 13388
rect 13596 13376 13602 13388
rect 13909 13379 13967 13385
rect 13909 13376 13921 13379
rect 13596 13348 13921 13376
rect 13596 13336 13602 13348
rect 13909 13345 13921 13348
rect 13955 13376 13967 13379
rect 14108 13376 14136 13404
rect 13955 13348 14136 13376
rect 13955 13345 13967 13348
rect 13909 13339 13967 13345
rect 14274 13336 14280 13388
rect 14332 13376 14338 13388
rect 14461 13379 14519 13385
rect 14461 13376 14473 13379
rect 14332 13348 14473 13376
rect 14332 13336 14338 13348
rect 14461 13345 14473 13348
rect 14507 13345 14519 13379
rect 14461 13339 14519 13345
rect 15378 13336 15384 13388
rect 15436 13376 15442 13388
rect 15749 13379 15807 13385
rect 15749 13376 15761 13379
rect 15436 13348 15761 13376
rect 15436 13336 15442 13348
rect 15749 13345 15761 13348
rect 15795 13345 15807 13379
rect 15749 13339 15807 13345
rect 13081 13311 13139 13317
rect 13081 13277 13093 13311
rect 13127 13308 13139 13311
rect 14093 13311 14151 13317
rect 13127 13280 13860 13308
rect 13127 13277 13139 13280
rect 13081 13271 13139 13277
rect 13722 13240 13728 13252
rect 11716 13212 13728 13240
rect 13722 13200 13728 13212
rect 13780 13200 13786 13252
rect 13832 13240 13860 13280
rect 14093 13277 14105 13311
rect 14139 13308 14151 13311
rect 14182 13308 14188 13320
rect 14139 13280 14188 13308
rect 14139 13277 14151 13280
rect 14093 13271 14151 13277
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 14918 13268 14924 13320
rect 14976 13308 14982 13320
rect 15841 13311 15899 13317
rect 15841 13308 15853 13311
rect 14976 13280 15853 13308
rect 14976 13268 14982 13280
rect 15841 13277 15853 13280
rect 15887 13277 15899 13311
rect 16224 13308 16252 13416
rect 16684 13416 20300 13444
rect 16298 13336 16304 13388
rect 16356 13376 16362 13388
rect 16485 13379 16543 13385
rect 16485 13376 16497 13379
rect 16356 13348 16497 13376
rect 16356 13336 16362 13348
rect 16485 13345 16497 13348
rect 16531 13345 16543 13379
rect 16684 13376 16712 13416
rect 16485 13339 16543 13345
rect 16592 13348 16712 13376
rect 16752 13379 16810 13385
rect 16592 13308 16620 13348
rect 16752 13345 16764 13379
rect 16798 13376 16810 13379
rect 16798 13348 17632 13376
rect 16798 13345 16810 13348
rect 16752 13339 16810 13345
rect 16224 13280 16620 13308
rect 15841 13271 15899 13277
rect 16022 13240 16028 13252
rect 13832 13212 16028 13240
rect 16022 13200 16028 13212
rect 16080 13240 16086 13252
rect 16390 13240 16396 13252
rect 16080 13212 16396 13240
rect 16080 13200 16086 13212
rect 16390 13200 16396 13212
rect 16448 13200 16454 13252
rect 17604 13240 17632 13348
rect 17862 13336 17868 13388
rect 17920 13376 17926 13388
rect 18509 13379 18567 13385
rect 18509 13376 18521 13379
rect 17920 13348 18521 13376
rect 17920 13336 17926 13348
rect 18509 13345 18521 13348
rect 18555 13376 18567 13379
rect 19150 13376 19156 13388
rect 18555 13348 19156 13376
rect 18555 13345 18567 13348
rect 18509 13339 18567 13345
rect 19150 13336 19156 13348
rect 19208 13336 19214 13388
rect 19334 13336 19340 13388
rect 19392 13376 19398 13388
rect 20272 13385 20300 13416
rect 19521 13379 19579 13385
rect 19521 13376 19533 13379
rect 19392 13348 19533 13376
rect 19392 13336 19398 13348
rect 19521 13345 19533 13348
rect 19567 13345 19579 13379
rect 19521 13339 19579 13345
rect 20257 13379 20315 13385
rect 20257 13345 20269 13379
rect 20303 13345 20315 13379
rect 20257 13339 20315 13345
rect 17678 13268 17684 13320
rect 17736 13308 17742 13320
rect 18601 13311 18659 13317
rect 18601 13308 18613 13311
rect 17736 13280 18613 13308
rect 17736 13268 17742 13280
rect 18601 13277 18613 13280
rect 18647 13277 18659 13311
rect 18601 13271 18659 13277
rect 18690 13268 18696 13320
rect 18748 13308 18754 13320
rect 19705 13311 19763 13317
rect 18748 13280 18793 13308
rect 18748 13268 18754 13280
rect 19705 13277 19717 13311
rect 19751 13277 19763 13311
rect 19705 13271 19763 13277
rect 18708 13240 18736 13268
rect 17604 13212 18736 13240
rect 19426 13200 19432 13252
rect 19484 13240 19490 13252
rect 19720 13240 19748 13271
rect 19484 13212 19748 13240
rect 19484 13200 19490 13212
rect 12986 13132 12992 13184
rect 13044 13172 13050 13184
rect 15289 13175 15347 13181
rect 15289 13172 15301 13175
rect 13044 13144 15301 13172
rect 13044 13132 13050 13144
rect 15289 13141 15301 13144
rect 15335 13141 15347 13175
rect 15289 13135 15347 13141
rect 16850 13132 16856 13184
rect 16908 13172 16914 13184
rect 19153 13175 19211 13181
rect 19153 13172 19165 13175
rect 16908 13144 19165 13172
rect 16908 13132 16914 13144
rect 19153 13141 19165 13144
rect 19199 13141 19211 13175
rect 19153 13135 19211 13141
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 12069 12971 12127 12977
rect 12069 12937 12081 12971
rect 12115 12968 12127 12971
rect 12158 12968 12164 12980
rect 12115 12940 12164 12968
rect 12115 12937 12127 12940
rect 12069 12931 12127 12937
rect 12158 12928 12164 12940
rect 12216 12928 12222 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 12492 12940 12537 12968
rect 12492 12928 12498 12940
rect 14458 12928 14464 12980
rect 14516 12968 14522 12980
rect 14516 12940 16344 12968
rect 14516 12928 14522 12940
rect 12894 12860 12900 12912
rect 12952 12900 12958 12912
rect 13262 12900 13268 12912
rect 12952 12872 13268 12900
rect 12952 12860 12958 12872
rect 13262 12860 13268 12872
rect 13320 12900 13326 12912
rect 13320 12872 13492 12900
rect 13320 12860 13326 12872
rect 9214 12792 9220 12844
rect 9272 12832 9278 12844
rect 9309 12835 9367 12841
rect 9309 12832 9321 12835
rect 9272 12804 9321 12832
rect 9272 12792 9278 12804
rect 9309 12801 9321 12804
rect 9355 12801 9367 12835
rect 9309 12795 9367 12801
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12801 11575 12835
rect 12986 12832 12992 12844
rect 11517 12795 11575 12801
rect 12912 12804 12992 12832
rect 9576 12767 9634 12773
rect 9576 12733 9588 12767
rect 9622 12764 9634 12767
rect 10594 12764 10600 12776
rect 9622 12736 10600 12764
rect 9622 12733 9634 12736
rect 9576 12727 9634 12733
rect 10594 12724 10600 12736
rect 10652 12764 10658 12776
rect 11532 12764 11560 12795
rect 10652 12736 11560 12764
rect 12253 12767 12311 12773
rect 10652 12724 10658 12736
rect 12253 12733 12265 12767
rect 12299 12764 12311 12767
rect 12434 12764 12440 12776
rect 12299 12736 12440 12764
rect 12299 12733 12311 12736
rect 12253 12727 12311 12733
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 12912 12773 12940 12804
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 13464 12841 13492 12872
rect 14642 12860 14648 12912
rect 14700 12900 14706 12912
rect 14700 12872 15148 12900
rect 14700 12860 14706 12872
rect 15120 12841 15148 12872
rect 13081 12835 13139 12841
rect 13081 12801 13093 12835
rect 13127 12801 13139 12835
rect 13081 12795 13139 12801
rect 13449 12835 13507 12841
rect 13449 12801 13461 12835
rect 13495 12801 13507 12835
rect 13449 12795 13507 12801
rect 15105 12835 15163 12841
rect 15105 12801 15117 12835
rect 15151 12801 15163 12835
rect 16316 12832 16344 12940
rect 16390 12928 16396 12980
rect 16448 12968 16454 12980
rect 16485 12971 16543 12977
rect 16485 12968 16497 12971
rect 16448 12940 16497 12968
rect 16448 12928 16454 12940
rect 16485 12937 16497 12940
rect 16531 12937 16543 12971
rect 18049 12971 18107 12977
rect 16485 12931 16543 12937
rect 17236 12940 17632 12968
rect 16761 12903 16819 12909
rect 16761 12869 16773 12903
rect 16807 12900 16819 12903
rect 17236 12900 17264 12940
rect 16807 12872 17264 12900
rect 17604 12900 17632 12940
rect 18049 12937 18061 12971
rect 18095 12968 18107 12971
rect 18506 12968 18512 12980
rect 18095 12940 18512 12968
rect 18095 12937 18107 12940
rect 18049 12931 18107 12937
rect 18506 12928 18512 12940
rect 18564 12928 18570 12980
rect 18690 12928 18696 12980
rect 18748 12968 18754 12980
rect 20441 12971 20499 12977
rect 20441 12968 20453 12971
rect 18748 12940 20453 12968
rect 18748 12928 18754 12940
rect 20441 12937 20453 12940
rect 20487 12937 20499 12971
rect 20898 12968 20904 12980
rect 20859 12940 20904 12968
rect 20441 12931 20499 12937
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 18598 12900 18604 12912
rect 17604 12872 18604 12900
rect 16807 12869 16819 12872
rect 16761 12863 16819 12869
rect 18598 12860 18604 12872
rect 18656 12860 18662 12912
rect 18708 12841 18736 12928
rect 17221 12835 17279 12841
rect 17221 12832 17233 12835
rect 16316 12804 17233 12832
rect 15105 12795 15163 12801
rect 17221 12801 17233 12804
rect 17267 12801 17279 12835
rect 17221 12795 17279 12801
rect 17405 12835 17463 12841
rect 17405 12801 17417 12835
rect 17451 12832 17463 12835
rect 18693 12835 18751 12841
rect 18693 12832 18705 12835
rect 17451 12804 18705 12832
rect 17451 12801 17463 12804
rect 17405 12795 17463 12801
rect 18693 12801 18705 12804
rect 18739 12801 18751 12835
rect 18693 12795 18751 12801
rect 12897 12767 12955 12773
rect 12897 12733 12909 12767
rect 12943 12733 12955 12767
rect 13096 12764 13124 12795
rect 15120 12764 15148 12795
rect 15194 12764 15200 12776
rect 13096 12736 14872 12764
rect 15120 12736 15200 12764
rect 12897 12727 12955 12733
rect 10502 12656 10508 12708
rect 10560 12696 10566 12708
rect 11333 12699 11391 12705
rect 11333 12696 11345 12699
rect 10560 12668 11345 12696
rect 10560 12656 10566 12668
rect 11333 12665 11345 12668
rect 11379 12696 11391 12699
rect 13078 12696 13084 12708
rect 11379 12668 13084 12696
rect 11379 12665 11391 12668
rect 11333 12659 11391 12665
rect 13078 12656 13084 12668
rect 13136 12656 13142 12708
rect 13716 12699 13774 12705
rect 13716 12665 13728 12699
rect 13762 12696 13774 12699
rect 14734 12696 14740 12708
rect 13762 12668 14740 12696
rect 13762 12665 13774 12668
rect 13716 12659 13774 12665
rect 14734 12656 14740 12668
rect 14792 12656 14798 12708
rect 10594 12588 10600 12640
rect 10652 12628 10658 12640
rect 10689 12631 10747 12637
rect 10689 12628 10701 12631
rect 10652 12600 10701 12628
rect 10652 12588 10658 12600
rect 10689 12597 10701 12600
rect 10735 12597 10747 12631
rect 10962 12628 10968 12640
rect 10923 12600 10968 12628
rect 10689 12591 10747 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 11425 12631 11483 12637
rect 11425 12597 11437 12631
rect 11471 12628 11483 12631
rect 11698 12628 11704 12640
rect 11471 12600 11704 12628
rect 11471 12597 11483 12600
rect 11425 12591 11483 12597
rect 11698 12588 11704 12600
rect 11756 12628 11762 12640
rect 12066 12628 12072 12640
rect 11756 12600 12072 12628
rect 11756 12588 11762 12600
rect 12066 12588 12072 12600
rect 12124 12588 12130 12640
rect 12805 12631 12863 12637
rect 12805 12597 12817 12631
rect 12851 12628 12863 12631
rect 14550 12628 14556 12640
rect 12851 12600 14556 12628
rect 12851 12597 12863 12600
rect 12805 12591 12863 12597
rect 14550 12588 14556 12600
rect 14608 12588 14614 12640
rect 14844 12637 14872 12736
rect 15194 12724 15200 12736
rect 15252 12724 15258 12776
rect 15372 12767 15430 12773
rect 15372 12733 15384 12767
rect 15418 12764 15430 12767
rect 15654 12764 15660 12776
rect 15418 12736 15660 12764
rect 15418 12733 15430 12736
rect 15372 12727 15430 12733
rect 14829 12631 14887 12637
rect 14829 12597 14841 12631
rect 14875 12628 14887 12631
rect 15387 12628 15415 12727
rect 15654 12724 15660 12736
rect 15712 12724 15718 12776
rect 15930 12724 15936 12776
rect 15988 12764 15994 12776
rect 17129 12767 17187 12773
rect 17129 12764 17141 12767
rect 15988 12736 17141 12764
rect 15988 12724 15994 12736
rect 17129 12733 17141 12736
rect 17175 12733 17187 12767
rect 17236 12764 17264 12795
rect 18046 12764 18052 12776
rect 17236 12736 18052 12764
rect 17129 12727 17187 12733
rect 18046 12724 18052 12736
rect 18104 12724 18110 12776
rect 18322 12724 18328 12776
rect 18380 12764 18386 12776
rect 19061 12767 19119 12773
rect 19061 12764 19073 12767
rect 18380 12736 19073 12764
rect 18380 12724 18386 12736
rect 19061 12733 19073 12736
rect 19107 12733 19119 12767
rect 20714 12764 20720 12776
rect 20675 12736 20720 12764
rect 19061 12727 19119 12733
rect 20714 12724 20720 12736
rect 20772 12724 20778 12776
rect 17678 12696 17684 12708
rect 17144 12668 17684 12696
rect 17144 12640 17172 12668
rect 17678 12656 17684 12668
rect 17736 12656 17742 12708
rect 18230 12656 18236 12708
rect 18288 12696 18294 12708
rect 18509 12699 18567 12705
rect 18509 12696 18521 12699
rect 18288 12668 18521 12696
rect 18288 12656 18294 12668
rect 18509 12665 18521 12668
rect 18555 12665 18567 12699
rect 18509 12659 18567 12665
rect 18690 12656 18696 12708
rect 18748 12696 18754 12708
rect 18874 12696 18880 12708
rect 18748 12668 18880 12696
rect 18748 12656 18754 12668
rect 18874 12656 18880 12668
rect 18932 12656 18938 12708
rect 19328 12699 19386 12705
rect 19328 12665 19340 12699
rect 19374 12696 19386 12699
rect 19610 12696 19616 12708
rect 19374 12668 19616 12696
rect 19374 12665 19386 12668
rect 19328 12659 19386 12665
rect 19610 12656 19616 12668
rect 19668 12656 19674 12708
rect 14875 12600 15415 12628
rect 14875 12597 14887 12600
rect 14829 12591 14887 12597
rect 17126 12588 17132 12640
rect 17184 12588 17190 12640
rect 17310 12588 17316 12640
rect 17368 12628 17374 12640
rect 18417 12631 18475 12637
rect 18417 12628 18429 12631
rect 17368 12600 18429 12628
rect 17368 12588 17374 12600
rect 18417 12597 18429 12600
rect 18463 12597 18475 12631
rect 18417 12591 18475 12597
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 10045 12427 10103 12433
rect 10045 12393 10057 12427
rect 10091 12424 10103 12427
rect 10226 12424 10232 12436
rect 10091 12396 10232 12424
rect 10091 12393 10103 12396
rect 10045 12387 10103 12393
rect 10226 12384 10232 12396
rect 10284 12384 10290 12436
rect 10505 12427 10563 12433
rect 10505 12393 10517 12427
rect 10551 12424 10563 12427
rect 10962 12424 10968 12436
rect 10551 12396 10968 12424
rect 10551 12393 10563 12396
rect 10505 12387 10563 12393
rect 10962 12384 10968 12396
rect 11020 12384 11026 12436
rect 11790 12384 11796 12436
rect 11848 12424 11854 12436
rect 13906 12424 13912 12436
rect 11848 12396 13912 12424
rect 11848 12384 11854 12396
rect 13906 12384 13912 12396
rect 13964 12384 13970 12436
rect 14550 12384 14556 12436
rect 14608 12424 14614 12436
rect 14737 12427 14795 12433
rect 14737 12424 14749 12427
rect 14608 12396 14749 12424
rect 14608 12384 14614 12396
rect 14737 12393 14749 12396
rect 14783 12393 14795 12427
rect 14737 12387 14795 12393
rect 15194 12384 15200 12436
rect 15252 12424 15258 12436
rect 15473 12427 15531 12433
rect 15473 12424 15485 12427
rect 15252 12396 15485 12424
rect 15252 12384 15258 12396
rect 15473 12393 15485 12396
rect 15519 12424 15531 12427
rect 15746 12424 15752 12436
rect 15519 12396 15752 12424
rect 15519 12393 15531 12396
rect 15473 12387 15531 12393
rect 15746 12384 15752 12396
rect 15804 12384 15810 12436
rect 16117 12427 16175 12433
rect 16117 12393 16129 12427
rect 16163 12424 16175 12427
rect 16850 12424 16856 12436
rect 16163 12396 16856 12424
rect 16163 12393 16175 12396
rect 16117 12387 16175 12393
rect 16850 12384 16856 12396
rect 16908 12384 16914 12436
rect 17221 12427 17279 12433
rect 17221 12424 17233 12427
rect 17144 12396 17233 12424
rect 8846 12316 8852 12368
rect 8904 12356 8910 12368
rect 16758 12356 16764 12368
rect 8904 12328 16764 12356
rect 8904 12316 8910 12328
rect 16758 12316 16764 12328
rect 16816 12316 16822 12368
rect 17034 12316 17040 12368
rect 17092 12356 17098 12368
rect 17144 12356 17172 12396
rect 17221 12393 17233 12396
rect 17267 12393 17279 12427
rect 17221 12387 17279 12393
rect 18046 12384 18052 12436
rect 18104 12424 18110 12436
rect 18966 12424 18972 12436
rect 18104 12396 18972 12424
rect 18104 12384 18110 12396
rect 18966 12384 18972 12396
rect 19024 12384 19030 12436
rect 19886 12384 19892 12436
rect 19944 12424 19950 12436
rect 20441 12427 20499 12433
rect 20441 12424 20453 12427
rect 19944 12396 20453 12424
rect 19944 12384 19950 12396
rect 20441 12393 20453 12396
rect 20487 12393 20499 12427
rect 20441 12387 20499 12393
rect 17092 12328 17172 12356
rect 17092 12316 17098 12328
rect 18506 12316 18512 12368
rect 18564 12356 18570 12368
rect 19150 12356 19156 12368
rect 18564 12328 19156 12356
rect 18564 12316 18570 12328
rect 19150 12316 19156 12328
rect 19208 12316 19214 12368
rect 19518 12316 19524 12368
rect 19576 12356 19582 12368
rect 20070 12356 20076 12368
rect 19576 12328 20076 12356
rect 19576 12316 19582 12328
rect 20070 12316 20076 12328
rect 20128 12316 20134 12368
rect 10410 12288 10416 12300
rect 10371 12260 10416 12288
rect 10410 12248 10416 12260
rect 10468 12248 10474 12300
rect 11692 12291 11750 12297
rect 11692 12257 11704 12291
rect 11738 12288 11750 12291
rect 12250 12288 12256 12300
rect 11738 12260 12256 12288
rect 11738 12257 11750 12260
rect 11692 12251 11750 12257
rect 12250 12248 12256 12260
rect 12308 12248 12314 12300
rect 13348 12291 13406 12297
rect 13348 12288 13360 12291
rect 13004 12260 13360 12288
rect 10594 12220 10600 12232
rect 10555 12192 10600 12220
rect 10594 12180 10600 12192
rect 10652 12180 10658 12232
rect 10870 12180 10876 12232
rect 10928 12220 10934 12232
rect 11425 12223 11483 12229
rect 11425 12220 11437 12223
rect 10928 12192 11437 12220
rect 10928 12180 10934 12192
rect 11425 12189 11437 12192
rect 11471 12189 11483 12223
rect 11425 12183 11483 12189
rect 8754 12112 8760 12164
rect 8812 12152 8818 12164
rect 9214 12152 9220 12164
rect 8812 12124 9220 12152
rect 8812 12112 8818 12124
rect 9214 12112 9220 12124
rect 9272 12152 9278 12164
rect 10888 12152 10916 12180
rect 9272 12124 10916 12152
rect 12805 12155 12863 12161
rect 9272 12112 9278 12124
rect 12805 12121 12817 12155
rect 12851 12152 12863 12155
rect 13004 12152 13032 12260
rect 13348 12257 13360 12260
rect 13394 12288 13406 12291
rect 14918 12288 14924 12300
rect 13394 12260 14924 12288
rect 13394 12257 13406 12260
rect 13348 12251 13406 12257
rect 14918 12248 14924 12260
rect 14976 12248 14982 12300
rect 15657 12291 15715 12297
rect 15657 12257 15669 12291
rect 15703 12288 15715 12291
rect 16942 12288 16948 12300
rect 15703 12260 16948 12288
rect 15703 12257 15715 12260
rect 15657 12251 15715 12257
rect 16942 12248 16948 12260
rect 17000 12248 17006 12300
rect 17129 12291 17187 12297
rect 17129 12288 17141 12291
rect 17052 12260 17141 12288
rect 13078 12180 13084 12232
rect 13136 12220 13142 12232
rect 16209 12223 16267 12229
rect 13136 12192 13181 12220
rect 13136 12180 13142 12192
rect 16209 12189 16221 12223
rect 16255 12189 16267 12223
rect 16209 12183 16267 12189
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12220 16451 12223
rect 16482 12220 16488 12232
rect 16439 12192 16488 12220
rect 16439 12189 16451 12192
rect 16393 12183 16451 12189
rect 12851 12124 13032 12152
rect 14461 12155 14519 12161
rect 12851 12121 12863 12124
rect 12805 12115 12863 12121
rect 14461 12121 14473 12155
rect 14507 12152 14519 12155
rect 15010 12152 15016 12164
rect 14507 12124 15016 12152
rect 14507 12121 14519 12124
rect 14461 12115 14519 12121
rect 15010 12112 15016 12124
rect 15068 12112 15074 12164
rect 16224 12152 16252 12183
rect 16482 12180 16488 12192
rect 16540 12180 16546 12232
rect 16666 12180 16672 12232
rect 16724 12220 16730 12232
rect 17052 12220 17080 12260
rect 17129 12257 17141 12260
rect 17175 12257 17187 12291
rect 17129 12251 17187 12257
rect 17678 12248 17684 12300
rect 17736 12288 17742 12300
rect 17773 12291 17831 12297
rect 17773 12288 17785 12291
rect 17736 12260 17785 12288
rect 17736 12248 17742 12260
rect 17773 12257 17785 12260
rect 17819 12257 17831 12291
rect 17773 12251 17831 12257
rect 18322 12248 18328 12300
rect 18380 12288 18386 12300
rect 18601 12291 18659 12297
rect 18601 12288 18613 12291
rect 18380 12260 18613 12288
rect 18380 12248 18386 12260
rect 18601 12257 18613 12260
rect 18647 12257 18659 12291
rect 18601 12251 18659 12257
rect 18868 12291 18926 12297
rect 18868 12257 18880 12291
rect 18914 12288 18926 12291
rect 19426 12288 19432 12300
rect 18914 12260 19432 12288
rect 18914 12257 18926 12260
rect 18868 12251 18926 12257
rect 19426 12248 19432 12260
rect 19484 12248 19490 12300
rect 20257 12291 20315 12297
rect 20257 12257 20269 12291
rect 20303 12257 20315 12291
rect 20257 12251 20315 12257
rect 16724 12192 17080 12220
rect 17405 12223 17463 12229
rect 16724 12180 16730 12192
rect 17405 12189 17417 12223
rect 17451 12220 17463 12223
rect 17494 12220 17500 12232
rect 17451 12192 17500 12220
rect 17451 12189 17463 12192
rect 17405 12183 17463 12189
rect 17494 12180 17500 12192
rect 17552 12180 17558 12232
rect 18046 12220 18052 12232
rect 18007 12192 18052 12220
rect 18046 12180 18052 12192
rect 18104 12180 18110 12232
rect 18598 12152 18604 12164
rect 16224 12124 18604 12152
rect 18598 12112 18604 12124
rect 18656 12112 18662 12164
rect 20272 12152 20300 12251
rect 19536 12124 20300 12152
rect 13998 12044 14004 12096
rect 14056 12084 14062 12096
rect 15378 12084 15384 12096
rect 14056 12056 15384 12084
rect 14056 12044 14062 12056
rect 15378 12044 15384 12056
rect 15436 12044 15442 12096
rect 15749 12087 15807 12093
rect 15749 12053 15761 12087
rect 15795 12084 15807 12087
rect 16114 12084 16120 12096
rect 15795 12056 16120 12084
rect 15795 12053 15807 12056
rect 15749 12047 15807 12053
rect 16114 12044 16120 12056
rect 16172 12044 16178 12096
rect 16761 12087 16819 12093
rect 16761 12053 16773 12087
rect 16807 12084 16819 12087
rect 17586 12084 17592 12096
rect 16807 12056 17592 12084
rect 16807 12053 16819 12056
rect 16761 12047 16819 12053
rect 17586 12044 17592 12056
rect 17644 12044 17650 12096
rect 18874 12044 18880 12096
rect 18932 12084 18938 12096
rect 19536 12084 19564 12124
rect 19978 12084 19984 12096
rect 18932 12056 19564 12084
rect 19939 12056 19984 12084
rect 18932 12044 18938 12056
rect 19978 12044 19984 12056
rect 20036 12044 20042 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 10134 11840 10140 11892
rect 10192 11880 10198 11892
rect 10413 11883 10471 11889
rect 10413 11880 10425 11883
rect 10192 11852 10425 11880
rect 10192 11840 10198 11852
rect 10413 11849 10425 11852
rect 10459 11849 10471 11883
rect 10413 11843 10471 11849
rect 11054 11840 11060 11892
rect 11112 11880 11118 11892
rect 12802 11880 12808 11892
rect 11112 11852 12808 11880
rect 11112 11840 11118 11852
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 13722 11840 13728 11892
rect 13780 11880 13786 11892
rect 14369 11883 14427 11889
rect 14369 11880 14381 11883
rect 13780 11852 14381 11880
rect 13780 11840 13786 11852
rect 14369 11849 14381 11852
rect 14415 11849 14427 11883
rect 16666 11880 16672 11892
rect 14369 11843 14427 11849
rect 14476 11852 16672 11880
rect 11698 11772 11704 11824
rect 11756 11812 11762 11824
rect 14476 11812 14504 11852
rect 16666 11840 16672 11852
rect 16724 11840 16730 11892
rect 18598 11880 18604 11892
rect 18559 11852 18604 11880
rect 18598 11840 18604 11852
rect 18656 11840 18662 11892
rect 19058 11840 19064 11892
rect 19116 11880 19122 11892
rect 19116 11852 20300 11880
rect 19116 11840 19122 11852
rect 11756 11784 14504 11812
rect 11756 11772 11762 11784
rect 19150 11772 19156 11824
rect 19208 11812 19214 11824
rect 19610 11812 19616 11824
rect 19208 11784 19616 11812
rect 19208 11772 19214 11784
rect 19610 11772 19616 11784
rect 19668 11812 19674 11824
rect 19978 11812 19984 11824
rect 19668 11784 19984 11812
rect 19668 11772 19674 11784
rect 19978 11772 19984 11784
rect 20036 11772 20042 11824
rect 8754 11744 8760 11756
rect 8715 11716 8760 11744
rect 8754 11704 8760 11716
rect 8812 11704 8818 11756
rect 10965 11747 11023 11753
rect 10965 11713 10977 11747
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 9024 11679 9082 11685
rect 9024 11645 9036 11679
rect 9070 11676 9082 11679
rect 10594 11676 10600 11688
rect 9070 11648 10600 11676
rect 9070 11645 9082 11648
rect 9024 11639 9082 11645
rect 10594 11636 10600 11648
rect 10652 11676 10658 11688
rect 10980 11676 11008 11707
rect 12250 11704 12256 11756
rect 12308 11744 12314 11756
rect 13173 11747 13231 11753
rect 13173 11744 13185 11747
rect 12308 11716 13185 11744
rect 12308 11704 12314 11716
rect 13173 11713 13185 11716
rect 13219 11744 13231 11747
rect 14093 11747 14151 11753
rect 14093 11744 14105 11747
rect 13219 11716 14105 11744
rect 13219 11713 13231 11716
rect 13173 11707 13231 11713
rect 14093 11713 14105 11716
rect 14139 11713 14151 11747
rect 14918 11744 14924 11756
rect 14879 11716 14924 11744
rect 14093 11707 14151 11713
rect 14918 11704 14924 11716
rect 14976 11704 14982 11756
rect 15746 11744 15752 11756
rect 15707 11716 15752 11744
rect 15746 11704 15752 11716
rect 15804 11704 15810 11756
rect 17405 11747 17463 11753
rect 17405 11713 17417 11747
rect 17451 11744 17463 11747
rect 17954 11744 17960 11756
rect 17451 11716 17960 11744
rect 17451 11713 17463 11716
rect 17405 11707 17463 11713
rect 17954 11704 17960 11716
rect 18012 11704 18018 11756
rect 19245 11747 19303 11753
rect 19245 11713 19257 11747
rect 19291 11744 19303 11747
rect 19426 11744 19432 11756
rect 19291 11716 19432 11744
rect 19291 11713 19303 11716
rect 19245 11707 19303 11713
rect 19426 11704 19432 11716
rect 19484 11704 19490 11756
rect 20162 11744 20168 11756
rect 20123 11716 20168 11744
rect 20162 11704 20168 11716
rect 20220 11704 20226 11756
rect 20272 11744 20300 11852
rect 20809 11747 20867 11753
rect 20809 11744 20821 11747
rect 20272 11716 20821 11744
rect 20809 11713 20821 11716
rect 20855 11713 20867 11747
rect 20809 11707 20867 11713
rect 16022 11685 16028 11688
rect 14829 11679 14887 11685
rect 14829 11676 14841 11679
rect 10652 11648 11008 11676
rect 12544 11648 14841 11676
rect 10652 11636 10658 11648
rect 10781 11611 10839 11617
rect 10781 11577 10793 11611
rect 10827 11608 10839 11611
rect 11425 11611 11483 11617
rect 11425 11608 11437 11611
rect 10827 11580 11437 11608
rect 10827 11577 10839 11580
rect 10781 11571 10839 11577
rect 11425 11577 11437 11580
rect 11471 11577 11483 11611
rect 11425 11571 11483 11577
rect 9858 11500 9864 11552
rect 9916 11540 9922 11552
rect 10137 11543 10195 11549
rect 10137 11540 10149 11543
rect 9916 11512 10149 11540
rect 9916 11500 9922 11512
rect 10137 11509 10149 11512
rect 10183 11540 10195 11543
rect 10318 11540 10324 11552
rect 10183 11512 10324 11540
rect 10183 11509 10195 11512
rect 10137 11503 10195 11509
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 10873 11543 10931 11549
rect 10873 11509 10885 11543
rect 10919 11540 10931 11543
rect 12342 11540 12348 11552
rect 10919 11512 12348 11540
rect 10919 11509 10931 11512
rect 10873 11503 10931 11509
rect 12342 11500 12348 11512
rect 12400 11500 12406 11552
rect 12544 11549 12572 11648
rect 14829 11645 14841 11648
rect 14875 11645 14887 11679
rect 14829 11639 14887 11645
rect 16016 11639 16028 11685
rect 16080 11676 16086 11688
rect 20625 11679 20683 11685
rect 20625 11676 20637 11679
rect 16080 11648 16116 11676
rect 17696 11648 20637 11676
rect 16022 11636 16028 11639
rect 16080 11636 16086 11648
rect 14737 11611 14795 11617
rect 14737 11608 14749 11611
rect 13556 11580 14749 11608
rect 12529 11543 12587 11549
rect 12529 11509 12541 11543
rect 12575 11509 12587 11543
rect 12894 11540 12900 11552
rect 12855 11512 12900 11540
rect 12529 11503 12587 11509
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 12986 11500 12992 11552
rect 13044 11540 13050 11552
rect 13556 11549 13584 11580
rect 14737 11577 14749 11580
rect 14783 11577 14795 11611
rect 14737 11571 14795 11577
rect 16114 11568 16120 11620
rect 16172 11608 16178 11620
rect 17696 11608 17724 11648
rect 20625 11645 20637 11648
rect 20671 11645 20683 11679
rect 20625 11639 20683 11645
rect 16172 11580 17724 11608
rect 18141 11611 18199 11617
rect 16172 11568 16178 11580
rect 18141 11577 18153 11611
rect 18187 11608 18199 11611
rect 19334 11608 19340 11620
rect 18187 11580 19340 11608
rect 18187 11577 18199 11580
rect 18141 11571 18199 11577
rect 19334 11568 19340 11580
rect 19392 11568 19398 11620
rect 19518 11568 19524 11620
rect 19576 11608 19582 11620
rect 19981 11611 20039 11617
rect 19576 11580 19748 11608
rect 19576 11568 19582 11580
rect 13541 11543 13599 11549
rect 13044 11512 13089 11540
rect 13044 11500 13050 11512
rect 13541 11509 13553 11543
rect 13587 11509 13599 11543
rect 13541 11503 13599 11509
rect 13630 11500 13636 11552
rect 13688 11540 13694 11552
rect 13909 11543 13967 11549
rect 13909 11540 13921 11543
rect 13688 11512 13921 11540
rect 13688 11500 13694 11512
rect 13909 11509 13921 11512
rect 13955 11509 13967 11543
rect 13909 11503 13967 11509
rect 13998 11500 14004 11552
rect 14056 11540 14062 11552
rect 17126 11540 17132 11552
rect 14056 11512 14101 11540
rect 17087 11512 17132 11540
rect 14056 11500 14062 11512
rect 17126 11500 17132 11512
rect 17184 11500 17190 11552
rect 18966 11540 18972 11552
rect 18927 11512 18972 11540
rect 18966 11500 18972 11512
rect 19024 11500 19030 11552
rect 19058 11500 19064 11552
rect 19116 11540 19122 11552
rect 19610 11540 19616 11552
rect 19116 11512 19161 11540
rect 19571 11512 19616 11540
rect 19116 11500 19122 11512
rect 19610 11500 19616 11512
rect 19668 11500 19674 11552
rect 19720 11540 19748 11580
rect 19981 11577 19993 11611
rect 20027 11608 20039 11611
rect 20806 11608 20812 11620
rect 20027 11580 20812 11608
rect 20027 11577 20039 11580
rect 19981 11571 20039 11577
rect 20806 11568 20812 11580
rect 20864 11568 20870 11620
rect 20073 11543 20131 11549
rect 20073 11540 20085 11543
rect 19720 11512 20085 11540
rect 20073 11509 20085 11512
rect 20119 11509 20131 11543
rect 20073 11503 20131 11509
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 12250 11336 12256 11348
rect 12211 11308 12256 11336
rect 12250 11296 12256 11308
rect 12308 11296 12314 11348
rect 12526 11296 12532 11348
rect 12584 11336 12590 11348
rect 13262 11336 13268 11348
rect 12584 11308 13268 11336
rect 12584 11296 12590 11308
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 13722 11296 13728 11348
rect 13780 11336 13786 11348
rect 15194 11336 15200 11348
rect 13780 11308 15200 11336
rect 13780 11296 13786 11308
rect 15194 11296 15200 11308
rect 15252 11296 15258 11348
rect 15289 11339 15347 11345
rect 15289 11305 15301 11339
rect 15335 11336 15347 11339
rect 15562 11336 15568 11348
rect 15335 11308 15568 11336
rect 15335 11305 15347 11308
rect 15289 11299 15347 11305
rect 15562 11296 15568 11308
rect 15620 11296 15626 11348
rect 15657 11339 15715 11345
rect 15657 11305 15669 11339
rect 15703 11336 15715 11339
rect 16114 11336 16120 11348
rect 15703 11308 16120 11336
rect 15703 11305 15715 11308
rect 15657 11299 15715 11305
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 18874 11336 18880 11348
rect 16316 11308 18880 11336
rect 8196 11271 8254 11277
rect 8196 11237 8208 11271
rect 8242 11268 8254 11271
rect 9858 11268 9864 11280
rect 8242 11240 9864 11268
rect 8242 11237 8254 11240
rect 8196 11231 8254 11237
rect 9858 11228 9864 11240
rect 9916 11228 9922 11280
rect 9953 11271 10011 11277
rect 9953 11237 9965 11271
rect 9999 11268 10011 11271
rect 16316 11268 16344 11308
rect 18874 11296 18880 11308
rect 18932 11296 18938 11348
rect 19426 11296 19432 11348
rect 19484 11336 19490 11348
rect 20533 11339 20591 11345
rect 20533 11336 20545 11339
rect 19484 11308 20545 11336
rect 19484 11296 19490 11308
rect 20533 11305 20545 11308
rect 20579 11305 20591 11339
rect 20533 11299 20591 11305
rect 9999 11240 16344 11268
rect 16844 11271 16902 11277
rect 9999 11237 10011 11240
rect 9953 11231 10011 11237
rect 16844 11237 16856 11271
rect 16890 11268 16902 11271
rect 17126 11268 17132 11280
rect 16890 11240 17132 11268
rect 16890 11237 16902 11240
rect 16844 11231 16902 11237
rect 17126 11228 17132 11240
rect 17184 11268 17190 11280
rect 17494 11268 17500 11280
rect 17184 11240 17500 11268
rect 17184 11228 17190 11240
rect 17494 11228 17500 11240
rect 17552 11228 17558 11280
rect 18690 11268 18696 11280
rect 18651 11240 18696 11268
rect 18690 11228 18696 11240
rect 18748 11228 18754 11280
rect 19702 11268 19708 11280
rect 18800 11240 19708 11268
rect 7929 11203 7987 11209
rect 7929 11169 7941 11203
rect 7975 11200 7987 11203
rect 8754 11200 8760 11212
rect 7975 11172 8760 11200
rect 7975 11169 7987 11172
rect 7929 11163 7987 11169
rect 8754 11160 8760 11172
rect 8812 11160 8818 11212
rect 9674 11200 9680 11212
rect 9635 11172 9680 11200
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 10870 11200 10876 11212
rect 10831 11172 10876 11200
rect 10870 11160 10876 11172
rect 10928 11160 10934 11212
rect 11140 11203 11198 11209
rect 11140 11169 11152 11203
rect 11186 11200 11198 11203
rect 11974 11200 11980 11212
rect 11186 11172 11980 11200
rect 11186 11169 11198 11172
rect 11140 11163 11198 11169
rect 11974 11160 11980 11172
rect 12032 11160 12038 11212
rect 12989 11203 13047 11209
rect 12989 11169 13001 11203
rect 13035 11200 13047 11203
rect 18417 11203 18475 11209
rect 13035 11172 17632 11200
rect 13035 11169 13047 11172
rect 12989 11163 13047 11169
rect 10410 11092 10416 11144
rect 10468 11132 10474 11144
rect 10778 11132 10784 11144
rect 10468 11104 10784 11132
rect 10468 11092 10474 11104
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 12618 11092 12624 11144
rect 12676 11132 12682 11144
rect 13722 11132 13728 11144
rect 12676 11104 13728 11132
rect 12676 11092 12682 11104
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 15746 11132 15752 11144
rect 15707 11104 15752 11132
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 15841 11135 15899 11141
rect 15841 11101 15853 11135
rect 15887 11101 15899 11135
rect 15841 11095 15899 11101
rect 12434 11024 12440 11076
rect 12492 11064 12498 11076
rect 13170 11064 13176 11076
rect 12492 11036 13176 11064
rect 12492 11024 12498 11036
rect 13170 11024 13176 11036
rect 13228 11064 13234 11076
rect 14277 11067 14335 11073
rect 14277 11064 14289 11067
rect 13228 11036 14289 11064
rect 13228 11024 13234 11036
rect 14277 11033 14289 11036
rect 14323 11033 14335 11067
rect 14277 11027 14335 11033
rect 15010 11024 15016 11076
rect 15068 11064 15074 11076
rect 15856 11064 15884 11095
rect 16298 11092 16304 11144
rect 16356 11132 16362 11144
rect 16577 11135 16635 11141
rect 16577 11132 16589 11135
rect 16356 11104 16589 11132
rect 16356 11092 16362 11104
rect 16577 11101 16589 11104
rect 16623 11101 16635 11135
rect 17604 11132 17632 11172
rect 18417 11169 18429 11203
rect 18463 11200 18475 11203
rect 18598 11200 18604 11212
rect 18463 11172 18604 11200
rect 18463 11169 18475 11172
rect 18417 11163 18475 11169
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 18800 11132 18828 11240
rect 19702 11228 19708 11240
rect 19760 11228 19766 11280
rect 19426 11209 19432 11212
rect 19420 11200 19432 11209
rect 19387 11172 19432 11200
rect 19420 11163 19432 11172
rect 19426 11160 19432 11163
rect 19484 11160 19490 11212
rect 17604 11104 18828 11132
rect 16577 11095 16635 11101
rect 18874 11092 18880 11144
rect 18932 11132 18938 11144
rect 19153 11135 19211 11141
rect 19153 11132 19165 11135
rect 18932 11104 19165 11132
rect 18932 11092 18938 11104
rect 19153 11101 19165 11104
rect 19199 11101 19211 11135
rect 19153 11095 19211 11101
rect 15068 11036 15884 11064
rect 15068 11024 15074 11036
rect 17586 11024 17592 11076
rect 17644 11064 17650 11076
rect 17644 11036 18819 11064
rect 17644 11024 17650 11036
rect 9306 10996 9312 11008
rect 9267 10968 9312 10996
rect 9306 10956 9312 10968
rect 9364 10956 9370 11008
rect 15286 10956 15292 11008
rect 15344 10996 15350 11008
rect 17678 10996 17684 11008
rect 15344 10968 17684 10996
rect 15344 10956 15350 10968
rect 17678 10956 17684 10968
rect 17736 10956 17742 11008
rect 17954 10996 17960 11008
rect 17915 10968 17960 10996
rect 17954 10956 17960 10968
rect 18012 10956 18018 11008
rect 18506 10956 18512 11008
rect 18564 10996 18570 11008
rect 18690 10996 18696 11008
rect 18564 10968 18696 10996
rect 18564 10956 18570 10968
rect 18690 10956 18696 10968
rect 18748 10956 18754 11008
rect 18791 10996 18819 11036
rect 19518 10996 19524 11008
rect 18791 10968 19524 10996
rect 19518 10956 19524 10968
rect 19576 10956 19582 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 8938 10752 8944 10804
rect 8996 10792 9002 10804
rect 9398 10792 9404 10804
rect 8996 10764 9404 10792
rect 8996 10752 9002 10764
rect 9398 10752 9404 10764
rect 9456 10792 9462 10804
rect 12437 10795 12495 10801
rect 12437 10792 12449 10795
rect 9456 10764 12449 10792
rect 9456 10752 9462 10764
rect 12437 10761 12449 10764
rect 12483 10761 12495 10795
rect 12437 10755 12495 10761
rect 12894 10752 12900 10804
rect 12952 10792 12958 10804
rect 13357 10795 13415 10801
rect 13357 10792 13369 10795
rect 12952 10764 13369 10792
rect 12952 10752 12958 10764
rect 13357 10761 13369 10764
rect 13403 10761 13415 10795
rect 13357 10755 13415 10761
rect 14461 10795 14519 10801
rect 14461 10761 14473 10795
rect 14507 10792 14519 10795
rect 15102 10792 15108 10804
rect 14507 10764 15108 10792
rect 14507 10761 14519 10764
rect 14461 10755 14519 10761
rect 15102 10752 15108 10764
rect 15160 10752 15166 10804
rect 15286 10792 15292 10804
rect 15247 10764 15292 10792
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 15930 10752 15936 10804
rect 15988 10752 15994 10804
rect 18049 10795 18107 10801
rect 18049 10792 18061 10795
rect 16224 10764 18061 10792
rect 12529 10727 12587 10733
rect 12529 10693 12541 10727
rect 12575 10724 12587 10727
rect 13998 10724 14004 10736
rect 12575 10696 14004 10724
rect 12575 10693 12587 10696
rect 12529 10687 12587 10693
rect 13998 10684 14004 10696
rect 14056 10684 14062 10736
rect 15948 10724 15976 10752
rect 15120 10696 15976 10724
rect 15120 10668 15148 10696
rect 9306 10616 9312 10668
rect 9364 10656 9370 10668
rect 10413 10659 10471 10665
rect 10413 10656 10425 10659
rect 9364 10628 10425 10656
rect 9364 10616 9370 10628
rect 10413 10625 10425 10628
rect 10459 10625 10471 10659
rect 11422 10656 11428 10668
rect 11383 10628 11428 10656
rect 10413 10619 10471 10625
rect 11422 10616 11428 10628
rect 11480 10616 11486 10668
rect 11974 10616 11980 10668
rect 12032 10656 12038 10668
rect 13081 10659 13139 10665
rect 13081 10656 13093 10659
rect 12032 10628 13093 10656
rect 12032 10616 12038 10628
rect 13081 10625 13093 10628
rect 13127 10656 13139 10659
rect 13354 10656 13360 10668
rect 13127 10628 13360 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 13354 10616 13360 10628
rect 13412 10656 13418 10668
rect 13909 10659 13967 10665
rect 13909 10656 13921 10659
rect 13412 10628 13921 10656
rect 13412 10616 13418 10628
rect 13909 10625 13921 10628
rect 13955 10625 13967 10659
rect 15010 10656 15016 10668
rect 14971 10628 15016 10656
rect 13909 10619 13967 10625
rect 15010 10616 15016 10628
rect 15068 10616 15074 10668
rect 15102 10616 15108 10668
rect 15160 10616 15166 10668
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10656 15991 10659
rect 16117 10659 16175 10665
rect 16117 10656 16129 10659
rect 15979 10628 16129 10656
rect 15979 10625 15991 10628
rect 15933 10619 15991 10625
rect 16117 10625 16129 10628
rect 16163 10625 16175 10659
rect 16117 10619 16175 10625
rect 7742 10548 7748 10600
rect 7800 10588 7806 10600
rect 8205 10591 8263 10597
rect 8205 10588 8217 10591
rect 7800 10560 8217 10588
rect 7800 10548 7806 10560
rect 8205 10557 8217 10560
rect 8251 10557 8263 10591
rect 8205 10551 8263 10557
rect 8472 10591 8530 10597
rect 8472 10557 8484 10591
rect 8518 10588 8530 10591
rect 9324 10588 9352 10616
rect 8518 10560 9352 10588
rect 10321 10591 10379 10597
rect 8518 10557 8530 10560
rect 8472 10551 8530 10557
rect 10321 10557 10333 10591
rect 10367 10588 10379 10591
rect 10502 10588 10508 10600
rect 10367 10560 10508 10588
rect 10367 10557 10379 10560
rect 10321 10551 10379 10557
rect 10502 10548 10508 10560
rect 10560 10588 10566 10600
rect 12069 10591 12127 10597
rect 10560 10560 12020 10588
rect 10560 10548 10566 10560
rect 9306 10480 9312 10532
rect 9364 10520 9370 10532
rect 10229 10523 10287 10529
rect 10229 10520 10241 10523
rect 9364 10492 10241 10520
rect 9364 10480 9370 10492
rect 10229 10489 10241 10492
rect 10275 10489 10287 10523
rect 10229 10483 10287 10489
rect 11054 10480 11060 10532
rect 11112 10520 11118 10532
rect 11241 10523 11299 10529
rect 11241 10520 11253 10523
rect 11112 10492 11253 10520
rect 11112 10480 11118 10492
rect 11241 10489 11253 10492
rect 11287 10489 11299 10523
rect 11992 10520 12020 10560
rect 12069 10557 12081 10591
rect 12115 10588 12127 10591
rect 13630 10588 13636 10600
rect 12115 10560 13636 10588
rect 12115 10557 12127 10560
rect 12069 10551 12127 10557
rect 13630 10548 13636 10560
rect 13688 10548 13694 10600
rect 13725 10591 13783 10597
rect 13725 10557 13737 10591
rect 13771 10588 13783 10591
rect 14458 10588 14464 10600
rect 13771 10560 14464 10588
rect 13771 10557 13783 10560
rect 13725 10551 13783 10557
rect 14458 10548 14464 10560
rect 14516 10588 14522 10600
rect 14642 10588 14648 10600
rect 14516 10560 14648 10588
rect 14516 10548 14522 10560
rect 14642 10548 14648 10560
rect 14700 10548 14706 10600
rect 14829 10591 14887 10597
rect 14829 10557 14841 10591
rect 14875 10588 14887 10591
rect 15378 10588 15384 10600
rect 14875 10560 15384 10588
rect 14875 10557 14887 10560
rect 14829 10551 14887 10557
rect 15378 10548 15384 10560
rect 15436 10548 15442 10600
rect 15657 10591 15715 10597
rect 15657 10557 15669 10591
rect 15703 10588 15715 10591
rect 16224 10588 16252 10764
rect 18049 10761 18061 10764
rect 18095 10761 18107 10795
rect 18049 10755 18107 10761
rect 18601 10659 18659 10665
rect 18601 10625 18613 10659
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 15703 10560 16252 10588
rect 15703 10557 15715 10560
rect 15657 10551 15715 10557
rect 16298 10548 16304 10600
rect 16356 10588 16362 10600
rect 16568 10591 16626 10597
rect 16356 10560 16401 10588
rect 16356 10548 16362 10560
rect 16568 10557 16580 10591
rect 16614 10588 16626 10591
rect 17954 10588 17960 10600
rect 16614 10560 17960 10588
rect 16614 10557 16626 10560
rect 16568 10551 16626 10557
rect 17954 10548 17960 10560
rect 18012 10588 18018 10600
rect 18506 10588 18512 10600
rect 18012 10560 18512 10588
rect 18012 10548 18018 10560
rect 18506 10548 18512 10560
rect 18564 10588 18570 10600
rect 18616 10588 18644 10619
rect 18564 10560 18644 10588
rect 18564 10548 18570 10560
rect 18874 10548 18880 10600
rect 18932 10588 18938 10600
rect 19705 10591 19763 10597
rect 19705 10588 19717 10591
rect 18932 10560 19717 10588
rect 18932 10548 18938 10560
rect 19705 10557 19717 10560
rect 19751 10557 19763 10591
rect 19705 10551 19763 10557
rect 12158 10520 12164 10532
rect 11992 10492 12164 10520
rect 11241 10483 11299 10489
rect 12158 10480 12164 10492
rect 12216 10480 12222 10532
rect 12437 10523 12495 10529
rect 12437 10489 12449 10523
rect 12483 10520 12495 10523
rect 16022 10520 16028 10532
rect 12483 10492 16028 10520
rect 12483 10489 12495 10492
rect 12437 10483 12495 10489
rect 16022 10480 16028 10492
rect 16080 10480 16086 10532
rect 16117 10523 16175 10529
rect 16117 10489 16129 10523
rect 16163 10520 16175 10523
rect 18417 10523 18475 10529
rect 16163 10492 17724 10520
rect 16163 10489 16175 10492
rect 16117 10483 16175 10489
rect 17696 10464 17724 10492
rect 18417 10489 18429 10523
rect 18463 10520 18475 10523
rect 19061 10523 19119 10529
rect 19061 10520 19073 10523
rect 18463 10492 19073 10520
rect 18463 10489 18475 10492
rect 18417 10483 18475 10489
rect 19061 10489 19073 10492
rect 19107 10489 19119 10523
rect 19061 10483 19119 10489
rect 19972 10523 20030 10529
rect 19972 10489 19984 10523
rect 20018 10520 20030 10523
rect 20438 10520 20444 10532
rect 20018 10492 20444 10520
rect 20018 10489 20030 10492
rect 19972 10483 20030 10489
rect 20438 10480 20444 10492
rect 20496 10480 20502 10532
rect 9582 10452 9588 10464
rect 9543 10424 9588 10452
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 9858 10452 9864 10464
rect 9819 10424 9864 10452
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 10873 10455 10931 10461
rect 10873 10421 10885 10455
rect 10919 10452 10931 10455
rect 11146 10452 11152 10464
rect 10919 10424 11152 10452
rect 10919 10421 10931 10424
rect 10873 10415 10931 10421
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 11333 10455 11391 10461
rect 11333 10421 11345 10455
rect 11379 10452 11391 10455
rect 11698 10452 11704 10464
rect 11379 10424 11704 10452
rect 11379 10421 11391 10424
rect 11333 10415 11391 10421
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 12526 10412 12532 10464
rect 12584 10452 12590 10464
rect 12894 10452 12900 10464
rect 12584 10424 12900 10452
rect 12584 10412 12590 10424
rect 12894 10412 12900 10424
rect 12952 10412 12958 10464
rect 12989 10455 13047 10461
rect 12989 10421 13001 10455
rect 13035 10452 13047 10455
rect 13078 10452 13084 10464
rect 13035 10424 13084 10452
rect 13035 10421 13047 10424
rect 12989 10415 13047 10421
rect 13078 10412 13084 10424
rect 13136 10452 13142 10464
rect 13538 10452 13544 10464
rect 13136 10424 13544 10452
rect 13136 10412 13142 10424
rect 13538 10412 13544 10424
rect 13596 10412 13602 10464
rect 13630 10412 13636 10464
rect 13688 10452 13694 10464
rect 13817 10455 13875 10461
rect 13817 10452 13829 10455
rect 13688 10424 13829 10452
rect 13688 10412 13694 10424
rect 13817 10421 13829 10424
rect 13863 10421 13875 10455
rect 13817 10415 13875 10421
rect 14921 10455 14979 10461
rect 14921 10421 14933 10455
rect 14967 10452 14979 10455
rect 15654 10452 15660 10464
rect 14967 10424 15660 10452
rect 14967 10421 14979 10424
rect 14921 10415 14979 10421
rect 15654 10412 15660 10424
rect 15712 10412 15718 10464
rect 15749 10455 15807 10461
rect 15749 10421 15761 10455
rect 15795 10452 15807 10455
rect 17586 10452 17592 10464
rect 15795 10424 17592 10452
rect 15795 10421 15807 10424
rect 15749 10415 15807 10421
rect 17586 10412 17592 10424
rect 17644 10412 17650 10464
rect 17678 10412 17684 10464
rect 17736 10452 17742 10464
rect 17736 10424 17829 10452
rect 17736 10412 17742 10424
rect 18322 10412 18328 10464
rect 18380 10452 18386 10464
rect 18509 10455 18567 10461
rect 18509 10452 18521 10455
rect 18380 10424 18521 10452
rect 18380 10412 18386 10424
rect 18509 10421 18521 10424
rect 18555 10421 18567 10455
rect 18509 10415 18567 10421
rect 19426 10412 19432 10464
rect 19484 10452 19490 10464
rect 21085 10455 21143 10461
rect 21085 10452 21097 10455
rect 19484 10424 21097 10452
rect 19484 10412 19490 10424
rect 21085 10421 21097 10424
rect 21131 10421 21143 10455
rect 21085 10415 21143 10421
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 9033 10251 9091 10257
rect 9033 10217 9045 10251
rect 9079 10248 9091 10251
rect 9858 10248 9864 10260
rect 9079 10220 9864 10248
rect 9079 10217 9091 10220
rect 9033 10211 9091 10217
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 11974 10248 11980 10260
rect 11935 10220 11980 10248
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 12986 10208 12992 10260
rect 13044 10248 13050 10260
rect 13173 10251 13231 10257
rect 13173 10248 13185 10251
rect 13044 10220 13185 10248
rect 13044 10208 13050 10220
rect 13173 10217 13185 10220
rect 13219 10217 13231 10251
rect 13173 10211 13231 10217
rect 14553 10251 14611 10257
rect 14553 10217 14565 10251
rect 14599 10248 14611 10251
rect 15289 10251 15347 10257
rect 15289 10248 15301 10251
rect 14599 10220 15301 10248
rect 14599 10217 14611 10220
rect 14553 10211 14611 10217
rect 15289 10217 15301 10220
rect 15335 10217 15347 10251
rect 15289 10211 15347 10217
rect 15378 10208 15384 10260
rect 15436 10248 15442 10260
rect 16758 10248 16764 10260
rect 15436 10220 16764 10248
rect 15436 10208 15442 10220
rect 16758 10208 16764 10220
rect 16816 10208 16822 10260
rect 16853 10251 16911 10257
rect 16853 10217 16865 10251
rect 16899 10248 16911 10251
rect 18233 10251 18291 10257
rect 18233 10248 18245 10251
rect 16899 10220 18245 10248
rect 16899 10217 16911 10220
rect 16853 10211 16911 10217
rect 18233 10217 18245 10220
rect 18279 10217 18291 10251
rect 18233 10211 18291 10217
rect 10864 10183 10922 10189
rect 10864 10149 10876 10183
rect 10910 10180 10922 10183
rect 11054 10180 11060 10192
rect 10910 10152 11060 10180
rect 10910 10149 10922 10152
rect 10864 10143 10922 10149
rect 11054 10140 11060 10152
rect 11112 10180 11118 10192
rect 11422 10180 11428 10192
rect 11112 10152 11428 10180
rect 11112 10140 11118 10152
rect 11422 10140 11428 10152
rect 11480 10140 11486 10192
rect 13633 10183 13691 10189
rect 13633 10180 13645 10183
rect 12443 10152 13645 10180
rect 8941 10115 8999 10121
rect 8941 10081 8953 10115
rect 8987 10112 8999 10115
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 8987 10084 9689 10112
rect 8987 10081 8999 10084
rect 8941 10075 8999 10081
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 10686 10072 10692 10124
rect 10744 10112 10750 10124
rect 12443 10112 12471 10152
rect 13633 10149 13645 10152
rect 13679 10180 13691 10183
rect 15746 10180 15752 10192
rect 13679 10152 15752 10180
rect 13679 10149 13691 10152
rect 13633 10143 13691 10149
rect 15746 10140 15752 10152
rect 15804 10140 15810 10192
rect 16022 10140 16028 10192
rect 16080 10180 16086 10192
rect 19613 10183 19671 10189
rect 19613 10180 19625 10183
rect 16080 10152 19625 10180
rect 16080 10140 16086 10152
rect 19613 10149 19625 10152
rect 19659 10149 19671 10183
rect 19613 10143 19671 10149
rect 10744 10084 12471 10112
rect 10744 10072 10750 10084
rect 12526 10072 12532 10124
rect 12584 10112 12590 10124
rect 13078 10112 13084 10124
rect 12584 10084 13084 10112
rect 12584 10072 12590 10084
rect 13078 10072 13084 10084
rect 13136 10072 13142 10124
rect 13538 10112 13544 10124
rect 13499 10084 13544 10112
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 14645 10115 14703 10121
rect 14645 10081 14657 10115
rect 14691 10112 14703 10115
rect 15286 10112 15292 10124
rect 14691 10084 15292 10112
rect 14691 10081 14703 10084
rect 14645 10075 14703 10081
rect 15286 10072 15292 10084
rect 15344 10072 15350 10124
rect 15378 10072 15384 10124
rect 15436 10112 15442 10124
rect 15654 10112 15660 10124
rect 15436 10084 15660 10112
rect 15436 10072 15442 10084
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 16850 10072 16856 10124
rect 16908 10112 16914 10124
rect 17221 10115 17279 10121
rect 17221 10112 17233 10115
rect 16908 10084 17233 10112
rect 16908 10072 16914 10084
rect 17221 10081 17233 10084
rect 17267 10081 17279 10115
rect 17862 10112 17868 10124
rect 17221 10075 17279 10081
rect 17328 10084 17868 10112
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10044 9275 10047
rect 9582 10044 9588 10056
rect 9263 10016 9588 10044
rect 9263 10013 9275 10016
rect 9217 10007 9275 10013
rect 9582 10004 9588 10016
rect 9640 10004 9646 10056
rect 10594 10044 10600 10056
rect 10555 10016 10600 10044
rect 10594 10004 10600 10016
rect 10652 10004 10658 10056
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10013 13783 10047
rect 13725 10007 13783 10013
rect 8573 9979 8631 9985
rect 8573 9945 8585 9979
rect 8619 9976 8631 9979
rect 9674 9976 9680 9988
rect 8619 9948 9680 9976
rect 8619 9945 8631 9948
rect 8573 9939 8631 9945
rect 9674 9936 9680 9948
rect 9732 9936 9738 9988
rect 13354 9936 13360 9988
rect 13412 9976 13418 9988
rect 13740 9976 13768 10007
rect 14458 10004 14464 10056
rect 14516 10044 14522 10056
rect 14737 10047 14795 10053
rect 14737 10044 14749 10047
rect 14516 10016 14749 10044
rect 14516 10004 14522 10016
rect 14737 10013 14749 10016
rect 14783 10013 14795 10047
rect 14737 10007 14795 10013
rect 15749 10047 15807 10053
rect 15749 10013 15761 10047
rect 15795 10013 15807 10047
rect 15930 10044 15936 10056
rect 15891 10016 15936 10044
rect 15749 10007 15807 10013
rect 13412 9948 13768 9976
rect 15764 9976 15792 10007
rect 15930 10004 15936 10016
rect 15988 10004 15994 10056
rect 17328 10053 17356 10084
rect 17862 10072 17868 10084
rect 17920 10072 17926 10124
rect 17313 10047 17371 10053
rect 17313 10013 17325 10047
rect 17359 10013 17371 10047
rect 17494 10044 17500 10056
rect 17455 10016 17500 10044
rect 17313 10007 17371 10013
rect 16022 9976 16028 9988
rect 15764 9948 16028 9976
rect 13412 9936 13418 9948
rect 16022 9936 16028 9948
rect 16080 9936 16086 9988
rect 16850 9936 16856 9988
rect 16908 9976 16914 9988
rect 17328 9976 17356 10007
rect 17494 10004 17500 10016
rect 17552 10004 17558 10056
rect 17954 10004 17960 10056
rect 18012 10044 18018 10056
rect 18325 10047 18383 10053
rect 18325 10044 18337 10047
rect 18012 10016 18337 10044
rect 18012 10004 18018 10016
rect 18325 10013 18337 10016
rect 18371 10013 18383 10047
rect 18506 10044 18512 10056
rect 18467 10016 18512 10044
rect 18325 10007 18383 10013
rect 18506 10004 18512 10016
rect 18564 10004 18570 10056
rect 19702 10044 19708 10056
rect 19663 10016 19708 10044
rect 19702 10004 19708 10016
rect 19760 10004 19766 10056
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10044 19947 10047
rect 20162 10044 20168 10056
rect 19935 10016 20168 10044
rect 19935 10013 19947 10016
rect 19889 10007 19947 10013
rect 20162 10004 20168 10016
rect 20220 10004 20226 10056
rect 16908 9948 17356 9976
rect 16908 9936 16914 9948
rect 17586 9936 17592 9988
rect 17644 9976 17650 9988
rect 17865 9979 17923 9985
rect 17865 9976 17877 9979
rect 17644 9948 17877 9976
rect 17644 9936 17650 9948
rect 17865 9945 17877 9948
rect 17911 9945 17923 9979
rect 17865 9939 17923 9945
rect 18046 9936 18052 9988
rect 18104 9936 18110 9988
rect 14182 9908 14188 9920
rect 14143 9880 14188 9908
rect 14182 9868 14188 9880
rect 14240 9868 14246 9920
rect 16574 9868 16580 9920
rect 16632 9908 16638 9920
rect 18064 9908 18092 9936
rect 16632 9880 18092 9908
rect 16632 9868 16638 9880
rect 18506 9868 18512 9920
rect 18564 9908 18570 9920
rect 19245 9911 19303 9917
rect 19245 9908 19257 9911
rect 18564 9880 19257 9908
rect 18564 9868 18570 9880
rect 19245 9877 19257 9880
rect 19291 9877 19303 9911
rect 19245 9871 19303 9877
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 9030 9664 9036 9716
rect 9088 9704 9094 9716
rect 9306 9704 9312 9716
rect 9088 9676 9312 9704
rect 9088 9664 9094 9676
rect 9306 9664 9312 9676
rect 9364 9664 9370 9716
rect 10594 9704 10600 9716
rect 9968 9676 10600 9704
rect 9766 9528 9772 9580
rect 9824 9568 9830 9580
rect 9968 9577 9996 9676
rect 10594 9664 10600 9676
rect 10652 9704 10658 9716
rect 10652 9676 10916 9704
rect 10652 9664 10658 9676
rect 10888 9636 10916 9676
rect 11054 9664 11060 9716
rect 11112 9704 11118 9716
rect 11333 9707 11391 9713
rect 11333 9704 11345 9707
rect 11112 9676 11345 9704
rect 11112 9664 11118 9676
rect 11333 9673 11345 9676
rect 11379 9673 11391 9707
rect 11333 9667 11391 9673
rect 15378 9664 15384 9716
rect 15436 9704 15442 9716
rect 15436 9676 16160 9704
rect 15436 9664 15442 9676
rect 16025 9639 16083 9645
rect 16025 9636 16037 9639
rect 10888 9608 12572 9636
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 9824 9540 9965 9568
rect 9824 9528 9830 9540
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 11882 9568 11888 9580
rect 11843 9540 11888 9568
rect 9953 9531 10011 9537
rect 11882 9528 11888 9540
rect 11940 9528 11946 9580
rect 12544 9577 12572 9608
rect 15672 9608 16037 9636
rect 12529 9571 12587 9577
rect 12529 9537 12541 9571
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 13722 9528 13728 9580
rect 13780 9568 13786 9580
rect 14645 9571 14703 9577
rect 14645 9568 14657 9571
rect 13780 9540 14657 9568
rect 13780 9528 13786 9540
rect 14645 9537 14657 9540
rect 14691 9537 14703 9571
rect 14645 9531 14703 9537
rect 7742 9500 7748 9512
rect 7703 9472 7748 9500
rect 7742 9460 7748 9472
rect 7800 9460 7806 9512
rect 8012 9503 8070 9509
rect 8012 9469 8024 9503
rect 8058 9500 8070 9503
rect 8570 9500 8576 9512
rect 8058 9472 8576 9500
rect 8058 9469 8070 9472
rect 8012 9463 8070 9469
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 9861 9503 9919 9509
rect 9861 9469 9873 9503
rect 9907 9469 9919 9503
rect 9861 9463 9919 9469
rect 9582 9432 9588 9444
rect 8956 9404 9588 9432
rect 8570 9324 8576 9376
rect 8628 9364 8634 9376
rect 8956 9364 8984 9404
rect 9582 9392 9588 9404
rect 9640 9392 9646 9444
rect 9122 9364 9128 9376
rect 8628 9336 8984 9364
rect 9083 9336 9128 9364
rect 8628 9324 8634 9336
rect 9122 9324 9128 9336
rect 9180 9324 9186 9376
rect 9677 9367 9735 9373
rect 9677 9333 9689 9367
rect 9723 9364 9735 9367
rect 9766 9364 9772 9376
rect 9723 9336 9772 9364
rect 9723 9333 9735 9336
rect 9677 9327 9735 9333
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 9876 9364 9904 9463
rect 11146 9460 11152 9512
rect 11204 9500 11210 9512
rect 11609 9503 11667 9509
rect 11609 9500 11621 9503
rect 11204 9472 11621 9500
rect 11204 9460 11210 9472
rect 11609 9469 11621 9472
rect 11655 9469 11667 9503
rect 11609 9463 11667 9469
rect 12796 9503 12854 9509
rect 12796 9469 12808 9503
rect 12842 9500 12854 9503
rect 14458 9500 14464 9512
rect 12842 9472 14464 9500
rect 12842 9469 12854 9472
rect 12796 9463 12854 9469
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 15672 9500 15700 9608
rect 16025 9605 16037 9608
rect 16071 9605 16083 9639
rect 16132 9636 16160 9676
rect 17954 9664 17960 9716
rect 18012 9704 18018 9716
rect 18049 9707 18107 9713
rect 18049 9704 18061 9707
rect 18012 9676 18061 9704
rect 18012 9664 18018 9676
rect 18049 9673 18061 9676
rect 18095 9673 18107 9707
rect 18049 9667 18107 9673
rect 18138 9636 18144 9648
rect 16132 9608 18144 9636
rect 16025 9599 16083 9605
rect 16040 9568 16068 9599
rect 18138 9596 18144 9608
rect 18196 9596 18202 9648
rect 18230 9596 18236 9648
rect 18288 9636 18294 9648
rect 18782 9636 18788 9648
rect 18288 9608 18788 9636
rect 18288 9596 18294 9608
rect 18782 9596 18788 9608
rect 18840 9596 18846 9648
rect 20162 9596 20168 9648
rect 20220 9596 20226 9648
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16040 9540 16865 9568
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 17494 9528 17500 9580
rect 17552 9568 17558 9580
rect 18601 9571 18659 9577
rect 18601 9568 18613 9571
rect 17552 9540 18613 9568
rect 17552 9528 17558 9540
rect 18601 9537 18613 9540
rect 18647 9537 18659 9571
rect 18601 9531 18659 9537
rect 18874 9528 18880 9580
rect 18932 9528 18938 9580
rect 14844 9472 15700 9500
rect 10220 9435 10278 9441
rect 10220 9401 10232 9435
rect 10266 9432 10278 9435
rect 10410 9432 10416 9444
rect 10266 9404 10416 9432
rect 10266 9401 10278 9404
rect 10220 9395 10278 9401
rect 10410 9392 10416 9404
rect 10468 9392 10474 9444
rect 10594 9392 10600 9444
rect 10652 9432 10658 9444
rect 14274 9432 14280 9444
rect 10652 9404 14280 9432
rect 10652 9392 10658 9404
rect 14274 9392 14280 9404
rect 14332 9392 14338 9444
rect 14476 9432 14504 9460
rect 14844 9432 14872 9472
rect 18322 9460 18328 9512
rect 18380 9500 18386 9512
rect 18892 9500 18920 9528
rect 19153 9503 19211 9509
rect 19153 9500 19165 9503
rect 18380 9472 18736 9500
rect 18380 9460 18386 9472
rect 14476 9404 14872 9432
rect 14912 9435 14970 9441
rect 14912 9401 14924 9435
rect 14958 9432 14970 9435
rect 15378 9432 15384 9444
rect 14958 9404 15384 9432
rect 14958 9401 14970 9404
rect 14912 9395 14970 9401
rect 15378 9392 15384 9404
rect 15436 9392 15442 9444
rect 16669 9435 16727 9441
rect 16669 9432 16681 9435
rect 15488 9404 16681 9432
rect 10870 9364 10876 9376
rect 9876 9336 10876 9364
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 13909 9367 13967 9373
rect 13909 9333 13921 9367
rect 13955 9364 13967 9367
rect 14090 9364 14096 9376
rect 13955 9336 14096 9364
rect 13955 9333 13967 9336
rect 13909 9327 13967 9333
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 14185 9367 14243 9373
rect 14185 9333 14197 9367
rect 14231 9364 14243 9367
rect 15488 9364 15516 9404
rect 16669 9401 16681 9404
rect 16715 9401 16727 9435
rect 16669 9395 16727 9401
rect 16758 9392 16764 9444
rect 16816 9432 16822 9444
rect 17402 9432 17408 9444
rect 16816 9404 17408 9432
rect 16816 9392 16822 9404
rect 17402 9392 17408 9404
rect 17460 9392 17466 9444
rect 17954 9392 17960 9444
rect 18012 9432 18018 9444
rect 18414 9432 18420 9444
rect 18012 9404 18420 9432
rect 18012 9392 18018 9404
rect 18414 9392 18420 9404
rect 18472 9392 18478 9444
rect 18708 9432 18736 9472
rect 18892 9472 19165 9500
rect 18892 9432 18920 9472
rect 19153 9469 19165 9472
rect 19199 9469 19211 9503
rect 19153 9463 19211 9469
rect 18708 9404 18920 9432
rect 19420 9435 19478 9441
rect 19420 9401 19432 9435
rect 19466 9432 19478 9435
rect 19518 9432 19524 9444
rect 19466 9404 19524 9432
rect 19466 9401 19478 9404
rect 19420 9395 19478 9401
rect 19518 9392 19524 9404
rect 19576 9432 19582 9444
rect 20180 9432 20208 9596
rect 20806 9568 20812 9580
rect 20767 9540 20812 9568
rect 20806 9528 20812 9540
rect 20864 9528 20870 9580
rect 19576 9404 20208 9432
rect 19576 9392 19582 9404
rect 16298 9364 16304 9376
rect 14231 9336 15516 9364
rect 16259 9336 16304 9364
rect 14231 9333 14243 9336
rect 14185 9327 14243 9333
rect 16298 9324 16304 9336
rect 16356 9324 16362 9376
rect 17586 9324 17592 9376
rect 17644 9364 17650 9376
rect 18509 9367 18567 9373
rect 18509 9364 18521 9367
rect 17644 9336 18521 9364
rect 17644 9324 17650 9336
rect 18509 9333 18521 9336
rect 18555 9333 18567 9367
rect 18509 9327 18567 9333
rect 19242 9324 19248 9376
rect 19300 9364 19306 9376
rect 19610 9364 19616 9376
rect 19300 9336 19616 9364
rect 19300 9324 19306 9336
rect 19610 9324 19616 9336
rect 19668 9324 19674 9376
rect 20438 9324 20444 9376
rect 20496 9364 20502 9376
rect 20533 9367 20591 9373
rect 20533 9364 20545 9367
rect 20496 9336 20545 9364
rect 20496 9324 20502 9336
rect 20533 9333 20545 9336
rect 20579 9333 20591 9367
rect 20533 9327 20591 9333
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 9861 9163 9919 9169
rect 9861 9129 9873 9163
rect 9907 9160 9919 9163
rect 11054 9160 11060 9172
rect 9907 9132 11060 9160
rect 9907 9129 9919 9132
rect 9861 9123 9919 9129
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 11333 9163 11391 9169
rect 11333 9129 11345 9163
rect 11379 9160 11391 9163
rect 11885 9163 11943 9169
rect 11885 9160 11897 9163
rect 11379 9132 11897 9160
rect 11379 9129 11391 9132
rect 11333 9123 11391 9129
rect 11885 9129 11897 9132
rect 11931 9129 11943 9163
rect 11885 9123 11943 9129
rect 12253 9163 12311 9169
rect 12253 9129 12265 9163
rect 12299 9160 12311 9163
rect 14001 9163 14059 9169
rect 12299 9132 13860 9160
rect 12299 9129 12311 9132
rect 12253 9123 12311 9129
rect 9033 9095 9091 9101
rect 9033 9061 9045 9095
rect 9079 9092 9091 9095
rect 10042 9092 10048 9104
rect 9079 9064 10048 9092
rect 9079 9061 9091 9064
rect 9033 9055 9091 9061
rect 10042 9052 10048 9064
rect 10100 9052 10106 9104
rect 10229 9095 10287 9101
rect 10229 9061 10241 9095
rect 10275 9092 10287 9095
rect 12897 9095 12955 9101
rect 12897 9092 12909 9095
rect 10275 9064 12909 9092
rect 10275 9061 10287 9064
rect 10229 9055 10287 9061
rect 12897 9061 12909 9064
rect 12943 9061 12955 9095
rect 12897 9055 12955 9061
rect 6914 8984 6920 9036
rect 6972 9024 6978 9036
rect 8941 9027 8999 9033
rect 8941 9024 8953 9027
rect 6972 8996 8953 9024
rect 6972 8984 6978 8996
rect 8941 8993 8953 8996
rect 8987 8993 8999 9027
rect 10594 9024 10600 9036
rect 8941 8987 8999 8993
rect 10336 8996 10600 9024
rect 9122 8916 9128 8968
rect 9180 8956 9186 8968
rect 9180 8928 9225 8956
rect 9180 8916 9186 8928
rect 9766 8916 9772 8968
rect 9824 8956 9830 8968
rect 10336 8965 10364 8996
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 11054 8984 11060 9036
rect 11112 9024 11118 9036
rect 11241 9027 11299 9033
rect 11241 9024 11253 9027
rect 11112 8996 11253 9024
rect 11112 8984 11118 8996
rect 11241 8993 11253 8996
rect 11287 8993 11299 9027
rect 11241 8987 11299 8993
rect 12345 9027 12403 9033
rect 12345 8993 12357 9027
rect 12391 9024 12403 9027
rect 13446 9024 13452 9036
rect 12391 8996 13452 9024
rect 12391 8993 12403 8996
rect 12345 8987 12403 8993
rect 13446 8984 13452 8996
rect 13504 8984 13510 9036
rect 13832 9024 13860 9132
rect 14001 9129 14013 9163
rect 14047 9160 14059 9163
rect 14182 9160 14188 9172
rect 14047 9132 14188 9160
rect 14047 9129 14059 9132
rect 14001 9123 14059 9129
rect 14182 9120 14188 9132
rect 14240 9120 14246 9172
rect 14274 9120 14280 9172
rect 14332 9160 14338 9172
rect 15102 9160 15108 9172
rect 14332 9132 15108 9160
rect 14332 9120 14338 9132
rect 15102 9120 15108 9132
rect 15160 9120 15166 9172
rect 15286 9160 15292 9172
rect 15247 9132 15292 9160
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 15378 9120 15384 9172
rect 15436 9160 15442 9172
rect 15930 9160 15936 9172
rect 15436 9132 15936 9160
rect 15436 9120 15442 9132
rect 15930 9120 15936 9132
rect 15988 9120 15994 9172
rect 18877 9163 18935 9169
rect 18877 9129 18889 9163
rect 18923 9129 18935 9163
rect 18877 9123 18935 9129
rect 13909 9095 13967 9101
rect 13909 9061 13921 9095
rect 13955 9092 13967 9095
rect 16298 9092 16304 9104
rect 13955 9064 16304 9092
rect 13955 9061 13967 9064
rect 13909 9055 13967 9061
rect 16298 9052 16304 9064
rect 16356 9052 16362 9104
rect 17678 9052 17684 9104
rect 17736 9101 17742 9104
rect 17736 9095 17800 9101
rect 17736 9061 17754 9095
rect 17788 9061 17800 9095
rect 17736 9055 17800 9061
rect 17736 9052 17742 9055
rect 18230 9052 18236 9104
rect 18288 9092 18294 9104
rect 18690 9092 18696 9104
rect 18288 9064 18696 9092
rect 18288 9052 18294 9064
rect 18690 9052 18696 9064
rect 18748 9052 18754 9104
rect 18892 9092 18920 9123
rect 19518 9120 19524 9172
rect 19576 9160 19582 9172
rect 20533 9163 20591 9169
rect 20533 9160 20545 9163
rect 19576 9132 20545 9160
rect 19576 9120 19582 9132
rect 20533 9129 20545 9132
rect 20579 9129 20591 9163
rect 20533 9123 20591 9129
rect 19398 9095 19456 9101
rect 19398 9092 19410 9095
rect 18892 9064 19410 9092
rect 19398 9061 19410 9064
rect 19444 9092 19456 9095
rect 19610 9092 19616 9104
rect 19444 9064 19616 9092
rect 19444 9061 19456 9064
rect 19398 9055 19456 9061
rect 19610 9052 19616 9064
rect 19668 9052 19674 9104
rect 14734 9024 14740 9036
rect 13832 8996 14228 9024
rect 14695 8996 14740 9024
rect 10321 8959 10379 8965
rect 10321 8956 10333 8959
rect 9824 8928 10333 8956
rect 9824 8916 9830 8928
rect 10321 8925 10333 8928
rect 10367 8925 10379 8959
rect 10321 8919 10379 8925
rect 10410 8916 10416 8968
rect 10468 8956 10474 8968
rect 11146 8956 11152 8968
rect 10468 8928 11152 8956
rect 10468 8916 10474 8928
rect 11146 8916 11152 8928
rect 11204 8956 11210 8968
rect 11425 8959 11483 8965
rect 11425 8956 11437 8959
rect 11204 8928 11437 8956
rect 11204 8916 11210 8928
rect 11425 8925 11437 8928
rect 11471 8925 11483 8959
rect 12437 8959 12495 8965
rect 12437 8956 12449 8959
rect 11425 8919 11483 8925
rect 11808 8928 12449 8956
rect 10873 8891 10931 8897
rect 10873 8857 10885 8891
rect 10919 8888 10931 8891
rect 11698 8888 11704 8900
rect 10919 8860 11704 8888
rect 10919 8857 10931 8860
rect 10873 8851 10931 8857
rect 11698 8848 11704 8860
rect 11756 8848 11762 8900
rect 8570 8820 8576 8832
rect 8531 8792 8576 8820
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 10778 8780 10784 8832
rect 10836 8820 10842 8832
rect 11808 8820 11836 8928
rect 12437 8925 12449 8928
rect 12483 8925 12495 8959
rect 12437 8919 12495 8925
rect 12710 8916 12716 8968
rect 12768 8956 12774 8968
rect 13354 8956 13360 8968
rect 12768 8928 13360 8956
rect 12768 8916 12774 8928
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 14090 8956 14096 8968
rect 14051 8928 14096 8956
rect 14090 8916 14096 8928
rect 14148 8916 14154 8968
rect 14200 8956 14228 8996
rect 14734 8984 14740 8996
rect 14792 8984 14798 9036
rect 15654 9024 15660 9036
rect 15615 8996 15660 9024
rect 15654 8984 15660 8996
rect 15712 8984 15718 9036
rect 15838 8984 15844 9036
rect 15896 9024 15902 9036
rect 16390 9024 16396 9036
rect 15896 8996 16396 9024
rect 15896 8984 15902 8996
rect 16390 8984 16396 8996
rect 16448 9024 16454 9036
rect 16761 9027 16819 9033
rect 16761 9024 16773 9027
rect 16448 8996 16773 9024
rect 16448 8984 16454 8996
rect 16761 8993 16773 8996
rect 16807 8993 16819 9027
rect 18322 9024 18328 9036
rect 16761 8987 16819 8993
rect 17512 8996 18328 9024
rect 15102 8956 15108 8968
rect 14200 8928 15108 8956
rect 15102 8916 15108 8928
rect 15160 8916 15166 8968
rect 15470 8916 15476 8968
rect 15528 8956 15534 8968
rect 15749 8959 15807 8965
rect 15749 8956 15761 8959
rect 15528 8928 15761 8956
rect 15528 8916 15534 8928
rect 15749 8925 15761 8928
rect 15795 8925 15807 8959
rect 15930 8956 15936 8968
rect 15891 8928 15936 8956
rect 15749 8919 15807 8925
rect 12802 8848 12808 8900
rect 12860 8888 12866 8900
rect 14550 8888 14556 8900
rect 12860 8860 14556 8888
rect 12860 8848 12866 8860
rect 14550 8848 14556 8860
rect 14608 8848 14614 8900
rect 15764 8888 15792 8919
rect 15930 8916 15936 8928
rect 15988 8916 15994 8968
rect 16298 8916 16304 8968
rect 16356 8956 16362 8968
rect 16482 8956 16488 8968
rect 16356 8928 16488 8956
rect 16356 8916 16362 8928
rect 16482 8916 16488 8928
rect 16540 8916 16546 8968
rect 17512 8965 17540 8996
rect 18322 8984 18328 8996
rect 18380 9024 18386 9036
rect 19153 9027 19211 9033
rect 19153 9024 19165 9027
rect 18380 8996 19165 9024
rect 18380 8984 18386 8996
rect 19153 8993 19165 8996
rect 19199 8993 19211 9027
rect 19153 8987 19211 8993
rect 17497 8959 17555 8965
rect 17497 8956 17509 8959
rect 17328 8928 17509 8956
rect 17218 8888 17224 8900
rect 15764 8860 17224 8888
rect 17218 8848 17224 8860
rect 17276 8848 17282 8900
rect 10836 8792 11836 8820
rect 10836 8780 10842 8792
rect 12710 8780 12716 8832
rect 12768 8820 12774 8832
rect 13541 8823 13599 8829
rect 13541 8820 13553 8823
rect 12768 8792 13553 8820
rect 12768 8780 12774 8792
rect 13541 8789 13553 8792
rect 13587 8789 13599 8823
rect 13541 8783 13599 8789
rect 15654 8780 15660 8832
rect 15712 8820 15718 8832
rect 16206 8820 16212 8832
rect 15712 8792 16212 8820
rect 15712 8780 15718 8792
rect 16206 8780 16212 8792
rect 16264 8820 16270 8832
rect 16577 8823 16635 8829
rect 16577 8820 16589 8823
rect 16264 8792 16589 8820
rect 16264 8780 16270 8792
rect 16577 8789 16589 8792
rect 16623 8820 16635 8823
rect 17328 8820 17356 8928
rect 17497 8925 17509 8928
rect 17543 8925 17555 8959
rect 17497 8919 17555 8925
rect 16623 8792 17356 8820
rect 16623 8789 16635 8792
rect 16577 8783 16635 8789
rect 18966 8780 18972 8832
rect 19024 8820 19030 8832
rect 19334 8820 19340 8832
rect 19024 8792 19340 8820
rect 19024 8780 19030 8792
rect 19334 8780 19340 8792
rect 19392 8780 19398 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 11146 8576 11152 8628
rect 11204 8616 11210 8628
rect 11241 8619 11299 8625
rect 11241 8616 11253 8619
rect 11204 8588 11253 8616
rect 11204 8576 11210 8588
rect 11241 8585 11253 8588
rect 11287 8585 11299 8619
rect 13722 8616 13728 8628
rect 11241 8579 11299 8585
rect 13096 8588 13728 8616
rect 10870 8508 10876 8560
rect 10928 8548 10934 8560
rect 12621 8551 12679 8557
rect 12621 8548 12633 8551
rect 10928 8520 12633 8548
rect 10928 8508 10934 8520
rect 12621 8517 12633 8520
rect 12667 8517 12679 8551
rect 12621 8511 12679 8517
rect 11606 8440 11612 8492
rect 11664 8480 11670 8492
rect 13096 8489 13124 8588
rect 13722 8576 13728 8588
rect 13780 8616 13786 8628
rect 15105 8619 15163 8625
rect 13780 8588 15056 8616
rect 13780 8576 13786 8588
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 11664 8452 11713 8480
rect 11664 8440 11670 8452
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8449 13139 8483
rect 15028 8480 15056 8588
rect 15105 8585 15117 8619
rect 15151 8616 15163 8619
rect 15838 8616 15844 8628
rect 15151 8588 15844 8616
rect 15151 8585 15163 8588
rect 15105 8579 15163 8585
rect 15838 8576 15844 8588
rect 15896 8576 15902 8628
rect 15930 8576 15936 8628
rect 15988 8616 15994 8628
rect 17313 8619 17371 8625
rect 17313 8616 17325 8619
rect 15988 8588 17325 8616
rect 15988 8576 15994 8588
rect 17313 8585 17325 8588
rect 17359 8585 17371 8619
rect 17313 8579 17371 8585
rect 18049 8619 18107 8625
rect 18049 8585 18061 8619
rect 18095 8616 18107 8619
rect 18598 8616 18604 8628
rect 18095 8588 18604 8616
rect 18095 8585 18107 8588
rect 18049 8579 18107 8585
rect 18598 8576 18604 8588
rect 18656 8576 18662 8628
rect 19061 8619 19119 8625
rect 19061 8585 19073 8619
rect 19107 8616 19119 8619
rect 19702 8616 19708 8628
rect 19107 8588 19708 8616
rect 19107 8585 19119 8588
rect 19061 8579 19119 8585
rect 19702 8576 19708 8588
rect 19760 8576 19766 8628
rect 20438 8548 20444 8560
rect 18708 8520 20444 8548
rect 15654 8480 15660 8492
rect 15028 8452 15660 8480
rect 13081 8443 13139 8449
rect 15654 8440 15660 8452
rect 15712 8480 15718 8492
rect 15933 8483 15991 8489
rect 15933 8480 15945 8483
rect 15712 8452 15945 8480
rect 15712 8440 15718 8452
rect 15933 8449 15945 8452
rect 15979 8449 15991 8483
rect 18506 8480 18512 8492
rect 18467 8452 18512 8480
rect 15933 8443 15991 8449
rect 18506 8440 18512 8452
rect 18564 8440 18570 8492
rect 18708 8489 18736 8520
rect 20438 8508 20444 8520
rect 20496 8508 20502 8560
rect 18693 8483 18751 8489
rect 18693 8449 18705 8483
rect 18739 8449 18751 8483
rect 18693 8443 18751 8449
rect 18969 8483 19027 8489
rect 18969 8449 18981 8483
rect 19015 8480 19027 8483
rect 19058 8480 19064 8492
rect 19015 8452 19064 8480
rect 19015 8449 19027 8452
rect 18969 8443 19027 8449
rect 19058 8440 19064 8452
rect 19116 8440 19122 8492
rect 19610 8480 19616 8492
rect 19571 8452 19616 8480
rect 19610 8440 19616 8452
rect 19668 8440 19674 8492
rect 20530 8480 20536 8492
rect 20491 8452 20536 8480
rect 20530 8440 20536 8452
rect 20588 8440 20594 8492
rect 20622 8440 20628 8492
rect 20680 8480 20686 8492
rect 20680 8452 20725 8480
rect 20680 8440 20686 8452
rect 7742 8372 7748 8424
rect 7800 8412 7806 8424
rect 8021 8415 8079 8421
rect 8021 8412 8033 8415
rect 7800 8384 8033 8412
rect 7800 8372 7806 8384
rect 8021 8381 8033 8384
rect 8067 8381 8079 8415
rect 8021 8375 8079 8381
rect 8288 8415 8346 8421
rect 8288 8381 8300 8415
rect 8334 8412 8346 8415
rect 9122 8412 9128 8424
rect 8334 8384 9128 8412
rect 8334 8381 8346 8384
rect 8288 8375 8346 8381
rect 8036 8344 8064 8375
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 9858 8372 9864 8424
rect 9916 8412 9922 8424
rect 9916 8384 9961 8412
rect 9916 8372 9922 8384
rect 11146 8372 11152 8424
rect 11204 8412 11210 8424
rect 11517 8415 11575 8421
rect 11517 8412 11529 8415
rect 11204 8384 11529 8412
rect 11204 8372 11210 8384
rect 11517 8381 11529 8384
rect 11563 8381 11575 8415
rect 12802 8412 12808 8424
rect 12763 8384 12808 8412
rect 11517 8375 11575 8381
rect 12802 8372 12808 8384
rect 12860 8372 12866 8424
rect 13348 8415 13406 8421
rect 13348 8381 13360 8415
rect 13394 8412 13406 8415
rect 14090 8412 14096 8424
rect 13394 8384 14096 8412
rect 13394 8381 13406 8384
rect 13348 8375 13406 8381
rect 14090 8372 14096 8384
rect 14148 8372 14154 8424
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 15289 8415 15347 8421
rect 15289 8412 15301 8415
rect 14608 8384 15301 8412
rect 14608 8372 14614 8384
rect 15289 8381 15301 8384
rect 15335 8381 15347 8415
rect 18046 8412 18052 8424
rect 15289 8375 15347 8381
rect 16040 8384 18052 8412
rect 9876 8344 9904 8372
rect 8036 8316 9904 8344
rect 10128 8347 10186 8353
rect 10128 8313 10140 8347
rect 10174 8344 10186 8347
rect 10778 8344 10784 8356
rect 10174 8316 10784 8344
rect 10174 8313 10186 8316
rect 10128 8307 10186 8313
rect 10778 8304 10784 8316
rect 10836 8304 10842 8356
rect 13170 8304 13176 8356
rect 13228 8344 13234 8356
rect 13630 8344 13636 8356
rect 13228 8316 13636 8344
rect 13228 8304 13234 8316
rect 13630 8304 13636 8316
rect 13688 8344 13694 8356
rect 16040 8344 16068 8384
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 18417 8415 18475 8421
rect 18417 8381 18429 8415
rect 18463 8412 18475 8415
rect 19242 8412 19248 8424
rect 18463 8384 19248 8412
rect 18463 8381 18475 8384
rect 18417 8375 18475 8381
rect 19242 8372 19248 8384
rect 19300 8372 19306 8424
rect 19429 8415 19487 8421
rect 19429 8381 19441 8415
rect 19475 8412 19487 8415
rect 20548 8412 20576 8440
rect 19475 8384 20576 8412
rect 19475 8381 19487 8384
rect 19429 8375 19487 8381
rect 13688 8316 16068 8344
rect 16200 8347 16258 8353
rect 13688 8304 13694 8316
rect 16200 8313 16212 8347
rect 16246 8344 16258 8347
rect 16482 8344 16488 8356
rect 16246 8316 16488 8344
rect 16246 8313 16258 8316
rect 16200 8307 16258 8313
rect 16482 8304 16488 8316
rect 16540 8304 16546 8356
rect 17402 8344 17408 8356
rect 16592 8316 17408 8344
rect 9214 8236 9220 8288
rect 9272 8276 9278 8288
rect 9401 8279 9459 8285
rect 9401 8276 9413 8279
rect 9272 8248 9413 8276
rect 9272 8236 9278 8248
rect 9401 8245 9413 8248
rect 9447 8245 9459 8279
rect 9401 8239 9459 8245
rect 10962 8236 10968 8288
rect 11020 8276 11026 8288
rect 13814 8276 13820 8288
rect 11020 8248 13820 8276
rect 11020 8236 11026 8248
rect 13814 8236 13820 8248
rect 13872 8236 13878 8288
rect 14458 8276 14464 8288
rect 14419 8248 14464 8276
rect 14458 8236 14464 8248
rect 14516 8236 14522 8288
rect 15746 8236 15752 8288
rect 15804 8276 15810 8288
rect 16592 8276 16620 8316
rect 17402 8304 17408 8316
rect 17460 8304 17466 8356
rect 18969 8347 19027 8353
rect 18969 8313 18981 8347
rect 19015 8344 19027 8347
rect 19058 8344 19064 8356
rect 19015 8316 19064 8344
rect 19015 8313 19027 8316
rect 18969 8307 19027 8313
rect 19058 8304 19064 8316
rect 19116 8304 19122 8356
rect 19521 8347 19579 8353
rect 19521 8313 19533 8347
rect 19567 8344 19579 8347
rect 19978 8344 19984 8356
rect 19567 8316 19984 8344
rect 19567 8313 19579 8316
rect 19521 8307 19579 8313
rect 19978 8304 19984 8316
rect 20036 8304 20042 8356
rect 20070 8276 20076 8288
rect 15804 8248 16620 8276
rect 20031 8248 20076 8276
rect 15804 8236 15810 8248
rect 20070 8236 20076 8248
rect 20128 8236 20134 8288
rect 20438 8276 20444 8288
rect 20399 8248 20444 8276
rect 20438 8236 20444 8248
rect 20496 8236 20502 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 8570 8032 8576 8084
rect 8628 8072 8634 8084
rect 9033 8075 9091 8081
rect 9033 8072 9045 8075
rect 8628 8044 9045 8072
rect 8628 8032 8634 8044
rect 9033 8041 9045 8044
rect 9079 8041 9091 8075
rect 9033 8035 9091 8041
rect 10137 8075 10195 8081
rect 10137 8041 10149 8075
rect 10183 8072 10195 8075
rect 11054 8072 11060 8084
rect 10183 8044 11060 8072
rect 10183 8041 10195 8044
rect 10137 8035 10195 8041
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 11790 8032 11796 8084
rect 11848 8072 11854 8084
rect 11848 8044 13860 8072
rect 11848 8032 11854 8044
rect 10597 8007 10655 8013
rect 10597 7973 10609 8007
rect 10643 8004 10655 8007
rect 12618 8004 12624 8016
rect 10643 7976 12624 8004
rect 10643 7973 10655 7976
rect 10597 7967 10655 7973
rect 12618 7964 12624 7976
rect 12676 7964 12682 8016
rect 13170 8004 13176 8016
rect 13131 7976 13176 8004
rect 13170 7964 13176 7976
rect 13228 7964 13234 8016
rect 13832 8004 13860 8044
rect 13906 8032 13912 8084
rect 13964 8072 13970 8084
rect 14277 8075 14335 8081
rect 14277 8072 14289 8075
rect 13964 8044 14289 8072
rect 13964 8032 13970 8044
rect 14277 8041 14289 8044
rect 14323 8072 14335 8075
rect 14550 8072 14556 8084
rect 14323 8044 14556 8072
rect 14323 8041 14335 8044
rect 14277 8035 14335 8041
rect 14550 8032 14556 8044
rect 14608 8032 14614 8084
rect 15102 8032 15108 8084
rect 15160 8072 15166 8084
rect 17862 8072 17868 8084
rect 15160 8044 17868 8072
rect 15160 8032 15166 8044
rect 17862 8032 17868 8044
rect 17920 8032 17926 8084
rect 17954 8032 17960 8084
rect 18012 8072 18018 8084
rect 18049 8075 18107 8081
rect 18049 8072 18061 8075
rect 18012 8044 18061 8072
rect 18012 8032 18018 8044
rect 18049 8041 18061 8044
rect 18095 8041 18107 8075
rect 18049 8035 18107 8041
rect 20438 8032 20444 8084
rect 20496 8072 20502 8084
rect 20901 8075 20959 8081
rect 20901 8072 20913 8075
rect 20496 8044 20913 8072
rect 20496 8032 20502 8044
rect 20901 8041 20913 8044
rect 20947 8041 20959 8075
rect 20901 8035 20959 8041
rect 19242 8004 19248 8016
rect 13832 7976 19248 8004
rect 19242 7964 19248 7976
rect 19300 7964 19306 8016
rect 8941 7939 8999 7945
rect 8941 7905 8953 7939
rect 8987 7936 8999 7939
rect 9677 7939 9735 7945
rect 9677 7936 9689 7939
rect 8987 7908 9689 7936
rect 8987 7905 8999 7908
rect 8941 7899 8999 7905
rect 9677 7905 9689 7908
rect 9723 7905 9735 7939
rect 9677 7899 9735 7905
rect 9858 7896 9864 7948
rect 9916 7936 9922 7948
rect 10505 7939 10563 7945
rect 10505 7936 10517 7939
rect 9916 7908 10517 7936
rect 9916 7896 9922 7908
rect 10505 7905 10517 7908
rect 10551 7936 10563 7939
rect 10962 7936 10968 7948
rect 10551 7908 10968 7936
rect 10551 7905 10563 7908
rect 10505 7899 10563 7905
rect 10962 7896 10968 7908
rect 11020 7896 11026 7948
rect 11416 7939 11474 7945
rect 11416 7905 11428 7939
rect 11462 7936 11474 7939
rect 12894 7936 12900 7948
rect 11462 7908 12900 7936
rect 11462 7905 11474 7908
rect 11416 7899 11474 7905
rect 12894 7896 12900 7908
rect 12952 7896 12958 7948
rect 13538 7936 13544 7948
rect 13280 7908 13544 7936
rect 9214 7868 9220 7880
rect 9175 7840 9220 7868
rect 9214 7828 9220 7840
rect 9272 7828 9278 7880
rect 10778 7868 10784 7880
rect 10739 7840 10784 7868
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 11149 7871 11207 7877
rect 11149 7837 11161 7871
rect 11195 7837 11207 7871
rect 11149 7831 11207 7837
rect 8573 7803 8631 7809
rect 8573 7769 8585 7803
rect 8619 7800 8631 7803
rect 8662 7800 8668 7812
rect 8619 7772 8668 7800
rect 8619 7769 8631 7772
rect 8573 7763 8631 7769
rect 8662 7760 8668 7772
rect 8720 7760 8726 7812
rect 9950 7760 9956 7812
rect 10008 7800 10014 7812
rect 11164 7800 11192 7831
rect 13170 7828 13176 7880
rect 13228 7868 13234 7880
rect 13280 7877 13308 7908
rect 13538 7896 13544 7908
rect 13596 7896 13602 7948
rect 14185 7939 14243 7945
rect 14185 7905 14197 7939
rect 14231 7936 14243 7939
rect 15194 7936 15200 7948
rect 14231 7908 15200 7936
rect 14231 7905 14243 7908
rect 14185 7899 14243 7905
rect 15194 7896 15200 7908
rect 15252 7896 15258 7948
rect 15565 7939 15623 7945
rect 15565 7905 15577 7939
rect 15611 7936 15623 7939
rect 15654 7936 15660 7948
rect 15611 7908 15660 7936
rect 15611 7905 15623 7908
rect 15565 7899 15623 7905
rect 15654 7896 15660 7908
rect 15712 7896 15718 7948
rect 15838 7945 15844 7948
rect 15832 7936 15844 7945
rect 15799 7908 15844 7936
rect 15832 7899 15844 7908
rect 15838 7896 15844 7899
rect 15896 7896 15902 7948
rect 16114 7896 16120 7948
rect 16172 7936 16178 7948
rect 17221 7939 17279 7945
rect 17221 7936 17233 7939
rect 16172 7908 17233 7936
rect 16172 7896 16178 7908
rect 17221 7905 17233 7908
rect 17267 7905 17279 7939
rect 17221 7899 17279 7905
rect 17586 7896 17592 7948
rect 17644 7936 17650 7948
rect 18141 7939 18199 7945
rect 18141 7936 18153 7939
rect 17644 7908 18153 7936
rect 17644 7896 17650 7908
rect 18141 7905 18153 7908
rect 18187 7936 18199 7939
rect 18874 7936 18880 7948
rect 18187 7908 18880 7936
rect 18187 7905 18199 7908
rect 18141 7899 18199 7905
rect 18874 7896 18880 7908
rect 18932 7896 18938 7948
rect 19978 7936 19984 7948
rect 19939 7908 19984 7936
rect 19978 7896 19984 7908
rect 20036 7896 20042 7948
rect 13265 7871 13323 7877
rect 13265 7868 13277 7871
rect 13228 7840 13277 7868
rect 13228 7828 13234 7840
rect 13265 7837 13277 7840
rect 13311 7837 13323 7871
rect 13265 7831 13323 7837
rect 13449 7871 13507 7877
rect 13449 7837 13461 7871
rect 13495 7837 13507 7871
rect 14458 7868 14464 7880
rect 14419 7840 14464 7868
rect 13449 7831 13507 7837
rect 10008 7772 11192 7800
rect 13464 7800 13492 7831
rect 14458 7828 14464 7840
rect 14516 7828 14522 7880
rect 13906 7800 13912 7812
rect 13464 7772 13912 7800
rect 10008 7760 10014 7772
rect 13906 7760 13912 7772
rect 13964 7800 13970 7812
rect 14476 7800 14504 7828
rect 13964 7772 14504 7800
rect 13964 7760 13970 7772
rect 3418 7692 3424 7744
rect 3476 7732 3482 7744
rect 11790 7732 11796 7744
rect 3476 7704 11796 7732
rect 3476 7692 3482 7704
rect 11790 7692 11796 7704
rect 11848 7692 11854 7744
rect 12066 7692 12072 7744
rect 12124 7732 12130 7744
rect 12529 7735 12587 7741
rect 12529 7732 12541 7735
rect 12124 7704 12541 7732
rect 12124 7692 12130 7704
rect 12529 7701 12541 7704
rect 12575 7701 12587 7735
rect 12529 7695 12587 7701
rect 12805 7735 12863 7741
rect 12805 7701 12817 7735
rect 12851 7732 12863 7735
rect 12986 7732 12992 7744
rect 12851 7704 12992 7732
rect 12851 7701 12863 7704
rect 12805 7695 12863 7701
rect 12986 7692 12992 7704
rect 13044 7692 13050 7744
rect 13078 7692 13084 7744
rect 13136 7732 13142 7744
rect 13817 7735 13875 7741
rect 13817 7732 13829 7735
rect 13136 7704 13829 7732
rect 13136 7692 13142 7704
rect 13817 7701 13829 7704
rect 13863 7701 13875 7735
rect 15212 7732 15240 7896
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7837 18291 7871
rect 18233 7831 18291 7837
rect 20073 7871 20131 7877
rect 20073 7837 20085 7871
rect 20119 7868 20131 7871
rect 20162 7868 20168 7880
rect 20119 7840 20168 7868
rect 20119 7837 20131 7840
rect 20073 7831 20131 7837
rect 16500 7772 17816 7800
rect 16500 7732 16528 7772
rect 15212 7704 16528 7732
rect 16945 7735 17003 7741
rect 13817 7695 13875 7701
rect 16945 7701 16957 7735
rect 16991 7732 17003 7735
rect 17126 7732 17132 7744
rect 16991 7704 17132 7732
rect 16991 7701 17003 7704
rect 16945 7695 17003 7701
rect 17126 7692 17132 7704
rect 17184 7692 17190 7744
rect 17678 7732 17684 7744
rect 17639 7704 17684 7732
rect 17678 7692 17684 7704
rect 17736 7692 17742 7744
rect 17788 7732 17816 7772
rect 17862 7760 17868 7812
rect 17920 7800 17926 7812
rect 18248 7800 18276 7831
rect 20162 7828 20168 7840
rect 20220 7828 20226 7880
rect 20257 7871 20315 7877
rect 20257 7837 20269 7871
rect 20303 7868 20315 7871
rect 20530 7868 20536 7880
rect 20303 7840 20536 7868
rect 20303 7837 20315 7840
rect 20257 7831 20315 7837
rect 20530 7828 20536 7840
rect 20588 7828 20594 7880
rect 20438 7800 20444 7812
rect 17920 7772 18276 7800
rect 18340 7772 20444 7800
rect 17920 7760 17926 7772
rect 18340 7732 18368 7772
rect 20438 7760 20444 7772
rect 20496 7760 20502 7812
rect 17788 7704 18368 7732
rect 19150 7692 19156 7744
rect 19208 7732 19214 7744
rect 19334 7732 19340 7744
rect 19208 7704 19340 7732
rect 19208 7692 19214 7704
rect 19334 7692 19340 7704
rect 19392 7692 19398 7744
rect 19610 7732 19616 7744
rect 19571 7704 19616 7732
rect 19610 7692 19616 7704
rect 19668 7692 19674 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 8205 7531 8263 7537
rect 8205 7497 8217 7531
rect 8251 7528 8263 7531
rect 11146 7528 11152 7540
rect 8251 7500 11152 7528
rect 8251 7497 8263 7500
rect 8205 7491 8263 7497
rect 11146 7488 11152 7500
rect 11204 7488 11210 7540
rect 15013 7531 15071 7537
rect 15013 7528 15025 7531
rect 13188 7500 15025 7528
rect 10597 7463 10655 7469
rect 10597 7429 10609 7463
rect 10643 7460 10655 7463
rect 10778 7460 10784 7472
rect 10643 7432 10784 7460
rect 10643 7429 10655 7432
rect 10597 7423 10655 7429
rect 10778 7420 10784 7432
rect 10836 7420 10842 7472
rect 12894 7420 12900 7472
rect 12952 7460 12958 7472
rect 13188 7460 13216 7500
rect 15013 7497 15025 7500
rect 15059 7497 15071 7531
rect 15013 7491 15071 7497
rect 12952 7432 13216 7460
rect 12952 7420 12958 7432
rect 8849 7395 8907 7401
rect 8849 7361 8861 7395
rect 8895 7392 8907 7395
rect 11977 7395 12035 7401
rect 8895 7364 9352 7392
rect 8895 7361 8907 7364
rect 8849 7355 8907 7361
rect 9324 7336 9352 7364
rect 11977 7361 11989 7395
rect 12023 7392 12035 7395
rect 12066 7392 12072 7404
rect 12023 7364 12072 7392
rect 12023 7361 12035 7364
rect 11977 7355 12035 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 13078 7392 13084 7404
rect 13039 7364 13084 7392
rect 13078 7352 13084 7364
rect 13136 7352 13142 7404
rect 13188 7401 13216 7432
rect 13262 7420 13268 7472
rect 13320 7460 13326 7472
rect 13538 7460 13544 7472
rect 13320 7432 13544 7460
rect 13320 7420 13326 7432
rect 13538 7420 13544 7432
rect 13596 7420 13602 7472
rect 13173 7395 13231 7401
rect 13173 7361 13185 7395
rect 13219 7361 13231 7395
rect 13173 7355 13231 7361
rect 15838 7352 15844 7404
rect 15896 7392 15902 7404
rect 15933 7395 15991 7401
rect 15933 7392 15945 7395
rect 15896 7364 15945 7392
rect 15896 7352 15902 7364
rect 15933 7361 15945 7364
rect 15979 7392 15991 7395
rect 15979 7364 16436 7392
rect 15979 7361 15991 7364
rect 15933 7355 15991 7361
rect 9217 7327 9275 7333
rect 9217 7293 9229 7327
rect 9263 7293 9275 7327
rect 9217 7287 9275 7293
rect 9232 7256 9260 7287
rect 9306 7284 9312 7336
rect 9364 7324 9370 7336
rect 9473 7327 9531 7333
rect 9473 7324 9485 7327
rect 9364 7296 9485 7324
rect 9364 7284 9370 7296
rect 9473 7293 9485 7296
rect 9519 7293 9531 7327
rect 12986 7324 12992 7336
rect 12947 7296 12992 7324
rect 9473 7287 9531 7293
rect 12986 7284 12992 7296
rect 13044 7284 13050 7336
rect 13446 7284 13452 7336
rect 13504 7324 13510 7336
rect 13906 7333 13912 7336
rect 13633 7327 13691 7333
rect 13633 7324 13645 7327
rect 13504 7296 13645 7324
rect 13504 7284 13510 7296
rect 13633 7293 13645 7296
rect 13679 7293 13691 7327
rect 13900 7324 13912 7333
rect 13867 7296 13912 7324
rect 13633 7287 13691 7293
rect 13900 7287 13912 7296
rect 13906 7284 13912 7287
rect 13964 7284 13970 7336
rect 15657 7327 15715 7333
rect 15657 7293 15669 7327
rect 15703 7324 15715 7327
rect 16114 7324 16120 7336
rect 15703 7296 16120 7324
rect 15703 7293 15715 7296
rect 15657 7287 15715 7293
rect 16114 7284 16120 7296
rect 16172 7284 16178 7336
rect 16301 7327 16359 7333
rect 16301 7293 16313 7327
rect 16347 7293 16359 7327
rect 16301 7287 16359 7293
rect 9582 7256 9588 7268
rect 9232 7228 9588 7256
rect 9582 7216 9588 7228
rect 9640 7216 9646 7268
rect 11701 7259 11759 7265
rect 11701 7225 11713 7259
rect 11747 7256 11759 7259
rect 13262 7256 13268 7268
rect 11747 7228 13268 7256
rect 11747 7225 11759 7228
rect 11701 7219 11759 7225
rect 13262 7216 13268 7228
rect 13320 7216 13326 7268
rect 16316 7256 16344 7287
rect 15672 7228 16344 7256
rect 15672 7200 15700 7228
rect 8570 7188 8576 7200
rect 8531 7160 8576 7188
rect 8570 7148 8576 7160
rect 8628 7148 8634 7200
rect 8665 7191 8723 7197
rect 8665 7157 8677 7191
rect 8711 7188 8723 7191
rect 9674 7188 9680 7200
rect 8711 7160 9680 7188
rect 8711 7157 8723 7160
rect 8665 7151 8723 7157
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 11333 7191 11391 7197
rect 11333 7157 11345 7191
rect 11379 7188 11391 7191
rect 11606 7188 11612 7200
rect 11379 7160 11612 7188
rect 11379 7157 11391 7160
rect 11333 7151 11391 7157
rect 11606 7148 11612 7160
rect 11664 7148 11670 7200
rect 11793 7191 11851 7197
rect 11793 7157 11805 7191
rect 11839 7188 11851 7191
rect 12621 7191 12679 7197
rect 12621 7188 12633 7191
rect 11839 7160 12633 7188
rect 11839 7157 11851 7160
rect 11793 7151 11851 7157
rect 12621 7157 12633 7160
rect 12667 7157 12679 7191
rect 15286 7188 15292 7200
rect 15247 7160 15292 7188
rect 12621 7151 12679 7157
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 15654 7148 15660 7200
rect 15712 7148 15718 7200
rect 15746 7148 15752 7200
rect 15804 7188 15810 7200
rect 16408 7188 16436 7364
rect 18782 7324 18788 7336
rect 18743 7296 18788 7324
rect 18782 7284 18788 7296
rect 18840 7284 18846 7336
rect 19886 7324 19892 7336
rect 18984 7296 19892 7324
rect 16568 7259 16626 7265
rect 16568 7225 16580 7259
rect 16614 7256 16626 7259
rect 16850 7256 16856 7268
rect 16614 7228 16856 7256
rect 16614 7225 16626 7228
rect 16568 7219 16626 7225
rect 16850 7216 16856 7228
rect 16908 7216 16914 7268
rect 17310 7216 17316 7268
rect 17368 7256 17374 7268
rect 18984 7256 19012 7296
rect 19886 7284 19892 7296
rect 19944 7284 19950 7336
rect 20254 7284 20260 7336
rect 20312 7324 20318 7336
rect 20441 7327 20499 7333
rect 20441 7324 20453 7327
rect 20312 7296 20453 7324
rect 20312 7284 20318 7296
rect 20441 7293 20453 7296
rect 20487 7293 20499 7327
rect 20441 7287 20499 7293
rect 17368 7228 19012 7256
rect 19052 7259 19110 7265
rect 17368 7216 17374 7228
rect 19052 7225 19064 7259
rect 19098 7256 19110 7259
rect 20530 7256 20536 7268
rect 19098 7228 20536 7256
rect 19098 7225 19110 7228
rect 19052 7219 19110 7225
rect 20530 7216 20536 7228
rect 20588 7216 20594 7268
rect 17494 7188 17500 7200
rect 15804 7160 15849 7188
rect 16408 7160 17500 7188
rect 15804 7148 15810 7160
rect 17494 7148 17500 7160
rect 17552 7188 17558 7200
rect 17681 7191 17739 7197
rect 17681 7188 17693 7191
rect 17552 7160 17693 7188
rect 17552 7148 17558 7160
rect 17681 7157 17693 7160
rect 17727 7157 17739 7191
rect 17681 7151 17739 7157
rect 19242 7148 19248 7200
rect 19300 7188 19306 7200
rect 19702 7188 19708 7200
rect 19300 7160 19708 7188
rect 19300 7148 19306 7160
rect 19702 7148 19708 7160
rect 19760 7188 19766 7200
rect 20165 7191 20223 7197
rect 20165 7188 20177 7191
rect 19760 7160 20177 7188
rect 19760 7148 19766 7160
rect 20165 7157 20177 7160
rect 20211 7157 20223 7191
rect 20622 7188 20628 7200
rect 20583 7160 20628 7188
rect 20165 7151 20223 7157
rect 20622 7148 20628 7160
rect 20680 7148 20686 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 9306 6984 9312 6996
rect 9267 6956 9312 6984
rect 9306 6944 9312 6956
rect 9364 6944 9370 6996
rect 9674 6984 9680 6996
rect 9635 6956 9680 6984
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 12618 6944 12624 6996
rect 12676 6984 12682 6996
rect 13078 6984 13084 6996
rect 12676 6956 13084 6984
rect 12676 6944 12682 6956
rect 13078 6944 13084 6956
rect 13136 6944 13142 6996
rect 15746 6944 15752 6996
rect 15804 6984 15810 6996
rect 16209 6987 16267 6993
rect 16209 6984 16221 6987
rect 15804 6956 16221 6984
rect 15804 6944 15810 6956
rect 16209 6953 16221 6956
rect 16255 6953 16267 6987
rect 16209 6947 16267 6953
rect 16669 6987 16727 6993
rect 16669 6953 16681 6987
rect 16715 6984 16727 6987
rect 16758 6984 16764 6996
rect 16715 6956 16764 6984
rect 16715 6953 16727 6956
rect 16669 6947 16727 6953
rect 16758 6944 16764 6956
rect 16816 6944 16822 6996
rect 17310 6944 17316 6996
rect 17368 6984 17374 6996
rect 17589 6987 17647 6993
rect 17589 6984 17601 6987
rect 17368 6956 17601 6984
rect 17368 6944 17374 6956
rect 17589 6953 17601 6956
rect 17635 6953 17647 6987
rect 17589 6947 17647 6953
rect 19153 6987 19211 6993
rect 19153 6953 19165 6987
rect 19199 6984 19211 6987
rect 20070 6984 20076 6996
rect 19199 6956 20076 6984
rect 19199 6953 19211 6956
rect 19153 6947 19211 6953
rect 20070 6944 20076 6956
rect 20128 6944 20134 6996
rect 10045 6919 10103 6925
rect 10045 6885 10057 6919
rect 10091 6916 10103 6919
rect 11146 6916 11152 6928
rect 10091 6888 11152 6916
rect 10091 6885 10103 6888
rect 10045 6879 10103 6885
rect 11146 6876 11152 6888
rect 11204 6876 11210 6928
rect 11508 6919 11566 6925
rect 11508 6885 11520 6919
rect 11554 6916 11566 6919
rect 12066 6916 12072 6928
rect 11554 6888 12072 6916
rect 11554 6885 11566 6888
rect 11508 6879 11566 6885
rect 12066 6876 12072 6888
rect 12124 6876 12130 6928
rect 12986 6876 12992 6928
rect 13044 6916 13050 6928
rect 14185 6919 14243 6925
rect 14185 6916 14197 6919
rect 13044 6888 14197 6916
rect 13044 6876 13050 6888
rect 14185 6885 14197 6888
rect 14231 6916 14243 6919
rect 16577 6919 16635 6925
rect 16577 6916 16589 6919
rect 14231 6888 16589 6916
rect 14231 6885 14243 6888
rect 14185 6879 14243 6885
rect 16577 6885 16589 6888
rect 16623 6885 16635 6919
rect 16577 6879 16635 6885
rect 17512 6888 17724 6916
rect 8196 6851 8254 6857
rect 8196 6817 8208 6851
rect 8242 6848 8254 6851
rect 8754 6848 8760 6860
rect 8242 6820 8760 6848
rect 8242 6817 8254 6820
rect 8196 6811 8254 6817
rect 8754 6808 8760 6820
rect 8812 6848 8818 6860
rect 10870 6848 10876 6860
rect 8812 6820 10272 6848
rect 10831 6820 10876 6848
rect 8812 6808 8818 6820
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6749 7987 6783
rect 10134 6780 10140 6792
rect 10095 6752 10140 6780
rect 7929 6743 7987 6749
rect 7466 6604 7472 6656
rect 7524 6644 7530 6656
rect 7944 6644 7972 6743
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10244 6789 10272 6820
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 10962 6808 10968 6860
rect 11020 6848 11026 6860
rect 15010 6848 15016 6860
rect 11020 6820 15016 6848
rect 11020 6808 11026 6820
rect 15010 6808 15016 6820
rect 15068 6808 15074 6860
rect 17512 6848 17540 6888
rect 16776 6820 17540 6848
rect 17696 6848 17724 6888
rect 18966 6876 18972 6928
rect 19024 6916 19030 6928
rect 20165 6919 20223 6925
rect 19024 6888 19748 6916
rect 19024 6876 19030 6888
rect 18233 6851 18291 6857
rect 18233 6848 18245 6851
rect 17696 6820 18245 6848
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 11054 6740 11060 6792
rect 11112 6780 11118 6792
rect 11241 6783 11299 6789
rect 11241 6780 11253 6783
rect 11112 6752 11253 6780
rect 11112 6740 11118 6752
rect 11241 6749 11253 6752
rect 11287 6749 11299 6783
rect 11241 6743 11299 6749
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6780 13415 6783
rect 13630 6780 13636 6792
rect 13403 6752 13636 6780
rect 13403 6749 13415 6752
rect 13357 6743 13415 6749
rect 13630 6740 13636 6752
rect 13688 6740 13694 6792
rect 14277 6783 14335 6789
rect 14277 6749 14289 6783
rect 14323 6749 14335 6783
rect 14458 6780 14464 6792
rect 14419 6752 14464 6780
rect 14277 6743 14335 6749
rect 14292 6712 14320 6743
rect 14458 6740 14464 6752
rect 14516 6740 14522 6792
rect 15562 6740 15568 6792
rect 15620 6780 15626 6792
rect 16776 6780 16804 6820
rect 18233 6817 18245 6820
rect 18279 6817 18291 6851
rect 18233 6811 18291 6817
rect 19245 6851 19303 6857
rect 19245 6817 19257 6851
rect 19291 6848 19303 6851
rect 19610 6848 19616 6860
rect 19291 6820 19616 6848
rect 19291 6817 19303 6820
rect 19245 6811 19303 6817
rect 19610 6808 19616 6820
rect 19668 6808 19674 6860
rect 19720 6848 19748 6888
rect 20165 6885 20177 6919
rect 20211 6916 20223 6919
rect 20898 6916 20904 6928
rect 20211 6888 20904 6916
rect 20211 6885 20223 6888
rect 20165 6879 20223 6885
rect 20898 6876 20904 6888
rect 20956 6876 20962 6928
rect 20257 6851 20315 6857
rect 20257 6848 20269 6851
rect 19720 6820 20269 6848
rect 20257 6817 20269 6820
rect 20303 6817 20315 6851
rect 20257 6811 20315 6817
rect 15620 6752 16804 6780
rect 15620 6740 15626 6752
rect 16850 6740 16856 6792
rect 16908 6780 16914 6792
rect 16908 6752 17001 6780
rect 16908 6740 16914 6752
rect 17034 6740 17040 6792
rect 17092 6780 17098 6792
rect 17681 6783 17739 6789
rect 17681 6780 17693 6783
rect 17092 6752 17693 6780
rect 17092 6740 17098 6752
rect 17681 6749 17693 6752
rect 17727 6749 17739 6783
rect 17862 6780 17868 6792
rect 17823 6752 17868 6780
rect 17681 6743 17739 6749
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 19429 6783 19487 6789
rect 18432 6752 19288 6780
rect 14366 6712 14372 6724
rect 14292 6684 14372 6712
rect 14366 6672 14372 6684
rect 14424 6672 14430 6724
rect 15286 6672 15292 6724
rect 15344 6712 15350 6724
rect 15930 6712 15936 6724
rect 15344 6684 15936 6712
rect 15344 6672 15350 6684
rect 15930 6672 15936 6684
rect 15988 6672 15994 6724
rect 16868 6712 16896 6740
rect 17880 6712 17908 6740
rect 18432 6721 18460 6752
rect 16868 6684 17908 6712
rect 18417 6715 18475 6721
rect 18417 6681 18429 6715
rect 18463 6681 18475 6715
rect 19260 6712 19288 6752
rect 19429 6749 19441 6783
rect 19475 6780 19487 6783
rect 19702 6780 19708 6792
rect 19475 6752 19708 6780
rect 19475 6749 19487 6752
rect 19429 6743 19487 6749
rect 19702 6740 19708 6752
rect 19760 6740 19766 6792
rect 20346 6740 20352 6792
rect 20404 6780 20410 6792
rect 20404 6752 20449 6780
rect 20404 6740 20410 6752
rect 21910 6712 21916 6724
rect 19260 6684 21916 6712
rect 18417 6675 18475 6681
rect 21910 6672 21916 6684
rect 21968 6672 21974 6724
rect 9582 6644 9588 6656
rect 7524 6616 9588 6644
rect 7524 6604 7530 6616
rect 9582 6604 9588 6616
rect 9640 6644 9646 6656
rect 10689 6647 10747 6653
rect 10689 6644 10701 6647
rect 9640 6616 10701 6644
rect 9640 6604 9646 6616
rect 10689 6613 10701 6616
rect 10735 6644 10747 6647
rect 11054 6644 11060 6656
rect 10735 6616 11060 6644
rect 10735 6613 10747 6616
rect 10689 6607 10747 6613
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 12618 6644 12624 6656
rect 12579 6616 12624 6644
rect 12618 6604 12624 6616
rect 12676 6604 12682 6656
rect 13722 6604 13728 6656
rect 13780 6644 13786 6656
rect 13817 6647 13875 6653
rect 13817 6644 13829 6647
rect 13780 6616 13829 6644
rect 13780 6604 13786 6616
rect 13817 6613 13829 6616
rect 13863 6613 13875 6647
rect 13817 6607 13875 6613
rect 15470 6604 15476 6656
rect 15528 6644 15534 6656
rect 17034 6644 17040 6656
rect 15528 6616 17040 6644
rect 15528 6604 15534 6616
rect 17034 6604 17040 6616
rect 17092 6604 17098 6656
rect 17221 6647 17279 6653
rect 17221 6613 17233 6647
rect 17267 6644 17279 6647
rect 17310 6644 17316 6656
rect 17267 6616 17316 6644
rect 17267 6613 17279 6616
rect 17221 6607 17279 6613
rect 17310 6604 17316 6616
rect 17368 6604 17374 6656
rect 18690 6604 18696 6656
rect 18748 6644 18754 6656
rect 18785 6647 18843 6653
rect 18785 6644 18797 6647
rect 18748 6616 18797 6644
rect 18748 6604 18754 6616
rect 18785 6613 18797 6616
rect 18831 6613 18843 6647
rect 18785 6607 18843 6613
rect 18966 6604 18972 6656
rect 19024 6644 19030 6656
rect 19797 6647 19855 6653
rect 19797 6644 19809 6647
rect 19024 6616 19809 6644
rect 19024 6604 19030 6616
rect 19797 6613 19809 6616
rect 19843 6613 19855 6647
rect 19797 6607 19855 6613
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 8570 6400 8576 6452
rect 8628 6440 8634 6452
rect 9125 6443 9183 6449
rect 9125 6440 9137 6443
rect 8628 6412 9137 6440
rect 8628 6400 8634 6412
rect 9125 6409 9137 6412
rect 9171 6409 9183 6443
rect 10134 6440 10140 6452
rect 10095 6412 10140 6440
rect 9125 6403 9183 6409
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 11146 6440 11152 6452
rect 11107 6412 11152 6440
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 13262 6440 13268 6452
rect 13223 6412 13268 6440
rect 13262 6400 13268 6412
rect 13320 6400 13326 6452
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 15841 6443 15899 6449
rect 15841 6440 15853 6443
rect 13872 6412 15853 6440
rect 13872 6400 13878 6412
rect 15841 6409 15853 6412
rect 15887 6409 15899 6443
rect 15841 6403 15899 6409
rect 18141 6443 18199 6449
rect 18141 6409 18153 6443
rect 18187 6440 18199 6443
rect 19058 6440 19064 6452
rect 18187 6412 19064 6440
rect 18187 6409 18199 6412
rect 18141 6403 18199 6409
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 19426 6440 19432 6452
rect 19168 6412 19432 6440
rect 8754 6332 8760 6384
rect 8812 6372 8818 6384
rect 8849 6375 8907 6381
rect 8849 6372 8861 6375
rect 8812 6344 8861 6372
rect 8812 6332 8818 6344
rect 8849 6341 8861 6344
rect 8895 6372 8907 6375
rect 8895 6344 9720 6372
rect 8895 6341 8907 6344
rect 8849 6335 8907 6341
rect 7466 6304 7472 6316
rect 7427 6276 7472 6304
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 9692 6313 9720 6344
rect 12894 6332 12900 6384
rect 12952 6372 12958 6384
rect 14829 6375 14887 6381
rect 12952 6344 13860 6372
rect 12952 6332 12958 6344
rect 9677 6307 9735 6313
rect 9677 6273 9689 6307
rect 9723 6273 9735 6307
rect 9677 6267 9735 6273
rect 10318 6264 10324 6316
rect 10376 6304 10382 6316
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 10376 6276 10793 6304
rect 10376 6264 10382 6276
rect 10781 6273 10793 6276
rect 10827 6304 10839 6307
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 10827 6276 11713 6304
rect 10827 6273 10839 6276
rect 10781 6267 10839 6273
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 12986 6264 12992 6316
rect 13044 6304 13050 6316
rect 13262 6304 13268 6316
rect 13044 6276 13268 6304
rect 13044 6264 13050 6276
rect 13262 6264 13268 6276
rect 13320 6264 13326 6316
rect 13832 6313 13860 6344
rect 14829 6341 14841 6375
rect 14875 6372 14887 6375
rect 15746 6372 15752 6384
rect 14875 6344 15752 6372
rect 14875 6341 14887 6344
rect 14829 6335 14887 6341
rect 15746 6332 15752 6344
rect 15804 6332 15810 6384
rect 16574 6372 16580 6384
rect 15847 6344 16580 6372
rect 13817 6307 13875 6313
rect 13817 6273 13829 6307
rect 13863 6273 13875 6307
rect 13817 6267 13875 6273
rect 15010 6264 15016 6316
rect 15068 6304 15074 6316
rect 15289 6307 15347 6313
rect 15289 6304 15301 6307
rect 15068 6276 15301 6304
rect 15068 6264 15074 6276
rect 15289 6273 15301 6276
rect 15335 6273 15347 6307
rect 15289 6267 15347 6273
rect 15378 6264 15384 6316
rect 15436 6304 15442 6316
rect 15436 6276 15481 6304
rect 15436 6264 15442 6276
rect 7742 6245 7748 6248
rect 7736 6236 7748 6245
rect 7655 6208 7748 6236
rect 7736 6199 7748 6208
rect 7800 6236 7806 6248
rect 10336 6236 10364 6264
rect 7800 6208 10364 6236
rect 10597 6239 10655 6245
rect 7742 6196 7748 6199
rect 7800 6196 7806 6208
rect 10597 6205 10609 6239
rect 10643 6236 10655 6239
rect 10686 6236 10692 6248
rect 10643 6208 10692 6236
rect 10643 6205 10655 6208
rect 10597 6199 10655 6205
rect 10686 6196 10692 6208
rect 10744 6196 10750 6248
rect 11517 6239 11575 6245
rect 11517 6205 11529 6239
rect 11563 6236 11575 6239
rect 15847 6236 15875 6344
rect 16574 6332 16580 6344
rect 16632 6332 16638 6384
rect 16666 6332 16672 6384
rect 16724 6372 16730 6384
rect 19168 6372 19196 6412
rect 19426 6400 19432 6412
rect 19484 6400 19490 6452
rect 20530 6440 20536 6452
rect 20491 6412 20536 6440
rect 20530 6400 20536 6412
rect 20588 6400 20594 6452
rect 16724 6344 18736 6372
rect 16724 6332 16730 6344
rect 16485 6307 16543 6313
rect 16485 6273 16497 6307
rect 16531 6304 16543 6307
rect 17126 6304 17132 6316
rect 16531 6276 17132 6304
rect 16531 6273 16543 6276
rect 16485 6267 16543 6273
rect 17126 6264 17132 6276
rect 17184 6264 17190 6316
rect 17310 6304 17316 6316
rect 17271 6276 17316 6304
rect 17310 6264 17316 6276
rect 17368 6264 17374 6316
rect 17494 6304 17500 6316
rect 17455 6276 17500 6304
rect 17494 6264 17500 6276
rect 17552 6264 17558 6316
rect 11563 6208 15875 6236
rect 11563 6205 11575 6208
rect 11517 6199 11575 6205
rect 15930 6196 15936 6248
rect 15988 6236 15994 6248
rect 16209 6239 16267 6245
rect 16209 6236 16221 6239
rect 15988 6208 16221 6236
rect 15988 6196 15994 6208
rect 16209 6205 16221 6208
rect 16255 6205 16267 6239
rect 16209 6199 16267 6205
rect 17221 6239 17279 6245
rect 17221 6205 17233 6239
rect 17267 6236 17279 6239
rect 17678 6236 17684 6248
rect 17267 6208 17684 6236
rect 17267 6205 17279 6208
rect 17221 6199 17279 6205
rect 17678 6196 17684 6208
rect 17736 6196 17742 6248
rect 10505 6171 10563 6177
rect 10505 6137 10517 6171
rect 10551 6168 10563 6171
rect 11698 6168 11704 6180
rect 10551 6140 11704 6168
rect 10551 6137 10563 6140
rect 10505 6131 10563 6137
rect 11698 6128 11704 6140
rect 11756 6128 11762 6180
rect 13630 6168 13636 6180
rect 13591 6140 13636 6168
rect 13630 6128 13636 6140
rect 13688 6128 13694 6180
rect 13722 6128 13728 6180
rect 13780 6168 13786 6180
rect 15197 6171 15255 6177
rect 13780 6140 13825 6168
rect 13780 6128 13786 6140
rect 15197 6137 15209 6171
rect 15243 6168 15255 6171
rect 16022 6168 16028 6180
rect 15243 6140 16028 6168
rect 15243 6137 15255 6140
rect 15197 6131 15255 6137
rect 16022 6128 16028 6140
rect 16080 6128 16086 6180
rect 16114 6128 16120 6180
rect 16172 6168 16178 6180
rect 18046 6168 18052 6180
rect 16172 6140 18052 6168
rect 16172 6128 16178 6140
rect 18046 6128 18052 6140
rect 18104 6128 18110 6180
rect 18414 6128 18420 6180
rect 18472 6168 18478 6180
rect 18509 6171 18567 6177
rect 18509 6168 18521 6171
rect 18472 6140 18521 6168
rect 18472 6128 18478 6140
rect 18509 6137 18521 6140
rect 18555 6137 18567 6171
rect 18708 6168 18736 6344
rect 18800 6344 19196 6372
rect 18800 6313 18828 6344
rect 18785 6307 18843 6313
rect 18785 6273 18797 6307
rect 18831 6273 18843 6307
rect 18785 6267 18843 6273
rect 19058 6196 19064 6248
rect 19116 6236 19122 6248
rect 19153 6239 19211 6245
rect 19153 6236 19165 6239
rect 19116 6208 19165 6236
rect 19116 6196 19122 6208
rect 19153 6205 19165 6208
rect 19199 6205 19211 6239
rect 20254 6236 20260 6248
rect 19153 6199 19211 6205
rect 19251 6208 20260 6236
rect 19251 6168 19279 6208
rect 20254 6196 20260 6208
rect 20312 6196 20318 6248
rect 20714 6196 20720 6248
rect 20772 6236 20778 6248
rect 20809 6239 20867 6245
rect 20809 6236 20821 6239
rect 20772 6208 20821 6236
rect 20772 6196 20778 6208
rect 20809 6205 20821 6208
rect 20855 6205 20867 6239
rect 20809 6199 20867 6205
rect 18708 6140 19279 6168
rect 18509 6131 18567 6137
rect 19334 6128 19340 6180
rect 19392 6177 19398 6180
rect 19392 6171 19456 6177
rect 19392 6137 19410 6171
rect 19444 6137 19456 6171
rect 19392 6131 19456 6137
rect 19392 6128 19398 6131
rect 9490 6100 9496 6112
rect 9451 6072 9496 6100
rect 9490 6060 9496 6072
rect 9548 6060 9554 6112
rect 9585 6103 9643 6109
rect 9585 6069 9597 6103
rect 9631 6100 9643 6103
rect 9674 6100 9680 6112
rect 9631 6072 9680 6100
rect 9631 6069 9643 6072
rect 9585 6063 9643 6069
rect 9674 6060 9680 6072
rect 9732 6060 9738 6112
rect 11609 6103 11667 6109
rect 11609 6069 11621 6103
rect 11655 6100 11667 6103
rect 11790 6100 11796 6112
rect 11655 6072 11796 6100
rect 11655 6069 11667 6072
rect 11609 6063 11667 6069
rect 11790 6060 11796 6072
rect 11848 6060 11854 6112
rect 12250 6060 12256 6112
rect 12308 6100 12314 6112
rect 12437 6103 12495 6109
rect 12437 6100 12449 6103
rect 12308 6072 12449 6100
rect 12308 6060 12314 6072
rect 12437 6069 12449 6072
rect 12483 6069 12495 6103
rect 12437 6063 12495 6069
rect 16301 6103 16359 6109
rect 16301 6069 16313 6103
rect 16347 6100 16359 6103
rect 16853 6103 16911 6109
rect 16853 6100 16865 6103
rect 16347 6072 16865 6100
rect 16347 6069 16359 6072
rect 16301 6063 16359 6069
rect 16853 6069 16865 6072
rect 16899 6069 16911 6103
rect 18598 6100 18604 6112
rect 18559 6072 18604 6100
rect 16853 6063 16911 6069
rect 18598 6060 18604 6072
rect 18656 6060 18662 6112
rect 18690 6060 18696 6112
rect 18748 6100 18754 6112
rect 19242 6100 19248 6112
rect 18748 6072 19248 6100
rect 18748 6060 18754 6072
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 20806 6060 20812 6112
rect 20864 6100 20870 6112
rect 20993 6103 21051 6109
rect 20993 6100 21005 6103
rect 20864 6072 21005 6100
rect 20864 6060 20870 6072
rect 20993 6069 21005 6072
rect 21039 6069 21051 6103
rect 20993 6063 21051 6069
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 7653 5899 7711 5905
rect 7653 5865 7665 5899
rect 7699 5896 7711 5899
rect 7742 5896 7748 5908
rect 7699 5868 7748 5896
rect 7699 5865 7711 5868
rect 7653 5859 7711 5865
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 9125 5899 9183 5905
rect 9125 5865 9137 5899
rect 9171 5896 9183 5899
rect 9490 5896 9496 5908
rect 9171 5868 9496 5896
rect 9171 5865 9183 5868
rect 9125 5859 9183 5865
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 9674 5896 9680 5908
rect 9635 5868 9680 5896
rect 9674 5856 9680 5868
rect 9732 5856 9738 5908
rect 10042 5896 10048 5908
rect 10003 5868 10048 5896
rect 10042 5856 10048 5868
rect 10100 5856 10106 5908
rect 12894 5856 12900 5908
rect 12952 5896 12958 5908
rect 13909 5899 13967 5905
rect 12952 5868 13032 5896
rect 12952 5856 12958 5868
rect 4062 5788 4068 5840
rect 4120 5828 4126 5840
rect 6518 5831 6576 5837
rect 6518 5828 6530 5831
rect 4120 5800 6530 5828
rect 4120 5788 4126 5800
rect 6518 5797 6530 5800
rect 6564 5797 6576 5831
rect 6518 5791 6576 5797
rect 7190 5788 7196 5840
rect 7248 5828 7254 5840
rect 12066 5828 12072 5840
rect 7248 5800 12072 5828
rect 7248 5788 7254 5800
rect 12066 5788 12072 5800
rect 12124 5788 12130 5840
rect 12250 5788 12256 5840
rect 12308 5828 12314 5840
rect 12802 5828 12808 5840
rect 12308 5800 12808 5828
rect 12308 5788 12314 5800
rect 12802 5788 12808 5800
rect 12860 5788 12866 5840
rect 13004 5837 13032 5868
rect 13909 5865 13921 5899
rect 13955 5896 13967 5899
rect 15102 5896 15108 5908
rect 13955 5868 15108 5896
rect 13955 5865 13967 5868
rect 13909 5859 13967 5865
rect 15102 5856 15108 5868
rect 15160 5856 15166 5908
rect 15562 5856 15568 5908
rect 15620 5896 15626 5908
rect 15657 5899 15715 5905
rect 15657 5896 15669 5899
rect 15620 5868 15669 5896
rect 15620 5856 15626 5868
rect 15657 5865 15669 5868
rect 15703 5865 15715 5899
rect 15657 5859 15715 5865
rect 15749 5899 15807 5905
rect 15749 5865 15761 5899
rect 15795 5896 15807 5899
rect 15838 5896 15844 5908
rect 15795 5868 15844 5896
rect 15795 5865 15807 5868
rect 15749 5859 15807 5865
rect 15838 5856 15844 5868
rect 15896 5856 15902 5908
rect 16761 5899 16819 5905
rect 16761 5865 16773 5899
rect 16807 5896 16819 5899
rect 16807 5868 16896 5896
rect 16807 5865 16819 5868
rect 16761 5859 16819 5865
rect 12989 5831 13047 5837
rect 12989 5797 13001 5831
rect 13035 5828 13047 5831
rect 14737 5831 14795 5837
rect 13035 5800 14412 5828
rect 13035 5797 13047 5800
rect 12989 5791 13047 5797
rect 6273 5763 6331 5769
rect 6273 5729 6285 5763
rect 6319 5760 6331 5763
rect 7466 5760 7472 5772
rect 6319 5732 7472 5760
rect 6319 5729 6331 5732
rect 6273 5723 6331 5729
rect 7466 5720 7472 5732
rect 7524 5720 7530 5772
rect 10962 5760 10968 5772
rect 10152 5732 10968 5760
rect 10152 5704 10180 5732
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 11140 5763 11198 5769
rect 11140 5729 11152 5763
rect 11186 5760 11198 5763
rect 12618 5760 12624 5772
rect 11186 5732 12624 5760
rect 11186 5729 11198 5732
rect 11140 5723 11198 5729
rect 12618 5720 12624 5732
rect 12676 5760 12682 5772
rect 12897 5763 12955 5769
rect 12676 5732 12839 5760
rect 12676 5720 12682 5732
rect 10134 5692 10140 5704
rect 10095 5664 10140 5692
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 10318 5692 10324 5704
rect 10279 5664 10324 5692
rect 10318 5652 10324 5664
rect 10376 5652 10382 5704
rect 10873 5695 10931 5701
rect 10873 5661 10885 5695
rect 10919 5661 10931 5695
rect 12811 5692 12839 5732
rect 12897 5729 12909 5763
rect 12943 5760 12955 5763
rect 13538 5760 13544 5772
rect 12943 5732 13544 5760
rect 12943 5729 12955 5732
rect 12897 5723 12955 5729
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 13078 5692 13084 5704
rect 12811 5664 13084 5692
rect 10873 5655 10931 5661
rect 10888 5556 10916 5655
rect 13078 5652 13084 5664
rect 13136 5652 13142 5704
rect 13998 5692 14004 5704
rect 13959 5664 14004 5692
rect 13998 5652 14004 5664
rect 14056 5652 14062 5704
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5661 14151 5695
rect 14093 5655 14151 5661
rect 13096 5624 13124 5652
rect 14108 5624 14136 5655
rect 13096 5596 14136 5624
rect 14384 5624 14412 5800
rect 14737 5797 14749 5831
rect 14783 5828 14795 5831
rect 16666 5828 16672 5840
rect 14783 5800 16672 5828
rect 14783 5797 14795 5800
rect 14737 5791 14795 5797
rect 16666 5788 16672 5800
rect 16724 5788 16730 5840
rect 16868 5828 16896 5868
rect 17862 5856 17868 5908
rect 17920 5896 17926 5908
rect 18509 5899 18567 5905
rect 18509 5896 18521 5899
rect 17920 5868 18521 5896
rect 17920 5856 17926 5868
rect 18509 5865 18521 5868
rect 18555 5865 18567 5899
rect 18509 5859 18567 5865
rect 19236 5831 19294 5837
rect 16868 5800 19196 5828
rect 15378 5720 15384 5772
rect 15436 5760 15442 5772
rect 15436 5732 16344 5760
rect 15436 5720 15442 5732
rect 15194 5652 15200 5704
rect 15252 5692 15258 5704
rect 15838 5692 15844 5704
rect 15252 5664 15844 5692
rect 15252 5652 15258 5664
rect 15838 5652 15844 5664
rect 15896 5652 15902 5704
rect 15933 5695 15991 5701
rect 15933 5661 15945 5695
rect 15979 5692 15991 5695
rect 16114 5692 16120 5704
rect 15979 5664 16120 5692
rect 15979 5661 15991 5664
rect 15933 5655 15991 5661
rect 16114 5652 16120 5664
rect 16172 5652 16178 5704
rect 16316 5692 16344 5732
rect 16390 5720 16396 5772
rect 16448 5760 16454 5772
rect 16485 5763 16543 5769
rect 16485 5760 16497 5763
rect 16448 5732 16497 5760
rect 16448 5720 16454 5732
rect 16485 5729 16497 5732
rect 16531 5729 16543 5763
rect 16485 5723 16543 5729
rect 16574 5720 16580 5772
rect 16632 5760 16638 5772
rect 17396 5763 17454 5769
rect 16632 5732 16677 5760
rect 16632 5720 16638 5732
rect 17396 5729 17408 5763
rect 17442 5760 17454 5763
rect 18874 5760 18880 5772
rect 17442 5732 18880 5760
rect 17442 5729 17454 5732
rect 17396 5723 17454 5729
rect 18874 5720 18880 5732
rect 18932 5720 18938 5772
rect 19058 5760 19064 5772
rect 18984 5732 19064 5760
rect 17034 5692 17040 5704
rect 16316 5664 17040 5692
rect 17034 5652 17040 5664
rect 17092 5652 17098 5704
rect 17129 5695 17187 5701
rect 17129 5661 17141 5695
rect 17175 5661 17187 5695
rect 18782 5692 18788 5704
rect 17129 5655 17187 5661
rect 18340 5664 18788 5692
rect 16850 5624 16856 5636
rect 14384 5596 16856 5624
rect 16850 5584 16856 5596
rect 16908 5584 16914 5636
rect 11054 5556 11060 5568
rect 10888 5528 11060 5556
rect 11054 5516 11060 5528
rect 11112 5556 11118 5568
rect 12066 5556 12072 5568
rect 11112 5528 12072 5556
rect 11112 5516 11118 5528
rect 12066 5516 12072 5528
rect 12124 5516 12130 5568
rect 12250 5556 12256 5568
rect 12211 5528 12256 5556
rect 12250 5516 12256 5528
rect 12308 5516 12314 5568
rect 12526 5556 12532 5568
rect 12487 5528 12532 5556
rect 12526 5516 12532 5528
rect 12584 5516 12590 5568
rect 13538 5556 13544 5568
rect 13499 5528 13544 5556
rect 13538 5516 13544 5528
rect 13596 5516 13602 5568
rect 15289 5559 15347 5565
rect 15289 5525 15301 5559
rect 15335 5556 15347 5559
rect 15654 5556 15660 5568
rect 15335 5528 15660 5556
rect 15335 5525 15347 5528
rect 15289 5519 15347 5525
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 15838 5516 15844 5568
rect 15896 5556 15902 5568
rect 16301 5559 16359 5565
rect 16301 5556 16313 5559
rect 15896 5528 16313 5556
rect 15896 5516 15902 5528
rect 16301 5525 16313 5528
rect 16347 5556 16359 5559
rect 17144 5556 17172 5655
rect 17862 5556 17868 5568
rect 16347 5528 17868 5556
rect 16347 5525 16359 5528
rect 16301 5519 16359 5525
rect 17862 5516 17868 5528
rect 17920 5556 17926 5568
rect 18340 5556 18368 5664
rect 18782 5652 18788 5664
rect 18840 5692 18846 5704
rect 18984 5701 19012 5732
rect 19058 5720 19064 5732
rect 19116 5720 19122 5772
rect 19168 5760 19196 5800
rect 19236 5797 19248 5831
rect 19282 5828 19294 5831
rect 19610 5828 19616 5840
rect 19282 5800 19616 5828
rect 19282 5797 19294 5800
rect 19236 5791 19294 5797
rect 19610 5788 19616 5800
rect 19668 5828 19674 5840
rect 20346 5828 20352 5840
rect 19668 5800 20352 5828
rect 19668 5788 19674 5800
rect 20346 5788 20352 5800
rect 20404 5788 20410 5840
rect 20530 5760 20536 5772
rect 19168 5732 20536 5760
rect 20530 5720 20536 5732
rect 20588 5720 20594 5772
rect 18969 5695 19027 5701
rect 18969 5692 18981 5695
rect 18840 5664 18981 5692
rect 18840 5652 18846 5664
rect 18969 5661 18981 5664
rect 19015 5661 19027 5695
rect 18969 5655 19027 5661
rect 18414 5584 18420 5636
rect 18472 5584 18478 5636
rect 17920 5528 18368 5556
rect 18432 5556 18460 5584
rect 19150 5556 19156 5568
rect 18432 5528 19156 5556
rect 17920 5516 17926 5528
rect 19150 5516 19156 5528
rect 19208 5516 19214 5568
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 20349 5559 20407 5565
rect 20349 5556 20361 5559
rect 19392 5528 20361 5556
rect 19392 5516 19398 5528
rect 20349 5525 20361 5528
rect 20395 5525 20407 5559
rect 20349 5519 20407 5525
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 11698 5312 11704 5364
rect 11756 5352 11762 5364
rect 16669 5355 16727 5361
rect 16669 5352 16681 5355
rect 11756 5324 16681 5352
rect 11756 5312 11762 5324
rect 16669 5321 16681 5324
rect 16715 5321 16727 5355
rect 16669 5315 16727 5321
rect 16758 5312 16764 5364
rect 16816 5352 16822 5364
rect 19426 5352 19432 5364
rect 16816 5324 19432 5352
rect 16816 5312 16822 5324
rect 19426 5312 19432 5324
rect 19484 5312 19490 5364
rect 19610 5352 19616 5364
rect 19571 5324 19616 5352
rect 19610 5312 19616 5324
rect 19668 5312 19674 5364
rect 9950 5244 9956 5296
rect 10008 5284 10014 5296
rect 12434 5284 12440 5296
rect 10008 5256 12440 5284
rect 10008 5244 10014 5256
rect 12434 5244 12440 5256
rect 12492 5244 12498 5296
rect 12986 5284 12992 5296
rect 12912 5256 12992 5284
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5216 12035 5219
rect 12250 5216 12256 5228
rect 12023 5188 12256 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 12250 5176 12256 5188
rect 12308 5176 12314 5228
rect 12912 5225 12940 5256
rect 12986 5244 12992 5256
rect 13044 5244 13050 5296
rect 12897 5219 12955 5225
rect 12897 5185 12909 5219
rect 12943 5185 12955 5219
rect 13078 5216 13084 5228
rect 13039 5188 13084 5216
rect 12897 5179 12955 5185
rect 13078 5176 13084 5188
rect 13136 5176 13142 5228
rect 13446 5216 13452 5228
rect 13407 5188 13452 5216
rect 13446 5176 13452 5188
rect 13504 5176 13510 5228
rect 16114 5176 16120 5228
rect 16172 5216 16178 5228
rect 17313 5219 17371 5225
rect 17313 5216 17325 5219
rect 16172 5188 17325 5216
rect 16172 5176 16178 5188
rect 17313 5185 17325 5188
rect 17359 5185 17371 5219
rect 17313 5179 17371 5185
rect 17862 5176 17868 5228
rect 17920 5216 17926 5228
rect 18233 5219 18291 5225
rect 18233 5216 18245 5219
rect 17920 5188 18245 5216
rect 17920 5176 17926 5188
rect 18233 5185 18245 5188
rect 18279 5185 18291 5219
rect 20438 5216 20444 5228
rect 20399 5188 20444 5216
rect 18233 5179 18291 5185
rect 20438 5176 20444 5188
rect 20496 5176 20502 5228
rect 20898 5216 20904 5228
rect 20859 5188 20904 5216
rect 20898 5176 20904 5188
rect 20956 5176 20962 5228
rect 11793 5151 11851 5157
rect 11793 5117 11805 5151
rect 11839 5148 11851 5151
rect 12526 5148 12532 5160
rect 11839 5120 12532 5148
rect 11839 5117 11851 5120
rect 11793 5111 11851 5117
rect 12526 5108 12532 5120
rect 12584 5108 12590 5160
rect 12805 5151 12863 5157
rect 12805 5117 12817 5151
rect 12851 5148 12863 5151
rect 12986 5148 12992 5160
rect 12851 5120 12992 5148
rect 12851 5117 12863 5120
rect 12805 5111 12863 5117
rect 12986 5108 12992 5120
rect 13044 5148 13050 5160
rect 13262 5148 13268 5160
rect 13044 5120 13268 5148
rect 13044 5108 13050 5120
rect 13262 5108 13268 5120
rect 13320 5108 13326 5160
rect 13464 5148 13492 5176
rect 15105 5151 15163 5157
rect 15105 5148 15117 5151
rect 13464 5120 15117 5148
rect 15105 5117 15117 5120
rect 15151 5148 15163 5151
rect 15194 5148 15200 5160
rect 15151 5120 15200 5148
rect 15151 5117 15163 5120
rect 15105 5111 15163 5117
rect 15194 5108 15200 5120
rect 15252 5108 15258 5160
rect 15372 5151 15430 5157
rect 15372 5117 15384 5151
rect 15418 5148 15430 5151
rect 16132 5148 16160 5176
rect 15418 5120 16160 5148
rect 17129 5151 17187 5157
rect 15418 5117 15430 5120
rect 15372 5111 15430 5117
rect 17129 5117 17141 5151
rect 17175 5148 17187 5151
rect 17586 5148 17592 5160
rect 17175 5120 17592 5148
rect 17175 5117 17187 5120
rect 17129 5111 17187 5117
rect 11701 5083 11759 5089
rect 11701 5049 11713 5083
rect 11747 5080 11759 5083
rect 13538 5080 13544 5092
rect 11747 5052 13544 5080
rect 11747 5049 11759 5052
rect 11701 5043 11759 5049
rect 13538 5040 13544 5052
rect 13596 5040 13602 5092
rect 13722 5089 13728 5092
rect 13716 5080 13728 5089
rect 13683 5052 13728 5080
rect 13716 5043 13728 5052
rect 13722 5040 13728 5043
rect 13780 5040 13786 5092
rect 11330 5012 11336 5024
rect 11291 4984 11336 5012
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 14829 5015 14887 5021
rect 12492 4984 12537 5012
rect 12492 4972 12498 4984
rect 14829 4981 14841 5015
rect 14875 5012 14887 5015
rect 15387 5012 15415 5111
rect 17586 5108 17592 5120
rect 17644 5108 17650 5160
rect 20254 5148 20260 5160
rect 20215 5120 20260 5148
rect 20254 5108 20260 5120
rect 20312 5108 20318 5160
rect 16669 5083 16727 5089
rect 16669 5049 16681 5083
rect 16715 5080 16727 5083
rect 18500 5083 18558 5089
rect 16715 5052 17264 5080
rect 16715 5049 16727 5052
rect 16669 5043 16727 5049
rect 16482 5012 16488 5024
rect 14875 4984 15415 5012
rect 16443 4984 16488 5012
rect 14875 4981 14887 4984
rect 14829 4975 14887 4981
rect 16482 4972 16488 4984
rect 16540 4972 16546 5024
rect 16574 4972 16580 5024
rect 16632 5012 16638 5024
rect 17236 5021 17264 5052
rect 18500 5049 18512 5083
rect 18546 5080 18558 5083
rect 18690 5080 18696 5092
rect 18546 5052 18696 5080
rect 18546 5049 18558 5052
rect 18500 5043 18558 5049
rect 18690 5040 18696 5052
rect 18748 5040 18754 5092
rect 19058 5040 19064 5092
rect 19116 5080 19122 5092
rect 20349 5083 20407 5089
rect 20349 5080 20361 5083
rect 19116 5052 20361 5080
rect 19116 5040 19122 5052
rect 20349 5049 20361 5052
rect 20395 5049 20407 5083
rect 20349 5043 20407 5049
rect 16761 5015 16819 5021
rect 16761 5012 16773 5015
rect 16632 4984 16773 5012
rect 16632 4972 16638 4984
rect 16761 4981 16773 4984
rect 16807 4981 16819 5015
rect 16761 4975 16819 4981
rect 17221 5015 17279 5021
rect 17221 4981 17233 5015
rect 17267 5012 17279 5015
rect 18782 5012 18788 5024
rect 17267 4984 18788 5012
rect 17267 4981 17279 4984
rect 17221 4975 17279 4981
rect 18782 4972 18788 4984
rect 18840 4972 18846 5024
rect 19886 5012 19892 5024
rect 19847 4984 19892 5012
rect 19886 4972 19892 4984
rect 19944 4972 19950 5024
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 11330 4768 11336 4820
rect 11388 4808 11394 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 11388 4780 14105 4808
rect 11388 4768 11394 4780
rect 14093 4777 14105 4780
rect 14139 4777 14151 4811
rect 14093 4771 14151 4777
rect 14182 4768 14188 4820
rect 14240 4808 14246 4820
rect 18046 4808 18052 4820
rect 14240 4780 18052 4808
rect 14240 4768 14246 4780
rect 18046 4768 18052 4780
rect 18104 4768 18110 4820
rect 18690 4808 18696 4820
rect 18603 4780 18696 4808
rect 18690 4768 18696 4780
rect 18748 4808 18754 4820
rect 20438 4808 20444 4820
rect 18748 4780 20444 4808
rect 18748 4768 18754 4780
rect 20438 4768 20444 4780
rect 20496 4768 20502 4820
rect 290 4700 296 4752
rect 348 4740 354 4752
rect 12986 4740 12992 4752
rect 348 4712 12992 4740
rect 348 4700 354 4712
rect 12986 4700 12992 4712
rect 13044 4700 13050 4752
rect 13170 4700 13176 4752
rect 13228 4740 13234 4752
rect 15924 4743 15982 4749
rect 13228 4712 14320 4740
rect 13228 4700 13234 4712
rect 11977 4675 12035 4681
rect 11977 4641 11989 4675
rect 12023 4672 12035 4675
rect 12066 4672 12072 4684
rect 12023 4644 12072 4672
rect 12023 4641 12035 4644
rect 11977 4635 12035 4641
rect 12066 4632 12072 4644
rect 12124 4632 12130 4684
rect 12250 4681 12256 4684
rect 12244 4672 12256 4681
rect 12211 4644 12256 4672
rect 12244 4635 12256 4644
rect 12250 4632 12256 4635
rect 12308 4632 12314 4684
rect 13998 4672 14004 4684
rect 13959 4644 14004 4672
rect 13998 4632 14004 4644
rect 14056 4632 14062 4684
rect 13722 4604 13728 4616
rect 13372 4576 13728 4604
rect 9674 4496 9680 4548
rect 9732 4536 9738 4548
rect 11974 4536 11980 4548
rect 9732 4508 11980 4536
rect 9732 4496 9738 4508
rect 11974 4496 11980 4508
rect 12032 4496 12038 4548
rect 13372 4545 13400 4576
rect 13722 4564 13728 4576
rect 13780 4604 13786 4616
rect 14185 4607 14243 4613
rect 14185 4604 14197 4607
rect 13780 4576 14197 4604
rect 13780 4564 13786 4576
rect 14185 4573 14197 4576
rect 14231 4573 14243 4607
rect 14185 4567 14243 4573
rect 13357 4539 13415 4545
rect 13357 4505 13369 4539
rect 13403 4505 13415 4539
rect 14292 4536 14320 4712
rect 15924 4709 15936 4743
rect 15970 4740 15982 4743
rect 16482 4740 16488 4752
rect 15970 4712 16488 4740
rect 15970 4709 15982 4712
rect 15924 4703 15982 4709
rect 16482 4700 16488 4712
rect 16540 4700 16546 4752
rect 17034 4700 17040 4752
rect 17092 4740 17098 4752
rect 17558 4743 17616 4749
rect 17558 4740 17570 4743
rect 17092 4712 17570 4740
rect 17092 4700 17098 4712
rect 17558 4709 17570 4712
rect 17604 4709 17616 4743
rect 17558 4703 17616 4709
rect 19150 4700 19156 4752
rect 19208 4740 19214 4752
rect 20165 4743 20223 4749
rect 20165 4740 20177 4743
rect 19208 4712 20177 4740
rect 19208 4700 19214 4712
rect 20165 4709 20177 4712
rect 20211 4709 20223 4743
rect 20165 4703 20223 4709
rect 14550 4632 14556 4684
rect 14608 4672 14614 4684
rect 14645 4675 14703 4681
rect 14645 4672 14657 4675
rect 14608 4644 14657 4672
rect 14608 4632 14614 4644
rect 14645 4641 14657 4644
rect 14691 4641 14703 4675
rect 14645 4635 14703 4641
rect 15194 4632 15200 4684
rect 15252 4672 15258 4684
rect 15657 4675 15715 4681
rect 15657 4672 15669 4675
rect 15252 4644 15669 4672
rect 15252 4632 15258 4644
rect 15657 4641 15669 4644
rect 15703 4672 15715 4675
rect 16758 4672 16764 4684
rect 15703 4644 16764 4672
rect 15703 4641 15715 4644
rect 15657 4635 15715 4641
rect 16758 4632 16764 4644
rect 16816 4672 16822 4684
rect 17313 4675 17371 4681
rect 17313 4672 17325 4675
rect 16816 4644 17325 4672
rect 16816 4632 16822 4644
rect 17313 4641 17325 4644
rect 17359 4641 17371 4675
rect 17313 4635 17371 4641
rect 17402 4632 17408 4684
rect 17460 4672 17466 4684
rect 18969 4675 19027 4681
rect 18969 4672 18981 4675
rect 17460 4644 18981 4672
rect 17460 4632 17466 4644
rect 18969 4641 18981 4644
rect 19015 4641 19027 4675
rect 18969 4635 19027 4641
rect 18598 4564 18604 4616
rect 18656 4604 18662 4616
rect 20257 4607 20315 4613
rect 20257 4604 20269 4607
rect 18656 4576 20269 4604
rect 18656 4564 18662 4576
rect 20257 4573 20269 4576
rect 20303 4573 20315 4607
rect 20438 4604 20444 4616
rect 20399 4576 20444 4604
rect 20257 4567 20315 4573
rect 17034 4536 17040 4548
rect 14292 4508 15332 4536
rect 16995 4508 17040 4536
rect 13357 4499 13415 4505
rect 7650 4428 7656 4480
rect 7708 4468 7714 4480
rect 13262 4468 13268 4480
rect 7708 4440 13268 4468
rect 7708 4428 7714 4440
rect 13262 4428 13268 4440
rect 13320 4428 13326 4480
rect 13446 4428 13452 4480
rect 13504 4468 13510 4480
rect 13633 4471 13691 4477
rect 13633 4468 13645 4471
rect 13504 4440 13645 4468
rect 13504 4428 13510 4440
rect 13633 4437 13645 4440
rect 13679 4437 13691 4471
rect 13633 4431 13691 4437
rect 14829 4471 14887 4477
rect 14829 4437 14841 4471
rect 14875 4468 14887 4471
rect 15194 4468 15200 4480
rect 14875 4440 15200 4468
rect 14875 4437 14887 4440
rect 14829 4431 14887 4437
rect 15194 4428 15200 4440
rect 15252 4428 15258 4480
rect 15304 4468 15332 4508
rect 17034 4496 17040 4508
rect 17092 4496 17098 4548
rect 18322 4496 18328 4548
rect 18380 4496 18386 4548
rect 19153 4539 19211 4545
rect 19153 4505 19165 4539
rect 19199 4536 19211 4539
rect 19702 4536 19708 4548
rect 19199 4508 19708 4536
rect 19199 4505 19211 4508
rect 19153 4499 19211 4505
rect 19702 4496 19708 4508
rect 19760 4496 19766 4548
rect 20272 4536 20300 4567
rect 20438 4564 20444 4576
rect 20496 4564 20502 4616
rect 20898 4604 20904 4616
rect 20859 4576 20904 4604
rect 20898 4564 20904 4576
rect 20956 4564 20962 4616
rect 20346 4536 20352 4548
rect 20272 4508 20352 4536
rect 20346 4496 20352 4508
rect 20404 4496 20410 4548
rect 18340 4468 18368 4496
rect 19794 4468 19800 4480
rect 15304 4440 18368 4468
rect 19755 4440 19800 4468
rect 19794 4428 19800 4440
rect 19852 4428 19858 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 13262 4224 13268 4276
rect 13320 4264 13326 4276
rect 19058 4264 19064 4276
rect 13320 4236 19064 4264
rect 13320 4224 13326 4236
rect 12250 4156 12256 4208
rect 12308 4196 12314 4208
rect 16482 4196 16488 4208
rect 12308 4168 13032 4196
rect 12308 4156 12314 4168
rect 5810 4088 5816 4140
rect 5868 4128 5874 4140
rect 8938 4128 8944 4140
rect 5868 4100 8944 4128
rect 5868 4088 5874 4100
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 12434 4088 12440 4140
rect 12492 4128 12498 4140
rect 13004 4137 13032 4168
rect 15856 4168 16488 4196
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12492 4100 12909 4128
rect 12492 4088 12498 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 12897 4091 12955 4097
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4097 13047 4131
rect 13998 4128 14004 4140
rect 12989 4091 13047 4097
rect 13188 4100 14004 4128
rect 9033 4063 9091 4069
rect 9033 4029 9045 4063
rect 9079 4060 9091 4063
rect 9122 4060 9128 4072
rect 9079 4032 9128 4060
rect 9079 4029 9091 4032
rect 9033 4023 9091 4029
rect 9122 4020 9128 4032
rect 9180 4020 9186 4072
rect 11606 4060 11612 4072
rect 11567 4032 11612 4060
rect 11606 4020 11612 4032
rect 11664 4020 11670 4072
rect 12618 4060 12624 4072
rect 11716 4032 12624 4060
rect 9214 3952 9220 4004
rect 9272 4001 9278 4004
rect 9272 3995 9336 4001
rect 9272 3961 9290 3995
rect 9324 3961 9336 3995
rect 11716 3992 11744 4032
rect 12618 4020 12624 4032
rect 12676 4020 12682 4072
rect 12802 4060 12808 4072
rect 12763 4032 12808 4060
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 9272 3955 9336 3961
rect 9416 3964 11744 3992
rect 11885 3995 11943 4001
rect 9272 3952 9278 3955
rect 3602 3884 3608 3936
rect 3660 3924 3666 3936
rect 9416 3924 9444 3964
rect 11885 3961 11897 3995
rect 11931 3992 11943 3995
rect 13078 3992 13084 4004
rect 11931 3964 13084 3992
rect 11931 3961 11943 3964
rect 11885 3955 11943 3961
rect 13078 3952 13084 3964
rect 13136 3952 13142 4004
rect 3660 3896 9444 3924
rect 3660 3884 3666 3896
rect 10318 3884 10324 3936
rect 10376 3924 10382 3936
rect 10413 3927 10471 3933
rect 10413 3924 10425 3927
rect 10376 3896 10425 3924
rect 10376 3884 10382 3896
rect 10413 3893 10425 3896
rect 10459 3893 10471 3927
rect 10413 3887 10471 3893
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3924 12495 3927
rect 13188 3924 13216 4100
rect 13998 4088 14004 4100
rect 14056 4088 14062 4140
rect 15470 4128 15476 4140
rect 14200 4100 15476 4128
rect 13446 4060 13452 4072
rect 13407 4032 13452 4060
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 14200 4069 14228 4100
rect 15470 4088 15476 4100
rect 15528 4088 15534 4140
rect 15654 4128 15660 4140
rect 15615 4100 15660 4128
rect 15654 4088 15660 4100
rect 15712 4088 15718 4140
rect 15856 4137 15884 4168
rect 16482 4156 16488 4168
rect 16540 4196 16546 4208
rect 16540 4168 16804 4196
rect 16540 4156 16546 4168
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4097 15899 4131
rect 15841 4091 15899 4097
rect 16390 4088 16396 4140
rect 16448 4128 16454 4140
rect 16776 4137 16804 4168
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 16448 4100 16681 4128
rect 16448 4088 16454 4100
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 16761 4131 16819 4137
rect 16761 4097 16773 4131
rect 16807 4097 16819 4131
rect 16761 4091 16819 4097
rect 14185 4063 14243 4069
rect 14185 4029 14197 4063
rect 14231 4029 14243 4063
rect 14185 4023 14243 4029
rect 14366 4020 14372 4072
rect 14424 4060 14430 4072
rect 14737 4063 14795 4069
rect 14737 4060 14749 4063
rect 14424 4032 14749 4060
rect 14424 4020 14430 4032
rect 14737 4029 14749 4032
rect 14783 4029 14795 4063
rect 14737 4023 14795 4029
rect 15565 4063 15623 4069
rect 15565 4029 15577 4063
rect 15611 4060 15623 4063
rect 16574 4060 16580 4072
rect 15611 4032 16580 4060
rect 15611 4029 15623 4032
rect 15565 4023 15623 4029
rect 16574 4020 16580 4032
rect 16632 4020 16638 4072
rect 16850 4020 16856 4072
rect 16908 4060 16914 4072
rect 18064 4069 18092 4236
rect 19058 4224 19064 4236
rect 19116 4224 19122 4276
rect 19334 4196 19340 4208
rect 19260 4168 19340 4196
rect 19260 4137 19288 4168
rect 19334 4156 19340 4168
rect 19392 4156 19398 4208
rect 19610 4156 19616 4208
rect 19668 4196 19674 4208
rect 19668 4168 20208 4196
rect 19668 4156 19674 4168
rect 19245 4131 19303 4137
rect 19245 4097 19257 4131
rect 19291 4097 19303 4131
rect 19245 4091 19303 4097
rect 19886 4088 19892 4140
rect 19944 4128 19950 4140
rect 20180 4137 20208 4168
rect 20073 4131 20131 4137
rect 20073 4128 20085 4131
rect 19944 4100 20085 4128
rect 19944 4088 19950 4100
rect 20073 4097 20085 4100
rect 20119 4097 20131 4131
rect 20073 4091 20131 4097
rect 20165 4131 20223 4137
rect 20165 4097 20177 4131
rect 20211 4097 20223 4131
rect 20165 4091 20223 4097
rect 20530 4088 20536 4140
rect 20588 4128 20594 4140
rect 22462 4128 22468 4140
rect 20588 4100 22468 4128
rect 20588 4088 20594 4100
rect 22462 4088 22468 4100
rect 22520 4088 22526 4140
rect 17221 4063 17279 4069
rect 17221 4060 17233 4063
rect 16908 4032 17233 4060
rect 16908 4020 16914 4032
rect 17221 4029 17233 4032
rect 17267 4029 17279 4063
rect 17221 4023 17279 4029
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4029 18107 4063
rect 18966 4060 18972 4072
rect 18927 4032 18972 4060
rect 18049 4023 18107 4029
rect 18966 4020 18972 4032
rect 19024 4020 19030 4072
rect 19794 4020 19800 4072
rect 19852 4060 19858 4072
rect 19981 4063 20039 4069
rect 19981 4060 19993 4063
rect 19852 4032 19993 4060
rect 19852 4020 19858 4032
rect 19981 4029 19993 4032
rect 20027 4029 20039 4063
rect 19981 4023 20039 4029
rect 20254 4020 20260 4072
rect 20312 4060 20318 4072
rect 20625 4063 20683 4069
rect 20625 4060 20637 4063
rect 20312 4032 20637 4060
rect 20312 4020 20318 4032
rect 20625 4029 20637 4032
rect 20671 4029 20683 4063
rect 20625 4023 20683 4029
rect 13262 3952 13268 4004
rect 13320 3992 13326 4004
rect 13725 3995 13783 4001
rect 13725 3992 13737 3995
rect 13320 3964 13737 3992
rect 13320 3952 13326 3964
rect 13725 3961 13737 3964
rect 13771 3961 13783 3995
rect 13725 3955 13783 3961
rect 15838 3952 15844 4004
rect 15896 3992 15902 4004
rect 15896 3964 17448 3992
rect 15896 3952 15902 3964
rect 12483 3896 13216 3924
rect 12483 3893 12495 3896
rect 12437 3887 12495 3893
rect 13906 3884 13912 3936
rect 13964 3924 13970 3936
rect 14369 3927 14427 3933
rect 14369 3924 14381 3927
rect 13964 3896 14381 3924
rect 13964 3884 13970 3896
rect 14369 3893 14381 3896
rect 14415 3893 14427 3927
rect 14369 3887 14427 3893
rect 15197 3927 15255 3933
rect 15197 3893 15209 3927
rect 15243 3924 15255 3927
rect 15286 3924 15292 3936
rect 15243 3896 15292 3924
rect 15243 3893 15255 3896
rect 15197 3887 15255 3893
rect 15286 3884 15292 3896
rect 15344 3884 15350 3936
rect 16022 3884 16028 3936
rect 16080 3924 16086 3936
rect 16209 3927 16267 3933
rect 16209 3924 16221 3927
rect 16080 3896 16221 3924
rect 16080 3884 16086 3896
rect 16209 3893 16221 3896
rect 16255 3893 16267 3927
rect 16574 3924 16580 3936
rect 16535 3896 16580 3924
rect 16209 3887 16267 3893
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 17420 3933 17448 3964
rect 17405 3927 17463 3933
rect 17405 3893 17417 3927
rect 17451 3893 17463 3927
rect 17405 3887 17463 3893
rect 17678 3884 17684 3936
rect 17736 3924 17742 3936
rect 18233 3927 18291 3933
rect 18233 3924 18245 3927
rect 17736 3896 18245 3924
rect 17736 3884 17742 3896
rect 18233 3893 18245 3896
rect 18279 3893 18291 3927
rect 18233 3887 18291 3893
rect 18601 3927 18659 3933
rect 18601 3893 18613 3927
rect 18647 3924 18659 3927
rect 18782 3924 18788 3936
rect 18647 3896 18788 3924
rect 18647 3893 18659 3896
rect 18601 3887 18659 3893
rect 18782 3884 18788 3896
rect 18840 3884 18846 3936
rect 19061 3927 19119 3933
rect 19061 3893 19073 3927
rect 19107 3924 19119 3927
rect 19613 3927 19671 3933
rect 19613 3924 19625 3927
rect 19107 3896 19625 3924
rect 19107 3893 19119 3896
rect 19061 3887 19119 3893
rect 19613 3893 19625 3896
rect 19659 3893 19671 3927
rect 19613 3887 19671 3893
rect 20254 3884 20260 3936
rect 20312 3924 20318 3936
rect 20809 3927 20867 3933
rect 20809 3924 20821 3927
rect 20312 3896 20821 3924
rect 20312 3884 20318 3896
rect 20809 3893 20821 3896
rect 20855 3893 20867 3927
rect 20809 3887 20867 3893
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 1394 3680 1400 3732
rect 1452 3720 1458 3732
rect 15841 3723 15899 3729
rect 15841 3720 15853 3723
rect 1452 3692 15853 3720
rect 1452 3680 1458 3692
rect 15841 3689 15853 3692
rect 15887 3689 15899 3723
rect 15841 3683 15899 3689
rect 15933 3723 15991 3729
rect 15933 3689 15945 3723
rect 15979 3720 15991 3723
rect 16942 3720 16948 3732
rect 15979 3692 16948 3720
rect 15979 3689 15991 3692
rect 15933 3683 15991 3689
rect 16942 3680 16948 3692
rect 17000 3720 17006 3732
rect 17862 3720 17868 3732
rect 17000 3692 17868 3720
rect 17000 3680 17006 3692
rect 17862 3680 17868 3692
rect 17920 3680 17926 3732
rect 18141 3723 18199 3729
rect 18141 3689 18153 3723
rect 18187 3689 18199 3723
rect 18141 3683 18199 3689
rect 7466 3612 7472 3664
rect 7524 3652 7530 3664
rect 10042 3652 10048 3664
rect 7524 3624 10048 3652
rect 7524 3612 7530 3624
rect 10042 3612 10048 3624
rect 10100 3612 10106 3664
rect 10226 3612 10232 3664
rect 10284 3652 10290 3664
rect 10413 3655 10471 3661
rect 10413 3652 10425 3655
rect 10284 3624 10425 3652
rect 10284 3612 10290 3624
rect 10413 3621 10425 3624
rect 10459 3621 10471 3655
rect 10413 3615 10471 3621
rect 10778 3612 10784 3664
rect 10836 3652 10842 3664
rect 13262 3652 13268 3664
rect 10836 3624 13268 3652
rect 10836 3612 10842 3624
rect 13262 3612 13268 3624
rect 13320 3612 13326 3664
rect 13817 3655 13875 3661
rect 13817 3652 13829 3655
rect 13731 3624 13829 3652
rect 9122 3544 9128 3596
rect 9180 3584 9186 3596
rect 10597 3587 10655 3593
rect 9180 3556 10272 3584
rect 9180 3544 9186 3556
rect 10244 3528 10272 3556
rect 10597 3553 10609 3587
rect 10643 3584 10655 3587
rect 11146 3584 11152 3596
rect 10643 3556 11152 3584
rect 10643 3553 10655 3556
rect 10597 3547 10655 3553
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 11324 3587 11382 3593
rect 11324 3553 11336 3587
rect 11370 3584 11382 3587
rect 11882 3584 11888 3596
rect 11370 3556 11888 3584
rect 11370 3553 11382 3556
rect 11324 3547 11382 3553
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 12713 3587 12771 3593
rect 12713 3553 12725 3587
rect 12759 3584 12771 3587
rect 13446 3584 13452 3596
rect 12759 3556 13452 3584
rect 12759 3553 12771 3556
rect 12713 3547 12771 3553
rect 13446 3544 13452 3556
rect 13504 3544 13510 3596
rect 1946 3476 1952 3528
rect 2004 3516 2010 3528
rect 10134 3516 10140 3528
rect 2004 3488 10140 3516
rect 2004 3476 2010 3488
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 10226 3476 10232 3528
rect 10284 3516 10290 3528
rect 10870 3516 10876 3528
rect 10284 3488 10876 3516
rect 10284 3476 10290 3488
rect 10870 3476 10876 3488
rect 10928 3516 10934 3528
rect 11057 3519 11115 3525
rect 11057 3516 11069 3519
rect 10928 3488 11069 3516
rect 10928 3476 10934 3488
rect 11057 3485 11069 3488
rect 11103 3485 11115 3519
rect 11057 3479 11115 3485
rect 12434 3476 12440 3528
rect 12492 3516 12498 3528
rect 12897 3519 12955 3525
rect 12897 3516 12909 3519
rect 12492 3488 12909 3516
rect 12492 3476 12498 3488
rect 12897 3485 12909 3488
rect 12943 3485 12955 3519
rect 12897 3479 12955 3485
rect 13078 3476 13084 3528
rect 13136 3516 13142 3528
rect 13630 3516 13636 3528
rect 13136 3488 13636 3516
rect 13136 3476 13142 3488
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 6362 3408 6368 3460
rect 6420 3448 6426 3460
rect 10413 3451 10471 3457
rect 10413 3448 10425 3451
rect 6420 3420 10425 3448
rect 6420 3408 6426 3420
rect 10413 3417 10425 3420
rect 10459 3417 10471 3451
rect 13731 3448 13759 3624
rect 13817 3621 13829 3624
rect 13863 3621 13875 3655
rect 13817 3615 13875 3621
rect 13909 3655 13967 3661
rect 13909 3621 13921 3655
rect 13955 3652 13967 3655
rect 16114 3652 16120 3664
rect 13955 3624 16120 3652
rect 13955 3621 13967 3624
rect 13909 3615 13967 3621
rect 16114 3612 16120 3624
rect 16172 3612 16178 3664
rect 18156 3652 18184 3683
rect 18874 3680 18880 3732
rect 18932 3720 18938 3732
rect 19150 3720 19156 3732
rect 18932 3692 19156 3720
rect 18932 3680 18938 3692
rect 19150 3680 19156 3692
rect 19208 3720 19214 3732
rect 19797 3723 19855 3729
rect 19797 3720 19809 3723
rect 19208 3692 19809 3720
rect 19208 3680 19214 3692
rect 19797 3689 19809 3692
rect 19843 3689 19855 3723
rect 19797 3683 19855 3689
rect 20622 3680 20628 3732
rect 20680 3720 20686 3732
rect 21358 3720 21364 3732
rect 20680 3692 21364 3720
rect 20680 3680 20686 3692
rect 21358 3680 21364 3692
rect 21416 3680 21422 3732
rect 18598 3652 18604 3664
rect 16776 3624 17724 3652
rect 18156 3624 18604 3652
rect 16776 3596 16804 3624
rect 14461 3587 14519 3593
rect 14461 3553 14473 3587
rect 14507 3553 14519 3587
rect 16758 3584 16764 3596
rect 16719 3556 16764 3584
rect 14461 3547 14519 3553
rect 13998 3516 14004 3528
rect 13959 3488 14004 3516
rect 13998 3476 14004 3488
rect 14056 3476 14062 3528
rect 10413 3411 10471 3417
rect 11992 3420 13759 3448
rect 2498 3340 2504 3392
rect 2556 3380 2562 3392
rect 11992 3380 12020 3420
rect 13814 3408 13820 3460
rect 13872 3448 13878 3460
rect 14476 3448 14504 3547
rect 16758 3544 16764 3556
rect 16816 3544 16822 3596
rect 17028 3587 17086 3593
rect 17028 3553 17040 3587
rect 17074 3584 17086 3587
rect 17586 3584 17592 3596
rect 17074 3556 17592 3584
rect 17074 3553 17086 3556
rect 17028 3547 17086 3553
rect 17586 3544 17592 3556
rect 17644 3544 17650 3596
rect 17696 3584 17724 3624
rect 18598 3612 18604 3624
rect 18656 3661 18662 3664
rect 18656 3655 18720 3661
rect 18656 3621 18674 3655
rect 18708 3621 18720 3655
rect 18656 3615 18720 3621
rect 18656 3612 18662 3615
rect 18966 3612 18972 3664
rect 19024 3652 19030 3664
rect 20901 3655 20959 3661
rect 20901 3652 20913 3655
rect 19024 3624 20913 3652
rect 19024 3612 19030 3624
rect 20901 3621 20913 3624
rect 20947 3621 20959 3655
rect 20901 3615 20959 3621
rect 18417 3587 18475 3593
rect 18417 3584 18429 3587
rect 17696 3556 18429 3584
rect 18417 3553 18429 3556
rect 18463 3553 18475 3587
rect 18417 3547 18475 3553
rect 19978 3544 19984 3596
rect 20036 3584 20042 3596
rect 20073 3587 20131 3593
rect 20073 3584 20085 3587
rect 20036 3556 20085 3584
rect 20036 3544 20042 3556
rect 20073 3553 20085 3556
rect 20119 3553 20131 3587
rect 20073 3547 20131 3553
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 16080 3488 16125 3516
rect 16080 3476 16086 3488
rect 20257 3451 20315 3457
rect 20257 3448 20269 3451
rect 13872 3420 14504 3448
rect 19343 3420 20269 3448
rect 13872 3408 13878 3420
rect 2556 3352 12020 3380
rect 12437 3383 12495 3389
rect 2556 3340 2562 3352
rect 12437 3349 12449 3383
rect 12483 3380 12495 3383
rect 12894 3380 12900 3392
rect 12483 3352 12900 3380
rect 12483 3349 12495 3352
rect 12437 3343 12495 3349
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 13449 3383 13507 3389
rect 13449 3349 13461 3383
rect 13495 3380 13507 3383
rect 14458 3380 14464 3392
rect 13495 3352 14464 3380
rect 13495 3349 13507 3352
rect 13449 3343 13507 3349
rect 14458 3340 14464 3352
rect 14516 3340 14522 3392
rect 14642 3380 14648 3392
rect 14603 3352 14648 3380
rect 14642 3340 14648 3352
rect 14700 3340 14706 3392
rect 15473 3383 15531 3389
rect 15473 3349 15485 3383
rect 15519 3380 15531 3383
rect 16942 3380 16948 3392
rect 15519 3352 16948 3380
rect 15519 3349 15531 3352
rect 15473 3343 15531 3349
rect 16942 3340 16948 3352
rect 17000 3340 17006 3392
rect 19058 3340 19064 3392
rect 19116 3380 19122 3392
rect 19343 3380 19371 3420
rect 20257 3417 20269 3420
rect 20303 3417 20315 3451
rect 20257 3411 20315 3417
rect 19116 3352 19371 3380
rect 19116 3340 19122 3352
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 842 3136 848 3188
rect 900 3176 906 3188
rect 12897 3179 12955 3185
rect 12897 3176 12909 3179
rect 900 3148 12909 3176
rect 900 3136 906 3148
rect 12897 3145 12909 3148
rect 12943 3145 12955 3179
rect 12897 3139 12955 3145
rect 13262 3136 13268 3188
rect 13320 3176 13326 3188
rect 14642 3176 14648 3188
rect 13320 3148 14648 3176
rect 13320 3136 13326 3148
rect 14642 3136 14648 3148
rect 14700 3136 14706 3188
rect 16022 3176 16028 3188
rect 15983 3148 16028 3176
rect 16022 3136 16028 3148
rect 16080 3136 16086 3188
rect 17586 3136 17592 3188
rect 17644 3176 17650 3188
rect 17681 3179 17739 3185
rect 17681 3176 17693 3179
rect 17644 3148 17693 3176
rect 17644 3136 17650 3148
rect 17681 3145 17693 3148
rect 17727 3145 17739 3179
rect 17681 3139 17739 3145
rect 8202 3068 8208 3120
rect 8260 3108 8266 3120
rect 9766 3108 9772 3120
rect 8260 3080 9772 3108
rect 8260 3068 8266 3080
rect 9766 3068 9772 3080
rect 9824 3068 9830 3120
rect 11974 3068 11980 3120
rect 12032 3108 12038 3120
rect 12621 3111 12679 3117
rect 12621 3108 12633 3111
rect 12032 3080 12633 3108
rect 12032 3068 12038 3080
rect 12621 3077 12633 3080
rect 12667 3077 12679 3111
rect 12621 3071 12679 3077
rect 14369 3111 14427 3117
rect 14369 3077 14381 3111
rect 14415 3077 14427 3111
rect 14369 3071 14427 3077
rect 10042 3040 10048 3052
rect 10003 3012 10048 3040
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 12066 3040 12072 3052
rect 11164 3012 12072 3040
rect 4154 2932 4160 2984
rect 4212 2972 4218 2984
rect 9674 2972 9680 2984
rect 4212 2944 9680 2972
rect 4212 2932 4218 2944
rect 9674 2932 9680 2944
rect 9732 2932 9738 2984
rect 10318 2981 10324 2984
rect 10312 2972 10324 2981
rect 10279 2944 10324 2972
rect 10312 2935 10324 2944
rect 10318 2932 10324 2935
rect 10376 2932 10382 2984
rect 10870 2932 10876 2984
rect 10928 2972 10934 2984
rect 11164 2972 11192 3012
rect 12066 3000 12072 3012
rect 12124 3040 12130 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12124 3012 13001 3040
rect 12124 3000 12130 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 10928 2944 11192 2972
rect 11793 2975 11851 2981
rect 10928 2932 10934 2944
rect 11793 2941 11805 2975
rect 11839 2941 11851 2975
rect 11793 2935 11851 2941
rect 8570 2864 8576 2916
rect 8628 2904 8634 2916
rect 9950 2904 9956 2916
rect 8628 2876 9956 2904
rect 8628 2864 8634 2876
rect 9950 2864 9956 2876
rect 10008 2864 10014 2916
rect 11808 2904 11836 2935
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 12492 2944 12537 2972
rect 12492 2932 12498 2944
rect 12894 2932 12900 2984
rect 12952 2972 12958 2984
rect 13245 2975 13303 2981
rect 13245 2972 13257 2975
rect 12952 2944 13257 2972
rect 12952 2932 12958 2944
rect 13245 2941 13257 2944
rect 13291 2972 13303 2975
rect 13998 2972 14004 2984
rect 13291 2944 14004 2972
rect 13291 2941 13303 2944
rect 13245 2935 13303 2941
rect 13998 2932 14004 2944
rect 14056 2932 14062 2984
rect 13078 2904 13084 2916
rect 11808 2876 13084 2904
rect 13078 2864 13084 2876
rect 13136 2864 13142 2916
rect 14384 2904 14412 3071
rect 16040 3040 16068 3136
rect 18598 3040 18604 3052
rect 16040 3012 16436 3040
rect 18559 3012 18604 3040
rect 14645 2975 14703 2981
rect 14645 2941 14657 2975
rect 14691 2972 14703 2975
rect 16301 2975 16359 2981
rect 16301 2972 16313 2975
rect 14691 2944 16313 2972
rect 14691 2941 14703 2944
rect 14645 2935 14703 2941
rect 15120 2916 15148 2944
rect 16301 2941 16313 2944
rect 16347 2941 16359 2975
rect 16408 2972 16436 3012
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 18877 3043 18935 3049
rect 18877 3040 18889 3043
rect 18708 3012 18889 3040
rect 16557 2975 16615 2981
rect 16557 2972 16569 2975
rect 16408 2944 16569 2972
rect 16301 2935 16359 2941
rect 16557 2941 16569 2944
rect 16603 2941 16615 2975
rect 16557 2935 16615 2941
rect 17865 2975 17923 2981
rect 17865 2941 17877 2975
rect 17911 2972 17923 2975
rect 18417 2975 18475 2981
rect 18417 2972 18429 2975
rect 17911 2944 18429 2972
rect 17911 2941 17923 2944
rect 17865 2935 17923 2941
rect 18417 2941 18429 2944
rect 18463 2972 18475 2975
rect 18708 2972 18736 3012
rect 18877 3009 18889 3012
rect 18923 3009 18935 3043
rect 18877 3003 18935 3009
rect 19337 3043 19395 3049
rect 19337 3009 19349 3043
rect 19383 3040 19395 3043
rect 19383 3012 20576 3040
rect 19383 3009 19395 3012
rect 19337 3003 19395 3009
rect 18463 2944 18736 2972
rect 18463 2941 18475 2944
rect 18417 2935 18475 2941
rect 18782 2932 18788 2984
rect 18840 2972 18846 2984
rect 19061 2975 19119 2981
rect 19061 2972 19073 2975
rect 18840 2944 19073 2972
rect 18840 2932 18846 2944
rect 19061 2941 19073 2944
rect 19107 2941 19119 2975
rect 19061 2935 19119 2941
rect 19242 2932 19248 2984
rect 19300 2972 19306 2984
rect 20548 2981 20576 3012
rect 19797 2975 19855 2981
rect 19797 2972 19809 2975
rect 19300 2944 19809 2972
rect 19300 2932 19306 2944
rect 19797 2941 19809 2944
rect 19843 2941 19855 2975
rect 19797 2935 19855 2941
rect 20533 2975 20591 2981
rect 20533 2941 20545 2975
rect 20579 2941 20591 2975
rect 20533 2935 20591 2941
rect 20714 2932 20720 2984
rect 20772 2932 20778 2984
rect 14550 2904 14556 2916
rect 14384 2876 14556 2904
rect 14550 2864 14556 2876
rect 14608 2904 14614 2916
rect 14890 2907 14948 2913
rect 14890 2904 14902 2907
rect 14608 2876 14902 2904
rect 14608 2864 14614 2876
rect 14890 2873 14902 2876
rect 14936 2873 14948 2907
rect 14890 2867 14948 2873
rect 15102 2864 15108 2916
rect 15160 2864 15166 2916
rect 18598 2864 18604 2916
rect 18656 2904 18662 2916
rect 20073 2907 20131 2913
rect 18656 2876 19012 2904
rect 18656 2864 18662 2876
rect 3050 2796 3056 2848
rect 3108 2836 3114 2848
rect 9858 2836 9864 2848
rect 3108 2808 9864 2836
rect 3108 2796 3114 2808
rect 9858 2796 9864 2808
rect 9916 2796 9922 2848
rect 11425 2839 11483 2845
rect 11425 2805 11437 2839
rect 11471 2836 11483 2839
rect 11882 2836 11888 2848
rect 11471 2808 11888 2836
rect 11471 2805 11483 2808
rect 11425 2799 11483 2805
rect 11882 2796 11888 2808
rect 11940 2796 11946 2848
rect 11977 2839 12035 2845
rect 11977 2805 11989 2839
rect 12023 2836 12035 2839
rect 12526 2836 12532 2848
rect 12023 2808 12532 2836
rect 12023 2805 12035 2808
rect 11977 2799 12035 2805
rect 12526 2796 12532 2808
rect 12584 2796 12590 2848
rect 12897 2839 12955 2845
rect 12897 2805 12909 2839
rect 12943 2836 12955 2839
rect 17865 2839 17923 2845
rect 17865 2836 17877 2839
rect 12943 2808 17877 2836
rect 12943 2805 12955 2808
rect 12897 2799 12955 2805
rect 17865 2805 17877 2808
rect 17911 2805 17923 2839
rect 18046 2836 18052 2848
rect 18007 2808 18052 2836
rect 17865 2799 17923 2805
rect 18046 2796 18052 2808
rect 18104 2796 18110 2848
rect 18414 2796 18420 2848
rect 18472 2836 18478 2848
rect 18509 2839 18567 2845
rect 18509 2836 18521 2839
rect 18472 2808 18521 2836
rect 18472 2796 18478 2808
rect 18509 2805 18521 2808
rect 18555 2805 18567 2839
rect 18984 2836 19012 2876
rect 20073 2873 20085 2907
rect 20119 2904 20131 2907
rect 20732 2904 20760 2932
rect 20119 2876 20760 2904
rect 20119 2873 20131 2876
rect 20073 2867 20131 2873
rect 20717 2839 20775 2845
rect 20717 2836 20729 2839
rect 18984 2808 20729 2836
rect 18509 2799 18567 2805
rect 20717 2805 20729 2808
rect 20763 2805 20775 2839
rect 20717 2799 20775 2805
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 4706 2592 4712 2644
rect 4764 2632 4770 2644
rect 10689 2635 10747 2641
rect 10689 2632 10701 2635
rect 4764 2604 10701 2632
rect 4764 2592 4770 2604
rect 10689 2601 10701 2604
rect 10735 2601 10747 2635
rect 10689 2595 10747 2601
rect 10781 2635 10839 2641
rect 10781 2601 10793 2635
rect 10827 2632 10839 2635
rect 10870 2632 10876 2644
rect 10827 2604 10876 2632
rect 10827 2601 10839 2604
rect 10781 2595 10839 2601
rect 10870 2592 10876 2604
rect 10928 2592 10934 2644
rect 11146 2592 11152 2644
rect 11204 2632 11210 2644
rect 11701 2635 11759 2641
rect 11701 2632 11713 2635
rect 11204 2604 11713 2632
rect 11204 2592 11210 2604
rect 11701 2601 11713 2604
rect 11747 2601 11759 2635
rect 11701 2595 11759 2601
rect 14001 2635 14059 2641
rect 14001 2601 14013 2635
rect 14047 2632 14059 2635
rect 14182 2632 14188 2644
rect 14047 2604 14188 2632
rect 14047 2601 14059 2604
rect 14001 2595 14059 2601
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 14366 2632 14372 2644
rect 14327 2604 14372 2632
rect 14366 2592 14372 2604
rect 14424 2592 14430 2644
rect 14458 2592 14464 2644
rect 14516 2632 14522 2644
rect 16485 2635 16543 2641
rect 14516 2604 14561 2632
rect 14516 2592 14522 2604
rect 16485 2601 16497 2635
rect 16531 2601 16543 2635
rect 16942 2632 16948 2644
rect 16903 2604 16948 2632
rect 16485 2595 16543 2601
rect 12710 2524 12716 2576
rect 12768 2564 12774 2576
rect 13170 2564 13176 2576
rect 12768 2536 12940 2564
rect 13131 2536 13176 2564
rect 12768 2524 12774 2536
rect 9769 2499 9827 2505
rect 9769 2465 9781 2499
rect 9815 2496 9827 2499
rect 10778 2496 10784 2508
rect 9815 2468 10784 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 12912 2505 12940 2536
rect 13170 2524 13176 2536
rect 13228 2524 13234 2576
rect 16500 2564 16528 2595
rect 16942 2592 16948 2604
rect 17000 2592 17006 2644
rect 18325 2635 18383 2641
rect 18325 2601 18337 2635
rect 18371 2632 18383 2635
rect 18506 2632 18512 2644
rect 18371 2604 18512 2632
rect 18371 2601 18383 2604
rect 18325 2595 18383 2601
rect 18506 2592 18512 2604
rect 18564 2592 18570 2644
rect 18690 2592 18696 2644
rect 18748 2632 18754 2644
rect 19521 2635 19579 2641
rect 19521 2632 19533 2635
rect 18748 2604 19533 2632
rect 18748 2592 18754 2604
rect 19521 2601 19533 2604
rect 19567 2601 19579 2635
rect 19521 2595 19579 2601
rect 17770 2564 17776 2576
rect 16500 2536 17776 2564
rect 17770 2524 17776 2536
rect 17828 2524 17834 2576
rect 20898 2564 20904 2576
rect 18892 2536 20904 2564
rect 12897 2499 12955 2505
rect 12897 2465 12909 2499
rect 12943 2465 12955 2499
rect 15746 2496 15752 2508
rect 15707 2468 15752 2496
rect 12897 2459 12955 2465
rect 15746 2456 15752 2468
rect 15804 2456 15810 2508
rect 16853 2499 16911 2505
rect 16853 2465 16865 2499
rect 16899 2465 16911 2499
rect 16853 2459 16911 2465
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10873 2431 10931 2437
rect 10873 2428 10885 2431
rect 10376 2400 10885 2428
rect 10376 2388 10382 2400
rect 10873 2397 10885 2400
rect 10919 2397 10931 2431
rect 10873 2391 10931 2397
rect 11054 2388 11060 2440
rect 11112 2428 11118 2440
rect 11793 2431 11851 2437
rect 11793 2428 11805 2431
rect 11112 2400 11805 2428
rect 11112 2388 11118 2400
rect 11793 2397 11805 2400
rect 11839 2397 11851 2431
rect 11793 2391 11851 2397
rect 11882 2388 11888 2440
rect 11940 2428 11946 2440
rect 14550 2428 14556 2440
rect 11940 2400 11985 2428
rect 14511 2400 14556 2428
rect 11940 2388 11946 2400
rect 14550 2388 14556 2400
rect 14608 2388 14614 2440
rect 16022 2428 16028 2440
rect 15983 2400 16028 2428
rect 16022 2388 16028 2400
rect 16080 2388 16086 2440
rect 16868 2428 16896 2459
rect 17218 2456 17224 2508
rect 17276 2496 17282 2508
rect 17497 2499 17555 2505
rect 17497 2496 17509 2499
rect 17276 2468 17509 2496
rect 17276 2456 17282 2468
rect 17497 2465 17509 2468
rect 17543 2465 17555 2499
rect 17497 2459 17555 2465
rect 18693 2499 18751 2505
rect 18693 2465 18705 2499
rect 18739 2496 18751 2499
rect 18892 2496 18920 2536
rect 20898 2524 20904 2536
rect 20956 2524 20962 2576
rect 19242 2496 19248 2508
rect 18739 2468 18920 2496
rect 18984 2468 19248 2496
rect 18739 2465 18751 2468
rect 18693 2459 18751 2465
rect 17034 2428 17040 2440
rect 16868 2400 17040 2428
rect 17034 2388 17040 2400
rect 17092 2388 17098 2440
rect 17129 2431 17187 2437
rect 17129 2397 17141 2431
rect 17175 2428 17187 2431
rect 17402 2428 17408 2440
rect 17175 2400 17408 2428
rect 17175 2397 17187 2400
rect 17129 2391 17187 2397
rect 17402 2388 17408 2400
rect 17460 2388 17466 2440
rect 18046 2388 18052 2440
rect 18104 2428 18110 2440
rect 18984 2437 19012 2468
rect 19242 2456 19248 2468
rect 19300 2456 19306 2508
rect 19337 2499 19395 2505
rect 19337 2465 19349 2499
rect 19383 2465 19395 2499
rect 19337 2459 19395 2465
rect 18785 2431 18843 2437
rect 18785 2428 18797 2431
rect 18104 2400 18797 2428
rect 18104 2388 18110 2400
rect 18785 2397 18797 2400
rect 18831 2397 18843 2431
rect 18785 2391 18843 2397
rect 18969 2431 19027 2437
rect 18969 2397 18981 2431
rect 19015 2397 19027 2431
rect 18969 2391 19027 2397
rect 19150 2388 19156 2440
rect 19208 2428 19214 2440
rect 19352 2428 19380 2459
rect 19426 2456 19432 2508
rect 19484 2496 19490 2508
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 19484 2468 19901 2496
rect 19484 2456 19490 2468
rect 19889 2465 19901 2468
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 20162 2456 20168 2508
rect 20220 2496 20226 2508
rect 20441 2499 20499 2505
rect 20441 2496 20453 2499
rect 20220 2468 20453 2496
rect 20220 2456 20226 2468
rect 20441 2465 20453 2468
rect 20487 2465 20499 2499
rect 20441 2459 20499 2465
rect 19208 2400 19380 2428
rect 19208 2388 19214 2400
rect 9953 2363 10011 2369
rect 9953 2329 9965 2363
rect 9999 2360 10011 2363
rect 11333 2363 11391 2369
rect 9999 2332 11192 2360
rect 9999 2329 10011 2332
rect 9953 2323 10011 2329
rect 10321 2295 10379 2301
rect 10321 2261 10333 2295
rect 10367 2292 10379 2295
rect 11054 2292 11060 2304
rect 10367 2264 11060 2292
rect 10367 2261 10379 2264
rect 10321 2255 10379 2261
rect 11054 2252 11060 2264
rect 11112 2252 11118 2304
rect 11164 2292 11192 2332
rect 11333 2329 11345 2363
rect 11379 2360 11391 2363
rect 14642 2360 14648 2372
rect 11379 2332 14648 2360
rect 11379 2329 11391 2332
rect 11333 2323 11391 2329
rect 14642 2320 14648 2332
rect 14700 2320 14706 2372
rect 14734 2320 14740 2372
rect 14792 2360 14798 2372
rect 17681 2363 17739 2369
rect 17681 2360 17693 2363
rect 14792 2332 17693 2360
rect 14792 2320 14798 2332
rect 17681 2329 17693 2332
rect 17727 2329 17739 2363
rect 17681 2323 17739 2329
rect 18506 2320 18512 2372
rect 18564 2360 18570 2372
rect 20625 2363 20683 2369
rect 20625 2360 20637 2363
rect 18564 2332 20637 2360
rect 18564 2320 18570 2332
rect 20625 2329 20637 2332
rect 20671 2329 20683 2363
rect 20625 2323 20683 2329
rect 14182 2292 14188 2304
rect 11164 2264 14188 2292
rect 14182 2252 14188 2264
rect 14240 2252 14246 2304
rect 16942 2252 16948 2304
rect 17000 2292 17006 2304
rect 20073 2295 20131 2301
rect 20073 2292 20085 2295
rect 17000 2264 20085 2292
rect 17000 2252 17006 2264
rect 20073 2261 20085 2264
rect 20119 2261 20131 2295
rect 20073 2255 20131 2261
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 9674 2048 9680 2100
rect 9732 2088 9738 2100
rect 16298 2088 16304 2100
rect 9732 2060 16304 2088
rect 9732 2048 9738 2060
rect 16298 2048 16304 2060
rect 16356 2048 16362 2100
rect 17034 2048 17040 2100
rect 17092 2088 17098 2100
rect 18966 2088 18972 2100
rect 17092 2060 18972 2088
rect 17092 2048 17098 2060
rect 18966 2048 18972 2060
rect 19024 2048 19030 2100
rect 16114 1980 16120 2032
rect 16172 2020 16178 2032
rect 18046 2020 18052 2032
rect 16172 1992 18052 2020
rect 16172 1980 16178 1992
rect 18046 1980 18052 1992
rect 18104 1980 18110 2032
rect 5258 1912 5264 1964
rect 5316 1952 5322 1964
rect 8846 1952 8852 1964
rect 5316 1924 8852 1952
rect 5316 1912 5322 1924
rect 8846 1912 8852 1924
rect 8904 1912 8910 1964
rect 14642 1912 14648 1964
rect 14700 1952 14706 1964
rect 19518 1952 19524 1964
rect 14700 1924 19524 1952
rect 14700 1912 14706 1924
rect 19518 1912 19524 1924
rect 19576 1912 19582 1964
rect 11330 1368 11336 1420
rect 11388 1408 11394 1420
rect 12342 1408 12348 1420
rect 11388 1380 12348 1408
rect 11388 1368 11394 1380
rect 12342 1368 12348 1380
rect 12400 1368 12406 1420
rect 16390 1164 16396 1216
rect 16448 1204 16454 1216
rect 18690 1204 18696 1216
rect 16448 1176 18696 1204
rect 16448 1164 16454 1176
rect 18690 1164 18696 1176
rect 18748 1164 18754 1216
<< via1 >>
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 13084 20000 13136 20052
rect 14188 20043 14240 20052
rect 14188 20009 14197 20043
rect 14197 20009 14231 20043
rect 14231 20009 14240 20043
rect 14188 20000 14240 20009
rect 14556 20000 14608 20052
rect 15844 20000 15896 20052
rect 17500 20000 17552 20052
rect 18052 20000 18104 20052
rect 18880 20000 18932 20052
rect 19064 20043 19116 20052
rect 19064 20009 19073 20043
rect 19073 20009 19107 20043
rect 19107 20009 19116 20043
rect 19064 20000 19116 20009
rect 19616 20043 19668 20052
rect 19616 20009 19625 20043
rect 19625 20009 19659 20043
rect 19659 20009 19668 20043
rect 19616 20000 19668 20009
rect 19156 19932 19208 19984
rect 12624 19907 12676 19916
rect 12624 19873 12633 19907
rect 12633 19873 12667 19907
rect 12667 19873 12676 19907
rect 12624 19864 12676 19873
rect 13360 19864 13412 19916
rect 14464 19864 14516 19916
rect 15476 19907 15528 19916
rect 15476 19873 15485 19907
rect 15485 19873 15519 19907
rect 15519 19873 15528 19907
rect 15476 19864 15528 19873
rect 16028 19864 16080 19916
rect 16580 19864 16632 19916
rect 16856 19864 16908 19916
rect 18696 19864 18748 19916
rect 19432 19907 19484 19916
rect 19432 19873 19441 19907
rect 19441 19873 19475 19907
rect 19475 19873 19484 19907
rect 19432 19864 19484 19873
rect 20536 19907 20588 19916
rect 20536 19873 20545 19907
rect 20545 19873 20579 19907
rect 20579 19873 20588 19907
rect 20536 19864 20588 19873
rect 20812 19796 20864 19848
rect 19708 19728 19760 19780
rect 17132 19660 17184 19712
rect 17960 19660 18012 19712
rect 20168 19703 20220 19712
rect 20168 19669 20177 19703
rect 20177 19669 20211 19703
rect 20211 19669 20220 19703
rect 20168 19660 20220 19669
rect 20628 19660 20680 19712
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 7748 19252 7800 19304
rect 9588 19456 9640 19508
rect 19156 19499 19208 19508
rect 1400 19184 1452 19236
rect 2688 19184 2740 19236
rect 8208 19184 8260 19236
rect 10048 19252 10100 19304
rect 11428 19252 11480 19304
rect 11796 19295 11848 19304
rect 11796 19261 11805 19295
rect 11805 19261 11839 19295
rect 11839 19261 11848 19295
rect 11796 19252 11848 19261
rect 8944 19227 8996 19236
rect 8944 19193 8978 19227
rect 8978 19193 8996 19227
rect 8944 19184 8996 19193
rect 9680 19184 9732 19236
rect 2504 19116 2556 19168
rect 9772 19116 9824 19168
rect 10140 19116 10192 19168
rect 10324 19184 10376 19236
rect 19156 19465 19165 19499
rect 19165 19465 19199 19499
rect 19199 19465 19208 19499
rect 19156 19456 19208 19465
rect 14280 19252 14332 19304
rect 14372 19252 14424 19304
rect 16304 19252 16356 19304
rect 16488 19295 16540 19304
rect 16488 19261 16497 19295
rect 16497 19261 16531 19295
rect 16531 19261 16540 19295
rect 16488 19252 16540 19261
rect 16764 19252 16816 19304
rect 17224 19252 17276 19304
rect 18972 19295 19024 19304
rect 18972 19261 18981 19295
rect 18981 19261 19015 19295
rect 19015 19261 19024 19295
rect 18972 19252 19024 19261
rect 19248 19252 19300 19304
rect 20812 19295 20864 19304
rect 20812 19261 20821 19295
rect 20821 19261 20855 19295
rect 20855 19261 20864 19295
rect 20812 19252 20864 19261
rect 12716 19227 12768 19236
rect 12716 19193 12750 19227
rect 12750 19193 12768 19227
rect 12716 19184 12768 19193
rect 12808 19184 12860 19236
rect 13636 19184 13688 19236
rect 10876 19116 10928 19168
rect 11888 19116 11940 19168
rect 12532 19116 12584 19168
rect 13084 19116 13136 19168
rect 17868 19184 17920 19236
rect 19708 19184 19760 19236
rect 16396 19116 16448 19168
rect 16948 19116 17000 19168
rect 18512 19116 18564 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 2688 18912 2740 18964
rect 8760 18912 8812 18964
rect 9128 18912 9180 18964
rect 11520 18912 11572 18964
rect 11612 18912 11664 18964
rect 15292 18912 15344 18964
rect 18788 18912 18840 18964
rect 8576 18844 8628 18896
rect 11980 18844 12032 18896
rect 4160 18776 4212 18828
rect 8852 18776 8904 18828
rect 8944 18776 8996 18828
rect 6368 18708 6420 18760
rect 10232 18776 10284 18828
rect 11060 18776 11112 18828
rect 11888 18776 11940 18828
rect 15384 18844 15436 18896
rect 17224 18887 17276 18896
rect 17224 18853 17233 18887
rect 17233 18853 17267 18887
rect 17267 18853 17276 18887
rect 17224 18844 17276 18853
rect 18696 18887 18748 18896
rect 18696 18853 18705 18887
rect 18705 18853 18739 18887
rect 18739 18853 18748 18887
rect 18696 18844 18748 18853
rect 19432 18844 19484 18896
rect 14096 18776 14148 18828
rect 15292 18819 15344 18828
rect 15292 18785 15301 18819
rect 15301 18785 15335 18819
rect 15335 18785 15344 18819
rect 15292 18776 15344 18785
rect 15844 18776 15896 18828
rect 17684 18776 17736 18828
rect 9680 18751 9732 18760
rect 3056 18640 3108 18692
rect 8760 18640 8812 18692
rect 9680 18717 9689 18751
rect 9689 18717 9723 18751
rect 9723 18717 9732 18751
rect 9680 18708 9732 18717
rect 10968 18708 11020 18760
rect 14004 18751 14056 18760
rect 10784 18640 10836 18692
rect 12716 18683 12768 18692
rect 3608 18572 3660 18624
rect 8484 18572 8536 18624
rect 10048 18572 10100 18624
rect 11060 18615 11112 18624
rect 11060 18581 11069 18615
rect 11069 18581 11103 18615
rect 11103 18581 11112 18615
rect 11060 18572 11112 18581
rect 12716 18649 12725 18683
rect 12725 18649 12759 18683
rect 12759 18649 12768 18683
rect 14004 18717 14013 18751
rect 14013 18717 14047 18751
rect 14047 18717 14056 18751
rect 14004 18708 14056 18717
rect 17316 18708 17368 18760
rect 18788 18776 18840 18828
rect 19800 18776 19852 18828
rect 19156 18751 19208 18760
rect 19156 18717 19165 18751
rect 19165 18717 19199 18751
rect 19199 18717 19208 18751
rect 19156 18708 19208 18717
rect 12716 18640 12768 18649
rect 12072 18572 12124 18624
rect 12348 18572 12400 18624
rect 12808 18572 12860 18624
rect 13268 18572 13320 18624
rect 13912 18572 13964 18624
rect 17960 18640 18012 18692
rect 18512 18640 18564 18692
rect 20260 18640 20312 18692
rect 16672 18615 16724 18624
rect 16672 18581 16681 18615
rect 16681 18581 16715 18615
rect 16715 18581 16724 18615
rect 16672 18572 16724 18581
rect 16856 18572 16908 18624
rect 19524 18572 19576 18624
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 7472 18368 7524 18420
rect 8944 18368 8996 18420
rect 11888 18368 11940 18420
rect 13912 18368 13964 18420
rect 15844 18411 15896 18420
rect 15844 18377 15853 18411
rect 15853 18377 15887 18411
rect 15887 18377 15896 18411
rect 15844 18368 15896 18377
rect 18604 18368 18656 18420
rect 10784 18300 10836 18352
rect 5816 18232 5868 18284
rect 7472 18232 7524 18284
rect 8852 18232 8904 18284
rect 9864 18232 9916 18284
rect 10048 18275 10100 18284
rect 10048 18241 10057 18275
rect 10057 18241 10091 18275
rect 10091 18241 10100 18275
rect 10048 18232 10100 18241
rect 10232 18275 10284 18284
rect 10232 18241 10241 18275
rect 10241 18241 10275 18275
rect 10275 18241 10284 18275
rect 10232 18232 10284 18241
rect 12808 18275 12860 18284
rect 12808 18241 12817 18275
rect 12817 18241 12851 18275
rect 12851 18241 12860 18275
rect 12808 18232 12860 18241
rect 15844 18232 15896 18284
rect 18604 18275 18656 18284
rect 18604 18241 18613 18275
rect 18613 18241 18647 18275
rect 18647 18241 18656 18275
rect 18604 18232 18656 18241
rect 4712 18096 4764 18148
rect 6828 18096 6880 18148
rect 5264 18028 5316 18080
rect 7196 18028 7248 18080
rect 7748 18164 7800 18216
rect 10324 18164 10376 18216
rect 10968 18164 11020 18216
rect 13084 18207 13136 18216
rect 13084 18173 13118 18207
rect 13118 18173 13136 18207
rect 8852 18096 8904 18148
rect 9864 18096 9916 18148
rect 8668 18028 8720 18080
rect 10048 18028 10100 18080
rect 10600 18071 10652 18080
rect 10600 18037 10609 18071
rect 10609 18037 10643 18071
rect 10643 18037 10652 18071
rect 10600 18028 10652 18037
rect 11152 18096 11204 18148
rect 13084 18164 13136 18173
rect 15200 18164 15252 18216
rect 16028 18164 16080 18216
rect 19156 18164 19208 18216
rect 19432 18207 19484 18216
rect 19432 18173 19441 18207
rect 19441 18173 19475 18207
rect 19475 18173 19484 18207
rect 19432 18164 19484 18173
rect 19984 18207 20036 18216
rect 19984 18173 19993 18207
rect 19993 18173 20027 18207
rect 20027 18173 20036 18207
rect 19984 18164 20036 18173
rect 20076 18164 20128 18216
rect 18880 18096 18932 18148
rect 11244 18028 11296 18080
rect 12716 18028 12768 18080
rect 14188 18071 14240 18080
rect 14188 18037 14197 18071
rect 14197 18037 14231 18071
rect 14231 18037 14240 18071
rect 14188 18028 14240 18037
rect 15292 18028 15344 18080
rect 15936 18028 15988 18080
rect 16120 18071 16172 18080
rect 16120 18037 16129 18071
rect 16129 18037 16163 18071
rect 16163 18037 16172 18071
rect 16120 18028 16172 18037
rect 16212 18028 16264 18080
rect 17960 18028 18012 18080
rect 18144 18028 18196 18080
rect 19248 18028 19300 18080
rect 20168 18071 20220 18080
rect 20168 18037 20177 18071
rect 20177 18037 20211 18071
rect 20211 18037 20220 18071
rect 20168 18028 20220 18037
rect 20720 18071 20772 18080
rect 20720 18037 20729 18071
rect 20729 18037 20763 18071
rect 20763 18037 20772 18071
rect 20720 18028 20772 18037
rect 21732 18003 21784 18012
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 21732 17969 21741 18003
rect 21741 17969 21775 18003
rect 21775 17969 21784 18003
rect 21732 17960 21784 17969
rect 6920 17824 6972 17876
rect 7472 17867 7524 17876
rect 7472 17833 7481 17867
rect 7481 17833 7515 17867
rect 7515 17833 7524 17867
rect 9864 17867 9916 17876
rect 7472 17824 7524 17833
rect 9864 17833 9873 17867
rect 9873 17833 9907 17867
rect 9907 17833 9916 17867
rect 9864 17824 9916 17833
rect 10600 17824 10652 17876
rect 10784 17867 10836 17876
rect 10784 17833 10793 17867
rect 10793 17833 10827 17867
rect 10827 17833 10836 17867
rect 10784 17824 10836 17833
rect 12348 17824 12400 17876
rect 13268 17824 13320 17876
rect 14004 17824 14056 17876
rect 14556 17824 14608 17876
rect 16212 17824 16264 17876
rect 9404 17756 9456 17808
rect 10508 17756 10560 17808
rect 20076 17824 20128 17876
rect 8576 17731 8628 17740
rect 8576 17697 8585 17731
rect 8585 17697 8619 17731
rect 8619 17697 8628 17731
rect 8576 17688 8628 17697
rect 16672 17756 16724 17808
rect 18604 17756 18656 17808
rect 19432 17756 19484 17808
rect 15660 17731 15712 17740
rect 15660 17697 15669 17731
rect 15669 17697 15703 17731
rect 15703 17697 15712 17731
rect 15660 17688 15712 17697
rect 15752 17731 15804 17740
rect 15752 17697 15761 17731
rect 15761 17697 15795 17731
rect 15795 17697 15804 17731
rect 15752 17688 15804 17697
rect 16396 17688 16448 17740
rect 7748 17620 7800 17672
rect 8300 17552 8352 17604
rect 8392 17552 8444 17604
rect 11060 17620 11112 17672
rect 13176 17620 13228 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 16028 17620 16080 17672
rect 9496 17484 9548 17536
rect 13268 17484 13320 17536
rect 13452 17484 13504 17536
rect 16212 17484 16264 17536
rect 17500 17552 17552 17604
rect 17868 17620 17920 17672
rect 19156 17688 19208 17740
rect 21916 17620 21968 17672
rect 17776 17484 17828 17536
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 7012 17144 7064 17196
rect 7840 17280 7892 17332
rect 8852 17323 8904 17332
rect 8852 17289 8861 17323
rect 8861 17289 8895 17323
rect 8895 17289 8904 17323
rect 8852 17280 8904 17289
rect 12256 17280 12308 17332
rect 15476 17280 15528 17332
rect 848 17076 900 17128
rect 8852 17144 8904 17196
rect 10876 17187 10928 17196
rect 10876 17153 10885 17187
rect 10885 17153 10919 17187
rect 10919 17153 10928 17187
rect 11888 17187 11940 17196
rect 10876 17144 10928 17153
rect 11888 17153 11897 17187
rect 11897 17153 11931 17187
rect 11931 17153 11940 17187
rect 11888 17144 11940 17153
rect 9496 17119 9548 17128
rect 9496 17085 9505 17119
rect 9505 17085 9539 17119
rect 9539 17085 9548 17119
rect 9496 17076 9548 17085
rect 9956 17076 10008 17128
rect 8392 17008 8444 17060
rect 9772 17008 9824 17060
rect 9128 16983 9180 16992
rect 9128 16949 9137 16983
rect 9137 16949 9171 16983
rect 9171 16949 9180 16983
rect 9128 16940 9180 16949
rect 9220 16940 9272 16992
rect 10508 16940 10560 16992
rect 10968 16940 11020 16992
rect 11612 16940 11664 16992
rect 12256 16940 12308 16992
rect 14556 17212 14608 17264
rect 16580 17280 16632 17332
rect 19156 17280 19208 17332
rect 13268 17144 13320 17196
rect 14188 17144 14240 17196
rect 16212 17187 16264 17196
rect 16212 17153 16221 17187
rect 16221 17153 16255 17187
rect 16255 17153 16264 17187
rect 16212 17144 16264 17153
rect 16672 17144 16724 17196
rect 17776 17144 17828 17196
rect 17868 17144 17920 17196
rect 18696 17187 18748 17196
rect 16028 17076 16080 17128
rect 16120 17119 16172 17128
rect 16120 17085 16129 17119
rect 16129 17085 16163 17119
rect 16163 17085 16172 17119
rect 16120 17076 16172 17085
rect 17960 17076 18012 17128
rect 18696 17153 18705 17187
rect 18705 17153 18739 17187
rect 18739 17153 18748 17187
rect 18696 17144 18748 17153
rect 19984 17187 20036 17196
rect 19984 17153 19993 17187
rect 19993 17153 20027 17187
rect 20027 17153 20036 17187
rect 19984 17144 20036 17153
rect 20812 17187 20864 17196
rect 20812 17153 20821 17187
rect 20821 17153 20855 17187
rect 20855 17153 20864 17187
rect 20812 17144 20864 17153
rect 13452 17051 13504 17060
rect 13452 17017 13461 17051
rect 13461 17017 13495 17051
rect 13495 17017 13504 17051
rect 13452 17008 13504 17017
rect 20076 17076 20128 17128
rect 14280 16940 14332 16992
rect 16396 16940 16448 16992
rect 18420 16940 18472 16992
rect 19432 16983 19484 16992
rect 19432 16949 19441 16983
rect 19441 16949 19475 16983
rect 19475 16949 19484 16983
rect 19432 16940 19484 16949
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 10324 16736 10376 16788
rect 18512 16736 18564 16788
rect 18604 16736 18656 16788
rect 21364 16736 21416 16788
rect 10876 16668 10928 16720
rect 7012 16643 7064 16652
rect 7012 16609 7021 16643
rect 7021 16609 7055 16643
rect 7055 16609 7064 16643
rect 7012 16600 7064 16609
rect 7748 16600 7800 16652
rect 9128 16600 9180 16652
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 10416 16643 10468 16652
rect 10416 16609 10425 16643
rect 10425 16609 10459 16643
rect 10459 16609 10468 16643
rect 10416 16600 10468 16609
rect 14188 16600 14240 16652
rect 15660 16643 15712 16652
rect 8392 16439 8444 16448
rect 8392 16405 8401 16439
rect 8401 16405 8435 16439
rect 8435 16405 8444 16439
rect 8392 16396 8444 16405
rect 13912 16532 13964 16584
rect 15660 16609 15669 16643
rect 15669 16609 15703 16643
rect 15703 16609 15712 16643
rect 15660 16600 15712 16609
rect 16396 16643 16448 16652
rect 16396 16609 16405 16643
rect 16405 16609 16439 16643
rect 16439 16609 16448 16643
rect 16396 16600 16448 16609
rect 14280 16464 14332 16516
rect 14924 16532 14976 16584
rect 15476 16532 15528 16584
rect 17040 16600 17092 16652
rect 17776 16643 17828 16652
rect 17776 16609 17810 16643
rect 17810 16609 17828 16643
rect 17776 16600 17828 16609
rect 18696 16600 18748 16652
rect 17500 16575 17552 16584
rect 17500 16541 17509 16575
rect 17509 16541 17543 16575
rect 17543 16541 17552 16575
rect 17500 16532 17552 16541
rect 18512 16532 18564 16584
rect 11980 16396 12032 16448
rect 13544 16439 13596 16448
rect 13544 16405 13553 16439
rect 13553 16405 13587 16439
rect 13587 16405 13596 16439
rect 13544 16396 13596 16405
rect 13636 16396 13688 16448
rect 15292 16439 15344 16448
rect 15292 16405 15301 16439
rect 15301 16405 15335 16439
rect 15335 16405 15344 16439
rect 15292 16396 15344 16405
rect 18604 16396 18656 16448
rect 19064 16396 19116 16448
rect 19248 16396 19300 16448
rect 20444 16439 20496 16448
rect 20444 16405 20453 16439
rect 20453 16405 20487 16439
rect 20487 16405 20496 16439
rect 20444 16396 20496 16405
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 7012 16192 7064 16244
rect 9220 16192 9272 16244
rect 8392 16056 8444 16108
rect 8300 15988 8352 16040
rect 10416 16192 10468 16244
rect 12716 16192 12768 16244
rect 13728 16192 13780 16244
rect 15660 16192 15712 16244
rect 15844 16192 15896 16244
rect 10324 15988 10376 16040
rect 11888 16056 11940 16108
rect 13544 16099 13596 16108
rect 13544 16065 13553 16099
rect 13553 16065 13587 16099
rect 13587 16065 13596 16099
rect 13544 16056 13596 16065
rect 15108 16124 15160 16176
rect 13268 16031 13320 16040
rect 13268 15997 13277 16031
rect 13277 15997 13311 16031
rect 13311 15997 13320 16031
rect 13268 15988 13320 15997
rect 13452 15988 13504 16040
rect 14924 16056 14976 16108
rect 16212 16099 16264 16108
rect 16212 16065 16221 16099
rect 16221 16065 16255 16099
rect 16255 16065 16264 16099
rect 17224 16099 17276 16108
rect 16212 16056 16264 16065
rect 17224 16065 17233 16099
rect 17233 16065 17267 16099
rect 17267 16065 17276 16099
rect 17224 16056 17276 16065
rect 17776 16031 17828 16040
rect 7472 15852 7524 15904
rect 11060 15920 11112 15972
rect 12348 15920 12400 15972
rect 10600 15852 10652 15904
rect 11152 15895 11204 15904
rect 11152 15861 11161 15895
rect 11161 15861 11195 15895
rect 11195 15861 11204 15895
rect 11152 15852 11204 15861
rect 11796 15852 11848 15904
rect 13544 15920 13596 15972
rect 17776 15997 17785 16031
rect 17785 15997 17819 16031
rect 17819 15997 17828 16031
rect 17776 15988 17828 15997
rect 20076 16192 20128 16244
rect 19156 16099 19208 16108
rect 19156 16065 19165 16099
rect 19165 16065 19199 16099
rect 19199 16065 19208 16099
rect 19156 16056 19208 16065
rect 19432 16056 19484 16108
rect 20536 16056 20588 16108
rect 19248 15988 19300 16040
rect 20628 16031 20680 16040
rect 20628 15997 20637 16031
rect 20637 15997 20671 16031
rect 20671 15997 20680 16031
rect 20628 15988 20680 15997
rect 14004 15920 14056 15972
rect 14924 15920 14976 15972
rect 16856 15920 16908 15972
rect 17868 15920 17920 15972
rect 15476 15852 15528 15904
rect 16580 15895 16632 15904
rect 16580 15861 16589 15895
rect 16589 15861 16623 15895
rect 16623 15861 16632 15895
rect 16580 15852 16632 15861
rect 17316 15852 17368 15904
rect 17500 15852 17552 15904
rect 17960 15852 18012 15904
rect 18236 15895 18288 15904
rect 18236 15861 18245 15895
rect 18245 15861 18279 15895
rect 18279 15861 18288 15895
rect 18236 15852 18288 15861
rect 18972 15895 19024 15904
rect 18972 15861 18981 15895
rect 18981 15861 19015 15895
rect 19015 15861 19024 15895
rect 18972 15852 19024 15861
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 7748 15691 7800 15700
rect 7748 15657 7757 15691
rect 7757 15657 7791 15691
rect 7791 15657 7800 15691
rect 7748 15648 7800 15657
rect 8576 15648 8628 15700
rect 10416 15648 10468 15700
rect 11152 15648 11204 15700
rect 11796 15691 11848 15700
rect 11796 15657 11805 15691
rect 11805 15657 11839 15691
rect 11839 15657 11848 15691
rect 11796 15648 11848 15657
rect 12440 15648 12492 15700
rect 12716 15648 12768 15700
rect 13912 15648 13964 15700
rect 14464 15648 14516 15700
rect 7012 15580 7064 15632
rect 10508 15580 10560 15632
rect 11612 15580 11664 15632
rect 15476 15580 15528 15632
rect 16672 15648 16724 15700
rect 17224 15648 17276 15700
rect 19432 15691 19484 15700
rect 19432 15657 19441 15691
rect 19441 15657 19475 15691
rect 19475 15657 19484 15691
rect 19432 15648 19484 15657
rect 20628 15648 20680 15700
rect 16948 15580 17000 15632
rect 17868 15580 17920 15632
rect 19156 15580 19208 15632
rect 8944 15555 8996 15564
rect 8944 15521 8953 15555
rect 8953 15521 8987 15555
rect 8987 15521 8996 15555
rect 8944 15512 8996 15521
rect 9772 15512 9824 15564
rect 9956 15512 10008 15564
rect 12716 15555 12768 15564
rect 12716 15521 12725 15555
rect 12725 15521 12759 15555
rect 12759 15521 12768 15555
rect 12716 15512 12768 15521
rect 9312 15444 9364 15496
rect 11060 15444 11112 15496
rect 11980 15487 12032 15496
rect 11980 15453 11989 15487
rect 11989 15453 12023 15487
rect 12023 15453 12032 15487
rect 11980 15444 12032 15453
rect 12808 15487 12860 15496
rect 12808 15453 12817 15487
rect 12817 15453 12851 15487
rect 12851 15453 12860 15487
rect 12808 15444 12860 15453
rect 8852 15308 8904 15360
rect 10324 15351 10376 15360
rect 10324 15317 10333 15351
rect 10333 15317 10367 15351
rect 10367 15317 10376 15351
rect 10324 15308 10376 15317
rect 11060 15308 11112 15360
rect 14280 15512 14332 15564
rect 17500 15512 17552 15564
rect 18144 15512 18196 15564
rect 19340 15512 19392 15564
rect 20076 15555 20128 15564
rect 20076 15521 20085 15555
rect 20085 15521 20119 15555
rect 20119 15521 20128 15555
rect 20076 15512 20128 15521
rect 13544 15487 13596 15496
rect 13544 15453 13553 15487
rect 13553 15453 13587 15487
rect 13587 15453 13596 15487
rect 13544 15444 13596 15453
rect 16212 15444 16264 15496
rect 14648 15376 14700 15428
rect 17960 15444 18012 15496
rect 20168 15487 20220 15496
rect 20168 15453 20177 15487
rect 20177 15453 20211 15487
rect 20211 15453 20220 15487
rect 20168 15444 20220 15453
rect 20260 15487 20312 15496
rect 20260 15453 20269 15487
rect 20269 15453 20303 15487
rect 20303 15453 20312 15487
rect 20260 15444 20312 15453
rect 14188 15308 14240 15360
rect 15016 15308 15068 15360
rect 15384 15351 15436 15360
rect 15384 15317 15393 15351
rect 15393 15317 15427 15351
rect 15427 15317 15436 15351
rect 15384 15308 15436 15317
rect 17960 15308 18012 15360
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 9312 15147 9364 15156
rect 9312 15113 9321 15147
rect 9321 15113 9355 15147
rect 9355 15113 9364 15147
rect 9312 15104 9364 15113
rect 9680 15104 9732 15156
rect 12716 15104 12768 15156
rect 9128 15036 9180 15088
rect 20168 15147 20220 15156
rect 6828 14968 6880 15020
rect 7472 15011 7524 15020
rect 7472 14977 7481 15011
rect 7481 14977 7515 15011
rect 7515 14977 7524 15011
rect 7472 14968 7524 14977
rect 10324 14968 10376 15020
rect 10600 15011 10652 15020
rect 10600 14977 10609 15011
rect 10609 14977 10643 15011
rect 10643 14977 10652 15011
rect 10600 14968 10652 14977
rect 7196 14943 7248 14952
rect 7196 14909 7205 14943
rect 7205 14909 7239 14943
rect 7239 14909 7248 14943
rect 7196 14900 7248 14909
rect 7748 14900 7800 14952
rect 11060 14900 11112 14952
rect 12348 14968 12400 15020
rect 12716 14968 12768 15020
rect 13452 15011 13504 15020
rect 13452 14977 13461 15011
rect 13461 14977 13495 15011
rect 13495 14977 13504 15011
rect 13452 14968 13504 14977
rect 15476 14968 15528 15020
rect 18512 15036 18564 15088
rect 20168 15113 20177 15147
rect 20177 15113 20211 15147
rect 20211 15113 20220 15147
rect 20168 15104 20220 15113
rect 18420 14968 18472 15020
rect 20352 14968 20404 15020
rect 11704 14900 11756 14952
rect 14004 14900 14056 14952
rect 14648 14900 14700 14952
rect 15384 14900 15436 14952
rect 16580 14900 16632 14952
rect 16856 14900 16908 14952
rect 17408 14943 17460 14952
rect 17408 14909 17417 14943
rect 17417 14909 17451 14943
rect 17451 14909 17460 14943
rect 17408 14900 17460 14909
rect 17960 14900 18012 14952
rect 18512 14943 18564 14952
rect 18512 14909 18521 14943
rect 18521 14909 18555 14943
rect 18555 14909 18564 14943
rect 18512 14900 18564 14909
rect 20536 14943 20588 14952
rect 20536 14909 20545 14943
rect 20545 14909 20579 14943
rect 20579 14909 20588 14943
rect 20536 14900 20588 14909
rect 8392 14832 8444 14884
rect 8576 14832 8628 14884
rect 6828 14807 6880 14816
rect 6828 14773 6837 14807
rect 6837 14773 6871 14807
rect 6871 14773 6880 14807
rect 6828 14764 6880 14773
rect 8484 14764 8536 14816
rect 11060 14807 11112 14816
rect 11060 14773 11069 14807
rect 11069 14773 11103 14807
rect 11103 14773 11112 14807
rect 11060 14764 11112 14773
rect 12164 14832 12216 14884
rect 15016 14832 15068 14884
rect 16304 14832 16356 14884
rect 19432 14832 19484 14884
rect 11796 14764 11848 14816
rect 13268 14807 13320 14816
rect 13268 14773 13277 14807
rect 13277 14773 13311 14807
rect 13311 14773 13320 14807
rect 13268 14764 13320 14773
rect 13360 14807 13412 14816
rect 13360 14773 13369 14807
rect 13369 14773 13403 14807
rect 13403 14773 13412 14807
rect 13360 14764 13412 14773
rect 13820 14764 13872 14816
rect 14004 14764 14056 14816
rect 15108 14764 15160 14816
rect 15660 14764 15712 14816
rect 16672 14764 16724 14816
rect 16948 14764 17000 14816
rect 22468 14832 22520 14884
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 6828 14560 6880 14612
rect 7472 14492 7524 14544
rect 9128 14535 9180 14544
rect 9128 14501 9137 14535
rect 9137 14501 9171 14535
rect 9171 14501 9180 14535
rect 9128 14492 9180 14501
rect 9772 14560 9824 14612
rect 10508 14560 10560 14612
rect 14188 14603 14240 14612
rect 11704 14492 11756 14544
rect 11980 14492 12032 14544
rect 14188 14569 14197 14603
rect 14197 14569 14231 14603
rect 14231 14569 14240 14603
rect 14188 14560 14240 14569
rect 15660 14603 15712 14612
rect 15660 14569 15669 14603
rect 15669 14569 15703 14603
rect 15703 14569 15712 14603
rect 15660 14560 15712 14569
rect 16028 14560 16080 14612
rect 18696 14560 18748 14612
rect 19984 14560 20036 14612
rect 13452 14492 13504 14544
rect 7748 14424 7800 14476
rect 8852 14467 8904 14476
rect 8852 14433 8861 14467
rect 8861 14433 8895 14467
rect 8895 14433 8904 14467
rect 8852 14424 8904 14433
rect 9312 14424 9364 14476
rect 12164 14424 12216 14476
rect 8392 14331 8444 14340
rect 8392 14297 8401 14331
rect 8401 14297 8435 14331
rect 8435 14297 8444 14331
rect 8392 14288 8444 14297
rect 8852 14288 8904 14340
rect 9956 14220 10008 14272
rect 12900 14424 12952 14476
rect 13820 14288 13872 14340
rect 15292 14492 15344 14544
rect 17132 14424 17184 14476
rect 17960 14424 18012 14476
rect 14740 14399 14792 14408
rect 14740 14365 14749 14399
rect 14749 14365 14783 14399
rect 14783 14365 14792 14399
rect 14740 14356 14792 14365
rect 15016 14356 15068 14408
rect 15660 14288 15712 14340
rect 16212 14356 16264 14408
rect 17868 14356 17920 14408
rect 18512 14492 18564 14544
rect 18420 14467 18472 14476
rect 18420 14433 18429 14467
rect 18429 14433 18463 14467
rect 18463 14433 18472 14467
rect 18420 14424 18472 14433
rect 20352 14492 20404 14544
rect 18512 14356 18564 14408
rect 20168 14356 20220 14408
rect 16120 14288 16172 14340
rect 18604 14331 18656 14340
rect 16856 14220 16908 14272
rect 17040 14220 17092 14272
rect 18604 14297 18613 14331
rect 18613 14297 18647 14331
rect 18647 14297 18656 14331
rect 18604 14288 18656 14297
rect 20260 14220 20312 14272
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 8944 14016 8996 14068
rect 12808 14016 12860 14068
rect 13360 14016 13412 14068
rect 14740 14016 14792 14068
rect 7748 13948 7800 14000
rect 8852 13923 8904 13932
rect 8852 13889 8861 13923
rect 8861 13889 8895 13923
rect 8895 13889 8904 13923
rect 8852 13880 8904 13889
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 8576 13855 8628 13864
rect 8576 13821 8585 13855
rect 8585 13821 8619 13855
rect 8619 13821 8628 13855
rect 8576 13812 8628 13821
rect 16120 13948 16172 14000
rect 20076 14016 20128 14068
rect 11060 13880 11112 13932
rect 11980 13923 12032 13932
rect 11980 13889 11989 13923
rect 11989 13889 12023 13923
rect 12023 13889 12032 13923
rect 11980 13880 12032 13889
rect 11704 13812 11756 13864
rect 14188 13880 14240 13932
rect 15108 13880 15160 13932
rect 15476 13880 15528 13932
rect 15660 13923 15712 13932
rect 15660 13889 15669 13923
rect 15669 13889 15703 13923
rect 15703 13889 15712 13923
rect 15660 13880 15712 13889
rect 17592 13880 17644 13932
rect 15568 13855 15620 13864
rect 15568 13821 15577 13855
rect 15577 13821 15611 13855
rect 15611 13821 15620 13855
rect 15568 13812 15620 13821
rect 15844 13812 15896 13864
rect 17868 13812 17920 13864
rect 20352 13923 20404 13932
rect 20352 13889 20361 13923
rect 20361 13889 20395 13923
rect 20395 13889 20404 13923
rect 20352 13880 20404 13889
rect 20628 13948 20680 14000
rect 20720 13812 20772 13864
rect 12992 13744 13044 13796
rect 13728 13744 13780 13796
rect 15016 13744 15068 13796
rect 16304 13744 16356 13796
rect 16672 13744 16724 13796
rect 20168 13787 20220 13796
rect 8852 13676 8904 13728
rect 10600 13719 10652 13728
rect 10600 13685 10609 13719
rect 10609 13685 10643 13719
rect 10643 13685 10652 13719
rect 10600 13676 10652 13685
rect 12808 13719 12860 13728
rect 12808 13685 12817 13719
rect 12817 13685 12851 13719
rect 12851 13685 12860 13719
rect 12808 13676 12860 13685
rect 13084 13676 13136 13728
rect 13820 13676 13872 13728
rect 14464 13719 14516 13728
rect 14464 13685 14473 13719
rect 14473 13685 14507 13719
rect 14507 13685 14516 13719
rect 14464 13676 14516 13685
rect 15108 13719 15160 13728
rect 15108 13685 15117 13719
rect 15117 13685 15151 13719
rect 15151 13685 15160 13719
rect 15108 13676 15160 13685
rect 15752 13676 15804 13728
rect 16212 13676 16264 13728
rect 17316 13676 17368 13728
rect 17500 13719 17552 13728
rect 17500 13685 17509 13719
rect 17509 13685 17543 13719
rect 17543 13685 17552 13719
rect 17500 13676 17552 13685
rect 20168 13753 20177 13787
rect 20177 13753 20211 13787
rect 20211 13753 20220 13787
rect 20168 13744 20220 13753
rect 18144 13676 18196 13728
rect 18604 13676 18656 13728
rect 19984 13676 20036 13728
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 9220 13472 9272 13524
rect 11152 13472 11204 13524
rect 12992 13472 13044 13524
rect 13268 13472 13320 13524
rect 13820 13515 13872 13524
rect 13820 13481 13829 13515
rect 13829 13481 13863 13515
rect 13863 13481 13872 13515
rect 13820 13472 13872 13481
rect 12624 13404 12676 13456
rect 15108 13472 15160 13524
rect 16120 13472 16172 13524
rect 16396 13472 16448 13524
rect 17868 13515 17920 13524
rect 17868 13481 17877 13515
rect 17877 13481 17911 13515
rect 17911 13481 17920 13515
rect 17868 13472 17920 13481
rect 17960 13472 18012 13524
rect 19340 13472 19392 13524
rect 20444 13515 20496 13524
rect 20444 13481 20453 13515
rect 20453 13481 20487 13515
rect 20487 13481 20496 13515
rect 20444 13472 20496 13481
rect 14096 13404 14148 13456
rect 9956 13336 10008 13388
rect 10140 13379 10192 13388
rect 10140 13345 10149 13379
rect 10149 13345 10183 13379
rect 10183 13345 10192 13379
rect 10140 13336 10192 13345
rect 10232 13311 10284 13320
rect 10232 13277 10241 13311
rect 10241 13277 10275 13311
rect 10275 13277 10284 13311
rect 10232 13268 10284 13277
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 12440 13336 12492 13388
rect 13544 13336 13596 13388
rect 14280 13336 14332 13388
rect 15384 13336 15436 13388
rect 13728 13200 13780 13252
rect 14188 13268 14240 13320
rect 14924 13268 14976 13320
rect 16304 13336 16356 13388
rect 16028 13200 16080 13252
rect 16396 13200 16448 13252
rect 17868 13336 17920 13388
rect 19156 13336 19208 13388
rect 19340 13336 19392 13388
rect 17684 13268 17736 13320
rect 18696 13311 18748 13320
rect 18696 13277 18705 13311
rect 18705 13277 18739 13311
rect 18739 13277 18748 13311
rect 18696 13268 18748 13277
rect 19432 13200 19484 13252
rect 12992 13132 13044 13184
rect 16856 13132 16908 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 12164 12928 12216 12980
rect 12440 12971 12492 12980
rect 12440 12937 12449 12971
rect 12449 12937 12483 12971
rect 12483 12937 12492 12971
rect 12440 12928 12492 12937
rect 14464 12928 14516 12980
rect 12900 12860 12952 12912
rect 13268 12860 13320 12912
rect 9220 12792 9272 12844
rect 10600 12724 10652 12776
rect 12440 12724 12492 12776
rect 12992 12792 13044 12844
rect 14648 12860 14700 12912
rect 16396 12928 16448 12980
rect 18512 12928 18564 12980
rect 18696 12928 18748 12980
rect 20904 12971 20956 12980
rect 20904 12937 20913 12971
rect 20913 12937 20947 12971
rect 20947 12937 20956 12971
rect 20904 12928 20956 12937
rect 18604 12860 18656 12912
rect 10508 12656 10560 12708
rect 13084 12656 13136 12708
rect 14740 12656 14792 12708
rect 10600 12588 10652 12640
rect 10968 12631 11020 12640
rect 10968 12597 10977 12631
rect 10977 12597 11011 12631
rect 11011 12597 11020 12631
rect 10968 12588 11020 12597
rect 11704 12588 11756 12640
rect 12072 12588 12124 12640
rect 14556 12588 14608 12640
rect 15200 12724 15252 12776
rect 15660 12724 15712 12776
rect 15936 12724 15988 12776
rect 18052 12724 18104 12776
rect 18328 12724 18380 12776
rect 20720 12767 20772 12776
rect 20720 12733 20729 12767
rect 20729 12733 20763 12767
rect 20763 12733 20772 12767
rect 20720 12724 20772 12733
rect 17684 12656 17736 12708
rect 18236 12656 18288 12708
rect 18696 12656 18748 12708
rect 18880 12656 18932 12708
rect 19616 12656 19668 12708
rect 17132 12588 17184 12640
rect 17316 12588 17368 12640
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 10232 12384 10284 12436
rect 10968 12384 11020 12436
rect 11796 12384 11848 12436
rect 13912 12384 13964 12436
rect 14556 12384 14608 12436
rect 15200 12384 15252 12436
rect 15752 12384 15804 12436
rect 16856 12384 16908 12436
rect 8852 12316 8904 12368
rect 16764 12316 16816 12368
rect 17040 12316 17092 12368
rect 18052 12384 18104 12436
rect 18972 12384 19024 12436
rect 19892 12384 19944 12436
rect 18512 12316 18564 12368
rect 19156 12316 19208 12368
rect 19524 12316 19576 12368
rect 20076 12316 20128 12368
rect 10416 12291 10468 12300
rect 10416 12257 10425 12291
rect 10425 12257 10459 12291
rect 10459 12257 10468 12291
rect 10416 12248 10468 12257
rect 12256 12248 12308 12300
rect 10600 12223 10652 12232
rect 10600 12189 10609 12223
rect 10609 12189 10643 12223
rect 10643 12189 10652 12223
rect 10600 12180 10652 12189
rect 10876 12180 10928 12232
rect 8760 12112 8812 12164
rect 9220 12112 9272 12164
rect 14924 12248 14976 12300
rect 16948 12248 17000 12300
rect 13084 12223 13136 12232
rect 13084 12189 13093 12223
rect 13093 12189 13127 12223
rect 13127 12189 13136 12223
rect 13084 12180 13136 12189
rect 15016 12112 15068 12164
rect 16488 12180 16540 12232
rect 16672 12180 16724 12232
rect 17684 12248 17736 12300
rect 18328 12248 18380 12300
rect 19432 12248 19484 12300
rect 17500 12180 17552 12232
rect 18052 12223 18104 12232
rect 18052 12189 18061 12223
rect 18061 12189 18095 12223
rect 18095 12189 18104 12223
rect 18052 12180 18104 12189
rect 18604 12112 18656 12164
rect 14004 12044 14056 12096
rect 15384 12044 15436 12096
rect 16120 12044 16172 12096
rect 17592 12044 17644 12096
rect 18880 12044 18932 12096
rect 19984 12087 20036 12096
rect 19984 12053 19993 12087
rect 19993 12053 20027 12087
rect 20027 12053 20036 12087
rect 19984 12044 20036 12053
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 10140 11840 10192 11892
rect 11060 11840 11112 11892
rect 12808 11840 12860 11892
rect 13728 11840 13780 11892
rect 11704 11772 11756 11824
rect 16672 11840 16724 11892
rect 18604 11883 18656 11892
rect 18604 11849 18613 11883
rect 18613 11849 18647 11883
rect 18647 11849 18656 11883
rect 18604 11840 18656 11849
rect 19064 11840 19116 11892
rect 19156 11772 19208 11824
rect 19616 11772 19668 11824
rect 19984 11772 20036 11824
rect 8760 11747 8812 11756
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 10600 11636 10652 11688
rect 12256 11704 12308 11756
rect 14924 11747 14976 11756
rect 14924 11713 14933 11747
rect 14933 11713 14967 11747
rect 14967 11713 14976 11747
rect 14924 11704 14976 11713
rect 15752 11747 15804 11756
rect 15752 11713 15761 11747
rect 15761 11713 15795 11747
rect 15795 11713 15804 11747
rect 15752 11704 15804 11713
rect 17960 11704 18012 11756
rect 19432 11704 19484 11756
rect 20168 11747 20220 11756
rect 20168 11713 20177 11747
rect 20177 11713 20211 11747
rect 20211 11713 20220 11747
rect 20168 11704 20220 11713
rect 9864 11500 9916 11552
rect 10324 11500 10376 11552
rect 12348 11500 12400 11552
rect 16028 11679 16080 11688
rect 16028 11645 16062 11679
rect 16062 11645 16080 11679
rect 16028 11636 16080 11645
rect 12900 11543 12952 11552
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 12900 11500 12952 11509
rect 12992 11543 13044 11552
rect 12992 11509 13001 11543
rect 13001 11509 13035 11543
rect 13035 11509 13044 11543
rect 16120 11568 16172 11620
rect 19340 11568 19392 11620
rect 19524 11568 19576 11620
rect 12992 11500 13044 11509
rect 13636 11500 13688 11552
rect 14004 11543 14056 11552
rect 14004 11509 14013 11543
rect 14013 11509 14047 11543
rect 14047 11509 14056 11543
rect 17132 11543 17184 11552
rect 14004 11500 14056 11509
rect 17132 11509 17141 11543
rect 17141 11509 17175 11543
rect 17175 11509 17184 11543
rect 17132 11500 17184 11509
rect 18972 11543 19024 11552
rect 18972 11509 18981 11543
rect 18981 11509 19015 11543
rect 19015 11509 19024 11543
rect 18972 11500 19024 11509
rect 19064 11543 19116 11552
rect 19064 11509 19073 11543
rect 19073 11509 19107 11543
rect 19107 11509 19116 11543
rect 19616 11543 19668 11552
rect 19064 11500 19116 11509
rect 19616 11509 19625 11543
rect 19625 11509 19659 11543
rect 19659 11509 19668 11543
rect 19616 11500 19668 11509
rect 20812 11568 20864 11620
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 12256 11339 12308 11348
rect 12256 11305 12265 11339
rect 12265 11305 12299 11339
rect 12299 11305 12308 11339
rect 12256 11296 12308 11305
rect 12532 11296 12584 11348
rect 13268 11296 13320 11348
rect 13728 11296 13780 11348
rect 15200 11296 15252 11348
rect 15568 11296 15620 11348
rect 16120 11296 16172 11348
rect 9864 11228 9916 11280
rect 18880 11296 18932 11348
rect 19432 11296 19484 11348
rect 17132 11228 17184 11280
rect 17500 11228 17552 11280
rect 18696 11271 18748 11280
rect 18696 11237 18705 11271
rect 18705 11237 18739 11271
rect 18739 11237 18748 11271
rect 18696 11228 18748 11237
rect 8760 11160 8812 11212
rect 9680 11203 9732 11212
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 9680 11160 9732 11169
rect 10876 11203 10928 11212
rect 10876 11169 10885 11203
rect 10885 11169 10919 11203
rect 10919 11169 10928 11203
rect 10876 11160 10928 11169
rect 11980 11160 12032 11212
rect 10416 11092 10468 11144
rect 10784 11092 10836 11144
rect 12624 11092 12676 11144
rect 13728 11092 13780 11144
rect 15752 11135 15804 11144
rect 15752 11101 15761 11135
rect 15761 11101 15795 11135
rect 15795 11101 15804 11135
rect 15752 11092 15804 11101
rect 12440 11024 12492 11076
rect 13176 11024 13228 11076
rect 15016 11024 15068 11076
rect 16304 11092 16356 11144
rect 18604 11160 18656 11212
rect 19708 11228 19760 11280
rect 19432 11203 19484 11212
rect 19432 11169 19466 11203
rect 19466 11169 19484 11203
rect 19432 11160 19484 11169
rect 18880 11092 18932 11144
rect 17592 11024 17644 11076
rect 9312 10999 9364 11008
rect 9312 10965 9321 10999
rect 9321 10965 9355 10999
rect 9355 10965 9364 10999
rect 9312 10956 9364 10965
rect 15292 10956 15344 11008
rect 17684 10956 17736 11008
rect 17960 10999 18012 11008
rect 17960 10965 17969 10999
rect 17969 10965 18003 10999
rect 18003 10965 18012 10999
rect 17960 10956 18012 10965
rect 18512 10956 18564 11008
rect 18696 10956 18748 11008
rect 19524 10956 19576 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 8944 10752 8996 10804
rect 9404 10752 9456 10804
rect 12900 10752 12952 10804
rect 15108 10752 15160 10804
rect 15292 10795 15344 10804
rect 15292 10761 15301 10795
rect 15301 10761 15335 10795
rect 15335 10761 15344 10795
rect 15292 10752 15344 10761
rect 15936 10752 15988 10804
rect 14004 10684 14056 10736
rect 9312 10616 9364 10668
rect 11428 10659 11480 10668
rect 11428 10625 11437 10659
rect 11437 10625 11471 10659
rect 11471 10625 11480 10659
rect 11428 10616 11480 10625
rect 11980 10616 12032 10668
rect 13360 10616 13412 10668
rect 15016 10659 15068 10668
rect 15016 10625 15025 10659
rect 15025 10625 15059 10659
rect 15059 10625 15068 10659
rect 15016 10616 15068 10625
rect 15108 10616 15160 10668
rect 7748 10548 7800 10600
rect 10508 10548 10560 10600
rect 9312 10480 9364 10532
rect 11060 10480 11112 10532
rect 13636 10548 13688 10600
rect 14464 10548 14516 10600
rect 14648 10548 14700 10600
rect 15384 10548 15436 10600
rect 16304 10591 16356 10600
rect 16304 10557 16313 10591
rect 16313 10557 16347 10591
rect 16347 10557 16356 10591
rect 16304 10548 16356 10557
rect 17960 10548 18012 10600
rect 18512 10548 18564 10600
rect 18880 10548 18932 10600
rect 12164 10480 12216 10532
rect 16028 10480 16080 10532
rect 20444 10480 20496 10532
rect 9588 10455 9640 10464
rect 9588 10421 9597 10455
rect 9597 10421 9631 10455
rect 9631 10421 9640 10455
rect 9588 10412 9640 10421
rect 9864 10455 9916 10464
rect 9864 10421 9873 10455
rect 9873 10421 9907 10455
rect 9907 10421 9916 10455
rect 9864 10412 9916 10421
rect 11152 10412 11204 10464
rect 11704 10412 11756 10464
rect 12532 10412 12584 10464
rect 12900 10455 12952 10464
rect 12900 10421 12909 10455
rect 12909 10421 12943 10455
rect 12943 10421 12952 10455
rect 12900 10412 12952 10421
rect 13084 10412 13136 10464
rect 13544 10412 13596 10464
rect 13636 10412 13688 10464
rect 15660 10412 15712 10464
rect 17592 10412 17644 10464
rect 17684 10455 17736 10464
rect 17684 10421 17693 10455
rect 17693 10421 17727 10455
rect 17727 10421 17736 10455
rect 17684 10412 17736 10421
rect 18328 10412 18380 10464
rect 19432 10412 19484 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 9864 10208 9916 10260
rect 11980 10251 12032 10260
rect 11980 10217 11989 10251
rect 11989 10217 12023 10251
rect 12023 10217 12032 10251
rect 11980 10208 12032 10217
rect 12992 10208 13044 10260
rect 15384 10208 15436 10260
rect 16764 10208 16816 10260
rect 11060 10140 11112 10192
rect 11428 10140 11480 10192
rect 10692 10072 10744 10124
rect 15752 10140 15804 10192
rect 16028 10140 16080 10192
rect 12532 10072 12584 10124
rect 13084 10072 13136 10124
rect 13544 10115 13596 10124
rect 13544 10081 13553 10115
rect 13553 10081 13587 10115
rect 13587 10081 13596 10115
rect 13544 10072 13596 10081
rect 15292 10072 15344 10124
rect 15384 10072 15436 10124
rect 15660 10115 15712 10124
rect 15660 10081 15669 10115
rect 15669 10081 15703 10115
rect 15703 10081 15712 10115
rect 15660 10072 15712 10081
rect 16856 10072 16908 10124
rect 9588 10004 9640 10056
rect 10600 10047 10652 10056
rect 10600 10013 10609 10047
rect 10609 10013 10643 10047
rect 10643 10013 10652 10047
rect 10600 10004 10652 10013
rect 9680 9936 9732 9988
rect 13360 9936 13412 9988
rect 14464 10004 14516 10056
rect 15936 10047 15988 10056
rect 15936 10013 15945 10047
rect 15945 10013 15979 10047
rect 15979 10013 15988 10047
rect 15936 10004 15988 10013
rect 17868 10072 17920 10124
rect 17500 10047 17552 10056
rect 16028 9936 16080 9988
rect 16856 9936 16908 9988
rect 17500 10013 17509 10047
rect 17509 10013 17543 10047
rect 17543 10013 17552 10047
rect 17500 10004 17552 10013
rect 17960 10004 18012 10056
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 19708 10047 19760 10056
rect 19708 10013 19717 10047
rect 19717 10013 19751 10047
rect 19751 10013 19760 10047
rect 19708 10004 19760 10013
rect 20168 10004 20220 10056
rect 17592 9936 17644 9988
rect 18052 9936 18104 9988
rect 14188 9911 14240 9920
rect 14188 9877 14197 9911
rect 14197 9877 14231 9911
rect 14231 9877 14240 9911
rect 14188 9868 14240 9877
rect 16580 9868 16632 9920
rect 18512 9868 18564 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 9036 9664 9088 9716
rect 9312 9664 9364 9716
rect 9772 9528 9824 9580
rect 10600 9664 10652 9716
rect 11060 9664 11112 9716
rect 15384 9664 15436 9716
rect 11888 9571 11940 9580
rect 11888 9537 11897 9571
rect 11897 9537 11931 9571
rect 11931 9537 11940 9571
rect 11888 9528 11940 9537
rect 13728 9528 13780 9580
rect 7748 9503 7800 9512
rect 7748 9469 7757 9503
rect 7757 9469 7791 9503
rect 7791 9469 7800 9503
rect 7748 9460 7800 9469
rect 8576 9460 8628 9512
rect 8576 9324 8628 9376
rect 9588 9392 9640 9444
rect 9128 9367 9180 9376
rect 9128 9333 9137 9367
rect 9137 9333 9171 9367
rect 9171 9333 9180 9367
rect 9128 9324 9180 9333
rect 9772 9324 9824 9376
rect 11152 9460 11204 9512
rect 14464 9460 14516 9512
rect 17960 9664 18012 9716
rect 18144 9596 18196 9648
rect 18236 9596 18288 9648
rect 18788 9596 18840 9648
rect 20168 9596 20220 9648
rect 17500 9528 17552 9580
rect 18880 9528 18932 9580
rect 10416 9392 10468 9444
rect 10600 9392 10652 9444
rect 14280 9392 14332 9444
rect 18328 9460 18380 9512
rect 15384 9392 15436 9444
rect 10876 9324 10928 9376
rect 14096 9324 14148 9376
rect 16764 9435 16816 9444
rect 16764 9401 16773 9435
rect 16773 9401 16807 9435
rect 16807 9401 16816 9435
rect 16764 9392 16816 9401
rect 17408 9392 17460 9444
rect 17960 9392 18012 9444
rect 18420 9435 18472 9444
rect 18420 9401 18429 9435
rect 18429 9401 18463 9435
rect 18463 9401 18472 9435
rect 18420 9392 18472 9401
rect 19524 9392 19576 9444
rect 20812 9571 20864 9580
rect 20812 9537 20821 9571
rect 20821 9537 20855 9571
rect 20855 9537 20864 9571
rect 20812 9528 20864 9537
rect 16304 9367 16356 9376
rect 16304 9333 16313 9367
rect 16313 9333 16347 9367
rect 16347 9333 16356 9367
rect 16304 9324 16356 9333
rect 17592 9324 17644 9376
rect 19248 9324 19300 9376
rect 19616 9324 19668 9376
rect 20444 9324 20496 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 11060 9120 11112 9172
rect 10048 9052 10100 9104
rect 6920 8984 6972 9036
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 9772 8916 9824 8968
rect 10600 8984 10652 9036
rect 11060 8984 11112 9036
rect 13452 8984 13504 9036
rect 14188 9120 14240 9172
rect 14280 9120 14332 9172
rect 15108 9120 15160 9172
rect 15292 9163 15344 9172
rect 15292 9129 15301 9163
rect 15301 9129 15335 9163
rect 15335 9129 15344 9163
rect 15292 9120 15344 9129
rect 15384 9120 15436 9172
rect 15936 9120 15988 9172
rect 16304 9052 16356 9104
rect 17684 9052 17736 9104
rect 18236 9052 18288 9104
rect 18696 9052 18748 9104
rect 19524 9120 19576 9172
rect 19616 9052 19668 9104
rect 14740 9027 14792 9036
rect 10416 8959 10468 8968
rect 10416 8925 10425 8959
rect 10425 8925 10459 8959
rect 10459 8925 10468 8959
rect 10416 8916 10468 8925
rect 11152 8916 11204 8968
rect 11704 8848 11756 8900
rect 8576 8823 8628 8832
rect 8576 8789 8585 8823
rect 8585 8789 8619 8823
rect 8619 8789 8628 8823
rect 8576 8780 8628 8789
rect 10784 8780 10836 8832
rect 12716 8916 12768 8968
rect 13360 8916 13412 8968
rect 14096 8959 14148 8968
rect 14096 8925 14105 8959
rect 14105 8925 14139 8959
rect 14139 8925 14148 8959
rect 14096 8916 14148 8925
rect 14740 8993 14749 9027
rect 14749 8993 14783 9027
rect 14783 8993 14792 9027
rect 14740 8984 14792 8993
rect 15660 9027 15712 9036
rect 15660 8993 15669 9027
rect 15669 8993 15703 9027
rect 15703 8993 15712 9027
rect 15660 8984 15712 8993
rect 15844 8984 15896 9036
rect 16396 8984 16448 9036
rect 15108 8916 15160 8968
rect 15476 8916 15528 8968
rect 15936 8959 15988 8968
rect 12808 8848 12860 8900
rect 14556 8891 14608 8900
rect 14556 8857 14565 8891
rect 14565 8857 14599 8891
rect 14599 8857 14608 8891
rect 14556 8848 14608 8857
rect 15936 8925 15945 8959
rect 15945 8925 15979 8959
rect 15979 8925 15988 8959
rect 15936 8916 15988 8925
rect 16304 8916 16356 8968
rect 16488 8916 16540 8968
rect 18328 8984 18380 9036
rect 17224 8848 17276 8900
rect 12716 8780 12768 8832
rect 15660 8780 15712 8832
rect 16212 8780 16264 8832
rect 18972 8780 19024 8832
rect 19340 8780 19392 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 11152 8576 11204 8628
rect 10876 8508 10928 8560
rect 11612 8440 11664 8492
rect 13728 8576 13780 8628
rect 15844 8576 15896 8628
rect 15936 8576 15988 8628
rect 18604 8576 18656 8628
rect 19708 8576 19760 8628
rect 15660 8440 15712 8492
rect 18512 8483 18564 8492
rect 18512 8449 18521 8483
rect 18521 8449 18555 8483
rect 18555 8449 18564 8483
rect 18512 8440 18564 8449
rect 20444 8508 20496 8560
rect 19064 8440 19116 8492
rect 19616 8483 19668 8492
rect 19616 8449 19625 8483
rect 19625 8449 19659 8483
rect 19659 8449 19668 8483
rect 19616 8440 19668 8449
rect 20536 8483 20588 8492
rect 20536 8449 20545 8483
rect 20545 8449 20579 8483
rect 20579 8449 20588 8483
rect 20536 8440 20588 8449
rect 20628 8483 20680 8492
rect 20628 8449 20637 8483
rect 20637 8449 20671 8483
rect 20671 8449 20680 8483
rect 20628 8440 20680 8449
rect 7748 8372 7800 8424
rect 9128 8372 9180 8424
rect 9864 8415 9916 8424
rect 9864 8381 9873 8415
rect 9873 8381 9907 8415
rect 9907 8381 9916 8415
rect 9864 8372 9916 8381
rect 11152 8372 11204 8424
rect 12808 8415 12860 8424
rect 12808 8381 12817 8415
rect 12817 8381 12851 8415
rect 12851 8381 12860 8415
rect 12808 8372 12860 8381
rect 14096 8372 14148 8424
rect 14556 8372 14608 8424
rect 10784 8304 10836 8356
rect 13176 8304 13228 8356
rect 13636 8304 13688 8356
rect 18052 8372 18104 8424
rect 19248 8372 19300 8424
rect 16488 8304 16540 8356
rect 9220 8236 9272 8288
rect 10968 8236 11020 8288
rect 13820 8236 13872 8288
rect 14464 8279 14516 8288
rect 14464 8245 14473 8279
rect 14473 8245 14507 8279
rect 14507 8245 14516 8279
rect 14464 8236 14516 8245
rect 15752 8236 15804 8288
rect 17408 8304 17460 8356
rect 19064 8304 19116 8356
rect 19984 8304 20036 8356
rect 20076 8279 20128 8288
rect 20076 8245 20085 8279
rect 20085 8245 20119 8279
rect 20119 8245 20128 8279
rect 20076 8236 20128 8245
rect 20444 8279 20496 8288
rect 20444 8245 20453 8279
rect 20453 8245 20487 8279
rect 20487 8245 20496 8279
rect 20444 8236 20496 8245
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 8576 8032 8628 8084
rect 11060 8032 11112 8084
rect 11796 8032 11848 8084
rect 12624 7964 12676 8016
rect 13176 8007 13228 8016
rect 13176 7973 13185 8007
rect 13185 7973 13219 8007
rect 13219 7973 13228 8007
rect 13176 7964 13228 7973
rect 13912 8032 13964 8084
rect 14556 8032 14608 8084
rect 15108 8032 15160 8084
rect 17868 8032 17920 8084
rect 17960 8032 18012 8084
rect 20444 8032 20496 8084
rect 19248 7964 19300 8016
rect 9864 7896 9916 7948
rect 10968 7896 11020 7948
rect 12900 7896 12952 7948
rect 9220 7871 9272 7880
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 8668 7760 8720 7812
rect 9956 7760 10008 7812
rect 13176 7828 13228 7880
rect 13544 7896 13596 7948
rect 15200 7896 15252 7948
rect 15660 7896 15712 7948
rect 15844 7939 15896 7948
rect 15844 7905 15878 7939
rect 15878 7905 15896 7939
rect 15844 7896 15896 7905
rect 16120 7896 16172 7948
rect 17592 7896 17644 7948
rect 18880 7896 18932 7948
rect 19984 7939 20036 7948
rect 19984 7905 19993 7939
rect 19993 7905 20027 7939
rect 20027 7905 20036 7939
rect 19984 7896 20036 7905
rect 14464 7871 14516 7880
rect 14464 7837 14473 7871
rect 14473 7837 14507 7871
rect 14507 7837 14516 7871
rect 14464 7828 14516 7837
rect 13912 7760 13964 7812
rect 3424 7692 3476 7744
rect 11796 7692 11848 7744
rect 12072 7692 12124 7744
rect 12992 7692 13044 7744
rect 13084 7692 13136 7744
rect 17132 7692 17184 7744
rect 17684 7735 17736 7744
rect 17684 7701 17693 7735
rect 17693 7701 17727 7735
rect 17727 7701 17736 7735
rect 17684 7692 17736 7701
rect 17868 7760 17920 7812
rect 20168 7828 20220 7880
rect 20536 7828 20588 7880
rect 20444 7760 20496 7812
rect 19156 7692 19208 7744
rect 19340 7692 19392 7744
rect 19616 7735 19668 7744
rect 19616 7701 19625 7735
rect 19625 7701 19659 7735
rect 19659 7701 19668 7735
rect 19616 7692 19668 7701
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 11152 7488 11204 7540
rect 10784 7420 10836 7472
rect 12900 7420 12952 7472
rect 12072 7352 12124 7404
rect 13084 7395 13136 7404
rect 13084 7361 13093 7395
rect 13093 7361 13127 7395
rect 13127 7361 13136 7395
rect 13084 7352 13136 7361
rect 13268 7420 13320 7472
rect 13544 7420 13596 7472
rect 15844 7352 15896 7404
rect 9312 7284 9364 7336
rect 12992 7327 13044 7336
rect 12992 7293 13001 7327
rect 13001 7293 13035 7327
rect 13035 7293 13044 7327
rect 12992 7284 13044 7293
rect 13452 7284 13504 7336
rect 13912 7327 13964 7336
rect 13912 7293 13946 7327
rect 13946 7293 13964 7327
rect 13912 7284 13964 7293
rect 16120 7284 16172 7336
rect 9588 7216 9640 7268
rect 13268 7216 13320 7268
rect 8576 7191 8628 7200
rect 8576 7157 8585 7191
rect 8585 7157 8619 7191
rect 8619 7157 8628 7191
rect 8576 7148 8628 7157
rect 9680 7148 9732 7200
rect 11612 7148 11664 7200
rect 15292 7191 15344 7200
rect 15292 7157 15301 7191
rect 15301 7157 15335 7191
rect 15335 7157 15344 7191
rect 15292 7148 15344 7157
rect 15660 7148 15712 7200
rect 15752 7191 15804 7200
rect 15752 7157 15761 7191
rect 15761 7157 15795 7191
rect 15795 7157 15804 7191
rect 18788 7327 18840 7336
rect 18788 7293 18797 7327
rect 18797 7293 18831 7327
rect 18831 7293 18840 7327
rect 18788 7284 18840 7293
rect 16856 7216 16908 7268
rect 17316 7216 17368 7268
rect 19892 7284 19944 7336
rect 20260 7284 20312 7336
rect 20536 7216 20588 7268
rect 15752 7148 15804 7157
rect 17500 7148 17552 7200
rect 19248 7148 19300 7200
rect 19708 7148 19760 7200
rect 20628 7191 20680 7200
rect 20628 7157 20637 7191
rect 20637 7157 20671 7191
rect 20671 7157 20680 7191
rect 20628 7148 20680 7157
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 9312 6987 9364 6996
rect 9312 6953 9321 6987
rect 9321 6953 9355 6987
rect 9355 6953 9364 6987
rect 9312 6944 9364 6953
rect 9680 6987 9732 6996
rect 9680 6953 9689 6987
rect 9689 6953 9723 6987
rect 9723 6953 9732 6987
rect 9680 6944 9732 6953
rect 12624 6944 12676 6996
rect 13084 6944 13136 6996
rect 15752 6944 15804 6996
rect 16764 6944 16816 6996
rect 17316 6944 17368 6996
rect 20076 6944 20128 6996
rect 11152 6876 11204 6928
rect 12072 6876 12124 6928
rect 12992 6876 13044 6928
rect 8760 6808 8812 6860
rect 10876 6851 10928 6860
rect 10140 6783 10192 6792
rect 7472 6604 7524 6656
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 10876 6817 10885 6851
rect 10885 6817 10919 6851
rect 10919 6817 10928 6851
rect 10876 6808 10928 6817
rect 10968 6808 11020 6860
rect 15016 6808 15068 6860
rect 18972 6876 19024 6928
rect 11060 6740 11112 6792
rect 13636 6740 13688 6792
rect 14464 6783 14516 6792
rect 14464 6749 14473 6783
rect 14473 6749 14507 6783
rect 14507 6749 14516 6783
rect 14464 6740 14516 6749
rect 15568 6740 15620 6792
rect 19616 6808 19668 6860
rect 20904 6876 20956 6928
rect 16856 6783 16908 6792
rect 16856 6749 16865 6783
rect 16865 6749 16899 6783
rect 16899 6749 16908 6783
rect 16856 6740 16908 6749
rect 17040 6740 17092 6792
rect 17868 6783 17920 6792
rect 17868 6749 17877 6783
rect 17877 6749 17911 6783
rect 17911 6749 17920 6783
rect 17868 6740 17920 6749
rect 14372 6672 14424 6724
rect 15292 6672 15344 6724
rect 15936 6672 15988 6724
rect 19708 6740 19760 6792
rect 20352 6783 20404 6792
rect 20352 6749 20361 6783
rect 20361 6749 20395 6783
rect 20395 6749 20404 6783
rect 20352 6740 20404 6749
rect 21916 6672 21968 6724
rect 9588 6604 9640 6656
rect 11060 6604 11112 6656
rect 12624 6647 12676 6656
rect 12624 6613 12633 6647
rect 12633 6613 12667 6647
rect 12667 6613 12676 6647
rect 12624 6604 12676 6613
rect 13728 6604 13780 6656
rect 15476 6604 15528 6656
rect 17040 6604 17092 6656
rect 17316 6604 17368 6656
rect 18696 6604 18748 6656
rect 18972 6604 19024 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 8576 6400 8628 6452
rect 10140 6443 10192 6452
rect 10140 6409 10149 6443
rect 10149 6409 10183 6443
rect 10183 6409 10192 6443
rect 10140 6400 10192 6409
rect 11152 6443 11204 6452
rect 11152 6409 11161 6443
rect 11161 6409 11195 6443
rect 11195 6409 11204 6443
rect 11152 6400 11204 6409
rect 13268 6443 13320 6452
rect 13268 6409 13277 6443
rect 13277 6409 13311 6443
rect 13311 6409 13320 6443
rect 13268 6400 13320 6409
rect 13820 6400 13872 6452
rect 19064 6400 19116 6452
rect 8760 6332 8812 6384
rect 7472 6307 7524 6316
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 12900 6332 12952 6384
rect 10324 6264 10376 6316
rect 12992 6264 13044 6316
rect 13268 6264 13320 6316
rect 15752 6332 15804 6384
rect 15016 6264 15068 6316
rect 15384 6307 15436 6316
rect 15384 6273 15393 6307
rect 15393 6273 15427 6307
rect 15427 6273 15436 6307
rect 15384 6264 15436 6273
rect 7748 6239 7800 6248
rect 7748 6205 7782 6239
rect 7782 6205 7800 6239
rect 7748 6196 7800 6205
rect 10692 6196 10744 6248
rect 16580 6332 16632 6384
rect 16672 6332 16724 6384
rect 19432 6400 19484 6452
rect 20536 6443 20588 6452
rect 20536 6409 20545 6443
rect 20545 6409 20579 6443
rect 20579 6409 20588 6443
rect 20536 6400 20588 6409
rect 17132 6264 17184 6316
rect 17316 6307 17368 6316
rect 17316 6273 17325 6307
rect 17325 6273 17359 6307
rect 17359 6273 17368 6307
rect 17316 6264 17368 6273
rect 17500 6307 17552 6316
rect 17500 6273 17509 6307
rect 17509 6273 17543 6307
rect 17543 6273 17552 6307
rect 17500 6264 17552 6273
rect 15936 6196 15988 6248
rect 17684 6196 17736 6248
rect 11704 6128 11756 6180
rect 13636 6171 13688 6180
rect 13636 6137 13645 6171
rect 13645 6137 13679 6171
rect 13679 6137 13688 6171
rect 13636 6128 13688 6137
rect 13728 6171 13780 6180
rect 13728 6137 13737 6171
rect 13737 6137 13771 6171
rect 13771 6137 13780 6171
rect 13728 6128 13780 6137
rect 16028 6128 16080 6180
rect 16120 6128 16172 6180
rect 18052 6128 18104 6180
rect 18420 6128 18472 6180
rect 19064 6196 19116 6248
rect 20260 6196 20312 6248
rect 20720 6196 20772 6248
rect 19340 6128 19392 6180
rect 9496 6103 9548 6112
rect 9496 6069 9505 6103
rect 9505 6069 9539 6103
rect 9539 6069 9548 6103
rect 9496 6060 9548 6069
rect 9680 6060 9732 6112
rect 11796 6060 11848 6112
rect 12256 6060 12308 6112
rect 18604 6103 18656 6112
rect 18604 6069 18613 6103
rect 18613 6069 18647 6103
rect 18647 6069 18656 6103
rect 18604 6060 18656 6069
rect 18696 6060 18748 6112
rect 19248 6060 19300 6112
rect 20812 6060 20864 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 7748 5856 7800 5908
rect 9496 5856 9548 5908
rect 9680 5899 9732 5908
rect 9680 5865 9689 5899
rect 9689 5865 9723 5899
rect 9723 5865 9732 5899
rect 9680 5856 9732 5865
rect 10048 5899 10100 5908
rect 10048 5865 10057 5899
rect 10057 5865 10091 5899
rect 10091 5865 10100 5899
rect 10048 5856 10100 5865
rect 12900 5856 12952 5908
rect 4068 5788 4120 5840
rect 7196 5788 7248 5840
rect 12072 5788 12124 5840
rect 12256 5788 12308 5840
rect 12808 5788 12860 5840
rect 15108 5856 15160 5908
rect 15568 5856 15620 5908
rect 15844 5856 15896 5908
rect 7472 5720 7524 5772
rect 10968 5720 11020 5772
rect 12624 5720 12676 5772
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 10324 5695 10376 5704
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 10324 5652 10376 5661
rect 13544 5720 13596 5772
rect 13084 5695 13136 5704
rect 13084 5661 13093 5695
rect 13093 5661 13127 5695
rect 13127 5661 13136 5695
rect 13084 5652 13136 5661
rect 14004 5695 14056 5704
rect 14004 5661 14013 5695
rect 14013 5661 14047 5695
rect 14047 5661 14056 5695
rect 14004 5652 14056 5661
rect 16672 5788 16724 5840
rect 17868 5856 17920 5908
rect 15384 5720 15436 5772
rect 15200 5652 15252 5704
rect 15844 5652 15896 5704
rect 16120 5652 16172 5704
rect 16396 5720 16448 5772
rect 16580 5763 16632 5772
rect 16580 5729 16589 5763
rect 16589 5729 16623 5763
rect 16623 5729 16632 5763
rect 16580 5720 16632 5729
rect 18880 5720 18932 5772
rect 17040 5652 17092 5704
rect 16856 5584 16908 5636
rect 11060 5516 11112 5568
rect 12072 5516 12124 5568
rect 12256 5559 12308 5568
rect 12256 5525 12265 5559
rect 12265 5525 12299 5559
rect 12299 5525 12308 5559
rect 12256 5516 12308 5525
rect 12532 5559 12584 5568
rect 12532 5525 12541 5559
rect 12541 5525 12575 5559
rect 12575 5525 12584 5559
rect 12532 5516 12584 5525
rect 13544 5559 13596 5568
rect 13544 5525 13553 5559
rect 13553 5525 13587 5559
rect 13587 5525 13596 5559
rect 13544 5516 13596 5525
rect 15660 5516 15712 5568
rect 15844 5516 15896 5568
rect 17868 5516 17920 5568
rect 18788 5652 18840 5704
rect 19064 5720 19116 5772
rect 19616 5788 19668 5840
rect 20352 5788 20404 5840
rect 20536 5720 20588 5772
rect 18420 5584 18472 5636
rect 19156 5516 19208 5568
rect 19340 5516 19392 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 11704 5312 11756 5364
rect 16764 5312 16816 5364
rect 19432 5312 19484 5364
rect 19616 5355 19668 5364
rect 19616 5321 19625 5355
rect 19625 5321 19659 5355
rect 19659 5321 19668 5355
rect 19616 5312 19668 5321
rect 9956 5244 10008 5296
rect 12440 5244 12492 5296
rect 12256 5176 12308 5228
rect 12992 5244 13044 5296
rect 13084 5219 13136 5228
rect 13084 5185 13093 5219
rect 13093 5185 13127 5219
rect 13127 5185 13136 5219
rect 13084 5176 13136 5185
rect 13452 5219 13504 5228
rect 13452 5185 13461 5219
rect 13461 5185 13495 5219
rect 13495 5185 13504 5219
rect 13452 5176 13504 5185
rect 16120 5176 16172 5228
rect 17868 5176 17920 5228
rect 20444 5219 20496 5228
rect 20444 5185 20453 5219
rect 20453 5185 20487 5219
rect 20487 5185 20496 5219
rect 20444 5176 20496 5185
rect 20904 5219 20956 5228
rect 20904 5185 20913 5219
rect 20913 5185 20947 5219
rect 20947 5185 20956 5219
rect 20904 5176 20956 5185
rect 12532 5108 12584 5160
rect 12992 5108 13044 5160
rect 13268 5108 13320 5160
rect 15200 5108 15252 5160
rect 13544 5040 13596 5092
rect 13728 5083 13780 5092
rect 13728 5049 13762 5083
rect 13762 5049 13780 5083
rect 13728 5040 13780 5049
rect 11336 5015 11388 5024
rect 11336 4981 11345 5015
rect 11345 4981 11379 5015
rect 11379 4981 11388 5015
rect 11336 4972 11388 4981
rect 12440 5015 12492 5024
rect 12440 4981 12449 5015
rect 12449 4981 12483 5015
rect 12483 4981 12492 5015
rect 12440 4972 12492 4981
rect 17592 5108 17644 5160
rect 20260 5151 20312 5160
rect 20260 5117 20269 5151
rect 20269 5117 20303 5151
rect 20303 5117 20312 5151
rect 20260 5108 20312 5117
rect 16488 5015 16540 5024
rect 16488 4981 16497 5015
rect 16497 4981 16531 5015
rect 16531 4981 16540 5015
rect 16488 4972 16540 4981
rect 16580 4972 16632 5024
rect 18696 5040 18748 5092
rect 19064 5040 19116 5092
rect 18788 4972 18840 5024
rect 19892 5015 19944 5024
rect 19892 4981 19901 5015
rect 19901 4981 19935 5015
rect 19935 4981 19944 5015
rect 19892 4972 19944 4981
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 11336 4768 11388 4820
rect 14188 4768 14240 4820
rect 18052 4768 18104 4820
rect 18696 4811 18748 4820
rect 18696 4777 18705 4811
rect 18705 4777 18739 4811
rect 18739 4777 18748 4811
rect 18696 4768 18748 4777
rect 20444 4768 20496 4820
rect 296 4700 348 4752
rect 12992 4700 13044 4752
rect 13176 4700 13228 4752
rect 12072 4632 12124 4684
rect 12256 4675 12308 4684
rect 12256 4641 12290 4675
rect 12290 4641 12308 4675
rect 12256 4632 12308 4641
rect 14004 4675 14056 4684
rect 14004 4641 14013 4675
rect 14013 4641 14047 4675
rect 14047 4641 14056 4675
rect 14004 4632 14056 4641
rect 9680 4496 9732 4548
rect 11980 4496 12032 4548
rect 13728 4564 13780 4616
rect 16488 4700 16540 4752
rect 17040 4700 17092 4752
rect 19156 4700 19208 4752
rect 14556 4632 14608 4684
rect 15200 4632 15252 4684
rect 16764 4632 16816 4684
rect 17408 4632 17460 4684
rect 18604 4564 18656 4616
rect 20444 4607 20496 4616
rect 17040 4539 17092 4548
rect 7656 4428 7708 4480
rect 13268 4428 13320 4480
rect 13452 4428 13504 4480
rect 15200 4428 15252 4480
rect 17040 4505 17049 4539
rect 17049 4505 17083 4539
rect 17083 4505 17092 4539
rect 17040 4496 17092 4505
rect 18328 4496 18380 4548
rect 19708 4496 19760 4548
rect 20444 4573 20453 4607
rect 20453 4573 20487 4607
rect 20487 4573 20496 4607
rect 20444 4564 20496 4573
rect 20904 4607 20956 4616
rect 20904 4573 20913 4607
rect 20913 4573 20947 4607
rect 20947 4573 20956 4607
rect 20904 4564 20956 4573
rect 20352 4496 20404 4548
rect 19800 4471 19852 4480
rect 19800 4437 19809 4471
rect 19809 4437 19843 4471
rect 19843 4437 19852 4471
rect 19800 4428 19852 4437
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 13268 4224 13320 4276
rect 12256 4156 12308 4208
rect 5816 4088 5868 4140
rect 8944 4088 8996 4140
rect 12440 4088 12492 4140
rect 9128 4020 9180 4072
rect 11612 4063 11664 4072
rect 11612 4029 11621 4063
rect 11621 4029 11655 4063
rect 11655 4029 11664 4063
rect 11612 4020 11664 4029
rect 9220 3952 9272 4004
rect 12624 4020 12676 4072
rect 12808 4063 12860 4072
rect 12808 4029 12817 4063
rect 12817 4029 12851 4063
rect 12851 4029 12860 4063
rect 12808 4020 12860 4029
rect 3608 3884 3660 3936
rect 13084 3952 13136 4004
rect 10324 3884 10376 3936
rect 14004 4088 14056 4140
rect 13452 4063 13504 4072
rect 13452 4029 13461 4063
rect 13461 4029 13495 4063
rect 13495 4029 13504 4063
rect 13452 4020 13504 4029
rect 15476 4088 15528 4140
rect 15660 4131 15712 4140
rect 15660 4097 15669 4131
rect 15669 4097 15703 4131
rect 15703 4097 15712 4131
rect 15660 4088 15712 4097
rect 16488 4156 16540 4208
rect 16396 4088 16448 4140
rect 14372 4020 14424 4072
rect 16580 4020 16632 4072
rect 16856 4020 16908 4072
rect 19064 4224 19116 4276
rect 19340 4156 19392 4208
rect 19616 4156 19668 4208
rect 19892 4088 19944 4140
rect 20536 4088 20588 4140
rect 22468 4088 22520 4140
rect 18972 4063 19024 4072
rect 18972 4029 18981 4063
rect 18981 4029 19015 4063
rect 19015 4029 19024 4063
rect 18972 4020 19024 4029
rect 19800 4020 19852 4072
rect 20260 4020 20312 4072
rect 13268 3952 13320 4004
rect 15844 3952 15896 4004
rect 13912 3884 13964 3936
rect 15292 3884 15344 3936
rect 16028 3884 16080 3936
rect 16580 3927 16632 3936
rect 16580 3893 16589 3927
rect 16589 3893 16623 3927
rect 16623 3893 16632 3927
rect 16580 3884 16632 3893
rect 17684 3884 17736 3936
rect 18788 3884 18840 3936
rect 20260 3884 20312 3936
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 1400 3680 1452 3732
rect 16948 3680 17000 3732
rect 17868 3680 17920 3732
rect 7472 3612 7524 3664
rect 10048 3612 10100 3664
rect 10232 3612 10284 3664
rect 10784 3612 10836 3664
rect 13268 3612 13320 3664
rect 9128 3544 9180 3596
rect 11152 3544 11204 3596
rect 11888 3544 11940 3596
rect 13452 3544 13504 3596
rect 1952 3476 2004 3528
rect 10140 3476 10192 3528
rect 10232 3476 10284 3528
rect 10876 3476 10928 3528
rect 12440 3476 12492 3528
rect 13084 3476 13136 3528
rect 13636 3476 13688 3528
rect 6368 3408 6420 3460
rect 16120 3612 16172 3664
rect 18880 3680 18932 3732
rect 19156 3680 19208 3732
rect 20628 3680 20680 3732
rect 21364 3680 21416 3732
rect 16764 3587 16816 3596
rect 14004 3519 14056 3528
rect 14004 3485 14013 3519
rect 14013 3485 14047 3519
rect 14047 3485 14056 3519
rect 14004 3476 14056 3485
rect 2504 3340 2556 3392
rect 13820 3408 13872 3460
rect 16764 3553 16773 3587
rect 16773 3553 16807 3587
rect 16807 3553 16816 3587
rect 16764 3544 16816 3553
rect 17592 3544 17644 3596
rect 18604 3612 18656 3664
rect 18972 3612 19024 3664
rect 19984 3544 20036 3596
rect 16028 3519 16080 3528
rect 16028 3485 16037 3519
rect 16037 3485 16071 3519
rect 16071 3485 16080 3519
rect 16028 3476 16080 3485
rect 12900 3340 12952 3392
rect 14464 3340 14516 3392
rect 14648 3383 14700 3392
rect 14648 3349 14657 3383
rect 14657 3349 14691 3383
rect 14691 3349 14700 3383
rect 14648 3340 14700 3349
rect 16948 3340 17000 3392
rect 19064 3340 19116 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 848 3136 900 3188
rect 13268 3136 13320 3188
rect 14648 3136 14700 3188
rect 16028 3179 16080 3188
rect 16028 3145 16037 3179
rect 16037 3145 16071 3179
rect 16071 3145 16080 3179
rect 16028 3136 16080 3145
rect 17592 3136 17644 3188
rect 8208 3068 8260 3120
rect 9772 3068 9824 3120
rect 11980 3068 12032 3120
rect 10048 3043 10100 3052
rect 10048 3009 10057 3043
rect 10057 3009 10091 3043
rect 10091 3009 10100 3043
rect 10048 3000 10100 3009
rect 4160 2932 4212 2984
rect 9680 2932 9732 2984
rect 10324 2975 10376 2984
rect 10324 2941 10358 2975
rect 10358 2941 10376 2975
rect 10324 2932 10376 2941
rect 10876 2932 10928 2984
rect 12072 3000 12124 3052
rect 8576 2864 8628 2916
rect 9956 2864 10008 2916
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 12440 2932 12492 2941
rect 12900 2932 12952 2984
rect 14004 2932 14056 2984
rect 13084 2864 13136 2916
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 18788 2932 18840 2984
rect 19248 2932 19300 2984
rect 20720 2932 20772 2984
rect 14556 2864 14608 2916
rect 15108 2864 15160 2916
rect 18604 2864 18656 2916
rect 3056 2796 3108 2848
rect 9864 2796 9916 2848
rect 11888 2796 11940 2848
rect 12532 2796 12584 2848
rect 18052 2839 18104 2848
rect 18052 2805 18061 2839
rect 18061 2805 18095 2839
rect 18095 2805 18104 2839
rect 18052 2796 18104 2805
rect 18420 2796 18472 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 4712 2592 4764 2644
rect 10876 2592 10928 2644
rect 11152 2592 11204 2644
rect 14188 2592 14240 2644
rect 14372 2635 14424 2644
rect 14372 2601 14381 2635
rect 14381 2601 14415 2635
rect 14415 2601 14424 2635
rect 14372 2592 14424 2601
rect 14464 2635 14516 2644
rect 14464 2601 14473 2635
rect 14473 2601 14507 2635
rect 14507 2601 14516 2635
rect 14464 2592 14516 2601
rect 16948 2635 17000 2644
rect 12716 2524 12768 2576
rect 13176 2567 13228 2576
rect 10784 2456 10836 2508
rect 13176 2533 13185 2567
rect 13185 2533 13219 2567
rect 13219 2533 13228 2567
rect 13176 2524 13228 2533
rect 16948 2601 16957 2635
rect 16957 2601 16991 2635
rect 16991 2601 17000 2635
rect 16948 2592 17000 2601
rect 18512 2592 18564 2644
rect 18696 2592 18748 2644
rect 17776 2524 17828 2576
rect 15752 2499 15804 2508
rect 15752 2465 15761 2499
rect 15761 2465 15795 2499
rect 15795 2465 15804 2499
rect 15752 2456 15804 2465
rect 10324 2388 10376 2440
rect 11060 2388 11112 2440
rect 11888 2431 11940 2440
rect 11888 2397 11897 2431
rect 11897 2397 11931 2431
rect 11931 2397 11940 2431
rect 14556 2431 14608 2440
rect 11888 2388 11940 2397
rect 14556 2397 14565 2431
rect 14565 2397 14599 2431
rect 14599 2397 14608 2431
rect 14556 2388 14608 2397
rect 16028 2431 16080 2440
rect 16028 2397 16037 2431
rect 16037 2397 16071 2431
rect 16071 2397 16080 2431
rect 16028 2388 16080 2397
rect 17224 2456 17276 2508
rect 20904 2524 20956 2576
rect 17040 2388 17092 2440
rect 17408 2388 17460 2440
rect 18052 2388 18104 2440
rect 19248 2456 19300 2508
rect 19156 2388 19208 2440
rect 19432 2456 19484 2508
rect 20168 2456 20220 2508
rect 11060 2252 11112 2304
rect 14648 2320 14700 2372
rect 14740 2320 14792 2372
rect 18512 2320 18564 2372
rect 14188 2252 14240 2304
rect 16948 2252 17000 2304
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 9680 2048 9732 2100
rect 16304 2048 16356 2100
rect 17040 2048 17092 2100
rect 18972 2048 19024 2100
rect 16120 1980 16172 2032
rect 18052 1980 18104 2032
rect 5264 1912 5316 1964
rect 8852 1912 8904 1964
rect 14648 1912 14700 1964
rect 19524 1912 19576 1964
rect 11336 1368 11388 1420
rect 12348 1368 12400 1420
rect 16396 1164 16448 1216
rect 18696 1164 18748 1216
<< metal2 >>
rect 294 22000 350 22800
rect 846 22000 902 22800
rect 1398 22000 1454 22800
rect 1950 22000 2006 22800
rect 2502 22000 2558 22800
rect 3054 22000 3110 22800
rect 3606 22000 3662 22800
rect 4158 22000 4214 22800
rect 4710 22000 4766 22800
rect 5262 22000 5318 22800
rect 5814 22000 5870 22800
rect 6366 22000 6422 22800
rect 6918 22000 6974 22800
rect 7470 22000 7526 22800
rect 8022 22000 8078 22800
rect 8574 22000 8630 22800
rect 9126 22000 9182 22800
rect 9678 22000 9734 22800
rect 10230 22000 10286 22800
rect 10782 22000 10838 22800
rect 11334 22000 11390 22800
rect 11978 22000 12034 22800
rect 12530 22000 12586 22800
rect 13082 22000 13138 22800
rect 13634 22000 13690 22800
rect 14186 22000 14242 22800
rect 14738 22000 14794 22800
rect 15290 22000 15346 22800
rect 15842 22000 15898 22800
rect 16394 22000 16450 22800
rect 16946 22000 17002 22800
rect 17498 22000 17554 22800
rect 18050 22000 18106 22800
rect 18602 22000 18658 22800
rect 18786 22128 18842 22137
rect 18786 22063 18842 22072
rect 308 18329 336 22000
rect 294 18320 350 18329
rect 294 18255 350 18264
rect 860 17134 888 22000
rect 1412 19242 1440 22000
rect 1400 19236 1452 19242
rect 1400 19178 1452 19184
rect 1964 18737 1992 22000
rect 2516 19174 2544 22000
rect 2688 19236 2740 19242
rect 2688 19178 2740 19184
rect 2504 19168 2556 19174
rect 2504 19110 2556 19116
rect 2700 18970 2728 19178
rect 2688 18964 2740 18970
rect 2688 18906 2740 18912
rect 1950 18728 2006 18737
rect 3068 18698 3096 22000
rect 1950 18663 2006 18672
rect 3056 18692 3108 18698
rect 3056 18634 3108 18640
rect 3620 18630 3648 22000
rect 4172 18834 4200 22000
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 3608 18624 3660 18630
rect 3608 18566 3660 18572
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4724 18154 4752 22000
rect 4712 18148 4764 18154
rect 4712 18090 4764 18096
rect 5276 18086 5304 22000
rect 5828 18290 5856 22000
rect 6380 18766 6408 22000
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 5816 18284 5868 18290
rect 5816 18226 5868 18232
rect 6828 18148 6880 18154
rect 6828 18090 6880 18096
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 3422 17232 3478 17241
rect 3422 17167 3478 17176
rect 848 17128 900 17134
rect 848 17070 900 17076
rect 3436 7750 3464 17167
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 6840 15026 6868 18090
rect 6932 17882 6960 22000
rect 7484 18426 7512 22000
rect 8036 20346 8064 22000
rect 8036 20318 8248 20346
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7196 18080 7248 18086
rect 7196 18022 7248 18028
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 7024 16658 7052 17138
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 7024 16250 7052 16594
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 7024 15638 7052 16186
rect 7012 15632 7064 15638
rect 7012 15574 7064 15580
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 7208 14958 7236 18022
rect 7484 17882 7512 18226
rect 7760 18222 7788 19246
rect 8220 19242 8248 20318
rect 8208 19236 8260 19242
rect 8208 19178 8260 19184
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 8588 18902 8616 22000
rect 8944 19236 8996 19242
rect 8944 19178 8996 19184
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8576 18896 8628 18902
rect 8772 18873 8800 18906
rect 8576 18838 8628 18844
rect 8758 18864 8814 18873
rect 8956 18834 8984 19178
rect 9140 18970 9168 22000
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9600 19122 9628 19450
rect 9692 19242 9720 22000
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 9680 19236 9732 19242
rect 9680 19178 9732 19184
rect 9772 19168 9824 19174
rect 9600 19094 9720 19122
rect 9772 19110 9824 19116
rect 9128 18964 9180 18970
rect 9128 18906 9180 18912
rect 8758 18799 8814 18808
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 8944 18828 8996 18834
rect 8944 18770 8996 18776
rect 8760 18692 8812 18698
rect 8760 18634 8812 18640
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7484 17354 7512 17818
rect 7760 17762 7788 18158
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 7760 17734 7880 17762
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7484 17326 7696 17354
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7484 15026 7512 15846
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6840 14618 6868 14758
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4068 5840 4120 5846
rect 4066 5808 4068 5817
rect 4120 5808 4122 5817
rect 4066 5743 4122 5752
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 296 4752 348 4758
rect 296 4694 348 4700
rect 308 800 336 4694
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 1400 3732 1452 3738
rect 1400 3674 1452 3680
rect 848 3188 900 3194
rect 848 3130 900 3136
rect 860 800 888 3130
rect 1412 800 1440 3674
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 1964 800 1992 3470
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2516 800 2544 3334
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 3068 800 3096 2790
rect 3620 800 3648 3878
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 4172 800 4200 2926
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4724 800 4752 2586
rect 5264 1964 5316 1970
rect 5264 1906 5316 1912
rect 5276 800 5304 1906
rect 5828 800 5856 4082
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 6380 800 6408 3402
rect 6932 800 6960 8978
rect 7208 5846 7236 14894
rect 7484 14550 7512 14962
rect 7472 14544 7524 14550
rect 7472 14486 7524 14492
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7484 6322 7512 6598
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7196 5840 7248 5846
rect 7196 5782 7248 5788
rect 7484 5778 7512 6258
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7668 4486 7696 17326
rect 7760 16658 7788 17614
rect 7852 17338 7880 17734
rect 8300 17604 8352 17610
rect 8300 17546 8352 17552
rect 8392 17604 8444 17610
rect 8392 17546 8444 17552
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7748 16652 7800 16658
rect 7748 16594 7800 16600
rect 7760 15706 7788 16594
rect 8312 16046 8340 17546
rect 8404 17066 8432 17546
rect 8392 17060 8444 17066
rect 8392 17002 8444 17008
rect 8404 16454 8432 17002
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8404 16114 8432 16390
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7760 14482 7788 14894
rect 8392 14884 8444 14890
rect 8392 14826 8444 14832
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7760 14006 7788 14418
rect 8404 14346 8432 14826
rect 8496 14822 8524 18566
rect 8772 18193 8800 18634
rect 8864 18290 8892 18770
rect 8956 18426 8984 18770
rect 9692 18766 9720 19094
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9692 18465 9720 18702
rect 9678 18456 9734 18465
rect 8944 18420 8996 18426
rect 9678 18391 9734 18400
rect 8944 18362 8996 18368
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 8758 18184 8814 18193
rect 8758 18119 8814 18128
rect 8852 18148 8904 18154
rect 8852 18090 8904 18096
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8588 15706 8616 17682
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8576 14884 8628 14890
rect 8576 14826 8628 14832
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8392 14340 8444 14346
rect 8392 14282 8444 14288
rect 7748 14000 7800 14006
rect 7748 13942 7800 13948
rect 8588 13870 8616 14826
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7760 9518 7788 10542
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 7760 8430 7788 9454
rect 8588 9382 8616 9454
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 8588 8090 8616 8774
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8680 7818 8708 18022
rect 8864 17338 8892 18090
rect 9404 17808 9456 17814
rect 9404 17750 9456 17756
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8864 17202 8892 17274
rect 8852 17196 8904 17202
rect 8852 17138 8904 17144
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 9140 16658 9168 16934
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 9232 16250 9260 16934
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8864 14482 8892 15302
rect 8852 14476 8904 14482
rect 8852 14418 8904 14424
rect 8852 14340 8904 14346
rect 8852 14282 8904 14288
rect 8864 13938 8892 14282
rect 8956 14074 8984 15506
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9324 15162 9352 15438
rect 9312 15156 9364 15162
rect 9312 15098 9364 15104
rect 9128 15088 9180 15094
rect 9128 15030 9180 15036
rect 9140 14550 9168 15030
rect 9128 14544 9180 14550
rect 9128 14486 9180 14492
rect 9312 14476 9364 14482
rect 9232 14436 9312 14464
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 9232 13938 9260 14436
rect 9312 14418 9364 14424
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8864 12374 8892 13670
rect 9232 13530 9260 13874
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9232 12850 9260 13466
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 8852 12368 8904 12374
rect 8852 12310 8904 12316
rect 8760 12164 8812 12170
rect 8760 12106 8812 12112
rect 8772 11762 8800 12106
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8772 11218 8800 11698
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8668 7812 8720 7818
rect 8668 7754 8720 7760
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 8588 6458 8616 7142
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8772 6390 8800 6802
rect 8760 6384 8812 6390
rect 8760 6326 8812 6332
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7760 5914 7788 6190
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7484 800 7512 3606
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 8220 1442 8248 3062
rect 8576 2916 8628 2922
rect 8576 2858 8628 2864
rect 8036 1414 8248 1442
rect 8036 800 8064 1414
rect 8588 800 8616 2858
rect 8864 1970 8892 12310
rect 9232 12170 9260 12786
rect 9220 12164 9272 12170
rect 9220 12106 9272 12112
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 8956 4146 8984 10746
rect 9324 10674 9352 10950
rect 9416 10810 9444 17750
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9508 17134 9536 17478
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9784 17066 9812 19110
rect 10060 18986 10088 19246
rect 10244 19224 10272 22000
rect 10506 19272 10562 19281
rect 10324 19236 10376 19242
rect 10244 19196 10324 19224
rect 10506 19207 10562 19216
rect 10324 19178 10376 19184
rect 10140 19168 10192 19174
rect 10192 19128 10272 19156
rect 10140 19110 10192 19116
rect 10060 18958 10180 18986
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 10060 18290 10088 18566
rect 9864 18284 9916 18290
rect 10048 18284 10100 18290
rect 9916 18244 9996 18272
rect 9864 18226 9916 18232
rect 9864 18148 9916 18154
rect 9864 18090 9916 18096
rect 9876 17882 9904 18090
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9968 17134 9996 18244
rect 10048 18226 10100 18232
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 9772 17060 9824 17066
rect 9772 17002 9824 17008
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9692 15162 9720 16594
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9784 14618 9812 15506
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9968 14278 9996 15506
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9968 13394 9996 14214
rect 10060 13705 10088 18022
rect 10152 17785 10180 18958
rect 10244 18834 10272 19128
rect 10232 18828 10284 18834
rect 10232 18770 10284 18776
rect 10244 18290 10272 18770
rect 10414 18456 10470 18465
rect 10414 18391 10470 18400
rect 10232 18284 10284 18290
rect 10232 18226 10284 18232
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10336 17921 10364 18158
rect 10322 17912 10378 17921
rect 10322 17847 10378 17856
rect 10138 17776 10194 17785
rect 10138 17711 10194 17720
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 10336 16697 10364 16730
rect 10322 16688 10378 16697
rect 10428 16658 10456 18391
rect 10520 17814 10548 19207
rect 10796 18698 10824 22000
rect 11348 20074 11376 22000
rect 11348 20046 11652 20074
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11428 19304 11480 19310
rect 11428 19246 11480 19252
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 10784 18692 10836 18698
rect 10784 18634 10836 18640
rect 10784 18352 10836 18358
rect 10690 18320 10746 18329
rect 10784 18294 10836 18300
rect 10690 18255 10746 18264
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 10612 17882 10640 18022
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10322 16623 10378 16632
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10428 16250 10456 16594
rect 10416 16244 10468 16250
rect 10416 16186 10468 16192
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10336 15450 10364 15982
rect 10428 15706 10456 16186
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10520 15638 10548 16934
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10508 15632 10560 15638
rect 10508 15574 10560 15580
rect 10336 15422 10456 15450
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10336 15026 10364 15302
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10046 13696 10102 13705
rect 10046 13631 10102 13640
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9876 11286 9904 11494
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9312 10532 9364 10538
rect 9312 10474 9364 10480
rect 9324 9722 9352 10474
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9600 10062 9628 10406
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 9048 3108 9076 9658
rect 9600 9450 9628 9998
rect 9692 9994 9720 11154
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9876 10266 9904 10406
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9784 9382 9812 9522
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 9772 9376 9824 9382
rect 9824 9336 9904 9364
rect 9772 9318 9824 9324
rect 9140 8974 9168 9318
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9140 8430 9168 8910
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9232 7886 9260 8230
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9140 3602 9168 4014
rect 9232 4010 9260 7822
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9324 7002 9352 7278
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9600 6662 9628 7210
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 7002 9720 7142
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9508 5914 9536 6054
rect 9692 5914 9720 6054
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 8956 3080 9076 3108
rect 8956 2666 8984 3080
rect 9692 2990 9720 4490
rect 9784 3126 9812 8910
rect 9876 8430 9904 9336
rect 10060 9110 10088 13631
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 10152 11898 10180 13330
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10244 12442 10272 13262
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10336 11558 10364 13262
rect 10428 12424 10456 15422
rect 10612 15026 10640 15846
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10520 12714 10548 14554
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10612 12782 10640 13670
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10508 12708 10560 12714
rect 10508 12650 10560 12656
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10428 12396 10548 12424
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10428 11370 10456 12242
rect 10336 11342 10456 11370
rect 10336 11121 10364 11342
rect 10416 11144 10468 11150
rect 10322 11112 10378 11121
rect 10416 11086 10468 11092
rect 10322 11047 10378 11056
rect 10230 9616 10286 9625
rect 10230 9551 10286 9560
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 9864 8424 9916 8430
rect 9916 8384 9996 8412
rect 9864 8366 9916 8372
rect 9864 7948 9916 7954
rect 9864 7890 9916 7896
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9876 2854 9904 7890
rect 9968 7818 9996 8384
rect 9956 7812 10008 7818
rect 9956 7754 10008 7760
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10152 6458 10180 6734
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10046 6352 10102 6361
rect 10046 6287 10102 6296
rect 10060 5914 10088 6287
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 9968 2922 9996 5238
rect 10060 3670 10088 5850
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 10152 3534 10180 5646
rect 10244 3670 10272 9551
rect 10336 6440 10364 11047
rect 10428 9625 10456 11086
rect 10520 10606 10548 12396
rect 10612 12238 10640 12582
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10612 11694 10640 12174
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10704 10130 10732 18255
rect 10796 17882 10824 18294
rect 10888 18057 10916 19110
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 10980 18465 11008 18702
rect 11072 18630 11100 18770
rect 11440 18680 11468 19246
rect 11518 19000 11574 19009
rect 11624 18970 11652 20046
rect 11796 19304 11848 19310
rect 11796 19246 11848 19252
rect 11518 18935 11520 18944
rect 11572 18935 11574 18944
rect 11612 18964 11664 18970
rect 11520 18906 11572 18912
rect 11612 18906 11664 18912
rect 11440 18652 11744 18680
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 10966 18456 11022 18465
rect 10966 18391 11022 18400
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 10874 18048 10930 18057
rect 10874 17983 10930 17992
rect 10784 17876 10836 17882
rect 10784 17818 10836 17824
rect 10980 17762 11008 18158
rect 10796 17734 11008 17762
rect 10796 15609 10824 17734
rect 11072 17678 11100 18566
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 11060 17672 11112 17678
rect 11060 17614 11112 17620
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 10888 16726 10916 17138
rect 10968 16992 11020 16998
rect 10968 16934 11020 16940
rect 10876 16720 10928 16726
rect 10876 16662 10928 16668
rect 10782 15600 10838 15609
rect 10782 15535 10838 15544
rect 10796 11150 10824 15535
rect 10980 13818 11008 16934
rect 11164 15994 11192 18090
rect 11244 18080 11296 18086
rect 11242 18048 11244 18057
rect 11296 18048 11298 18057
rect 11242 17983 11298 17992
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11060 15972 11112 15978
rect 11164 15966 11284 15994
rect 11060 15914 11112 15920
rect 11072 15502 11100 15914
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11164 15706 11192 15846
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11060 15496 11112 15502
rect 11256 15450 11284 15966
rect 11624 15638 11652 16934
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11060 15438 11112 15444
rect 11164 15422 11284 15450
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 11072 14958 11100 15302
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 11072 13938 11100 14758
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10980 13790 11100 13818
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10980 12442 11008 12582
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10888 11218 10916 12174
rect 11072 11898 11100 13790
rect 11164 13530 11192 15422
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11716 15042 11744 18652
rect 11808 15994 11836 19246
rect 11888 19168 11940 19174
rect 11992 19156 12020 22000
rect 12544 19174 12572 22000
rect 13096 20058 13124 22000
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 11940 19128 12020 19156
rect 12532 19168 12584 19174
rect 11888 19110 11940 19116
rect 12532 19110 12584 19116
rect 11980 18896 12032 18902
rect 11980 18838 12032 18844
rect 12070 18864 12126 18873
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 11900 18426 11928 18770
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11900 16114 11928 17138
rect 11992 17105 12020 18838
rect 12126 18822 12204 18850
rect 12070 18799 12126 18808
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 11978 17096 12034 17105
rect 11978 17031 12034 17040
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11808 15966 11928 15994
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11808 15706 11836 15846
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 11624 15014 11744 15042
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11428 10668 11480 10674
rect 11428 10610 11480 10616
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 11072 10282 11100 10474
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 10980 10254 11100 10282
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10612 9722 10640 9998
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10414 9616 10470 9625
rect 10414 9551 10470 9560
rect 10416 9444 10468 9450
rect 10416 9386 10468 9392
rect 10600 9444 10652 9450
rect 10600 9386 10652 9392
rect 10428 8974 10456 9386
rect 10612 9042 10640 9386
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10336 6412 10456 6440
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10336 5710 10364 6258
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10232 3664 10284 3670
rect 10232 3606 10284 3612
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10244 3074 10272 3470
rect 10060 3058 10272 3074
rect 10048 3052 10272 3058
rect 10100 3046 10272 3052
rect 10048 2994 10100 3000
rect 10336 2990 10364 3878
rect 10324 2984 10376 2990
rect 10230 2952 10286 2961
rect 9956 2916 10008 2922
rect 10324 2926 10376 2932
rect 10230 2887 10286 2896
rect 9956 2858 10008 2864
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 8956 2638 9168 2666
rect 8852 1964 8904 1970
rect 8852 1906 8904 1912
rect 9140 800 9168 2638
rect 9680 2100 9732 2106
rect 9680 2042 9732 2048
rect 9692 800 9720 2042
rect 10244 800 10272 2887
rect 10336 2446 10364 2926
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10428 2122 10456 6412
rect 10704 6254 10732 10066
rect 10980 9602 11008 10254
rect 11060 10192 11112 10198
rect 11060 10134 11112 10140
rect 11072 9722 11100 10134
rect 11060 9716 11112 9722
rect 11060 9658 11112 9664
rect 10980 9574 11100 9602
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10796 8362 10824 8774
rect 10888 8566 10916 9318
rect 11072 9178 11100 9574
rect 11164 9518 11192 10406
rect 11440 10198 11468 10610
rect 11428 10192 11480 10198
rect 11428 10134 11480 10140
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 10876 8560 10928 8566
rect 10876 8502 10928 8508
rect 10784 8356 10836 8362
rect 10784 8298 10836 8304
rect 10796 7886 10824 8298
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10796 7478 10824 7822
rect 10784 7472 10836 7478
rect 10784 7414 10836 7420
rect 10888 6866 10916 8502
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10980 7954 11008 8230
rect 11072 8090 11100 8978
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11164 8634 11192 8910
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11624 8498 11652 15014
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11716 14550 11744 14894
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11704 14544 11756 14550
rect 11704 14486 11756 14492
rect 11716 13870 11744 14486
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11716 11830 11744 12582
rect 11808 12442 11836 14758
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11716 8906 11744 10406
rect 11900 9586 11928 15966
rect 11992 15502 12020 16390
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 11992 13938 12020 14486
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 12084 12646 12112 18566
rect 12176 14890 12204 18822
rect 12348 18624 12400 18630
rect 12348 18566 12400 18572
rect 12360 18329 12388 18566
rect 12346 18320 12402 18329
rect 12346 18255 12402 18264
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 12268 16998 12296 17274
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12164 14884 12216 14890
rect 12164 14826 12216 14832
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12176 12986 12204 14418
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12268 12866 12296 16934
rect 12360 15978 12388 17818
rect 12348 15972 12400 15978
rect 12348 15914 12400 15920
rect 12360 15026 12388 15914
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12452 14906 12480 15642
rect 12452 14878 12572 14906
rect 12544 13954 12572 14878
rect 12452 13926 12572 13954
rect 12452 13512 12480 13926
rect 12452 13484 12572 13512
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12452 12986 12480 13330
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12176 12838 12296 12866
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 12070 12336 12126 12345
rect 12176 12322 12204 12838
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12126 12294 12204 12322
rect 12256 12300 12308 12306
rect 12070 12271 12126 12280
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11992 10674 12020 11154
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 11992 10266 12020 10610
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11152 8424 11204 8430
rect 11152 8366 11204 8372
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 11164 7546 11192 8366
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11808 7750 11836 8026
rect 12084 7834 12112 12271
rect 12256 12242 12308 12248
rect 12268 11762 12296 12242
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12268 11354 12296 11698
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12164 10532 12216 10538
rect 12164 10474 12216 10480
rect 11992 7806 12112 7834
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10980 5778 11008 6802
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11072 6662 11100 6734
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 11072 5574 11100 6598
rect 11164 6458 11192 6870
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11348 4826 11376 4966
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11624 4078 11652 7142
rect 11794 6216 11850 6225
rect 11704 6180 11756 6186
rect 11794 6151 11850 6160
rect 11704 6122 11756 6128
rect 11716 5370 11744 6122
rect 11808 6118 11836 6151
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11992 4554 12020 7806
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 12084 7410 12112 7686
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12084 6934 12112 7346
rect 12072 6928 12124 6934
rect 12072 6870 12124 6876
rect 12072 5840 12124 5846
rect 12070 5808 12072 5817
rect 12124 5808 12126 5817
rect 12070 5743 12126 5752
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 12084 4690 12112 5510
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 11980 4548 12032 4554
rect 11980 4490 12032 4496
rect 11612 4072 11664 4078
rect 11612 4014 11664 4020
rect 10784 3664 10836 3670
rect 10784 3606 10836 3612
rect 10796 2514 10824 3606
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10888 2990 10916 3470
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 11164 2650 11192 3538
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11900 2854 11928 3538
rect 11980 3120 12032 3126
rect 11980 3062 12032 3068
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10428 2094 10824 2122
rect 10796 800 10824 2094
rect 10888 1601 10916 2586
rect 11900 2446 11928 2790
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 11072 2310 11100 2382
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 10874 1592 10930 1601
rect 10874 1527 10930 1536
rect 11336 1420 11388 1426
rect 11336 1362 11388 1368
rect 11348 800 11376 1362
rect 11992 800 12020 3062
rect 12084 3058 12112 4626
rect 12072 3052 12124 3058
rect 12072 2994 12124 3000
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 1950 0 2006 800
rect 2502 0 2558 800
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4158 0 4214 800
rect 4710 0 4766 800
rect 5262 0 5318 800
rect 5814 0 5870 800
rect 6366 0 6422 800
rect 6918 0 6974 800
rect 7470 0 7526 800
rect 8022 0 8078 800
rect 8574 0 8630 800
rect 9126 0 9182 800
rect 9678 0 9734 800
rect 10230 0 10286 800
rect 10782 0 10838 800
rect 11334 0 11390 800
rect 11978 0 12034 800
rect 12176 649 12204 10474
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12268 5846 12296 6054
rect 12256 5840 12308 5846
rect 12256 5782 12308 5788
rect 12256 5568 12308 5574
rect 12256 5510 12308 5516
rect 12268 5234 12296 5510
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12268 4690 12296 5170
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12268 4214 12296 4626
rect 12256 4208 12308 4214
rect 12256 4150 12308 4156
rect 12360 1426 12388 11494
rect 12452 11082 12480 12718
rect 12544 11354 12572 13484
rect 12636 13462 12664 19858
rect 12716 19236 12768 19242
rect 12716 19178 12768 19184
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12728 18698 12756 19178
rect 12716 18692 12768 18698
rect 12716 18634 12768 18640
rect 12820 18630 12848 19178
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12820 18290 12848 18566
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 13096 18222 13124 19110
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13084 18216 13136 18222
rect 13136 18176 13216 18204
rect 13084 18158 13136 18164
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12728 16250 12756 18022
rect 13188 17678 13216 18176
rect 13280 17882 13308 18566
rect 13268 17876 13320 17882
rect 13268 17818 13320 17824
rect 13176 17672 13228 17678
rect 13176 17614 13228 17620
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13280 17202 13308 17478
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12728 15706 12756 16186
rect 13268 16040 13320 16046
rect 13266 16008 13268 16017
rect 13320 16008 13322 16017
rect 13266 15943 13322 15952
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12728 15162 12756 15506
rect 12808 15496 12860 15502
rect 12808 15438 12860 15444
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12624 13456 12676 13462
rect 12624 13398 12676 13404
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12532 10464 12584 10470
rect 12452 10424 12532 10452
rect 12452 5302 12480 10424
rect 12532 10406 12584 10412
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12544 5658 12572 10066
rect 12636 8022 12664 11086
rect 12728 8974 12756 14962
rect 12820 14074 12848 15438
rect 13372 15348 13400 19858
rect 13648 19242 13676 22000
rect 14200 20058 14228 22000
rect 14752 20346 14780 22000
rect 14568 20318 14780 20346
rect 14568 20058 14596 20318
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 13636 19236 13688 19242
rect 13636 19178 13688 19184
rect 14096 18828 14148 18834
rect 14096 18770 14148 18776
rect 14004 18760 14056 18766
rect 14004 18702 14056 18708
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13924 18426 13952 18566
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 13910 18184 13966 18193
rect 13910 18119 13966 18128
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13464 17066 13492 17478
rect 13452 17060 13504 17066
rect 13452 17002 13504 17008
rect 13924 16590 13952 18119
rect 14016 17882 14044 18702
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 13912 16584 13964 16590
rect 13832 16544 13912 16572
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13450 16144 13506 16153
rect 13556 16114 13584 16390
rect 13450 16079 13506 16088
rect 13544 16108 13596 16114
rect 13464 16046 13492 16079
rect 13544 16050 13596 16056
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 13556 15502 13584 15914
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 13372 15320 13584 15348
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12808 13728 12860 13734
rect 12806 13696 12808 13705
rect 12860 13696 12862 13705
rect 12806 13631 12862 13640
rect 12820 12889 12848 13631
rect 12912 12918 12940 14418
rect 12992 13796 13044 13802
rect 12992 13738 13044 13744
rect 13004 13530 13032 13738
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 13096 13433 13124 13670
rect 13280 13530 13308 14758
rect 13372 14074 13400 14758
rect 13464 14550 13492 14962
rect 13452 14544 13504 14550
rect 13556 14521 13584 15320
rect 13452 14486 13504 14492
rect 13542 14512 13598 14521
rect 13542 14447 13598 14456
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13268 13524 13320 13530
rect 13648 13512 13676 16390
rect 13726 16280 13782 16289
rect 13726 16215 13728 16224
rect 13780 16215 13782 16224
rect 13728 16186 13780 16192
rect 13832 14822 13860 16544
rect 13912 16526 13964 16532
rect 14004 15972 14056 15978
rect 14004 15914 14056 15920
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13820 14340 13872 14346
rect 13820 14282 13872 14288
rect 13832 13818 13860 14282
rect 13740 13802 13860 13818
rect 13728 13796 13860 13802
rect 13780 13790 13860 13796
rect 13728 13738 13780 13744
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13832 13530 13860 13670
rect 13268 13466 13320 13472
rect 13464 13484 13676 13512
rect 13820 13524 13872 13530
rect 13082 13424 13138 13433
rect 13082 13359 13138 13368
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 12900 12912 12952 12918
rect 12806 12880 12862 12889
rect 12900 12854 12952 12860
rect 13004 12850 13032 13126
rect 12806 12815 12862 12824
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13096 12714 13124 13359
rect 13266 13016 13322 13025
rect 13266 12951 13322 12960
rect 13280 12918 13308 12951
rect 13268 12912 13320 12918
rect 13268 12854 13320 12860
rect 13084 12708 13136 12714
rect 13084 12650 13136 12656
rect 13084 12232 13136 12238
rect 13280 12220 13308 12854
rect 13136 12192 13308 12220
rect 13084 12174 13136 12180
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12820 9704 12848 11834
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 12912 10810 12940 11494
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12898 10568 12954 10577
rect 12898 10503 12954 10512
rect 12912 10470 12940 10503
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 13004 10266 13032 11494
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 13096 10130 13124 10406
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 12811 9676 12848 9704
rect 12811 9636 12839 9676
rect 12811 9608 12848 9636
rect 12820 9024 12848 9608
rect 13188 9081 13216 11018
rect 13174 9072 13230 9081
rect 12820 8996 12940 9024
rect 13174 9007 13230 9016
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12636 7002 12664 7958
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12636 5778 12664 6598
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12544 5630 12664 5658
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 12544 5166 12572 5510
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12452 4146 12480 4966
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12636 4078 12664 5630
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12452 2990 12480 3470
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12532 2848 12584 2854
rect 12532 2790 12584 2796
rect 12348 1420 12400 1426
rect 12348 1362 12400 1368
rect 12544 800 12572 2790
rect 12728 2582 12756 8774
rect 12820 8430 12848 8842
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12912 8276 12940 8996
rect 13176 8356 13228 8362
rect 13176 8298 13228 8304
rect 12820 8248 12940 8276
rect 12820 6236 12848 8248
rect 13188 8022 13216 8298
rect 13176 8016 13228 8022
rect 13176 7958 13228 7964
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12912 7478 12940 7890
rect 13176 7880 13228 7886
rect 13280 7857 13308 11290
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13372 9994 13400 10610
rect 13464 10577 13492 13484
rect 13820 13466 13872 13472
rect 13924 13410 13952 15642
rect 14016 14958 14044 15914
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13832 13382 13952 13410
rect 13450 10568 13506 10577
rect 13450 10503 13506 10512
rect 13556 10470 13584 13330
rect 13728 13252 13780 13258
rect 13728 13194 13780 13200
rect 13740 11898 13768 13194
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13648 10606 13676 11494
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13740 11150 13768 11290
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13360 9988 13412 9994
rect 13360 9930 13412 9936
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13176 7822 13228 7828
rect 13266 7848 13322 7857
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12912 6390 12940 7414
rect 13004 7342 13032 7686
rect 13096 7410 13124 7686
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 12992 6928 13044 6934
rect 12992 6870 13044 6876
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 13004 6322 13032 6870
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 12820 6208 12940 6236
rect 12912 5914 12940 6208
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 12808 5840 12860 5846
rect 13096 5794 13124 6938
rect 12808 5782 12860 5788
rect 12820 4078 12848 5782
rect 13004 5766 13124 5794
rect 13004 5302 13032 5766
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 12992 5296 13044 5302
rect 12992 5238 13044 5244
rect 13096 5234 13124 5646
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 13004 4758 13032 5102
rect 13188 4758 13216 7822
rect 13266 7783 13322 7792
rect 13280 7478 13308 7783
rect 13268 7472 13320 7478
rect 13268 7414 13320 7420
rect 13268 7268 13320 7274
rect 13268 7210 13320 7216
rect 13280 6458 13308 7210
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 13280 5166 13308 6258
rect 13268 5160 13320 5166
rect 13268 5102 13320 5108
rect 12992 4752 13044 4758
rect 12992 4694 13044 4700
rect 13176 4752 13228 4758
rect 13176 4694 13228 4700
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 13280 4282 13308 4422
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 13084 4004 13136 4010
rect 13084 3946 13136 3952
rect 13268 4004 13320 4010
rect 13268 3946 13320 3952
rect 13096 3534 13124 3946
rect 13280 3670 13308 3946
rect 13268 3664 13320 3670
rect 13268 3606 13320 3612
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12912 2990 12940 3334
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 13096 2922 13216 2938
rect 13084 2916 13216 2922
rect 13136 2910 13216 2916
rect 13084 2858 13136 2864
rect 13188 2582 13216 2910
rect 12716 2576 12768 2582
rect 12716 2518 12768 2524
rect 13176 2576 13228 2582
rect 13176 2518 13228 2524
rect 13280 1714 13308 3130
rect 13096 1686 13308 1714
rect 13096 800 13124 1686
rect 13372 1601 13400 8910
rect 13464 7834 13492 8978
rect 13556 7954 13584 10066
rect 13648 8362 13676 10406
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13740 8634 13768 9522
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13832 8294 13860 13382
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13924 8090 13952 12378
rect 14016 12102 14044 14758
rect 14108 13462 14136 18770
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14200 17202 14228 18022
rect 14292 17241 14320 19246
rect 14278 17232 14334 17241
rect 14188 17196 14240 17202
rect 14278 17167 14334 17176
rect 14188 17138 14240 17144
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14200 15366 14228 16594
rect 14292 16522 14320 16934
rect 14280 16516 14332 16522
rect 14280 16458 14332 16464
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14200 14618 14228 15302
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14096 13456 14148 13462
rect 14096 13398 14148 13404
rect 14200 13326 14228 13874
rect 14292 13394 14320 15506
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14278 13288 14334 13297
rect 14278 13223 14334 13232
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 14016 10742 14044 11494
rect 14004 10736 14056 10742
rect 14004 10678 14056 10684
rect 14292 10010 14320 13223
rect 14016 9982 14320 10010
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13464 7806 13860 7834
rect 13544 7472 13596 7478
rect 13544 7414 13596 7420
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13464 5234 13492 7278
rect 13556 5778 13584 7414
rect 13832 7154 13860 7806
rect 13912 7812 13964 7818
rect 13912 7754 13964 7760
rect 13924 7342 13952 7754
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 13832 7126 13952 7154
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13648 6186 13676 6734
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13740 6186 13768 6598
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13452 5228 13504 5234
rect 13452 5170 13504 5176
rect 13556 5098 13584 5510
rect 13544 5092 13596 5098
rect 13544 5034 13596 5040
rect 13728 5092 13780 5098
rect 13728 5034 13780 5040
rect 13740 4622 13768 5034
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13452 4480 13504 4486
rect 13452 4422 13504 4428
rect 13464 4078 13492 4422
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13832 3754 13860 6394
rect 13924 6066 13952 7126
rect 14016 6361 14044 9982
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14108 8974 14136 9318
rect 14200 9178 14228 9862
rect 14280 9444 14332 9450
rect 14280 9386 14332 9392
rect 14292 9178 14320 9386
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14280 9172 14332 9178
rect 14280 9114 14332 9120
rect 14384 9058 14412 19246
rect 14476 15706 14504 19858
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 15304 18970 15332 22000
rect 15856 20058 15884 22000
rect 15844 20052 15896 20058
rect 15844 19994 15896 20000
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 15384 18896 15436 18902
rect 15384 18838 15436 18844
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 15200 18216 15252 18222
rect 15200 18158 15252 18164
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14568 17270 14596 17818
rect 14556 17264 14608 17270
rect 14556 17206 14608 17212
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14476 12986 14504 13670
rect 14568 13297 14596 17206
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 15106 16688 15162 16697
rect 15106 16623 15162 16632
rect 14924 16584 14976 16590
rect 14924 16526 14976 16532
rect 14936 16114 14964 16526
rect 15120 16182 15148 16623
rect 15108 16176 15160 16182
rect 15108 16118 15160 16124
rect 14924 16108 14976 16114
rect 14924 16050 14976 16056
rect 14936 15978 14964 16050
rect 14924 15972 14976 15978
rect 14924 15914 14976 15920
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 14648 15428 14700 15434
rect 14648 15370 14700 15376
rect 14660 14958 14688 15370
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 15028 14890 15056 15302
rect 15016 14884 15068 14890
rect 15016 14826 15068 14832
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 15028 14414 15056 14826
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 14752 14074 14780 14350
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 15120 13938 15148 14758
rect 15212 14396 15240 18158
rect 15304 18086 15332 18770
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 15304 14550 15332 16390
rect 15396 15473 15424 18838
rect 15488 17338 15516 19858
rect 15844 18828 15896 18834
rect 15844 18770 15896 18776
rect 15856 18426 15884 18770
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 15856 18290 15884 18362
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15750 17776 15806 17785
rect 15660 17740 15712 17746
rect 15750 17711 15752 17720
rect 15660 17682 15712 17688
rect 15804 17711 15806 17720
rect 15752 17682 15804 17688
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 15672 16776 15700 17682
rect 15764 16946 15792 17682
rect 15856 17678 15884 18226
rect 16040 18222 16068 19858
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 15936 18080 15988 18086
rect 15936 18022 15988 18028
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 15844 17672 15896 17678
rect 15948 17660 15976 18022
rect 16028 17672 16080 17678
rect 15948 17632 16028 17660
rect 15844 17614 15896 17620
rect 16028 17614 16080 17620
rect 16132 17134 16160 18022
rect 16224 17882 16252 18022
rect 16212 17876 16264 17882
rect 16212 17818 16264 17824
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 16224 17202 16252 17478
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 15764 16918 15976 16946
rect 15672 16748 15792 16776
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 15488 15910 15516 16526
rect 15672 16250 15700 16594
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15488 15638 15516 15846
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 15382 15464 15438 15473
rect 15382 15399 15438 15408
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15396 14958 15424 15302
rect 15488 15026 15516 15574
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15672 14618 15700 14758
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15292 14544 15344 14550
rect 15292 14486 15344 14492
rect 15212 14368 15332 14396
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15016 13796 15068 13802
rect 15016 13738 15068 13744
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 14924 13320 14976 13326
rect 14554 13288 14610 13297
rect 14924 13262 14976 13268
rect 14554 13223 14610 13232
rect 14646 13016 14702 13025
rect 14464 12980 14516 12986
rect 14646 12951 14702 12960
rect 14464 12922 14516 12928
rect 14660 12918 14688 12951
rect 14648 12912 14700 12918
rect 14936 12866 14964 13262
rect 15028 13138 15056 13738
rect 15108 13728 15160 13734
rect 15108 13670 15160 13676
rect 15120 13530 15148 13670
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15028 13110 15148 13138
rect 14648 12854 14700 12860
rect 14844 12838 15056 12866
rect 14844 12730 14872 12838
rect 14752 12714 14872 12730
rect 14740 12708 14872 12714
rect 14792 12702 14872 12708
rect 14740 12650 14792 12656
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14568 12442 14596 12582
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14556 12436 14608 12442
rect 14556 12378 14608 12384
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 14554 11792 14610 11801
rect 14936 11762 14964 12242
rect 15028 12170 15056 12838
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 14554 11727 14610 11736
rect 14924 11756 14976 11762
rect 14568 11234 14596 11727
rect 14924 11698 14976 11704
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 14568 11206 14688 11234
rect 14660 10606 14688 11206
rect 15028 11082 15056 12106
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 15028 10674 15056 11018
rect 15120 10810 15148 13110
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15212 12442 15240 12718
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15198 11384 15254 11393
rect 15198 11319 15200 11328
rect 15252 11319 15254 11328
rect 15200 11290 15252 11296
rect 15304 11234 15332 14368
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 15672 14226 15700 14282
rect 15396 14198 15700 14226
rect 15396 13818 15424 14198
rect 15764 14056 15792 16748
rect 15842 16280 15898 16289
rect 15842 16215 15844 16224
rect 15896 16215 15898 16224
rect 15844 16186 15896 16192
rect 15488 14028 15792 14056
rect 15488 13938 15516 14028
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15568 13864 15620 13870
rect 15396 13790 15516 13818
rect 15568 13806 15620 13812
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15396 12345 15424 13330
rect 15382 12336 15438 12345
rect 15382 12271 15438 12280
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15212 11206 15332 11234
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 14476 10146 14504 10542
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 14922 10160 14978 10169
rect 14476 10118 14688 10146
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14476 9518 14504 9998
rect 14464 9512 14516 9518
rect 14660 9466 14688 10118
rect 14922 10095 14978 10104
rect 14936 9489 14964 10095
rect 14464 9454 14516 9460
rect 14568 9438 14688 9466
rect 14922 9480 14978 9489
rect 14568 9058 14596 9438
rect 14922 9415 14978 9424
rect 15120 9330 15148 10610
rect 15028 9302 15148 9330
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 14292 9030 14412 9058
rect 14476 9030 14596 9058
rect 14738 9072 14794 9081
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 14108 8430 14136 8910
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14002 6352 14058 6361
rect 14002 6287 14058 6296
rect 13924 6038 14044 6066
rect 14016 5710 14044 6038
rect 14004 5704 14056 5710
rect 14056 5652 14228 5658
rect 14004 5646 14228 5652
rect 14016 5630 14228 5646
rect 14200 4826 14228 5630
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 14016 4146 14044 4626
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 13912 3936 13964 3942
rect 13912 3878 13964 3884
rect 13464 3726 13860 3754
rect 13464 3602 13492 3726
rect 13452 3596 13504 3602
rect 13452 3538 13504 3544
rect 13636 3528 13688 3534
rect 13688 3476 13860 3482
rect 13636 3470 13860 3476
rect 13648 3466 13860 3470
rect 13648 3460 13872 3466
rect 13648 3454 13820 3460
rect 13820 3402 13872 3408
rect 13924 3346 13952 3878
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 13556 3318 13952 3346
rect 13358 1592 13414 1601
rect 13358 1527 13414 1536
rect 13556 1442 13584 3318
rect 14016 2990 14044 3470
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 14292 2666 14320 9030
rect 14476 8378 14504 9030
rect 14738 9007 14740 9016
rect 14792 9007 14794 9016
rect 14740 8978 14792 8984
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 14568 8430 14596 8842
rect 14384 8350 14504 8378
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14384 6730 14412 8350
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 14476 7886 14504 8230
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14476 6798 14504 7822
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14372 6724 14424 6730
rect 14372 6666 14424 6672
rect 14568 4690 14596 8026
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 15028 6866 15056 9302
rect 15212 9194 15240 11206
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15304 10810 15332 10950
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15396 10724 15424 12038
rect 15488 10826 15516 13790
rect 15580 11354 15608 13806
rect 15672 12782 15700 13874
rect 15764 13734 15792 14028
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 15856 13274 15884 13806
rect 15764 13246 15884 13274
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15764 12442 15792 13246
rect 15948 13172 15976 16918
rect 16040 14618 16068 17070
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16224 15502 16252 16050
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16316 14890 16344 19246
rect 16408 19174 16436 22000
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 16856 19916 16908 19922
rect 16856 19858 16908 19864
rect 16488 19304 16540 19310
rect 16488 19246 16540 19252
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16408 16998 16436 17682
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16408 16561 16436 16594
rect 16394 16552 16450 16561
rect 16394 16487 16450 16496
rect 16304 14884 16356 14890
rect 16304 14826 16356 14832
rect 16028 14612 16080 14618
rect 16028 14554 16080 14560
rect 16316 14498 16344 14826
rect 16224 14470 16344 14498
rect 16224 14414 16252 14470
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16120 14340 16172 14346
rect 16120 14282 16172 14288
rect 16132 14006 16160 14282
rect 16120 14000 16172 14006
rect 16120 13942 16172 13948
rect 16304 13796 16356 13802
rect 16304 13738 16356 13744
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 16028 13252 16080 13258
rect 16028 13194 16080 13200
rect 15856 13144 15976 13172
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15764 11762 15792 12378
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15488 10798 15608 10826
rect 15396 10696 15516 10724
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15396 10266 15424 10542
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15120 9178 15240 9194
rect 15304 9178 15332 10066
rect 15396 9722 15424 10066
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15384 9444 15436 9450
rect 15384 9386 15436 9392
rect 15396 9178 15424 9386
rect 15108 9172 15240 9178
rect 15160 9166 15240 9172
rect 15292 9172 15344 9178
rect 15108 9114 15160 9120
rect 15292 9114 15344 9120
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15198 9072 15254 9081
rect 15198 9007 15254 9016
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15120 8090 15148 8910
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 15028 5794 15056 6258
rect 15120 5914 15148 8026
rect 15212 7954 15240 9007
rect 15488 8974 15516 10696
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15200 7948 15252 7954
rect 15200 7890 15252 7896
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15304 6730 15332 7142
rect 15580 6798 15608 10798
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15672 10130 15700 10406
rect 15764 10198 15792 11086
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15856 10044 15884 13144
rect 15934 13016 15990 13025
rect 15934 12951 15990 12960
rect 15948 12782 15976 12951
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 15948 10810 15976 12718
rect 16040 11694 16068 13194
rect 16132 12209 16160 13466
rect 16118 12200 16174 12209
rect 16118 12135 16174 12144
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 16132 11626 16160 12038
rect 16120 11620 16172 11626
rect 16120 11562 16172 11568
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 15936 10804 15988 10810
rect 15936 10746 15988 10752
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 16040 10198 16068 10474
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 15764 10016 15884 10044
rect 15936 10056 15988 10062
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15672 8922 15700 8978
rect 15764 8922 15792 10016
rect 16132 10010 16160 11290
rect 15936 9998 15988 10004
rect 15948 9178 15976 9998
rect 16040 9994 16160 10010
rect 16028 9988 16160 9994
rect 16080 9982 16160 9988
rect 16028 9930 16080 9936
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15844 9036 15896 9042
rect 15844 8978 15896 8984
rect 15672 8894 15792 8922
rect 15660 8832 15712 8838
rect 15660 8774 15712 8780
rect 15672 8498 15700 8774
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15672 7954 15700 8434
rect 15764 8294 15792 8894
rect 15856 8634 15884 8978
rect 15948 8974 15976 9114
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 15948 8634 15976 8910
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 15934 8528 15990 8537
rect 15934 8463 15990 8472
rect 15752 8288 15804 8294
rect 15752 8230 15804 8236
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 15672 7206 15700 7890
rect 15856 7410 15884 7890
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15764 7002 15792 7142
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 15948 6882 15976 8463
rect 16040 7154 16068 9930
rect 16224 9602 16252 13670
rect 16316 13394 16344 13738
rect 16408 13530 16436 16487
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16316 13025 16344 13330
rect 16396 13252 16448 13258
rect 16396 13194 16448 13200
rect 16302 13016 16358 13025
rect 16408 12986 16436 13194
rect 16302 12951 16358 12960
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16500 12345 16528 19246
rect 16592 17338 16620 19858
rect 16764 19304 16816 19310
rect 16868 19281 16896 19858
rect 16764 19246 16816 19252
rect 16854 19272 16910 19281
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 16684 17814 16712 18566
rect 16672 17808 16724 17814
rect 16672 17750 16724 17756
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16684 17202 16712 17750
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16580 15904 16632 15910
rect 16580 15846 16632 15852
rect 16592 14958 16620 15846
rect 16672 15700 16724 15706
rect 16672 15642 16724 15648
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16684 14822 16712 15642
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16672 13796 16724 13802
rect 16672 13738 16724 13744
rect 16486 12336 16542 12345
rect 16486 12271 16542 12280
rect 16684 12238 16712 13738
rect 16776 12374 16804 19246
rect 16854 19207 16910 19216
rect 16960 19174 16988 22000
rect 17512 20058 17540 22000
rect 17866 20632 17922 20641
rect 17866 20567 17922 20576
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 17132 19712 17184 19718
rect 17132 19654 17184 19660
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16854 18864 16910 18873
rect 16854 18799 16910 18808
rect 16868 18630 16896 18799
rect 16856 18624 16908 18630
rect 16856 18566 16908 18572
rect 17038 17776 17094 17785
rect 17038 17711 17094 17720
rect 17052 16658 17080 17711
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 16854 16144 16910 16153
rect 16854 16079 16910 16088
rect 16868 15978 16896 16079
rect 16856 15972 16908 15978
rect 16856 15914 16908 15920
rect 16868 15745 16896 15914
rect 16854 15736 16910 15745
rect 16854 15671 16910 15680
rect 16948 15632 17000 15638
rect 16948 15574 17000 15580
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16868 14278 16896 14894
rect 16960 14822 16988 15574
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 16856 13184 16908 13190
rect 16856 13126 16908 13132
rect 16868 12442 16896 13126
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 16764 12368 16816 12374
rect 16764 12310 16816 12316
rect 16488 12232 16540 12238
rect 16394 12200 16450 12209
rect 16488 12174 16540 12180
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16394 12135 16450 12144
rect 16408 11370 16436 12135
rect 16500 11529 16528 12174
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 16486 11520 16542 11529
rect 16486 11455 16542 11464
rect 16408 11342 16528 11370
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 16316 10606 16344 11086
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 16394 10568 16450 10577
rect 16132 9574 16252 9602
rect 16132 8650 16160 9574
rect 16316 9466 16344 10542
rect 16394 10503 16450 10512
rect 16224 9438 16344 9466
rect 16224 8838 16252 9438
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16316 9110 16344 9318
rect 16408 9217 16436 10503
rect 16394 9208 16450 9217
rect 16394 9143 16450 9152
rect 16304 9104 16356 9110
rect 16304 9046 16356 9052
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16132 8622 16252 8650
rect 16120 7948 16172 7954
rect 16120 7890 16172 7896
rect 16132 7342 16160 7890
rect 16120 7336 16172 7342
rect 16120 7278 16172 7284
rect 16040 7126 16160 7154
rect 15672 6854 15976 6882
rect 15568 6792 15620 6798
rect 15568 6734 15620 6740
rect 15292 6724 15344 6730
rect 15292 6666 15344 6672
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15028 5766 15332 5794
rect 15396 5778 15424 6258
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15212 5166 15240 5646
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 15212 4690 15240 5102
rect 14556 4684 14608 4690
rect 15200 4684 15252 4690
rect 14556 4626 14608 4632
rect 15120 4644 15200 4672
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14200 2650 14320 2666
rect 14384 2650 14412 4014
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14476 2650 14504 3334
rect 14660 3194 14688 3334
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 15120 2922 15148 4644
rect 15200 4626 15252 4632
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 14556 2916 14608 2922
rect 14556 2858 14608 2864
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 14188 2644 14320 2650
rect 14240 2638 14320 2644
rect 14372 2644 14424 2650
rect 14188 2586 14240 2592
rect 14372 2586 14424 2592
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 14568 2446 14596 2858
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14648 2372 14700 2378
rect 14648 2314 14700 2320
rect 14740 2372 14792 2378
rect 14740 2314 14792 2320
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 13556 1414 13676 1442
rect 13648 800 13676 1414
rect 14200 800 14228 2246
rect 14660 1970 14688 2314
rect 14648 1964 14700 1970
rect 14648 1906 14700 1912
rect 14752 800 14780 2314
rect 15212 1442 15240 4422
rect 15304 3942 15332 5766
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15488 4146 15516 6598
rect 15580 5914 15608 6734
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15672 5794 15700 6854
rect 15936 6724 15988 6730
rect 15936 6666 15988 6672
rect 15752 6384 15804 6390
rect 15752 6326 15804 6332
rect 15580 5766 15700 5794
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15580 2961 15608 5766
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15672 4146 15700 5510
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 15566 2952 15622 2961
rect 15566 2887 15622 2896
rect 15764 2514 15792 6326
rect 15948 6254 15976 6666
rect 15936 6248 15988 6254
rect 15936 6190 15988 6196
rect 16132 6186 16160 7126
rect 16028 6180 16080 6186
rect 16028 6122 16080 6128
rect 16120 6180 16172 6186
rect 16120 6122 16172 6128
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15856 5817 15884 5850
rect 15842 5808 15898 5817
rect 15842 5743 15898 5752
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15856 5574 15884 5646
rect 15844 5568 15896 5574
rect 15844 5510 15896 5516
rect 15844 4004 15896 4010
rect 15844 3946 15896 3952
rect 15752 2508 15804 2514
rect 15752 2450 15804 2456
rect 15212 1414 15332 1442
rect 15304 800 15332 1414
rect 15856 800 15884 3946
rect 16040 3942 16068 6122
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 16132 5234 16160 5646
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 16224 5114 16252 8622
rect 16132 5086 16252 5114
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 16132 3670 16160 5086
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 16040 3194 16068 3470
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 16028 2440 16080 2446
rect 16026 2408 16028 2417
rect 16080 2408 16082 2417
rect 16026 2343 16082 2352
rect 16132 2038 16160 3606
rect 16316 2106 16344 8910
rect 16408 5778 16436 8978
rect 16500 8974 16528 11342
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 16500 8265 16528 8298
rect 16486 8256 16542 8265
rect 16486 8191 16542 8200
rect 16592 6390 16620 9862
rect 16684 6390 16712 11834
rect 16776 10418 16804 12310
rect 16960 12306 16988 14758
rect 17144 14482 17172 19654
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17236 18902 17264 19246
rect 17880 19242 17908 20567
rect 18064 20058 18092 22000
rect 18510 21176 18566 21185
rect 18510 21111 18566 21120
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 17868 19236 17920 19242
rect 17868 19178 17920 19184
rect 17224 18896 17276 18902
rect 17224 18838 17276 18844
rect 17684 18828 17736 18834
rect 17684 18770 17736 18776
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17590 18728 17646 18737
rect 17224 16108 17276 16114
rect 17224 16050 17276 16056
rect 17236 15706 17264 16050
rect 17328 16017 17356 18702
rect 17590 18663 17646 18672
rect 17498 17640 17554 17649
rect 17498 17575 17500 17584
rect 17552 17575 17554 17584
rect 17500 17546 17552 17552
rect 17512 16590 17540 17546
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17314 16008 17370 16017
rect 17314 15943 17370 15952
rect 17328 15910 17356 15943
rect 17512 15910 17540 16526
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17500 15904 17552 15910
rect 17500 15846 17552 15852
rect 17224 15700 17276 15706
rect 17224 15642 17276 15648
rect 17222 15464 17278 15473
rect 17222 15399 17278 15408
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 17052 12374 17080 14214
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 17040 12368 17092 12374
rect 17040 12310 17092 12316
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 17144 12220 17172 12582
rect 16946 12200 17002 12209
rect 16946 12135 17002 12144
rect 17052 12192 17172 12220
rect 16776 10390 16896 10418
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 16776 9450 16804 10202
rect 16868 10130 16896 10390
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 16764 9444 16816 9450
rect 16764 9386 16816 9392
rect 16868 7562 16896 9930
rect 16776 7534 16896 7562
rect 16776 7002 16804 7534
rect 16856 7268 16908 7274
rect 16856 7210 16908 7216
rect 16764 6996 16816 7002
rect 16764 6938 16816 6944
rect 16868 6798 16896 7210
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16580 6384 16632 6390
rect 16580 6326 16632 6332
rect 16672 6384 16724 6390
rect 16672 6326 16724 6332
rect 16592 6168 16620 6326
rect 16500 6140 16620 6168
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 16500 5114 16528 6140
rect 16684 6100 16712 6326
rect 16592 6072 16712 6100
rect 16592 5778 16620 6072
rect 16672 5840 16724 5846
rect 16672 5782 16724 5788
rect 16762 5808 16818 5817
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 16408 5086 16528 5114
rect 16408 4146 16436 5086
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16500 4758 16528 4966
rect 16488 4752 16540 4758
rect 16488 4694 16540 4700
rect 16500 4214 16528 4694
rect 16488 4208 16540 4214
rect 16488 4150 16540 4156
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16592 4078 16620 4966
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16580 3936 16632 3942
rect 16684 3890 16712 5782
rect 16762 5743 16818 5752
rect 16776 5370 16804 5743
rect 16856 5636 16908 5642
rect 16856 5578 16908 5584
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 16632 3884 16712 3890
rect 16580 3878 16712 3884
rect 16592 3862 16712 3878
rect 16776 3602 16804 4626
rect 16868 4078 16896 5578
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 16960 3738 16988 12135
rect 17052 6798 17080 12192
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17144 11286 17172 11494
rect 17132 11280 17184 11286
rect 17132 11222 17184 11228
rect 17236 9058 17264 15399
rect 17328 14793 17356 15846
rect 17500 15564 17552 15570
rect 17500 15506 17552 15512
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17314 14784 17370 14793
rect 17314 14719 17370 14728
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17328 12646 17356 13670
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17420 12424 17448 14894
rect 17512 13734 17540 15506
rect 17604 14056 17632 18663
rect 17696 15586 17724 18770
rect 17972 18698 18000 19654
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 18524 19174 18552 21111
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 17960 18692 18012 18698
rect 17960 18634 18012 18640
rect 18512 18692 18564 18698
rect 18512 18634 18564 18640
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 17960 18080 18012 18086
rect 17960 18022 18012 18028
rect 18144 18080 18196 18086
rect 18144 18022 18196 18028
rect 17868 17672 17920 17678
rect 17866 17640 17868 17649
rect 17920 17640 17922 17649
rect 17866 17575 17922 17584
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 17788 17202 17816 17478
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 17788 16658 17816 17138
rect 17776 16652 17828 16658
rect 17776 16594 17828 16600
rect 17776 16040 17828 16046
rect 17776 15982 17828 15988
rect 17788 15722 17816 15982
rect 17880 15978 17908 17138
rect 17972 17134 18000 18022
rect 18156 17785 18184 18022
rect 18142 17776 18198 17785
rect 18142 17711 18198 17720
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 18418 17096 18474 17105
rect 18418 17031 18474 17040
rect 18432 16998 18460 17031
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18524 16794 18552 18634
rect 18616 18426 18644 22000
rect 18696 19916 18748 19922
rect 18696 19858 18748 19864
rect 18708 18902 18736 19858
rect 18800 18970 18828 22063
rect 19154 22000 19210 22800
rect 19246 22536 19302 22545
rect 19246 22471 19302 22480
rect 19062 21584 19118 21593
rect 19062 21519 19118 21528
rect 19076 20058 19104 21519
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 19064 20052 19116 20058
rect 19064 19994 19116 20000
rect 18892 19938 18920 19994
rect 19168 19990 19196 22000
rect 19156 19984 19208 19990
rect 18892 19910 19104 19938
rect 19156 19926 19208 19932
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18788 18964 18840 18970
rect 18788 18906 18840 18912
rect 18696 18896 18748 18902
rect 18696 18838 18748 18844
rect 18788 18828 18840 18834
rect 18788 18770 18840 18776
rect 18604 18420 18656 18426
rect 18604 18362 18656 18368
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18616 17814 18644 18226
rect 18604 17808 18656 17814
rect 18604 17750 18656 17756
rect 18616 17184 18644 17750
rect 18696 17196 18748 17202
rect 18616 17156 18696 17184
rect 18696 17138 18748 17144
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18512 16584 18564 16590
rect 18510 16552 18512 16561
rect 18564 16552 18566 16561
rect 18510 16487 18566 16496
rect 18616 16454 18644 16730
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 17868 15972 17920 15978
rect 17868 15914 17920 15920
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 18236 15904 18288 15910
rect 18236 15846 18288 15852
rect 17788 15694 17908 15722
rect 17880 15638 17908 15694
rect 17868 15632 17920 15638
rect 17696 15558 17816 15586
rect 17868 15574 17920 15580
rect 17604 14028 17724 14056
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17328 12396 17448 12424
rect 17328 11121 17356 12396
rect 17406 12336 17462 12345
rect 17406 12271 17462 12280
rect 17314 11112 17370 11121
rect 17314 11047 17370 11056
rect 17420 9450 17448 12271
rect 17512 12238 17540 13670
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17604 12102 17632 13874
rect 17696 13326 17724 14028
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17696 12714 17724 13262
rect 17684 12708 17736 12714
rect 17684 12650 17736 12656
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17500 11280 17552 11286
rect 17500 11222 17552 11228
rect 17512 10062 17540 11222
rect 17590 11112 17646 11121
rect 17590 11047 17592 11056
rect 17644 11047 17646 11056
rect 17592 11018 17644 11024
rect 17696 11014 17724 12242
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17512 9586 17540 9998
rect 17604 9994 17632 10406
rect 17592 9988 17644 9994
rect 17592 9930 17644 9936
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17236 9030 17356 9058
rect 17224 8900 17276 8906
rect 17224 8842 17276 8848
rect 17130 8256 17186 8265
rect 17130 8191 17186 8200
rect 17144 7750 17172 8191
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 17052 6662 17080 6734
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 17144 6322 17172 7686
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 17040 5704 17092 5710
rect 17040 5646 17092 5652
rect 17052 4758 17080 5646
rect 17040 4752 17092 4758
rect 17040 4694 17092 4700
rect 17052 4554 17080 4694
rect 17040 4548 17092 4554
rect 17040 4490 17092 4496
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 16960 2650 16988 3334
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 17236 2514 17264 8842
rect 17328 7274 17356 9030
rect 17408 8356 17460 8362
rect 17408 8298 17460 8304
rect 17316 7268 17368 7274
rect 17316 7210 17368 7216
rect 17328 7002 17356 7210
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 17328 6322 17356 6598
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17420 4690 17448 8298
rect 17604 7954 17632 9318
rect 17696 9110 17724 10406
rect 17684 9104 17736 9110
rect 17684 9046 17736 9052
rect 17592 7948 17644 7954
rect 17592 7890 17644 7896
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17590 7440 17646 7449
rect 17590 7375 17646 7384
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17512 6322 17540 7142
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17604 6225 17632 7375
rect 17696 6254 17724 7686
rect 17684 6248 17736 6254
rect 17590 6216 17646 6225
rect 17684 6190 17736 6196
rect 17590 6151 17646 6160
rect 17604 5166 17632 6151
rect 17592 5160 17644 5166
rect 17592 5102 17644 5108
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17592 3596 17644 3602
rect 17592 3538 17644 3544
rect 17604 3194 17632 3538
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17604 3074 17632 3130
rect 17512 3046 17632 3074
rect 17512 2530 17540 3046
rect 17696 2938 17724 3878
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 17420 2502 17540 2530
rect 17604 2910 17724 2938
rect 17420 2446 17448 2502
rect 17040 2440 17092 2446
rect 17040 2382 17092 2388
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 16304 2100 16356 2106
rect 16304 2042 16356 2048
rect 16120 2032 16172 2038
rect 16120 1974 16172 1980
rect 16396 1216 16448 1222
rect 16396 1158 16448 1164
rect 16408 800 16436 1158
rect 16960 800 16988 2246
rect 17052 2106 17080 2382
rect 17040 2100 17092 2106
rect 17040 2042 17092 2048
rect 17604 1034 17632 2910
rect 17788 2582 17816 15558
rect 17972 15502 18000 15846
rect 18248 15609 18276 15846
rect 18050 15600 18106 15609
rect 18234 15600 18290 15609
rect 18144 15564 18196 15570
rect 18106 15544 18144 15552
rect 18050 15535 18144 15544
rect 18064 15524 18144 15535
rect 18234 15535 18290 15544
rect 18144 15506 18196 15512
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17972 15366 18000 15438
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17972 14958 18000 15302
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18708 15178 18736 16594
rect 18524 15150 18736 15178
rect 18524 15094 18552 15150
rect 18512 15088 18564 15094
rect 18512 15030 18564 15036
rect 18602 15056 18658 15065
rect 18420 15020 18472 15026
rect 18602 14991 18658 15000
rect 18420 14962 18472 14968
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 18432 14482 18460 14962
rect 18512 14952 18564 14958
rect 18512 14894 18564 14900
rect 18524 14550 18552 14894
rect 18512 14544 18564 14550
rect 18512 14486 18564 14492
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 18420 14476 18472 14482
rect 18420 14418 18472 14424
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17880 13870 17908 14350
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17880 13530 17908 13806
rect 17972 13530 18000 14418
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 17866 13424 17922 13433
rect 17866 13359 17868 13368
rect 17920 13359 17922 13368
rect 17868 13330 17920 13336
rect 18156 13274 18184 13670
rect 17972 13246 18184 13274
rect 17866 12744 17922 12753
rect 17866 12679 17922 12688
rect 17880 10130 17908 12679
rect 17972 11762 18000 13246
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18524 12986 18552 14350
rect 18616 14346 18644 14991
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 18604 14340 18656 14346
rect 18604 14282 18656 14288
rect 18604 13728 18656 13734
rect 18604 13670 18656 13676
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18616 12918 18644 13670
rect 18708 13433 18736 14554
rect 18694 13424 18750 13433
rect 18694 13359 18750 13368
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18708 12986 18736 13262
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18604 12912 18656 12918
rect 18326 12880 18382 12889
rect 18604 12854 18656 12860
rect 18326 12815 18382 12824
rect 18340 12782 18368 12815
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18064 12442 18092 12718
rect 18236 12708 18288 12714
rect 18236 12650 18288 12656
rect 18248 12481 18276 12650
rect 18234 12472 18290 12481
rect 18052 12436 18104 12442
rect 18234 12407 18290 12416
rect 18052 12378 18104 12384
rect 18340 12306 18368 12718
rect 18696 12708 18748 12714
rect 18696 12650 18748 12656
rect 18512 12368 18564 12374
rect 18512 12310 18564 12316
rect 18328 12300 18380 12306
rect 18328 12242 18380 12248
rect 18052 12232 18104 12238
rect 18050 12200 18052 12209
rect 18104 12200 18106 12209
rect 18050 12135 18106 12144
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 18524 11014 18552 12310
rect 18604 12164 18656 12170
rect 18604 12106 18656 12112
rect 18616 11898 18644 12106
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18708 11286 18736 12650
rect 18696 11280 18748 11286
rect 18696 11222 18748 11228
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 17972 10606 18000 10950
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18050 10704 18106 10713
rect 18050 10639 18106 10648
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17972 9722 18000 9998
rect 18064 9994 18092 10639
rect 18512 10600 18564 10606
rect 18326 10568 18382 10577
rect 18512 10542 18564 10548
rect 18326 10503 18382 10512
rect 18340 10470 18368 10503
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18524 10062 18552 10542
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18052 9988 18104 9994
rect 18052 9930 18104 9936
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18236 9648 18288 9654
rect 18524 9602 18552 9862
rect 18236 9590 18288 9596
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 17866 8120 17922 8129
rect 17972 8090 18000 9386
rect 18156 9081 18184 9590
rect 18248 9110 18276 9590
rect 18515 9574 18552 9602
rect 18328 9512 18380 9518
rect 18515 9500 18543 9574
rect 18328 9454 18380 9460
rect 18418 9480 18474 9489
rect 18236 9104 18288 9110
rect 18142 9072 18198 9081
rect 18236 9046 18288 9052
rect 18340 9042 18368 9454
rect 18515 9472 18552 9500
rect 18418 9415 18420 9424
rect 18472 9415 18474 9424
rect 18420 9386 18472 9392
rect 18142 9007 18198 9016
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 18050 8528 18106 8537
rect 18524 8498 18552 9472
rect 18616 8634 18644 11154
rect 18696 11008 18748 11014
rect 18696 10950 18748 10956
rect 18708 9636 18736 10950
rect 18800 9654 18828 18770
rect 18984 18193 19012 19246
rect 18970 18184 19026 18193
rect 18880 18148 18932 18154
rect 18970 18119 19026 18128
rect 18880 18090 18932 18096
rect 18892 12714 18920 18090
rect 19076 16538 19104 19910
rect 19154 19816 19210 19825
rect 19154 19751 19210 19760
rect 19168 19514 19196 19751
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 19260 19310 19288 22471
rect 19706 22000 19762 22800
rect 20258 22000 20314 22800
rect 20810 22000 20866 22800
rect 21362 22000 21418 22800
rect 21914 22000 21970 22800
rect 22466 22000 22522 22800
rect 19614 20224 19670 20233
rect 19614 20159 19670 20168
rect 19628 20058 19656 20159
rect 19616 20052 19668 20058
rect 19616 19994 19668 20000
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 19444 18902 19472 19858
rect 19720 19786 19748 22000
rect 19708 19780 19760 19786
rect 19708 19722 19760 19728
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 19890 19272 19946 19281
rect 19708 19236 19760 19242
rect 19890 19207 19946 19216
rect 19708 19178 19760 19184
rect 19432 18896 19484 18902
rect 19432 18838 19484 18844
rect 19156 18760 19208 18766
rect 19156 18702 19208 18708
rect 19168 18222 19196 18702
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19156 18216 19208 18222
rect 19156 18158 19208 18164
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19156 17740 19208 17746
rect 19156 17682 19208 17688
rect 19168 17338 19196 17682
rect 19260 17377 19288 18022
rect 19444 17814 19472 18158
rect 19432 17808 19484 17814
rect 19432 17750 19484 17756
rect 19246 17368 19302 17377
rect 19156 17332 19208 17338
rect 19246 17303 19302 17312
rect 19156 17274 19208 17280
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 19444 16561 19472 16934
rect 19430 16552 19486 16561
rect 19076 16510 19380 16538
rect 19064 16448 19116 16454
rect 19248 16448 19300 16454
rect 19116 16396 19196 16402
rect 19064 16390 19196 16396
rect 19248 16390 19300 16396
rect 19076 16374 19196 16390
rect 19168 16114 19196 16374
rect 19156 16108 19208 16114
rect 19156 16050 19208 16056
rect 18972 15904 19024 15910
rect 18972 15846 19024 15852
rect 18880 12708 18932 12714
rect 18880 12650 18932 12656
rect 18984 12442 19012 15846
rect 19168 15638 19196 16050
rect 19260 16046 19288 16390
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 19156 15632 19208 15638
rect 19156 15574 19208 15580
rect 19352 15570 19380 16510
rect 19430 16487 19486 16496
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 19444 15706 19472 16050
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19062 14512 19118 14521
rect 19062 14447 19118 14456
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18892 11354 18920 12038
rect 18984 11665 19012 12378
rect 19076 11898 19104 14447
rect 19352 13530 19380 15506
rect 19444 14890 19472 15642
rect 19432 14884 19484 14890
rect 19432 14826 19484 14832
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19168 12374 19196 13330
rect 19156 12368 19208 12374
rect 19156 12310 19208 12316
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 19156 11824 19208 11830
rect 19156 11766 19208 11772
rect 18970 11656 19026 11665
rect 18970 11591 19026 11600
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 19064 11552 19116 11558
rect 19168 11529 19196 11766
rect 19352 11626 19380 13330
rect 19432 13252 19484 13258
rect 19432 13194 19484 13200
rect 19444 12306 19472 13194
rect 19536 12374 19564 18566
rect 19616 12708 19668 12714
rect 19616 12650 19668 12656
rect 19524 12368 19576 12374
rect 19524 12310 19576 12316
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19444 11762 19472 12242
rect 19628 11830 19656 12650
rect 19616 11824 19668 11830
rect 19616 11766 19668 11772
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 19064 11494 19116 11500
rect 19154 11520 19210 11529
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18892 10606 18920 11086
rect 18880 10600 18932 10606
rect 18880 10542 18932 10548
rect 18677 9608 18736 9636
rect 18788 9648 18840 9654
rect 18677 9353 18705 9608
rect 18788 9590 18840 9596
rect 18892 9586 18920 10542
rect 18984 10441 19012 11494
rect 18970 10432 19026 10441
rect 18970 10367 19026 10376
rect 19076 9976 19104 11494
rect 19154 11455 19210 11464
rect 19444 11354 19472 11698
rect 19524 11620 19576 11626
rect 19524 11562 19576 11568
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19444 10470 19472 11154
rect 19536 11014 19564 11562
rect 19616 11552 19668 11558
rect 19616 11494 19668 11500
rect 19524 11008 19576 11014
rect 19524 10950 19576 10956
rect 19432 10464 19484 10470
rect 19338 10432 19394 10441
rect 19432 10406 19484 10412
rect 19338 10367 19394 10376
rect 19076 9948 19196 9976
rect 19168 9602 19196 9948
rect 19352 9636 19380 10367
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 19076 9574 19196 9602
rect 19343 9608 19380 9636
rect 18677 9344 18750 9353
rect 18677 9302 18694 9344
rect 18694 9279 18750 9288
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18050 8463 18106 8472
rect 18512 8492 18564 8498
rect 18064 8430 18092 8463
rect 18512 8434 18564 8440
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 17866 8055 17868 8064
rect 17920 8055 17922 8064
rect 17960 8084 18012 8090
rect 17868 8026 17920 8032
rect 17960 8026 18012 8032
rect 17868 7812 17920 7818
rect 17868 7754 17920 7760
rect 17880 6798 17908 7754
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 17868 6792 17920 6798
rect 18708 6746 18736 9046
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 18880 7948 18932 7954
rect 18880 7890 18932 7896
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 17868 6734 17920 6740
rect 17880 5914 17908 6734
rect 18524 6718 18736 6746
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 18052 6180 18104 6186
rect 18052 6122 18104 6128
rect 18420 6180 18472 6186
rect 18420 6122 18472 6128
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 18064 5817 18092 6122
rect 18050 5808 18106 5817
rect 18050 5743 18106 5752
rect 18432 5642 18460 6122
rect 18420 5636 18472 5642
rect 18420 5578 18472 5584
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17880 5234 17908 5510
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 18326 5264 18382 5273
rect 17868 5228 17920 5234
rect 18326 5199 18382 5208
rect 17868 5170 17920 5176
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 18064 4593 18092 4762
rect 18050 4584 18106 4593
rect 18340 4554 18368 5199
rect 18050 4519 18106 4528
rect 18328 4548 18380 4554
rect 18328 4490 18380 4496
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 17776 2576 17828 2582
rect 17880 2553 17908 3674
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18418 2952 18474 2961
rect 18418 2887 18474 2896
rect 18432 2854 18460 2887
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 17776 2518 17828 2524
rect 17866 2544 17922 2553
rect 17866 2479 17922 2488
rect 18064 2446 18092 2790
rect 18524 2650 18552 6718
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18708 6118 18736 6598
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18616 4622 18644 6054
rect 18800 5710 18828 7278
rect 18892 6225 18920 7890
rect 18984 6934 19012 8774
rect 19076 8498 19104 9574
rect 19343 9500 19371 9608
rect 19343 9472 19380 9500
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 19260 8430 19288 9318
rect 19352 8838 19380 9472
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 19064 8356 19116 8362
rect 19064 8298 19116 8304
rect 18972 6928 19024 6934
rect 18972 6870 19024 6876
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 18878 6216 18934 6225
rect 18878 6151 18934 6160
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18696 5092 18748 5098
rect 18696 5034 18748 5040
rect 18708 4826 18736 5034
rect 18788 5024 18840 5030
rect 18788 4966 18840 4972
rect 18696 4820 18748 4826
rect 18696 4762 18748 4768
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18800 4321 18828 4966
rect 18786 4312 18842 4321
rect 18786 4247 18842 4256
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18604 3664 18656 3670
rect 18604 3606 18656 3612
rect 18616 3058 18644 3606
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18800 2990 18828 3878
rect 18892 3738 18920 5714
rect 18984 4078 19012 6598
rect 19076 6458 19104 8298
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 19154 7848 19210 7857
rect 19154 7783 19210 7792
rect 19168 7750 19196 7783
rect 19156 7744 19208 7750
rect 19156 7686 19208 7692
rect 19260 7206 19288 7958
rect 19340 7744 19392 7750
rect 19338 7712 19340 7721
rect 19392 7712 19394 7721
rect 19338 7647 19394 7656
rect 19248 7200 19300 7206
rect 19154 7168 19210 7177
rect 19248 7142 19300 7148
rect 19154 7103 19210 7112
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 19064 6248 19116 6254
rect 19064 6190 19116 6196
rect 19076 5778 19104 6190
rect 19064 5772 19116 5778
rect 19064 5714 19116 5720
rect 19168 5574 19196 7103
rect 19444 6458 19472 10406
rect 19524 9444 19576 9450
rect 19524 9386 19576 9392
rect 19536 9178 19564 9386
rect 19628 9382 19656 11494
rect 19720 11286 19748 19178
rect 19800 18828 19852 18834
rect 19800 18770 19852 18776
rect 19708 11280 19760 11286
rect 19708 11222 19760 11228
rect 19708 10056 19760 10062
rect 19708 9998 19760 10004
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 19628 8498 19656 9046
rect 19720 8634 19748 9998
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19616 7744 19668 7750
rect 19616 7686 19668 7692
rect 19628 6866 19656 7686
rect 19708 7200 19760 7206
rect 19708 7142 19760 7148
rect 19616 6860 19668 6866
rect 19616 6802 19668 6808
rect 19720 6798 19748 7142
rect 19708 6792 19760 6798
rect 19708 6734 19760 6740
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19340 6180 19392 6186
rect 19340 6122 19392 6128
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19156 5568 19208 5574
rect 19156 5510 19208 5516
rect 19064 5092 19116 5098
rect 19064 5034 19116 5040
rect 19076 4282 19104 5034
rect 19168 4758 19196 5510
rect 19156 4752 19208 4758
rect 19156 4694 19208 4700
rect 19064 4276 19116 4282
rect 19064 4218 19116 4224
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 19156 3732 19208 3738
rect 19156 3674 19208 3680
rect 18972 3664 19024 3670
rect 18972 3606 19024 3612
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 18604 2916 18656 2922
rect 18604 2858 18656 2864
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 18512 2372 18564 2378
rect 18512 2314 18564 2320
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 18052 2032 18104 2038
rect 18050 2000 18052 2009
rect 18104 2000 18106 2009
rect 18050 1935 18106 1944
rect 18524 1170 18552 2314
rect 17512 1006 17632 1034
rect 18064 1142 18552 1170
rect 17512 800 17540 1006
rect 18064 800 18092 1142
rect 18616 800 18644 2858
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 18708 1222 18736 2586
rect 18984 2106 19012 3606
rect 19064 3392 19116 3398
rect 19064 3334 19116 3340
rect 18972 2100 19024 2106
rect 18972 2042 19024 2048
rect 19076 1442 19104 3334
rect 19168 2530 19196 3674
rect 19260 2990 19288 6054
rect 19352 5574 19380 6122
rect 19812 5930 19840 18770
rect 19904 12442 19932 19207
rect 20180 18873 20208 19654
rect 20166 18864 20222 18873
rect 20166 18799 20222 18808
rect 20272 18698 20300 22000
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20260 18692 20312 18698
rect 20260 18634 20312 18640
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19996 17202 20024 18158
rect 20088 17882 20116 18158
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 19984 17196 20036 17202
rect 19984 17138 20036 17144
rect 20076 17128 20128 17134
rect 20076 17070 20128 17076
rect 20088 16250 20116 17070
rect 20180 16969 20208 18022
rect 20166 16960 20222 16969
rect 20166 16895 20222 16904
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 20076 16244 20128 16250
rect 20076 16186 20128 16192
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19996 13734 20024 14554
rect 20088 14074 20116 15506
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20180 15162 20208 15438
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 20180 13802 20208 14350
rect 20272 14278 20300 15438
rect 20352 15020 20404 15026
rect 20352 14962 20404 14968
rect 20364 14550 20392 14962
rect 20456 14657 20484 16390
rect 20548 16114 20576 19858
rect 20824 19854 20852 22000
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20640 18329 20668 19654
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20626 18320 20682 18329
rect 20626 18255 20682 18264
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20628 16040 20680 16046
rect 20732 16017 20760 18022
rect 20824 17202 20852 19246
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 21376 16794 21404 22000
rect 21732 18012 21784 18018
rect 21732 17954 21784 17960
rect 21744 17921 21772 17954
rect 21730 17912 21786 17921
rect 21730 17847 21786 17856
rect 21928 17678 21956 22000
rect 21916 17672 21968 17678
rect 21916 17614 21968 17620
rect 21364 16788 21416 16794
rect 21364 16730 21416 16736
rect 20628 15982 20680 15988
rect 20718 16008 20774 16017
rect 20640 15706 20668 15982
rect 20718 15943 20774 15952
rect 20628 15700 20680 15706
rect 20628 15642 20680 15648
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20548 14793 20576 14894
rect 22480 14890 22508 22000
rect 22468 14884 22520 14890
rect 22468 14826 22520 14832
rect 20534 14784 20590 14793
rect 20534 14719 20590 14728
rect 20442 14648 20498 14657
rect 20442 14583 20498 14592
rect 20352 14544 20404 14550
rect 20352 14486 20404 14492
rect 20260 14272 20312 14278
rect 20260 14214 20312 14220
rect 20364 13938 20392 14486
rect 20442 14104 20498 14113
rect 20442 14039 20498 14048
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20168 13796 20220 13802
rect 20168 13738 20220 13744
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 20456 13530 20484 14039
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20640 13705 20668 13942
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20626 13696 20682 13705
rect 20626 13631 20682 13640
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20732 12782 20760 13806
rect 20902 13288 20958 13297
rect 20902 13223 20958 13232
rect 20916 12986 20944 13223
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 19892 12436 19944 12442
rect 19892 12378 19944 12384
rect 20076 12368 20128 12374
rect 20076 12310 20128 12316
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19996 11830 20024 12038
rect 19984 11824 20036 11830
rect 19984 11766 20036 11772
rect 20088 8378 20116 12310
rect 20168 11756 20220 11762
rect 20168 11698 20220 11704
rect 20180 10062 20208 11698
rect 20812 11620 20864 11626
rect 20812 11562 20864 11568
rect 20444 10532 20496 10538
rect 20444 10474 20496 10480
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 20180 9654 20208 9998
rect 20168 9648 20220 9654
rect 20168 9590 20220 9596
rect 20456 9382 20484 10474
rect 20534 10024 20590 10033
rect 20534 9959 20590 9968
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20456 8566 20484 9318
rect 20444 8560 20496 8566
rect 20444 8502 20496 8508
rect 20548 8498 20576 9959
rect 20824 9586 20852 11562
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 19984 8356 20036 8362
rect 20088 8350 20208 8378
rect 19984 8298 20036 8304
rect 19996 7954 20024 8298
rect 20076 8288 20128 8294
rect 20076 8230 20128 8236
rect 19984 7948 20036 7954
rect 19984 7890 20036 7896
rect 19892 7336 19944 7342
rect 19892 7278 19944 7284
rect 19536 5902 19840 5930
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19352 4214 19380 5510
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19340 4208 19392 4214
rect 19340 4150 19392 4156
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 19168 2514 19288 2530
rect 19444 2514 19472 5306
rect 19168 2508 19300 2514
rect 19168 2502 19248 2508
rect 19248 2450 19300 2456
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 19156 2440 19208 2446
rect 19154 2408 19156 2417
rect 19208 2408 19210 2417
rect 19154 2343 19210 2352
rect 19536 1970 19564 5902
rect 19616 5840 19668 5846
rect 19616 5782 19668 5788
rect 19628 5370 19656 5782
rect 19616 5364 19668 5370
rect 19616 5306 19668 5312
rect 19628 4214 19656 5306
rect 19904 5114 19932 7278
rect 19996 6769 20024 7890
rect 20088 7002 20116 8230
rect 20180 7886 20208 8350
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 20456 8090 20484 8230
rect 20444 8084 20496 8090
rect 20444 8026 20496 8032
rect 20640 7970 20668 8434
rect 20548 7942 20668 7970
rect 20548 7886 20576 7942
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20076 6996 20128 7002
rect 20076 6938 20128 6944
rect 19982 6760 20038 6769
rect 19982 6695 20038 6704
rect 19904 5086 20024 5114
rect 19892 5024 19944 5030
rect 19892 4966 19944 4972
rect 19708 4548 19760 4554
rect 19708 4490 19760 4496
rect 19616 4208 19668 4214
rect 19616 4150 19668 4156
rect 19524 1964 19576 1970
rect 19524 1906 19576 1912
rect 19076 1414 19196 1442
rect 18696 1216 18748 1222
rect 18696 1158 18748 1164
rect 19168 800 19196 1414
rect 19720 800 19748 4490
rect 19800 4480 19852 4486
rect 19800 4422 19852 4428
rect 19812 4078 19840 4422
rect 19904 4146 19932 4966
rect 19892 4140 19944 4146
rect 19892 4082 19944 4088
rect 19800 4072 19852 4078
rect 19800 4014 19852 4020
rect 19996 3602 20024 5086
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 20180 2514 20208 7822
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 20258 7712 20314 7721
rect 20258 7647 20314 7656
rect 20272 7342 20300 7647
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 20352 6792 20404 6798
rect 20352 6734 20404 6740
rect 20260 6248 20312 6254
rect 20260 6190 20312 6196
rect 20272 5166 20300 6190
rect 20364 5846 20392 6734
rect 20352 5840 20404 5846
rect 20352 5782 20404 5788
rect 20456 5658 20484 7754
rect 20548 7274 20576 7822
rect 20536 7268 20588 7274
rect 20536 7210 20588 7216
rect 20548 6458 20576 7210
rect 20628 7200 20680 7206
rect 20628 7142 20680 7148
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 20536 5772 20588 5778
rect 20536 5714 20588 5720
rect 20364 5630 20484 5658
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20364 4978 20392 5630
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 20272 4950 20392 4978
rect 20272 4078 20300 4950
rect 20456 4826 20484 5170
rect 20444 4820 20496 4826
rect 20444 4762 20496 4768
rect 20456 4622 20484 4762
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 20352 4548 20404 4554
rect 20352 4490 20404 4496
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 20260 3936 20312 3942
rect 20364 3913 20392 4490
rect 20548 4146 20576 5714
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20260 3878 20312 3884
rect 20350 3904 20406 3913
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 20272 800 20300 3878
rect 20350 3839 20406 3848
rect 20640 3738 20668 7142
rect 20904 6928 20956 6934
rect 20904 6870 20956 6876
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20732 2990 20760 6190
rect 20812 6112 20864 6118
rect 20812 6054 20864 6060
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20824 800 20852 6054
rect 20916 5234 20944 6870
rect 21916 6724 21968 6730
rect 21916 6666 21968 6672
rect 20904 5228 20956 5234
rect 20904 5170 20956 5176
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20916 2582 20944 4558
rect 21364 3732 21416 3738
rect 21364 3674 21416 3680
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 21376 800 21404 3674
rect 21928 800 21956 6666
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 22480 800 22508 4082
rect 12162 640 12218 649
rect 12162 575 12218 584
rect 12530 0 12586 800
rect 13082 0 13138 800
rect 13634 0 13690 800
rect 14186 0 14242 800
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15842 0 15898 800
rect 16394 0 16450 800
rect 16946 0 17002 800
rect 17498 0 17554 800
rect 18050 0 18106 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21914 0 21970 800
rect 22466 0 22522 800
<< via2 >>
rect 18786 22072 18842 22128
rect 294 18264 350 18320
rect 1950 18672 2006 18728
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 3422 17176 3478 17232
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 8758 18808 8814 18864
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4066 5788 4068 5808
rect 4068 5788 4120 5808
rect 4120 5788 4122 5808
rect 4066 5752 4122 5788
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 9678 18400 9734 18456
rect 8758 18128 8814 18184
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 10506 19216 10562 19272
rect 10414 18400 10470 18456
rect 10322 17856 10378 17912
rect 10138 17720 10194 17776
rect 10322 16632 10378 16688
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 10690 18264 10746 18320
rect 10046 13640 10102 13696
rect 10322 11056 10378 11112
rect 10230 9560 10286 9616
rect 10046 6296 10102 6352
rect 11518 18964 11574 19000
rect 11518 18944 11520 18964
rect 11520 18944 11572 18964
rect 11572 18944 11574 18964
rect 10966 18400 11022 18456
rect 10874 17992 10930 18048
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 10782 15544 10838 15600
rect 11242 18028 11244 18048
rect 11244 18028 11296 18048
rect 11296 18028 11298 18048
rect 11242 17992 11298 18028
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 12070 18808 12126 18864
rect 11978 17040 12034 17096
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 10414 9560 10470 9616
rect 10230 2896 10286 2952
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 12346 18264 12402 18320
rect 12070 12280 12126 12336
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11794 6160 11850 6216
rect 12070 5788 12072 5808
rect 12072 5788 12124 5808
rect 12124 5788 12126 5808
rect 12070 5752 12126 5788
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 10874 1536 10930 1592
rect 13266 15988 13268 16008
rect 13268 15988 13320 16008
rect 13320 15988 13322 16008
rect 13266 15952 13322 15988
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 13910 18128 13966 18184
rect 13450 16088 13506 16144
rect 12806 13676 12808 13696
rect 12808 13676 12860 13696
rect 12860 13676 12862 13696
rect 12806 13640 12862 13676
rect 13542 14456 13598 14512
rect 13726 16244 13782 16280
rect 13726 16224 13728 16244
rect 13728 16224 13780 16244
rect 13780 16224 13782 16244
rect 13082 13368 13138 13424
rect 12806 12824 12862 12880
rect 13266 12960 13322 13016
rect 12898 10512 12954 10568
rect 13174 9016 13230 9072
rect 13450 10512 13506 10568
rect 13266 7792 13322 7848
rect 14278 17176 14334 17232
rect 14278 13232 14334 13288
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 15106 16632 15162 16688
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 15750 17740 15806 17776
rect 15750 17720 15752 17740
rect 15752 17720 15804 17740
rect 15804 17720 15806 17740
rect 15382 15408 15438 15464
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14554 13232 14610 13288
rect 14646 12960 14702 13016
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 14554 11736 14610 11792
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 15198 11348 15254 11384
rect 15198 11328 15200 11348
rect 15200 11328 15252 11348
rect 15252 11328 15254 11348
rect 15842 16244 15898 16280
rect 15842 16224 15844 16244
rect 15844 16224 15896 16244
rect 15896 16224 15898 16244
rect 15382 12280 15438 12336
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14922 10104 14978 10160
rect 14922 9424 14978 9480
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14738 9036 14794 9072
rect 14002 6296 14058 6352
rect 13358 1536 13414 1592
rect 14738 9016 14740 9036
rect 14740 9016 14792 9036
rect 14792 9016 14794 9036
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 16394 16496 16450 16552
rect 15198 9016 15254 9072
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 15934 12960 15990 13016
rect 16118 12144 16174 12200
rect 15934 8472 15990 8528
rect 16302 12960 16358 13016
rect 16486 12280 16542 12336
rect 16854 19216 16910 19272
rect 17866 20576 17922 20632
rect 16854 18808 16910 18864
rect 17038 17720 17094 17776
rect 16854 16088 16910 16144
rect 16854 15680 16910 15736
rect 16394 12144 16450 12200
rect 16486 11464 16542 11520
rect 16394 10512 16450 10568
rect 16394 9152 16450 9208
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 15566 2896 15622 2952
rect 15842 5752 15898 5808
rect 16026 2388 16028 2408
rect 16028 2388 16080 2408
rect 16080 2388 16082 2408
rect 16026 2352 16082 2388
rect 16486 8200 16542 8256
rect 18510 21120 18566 21176
rect 17590 18672 17646 18728
rect 17498 17604 17554 17640
rect 17498 17584 17500 17604
rect 17500 17584 17552 17604
rect 17552 17584 17554 17604
rect 17314 15952 17370 16008
rect 17222 15408 17278 15464
rect 16946 12144 17002 12200
rect 16762 5752 16818 5808
rect 17314 14728 17370 14784
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 17866 17620 17868 17640
rect 17868 17620 17920 17640
rect 17920 17620 17922 17640
rect 17866 17584 17922 17620
rect 18142 17720 18198 17776
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18418 17040 18474 17096
rect 19246 22480 19302 22536
rect 19062 21528 19118 21584
rect 18510 16532 18512 16552
rect 18512 16532 18564 16552
rect 18564 16532 18566 16552
rect 18510 16496 18566 16532
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 17406 12280 17462 12336
rect 17314 11056 17370 11112
rect 17590 11076 17646 11112
rect 17590 11056 17592 11076
rect 17592 11056 17644 11076
rect 17644 11056 17646 11076
rect 17130 8200 17186 8256
rect 17590 7384 17646 7440
rect 17590 6160 17646 6216
rect 18050 15544 18106 15600
rect 18234 15544 18290 15600
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18602 15000 18658 15056
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 17866 13388 17922 13424
rect 17866 13368 17868 13388
rect 17868 13368 17920 13388
rect 17920 13368 17922 13388
rect 17866 12688 17922 12744
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18694 13368 18750 13424
rect 18326 12824 18382 12880
rect 18234 12416 18290 12472
rect 18050 12180 18052 12200
rect 18052 12180 18104 12200
rect 18104 12180 18106 12200
rect 18050 12144 18106 12180
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18050 10648 18106 10704
rect 18326 10512 18382 10568
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 17866 8084 17922 8120
rect 18142 9016 18198 9072
rect 18418 9444 18474 9480
rect 18418 9424 18420 9444
rect 18420 9424 18472 9444
rect 18472 9424 18474 9444
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18050 8472 18106 8528
rect 18970 18128 19026 18184
rect 19154 19760 19210 19816
rect 19614 20168 19670 20224
rect 19890 19216 19946 19272
rect 19246 17312 19302 17368
rect 19430 16496 19486 16552
rect 19062 14456 19118 14512
rect 18970 11600 19026 11656
rect 18970 10376 19026 10432
rect 19154 11464 19210 11520
rect 19338 10376 19394 10432
rect 18694 9288 18750 9344
rect 17866 8064 17868 8084
rect 17868 8064 17920 8084
rect 17920 8064 17922 8084
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 18050 5752 18106 5808
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18326 5208 18382 5264
rect 18050 4528 18106 4584
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18418 2896 18474 2952
rect 17866 2488 17922 2544
rect 18878 6160 18934 6216
rect 18786 4256 18842 4312
rect 19154 7792 19210 7848
rect 19338 7692 19340 7712
rect 19340 7692 19392 7712
rect 19392 7692 19394 7712
rect 19338 7656 19394 7692
rect 19154 7112 19210 7168
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 18050 1980 18052 2000
rect 18052 1980 18104 2000
rect 18104 1980 18106 2000
rect 18050 1944 18106 1980
rect 20166 18808 20222 18864
rect 20166 16904 20222 16960
rect 20626 18264 20682 18320
rect 21730 17856 21786 17912
rect 20718 15952 20774 16008
rect 20534 14728 20590 14784
rect 20442 14592 20498 14648
rect 20442 14048 20498 14104
rect 20626 13640 20682 13696
rect 20902 13232 20958 13288
rect 20534 9968 20590 10024
rect 19154 2388 19156 2408
rect 19156 2388 19208 2408
rect 19208 2388 19210 2408
rect 19154 2352 19210 2388
rect 19982 6704 20038 6760
rect 20258 7656 20314 7712
rect 20350 3848 20406 3904
rect 12162 584 12218 640
<< metal3 >>
rect 19241 22538 19307 22541
rect 22000 22538 22800 22568
rect 19241 22536 22800 22538
rect 19241 22480 19246 22536
rect 19302 22480 22800 22536
rect 19241 22478 22800 22480
rect 19241 22475 19307 22478
rect 22000 22448 22800 22478
rect 18781 22130 18847 22133
rect 22000 22130 22800 22160
rect 18781 22128 22800 22130
rect 18781 22072 18786 22128
rect 18842 22072 22800 22128
rect 18781 22070 22800 22072
rect 18781 22067 18847 22070
rect 22000 22040 22800 22070
rect 19057 21586 19123 21589
rect 22000 21586 22800 21616
rect 19057 21584 22800 21586
rect 19057 21528 19062 21584
rect 19118 21528 22800 21584
rect 19057 21526 22800 21528
rect 19057 21523 19123 21526
rect 22000 21496 22800 21526
rect 18505 21178 18571 21181
rect 22000 21178 22800 21208
rect 18505 21176 22800 21178
rect 18505 21120 18510 21176
rect 18566 21120 22800 21176
rect 18505 21118 22800 21120
rect 18505 21115 18571 21118
rect 22000 21088 22800 21118
rect 17861 20634 17927 20637
rect 22000 20634 22800 20664
rect 17861 20632 22800 20634
rect 17861 20576 17866 20632
rect 17922 20576 22800 20632
rect 17861 20574 22800 20576
rect 17861 20571 17927 20574
rect 22000 20544 22800 20574
rect 19609 20226 19675 20229
rect 22000 20226 22800 20256
rect 19609 20224 22800 20226
rect 19609 20168 19614 20224
rect 19670 20168 22800 20224
rect 19609 20166 22800 20168
rect 19609 20163 19675 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22000 20136 22800 20166
rect 14672 20095 14992 20096
rect 19149 19818 19215 19821
rect 22000 19818 22800 19848
rect 19149 19816 22800 19818
rect 19149 19760 19154 19816
rect 19210 19760 22800 19816
rect 19149 19758 22800 19760
rect 19149 19755 19215 19758
rect 22000 19728 22800 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 10501 19274 10567 19277
rect 16849 19274 16915 19277
rect 10501 19272 16915 19274
rect 10501 19216 10506 19272
rect 10562 19216 16854 19272
rect 16910 19216 16915 19272
rect 10501 19214 16915 19216
rect 10501 19211 10567 19214
rect 16849 19211 16915 19214
rect 19885 19274 19951 19277
rect 22000 19274 22800 19304
rect 19885 19272 22800 19274
rect 19885 19216 19890 19272
rect 19946 19216 22800 19272
rect 19885 19214 22800 19216
rect 19885 19211 19951 19214
rect 22000 19184 22800 19214
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 11513 19002 11579 19005
rect 11513 19000 12266 19002
rect 11513 18944 11518 19000
rect 11574 18944 12266 19000
rect 11513 18942 12266 18944
rect 11513 18939 11579 18942
rect 8753 18866 8819 18869
rect 12065 18866 12131 18869
rect 8753 18864 12131 18866
rect 8753 18808 8758 18864
rect 8814 18808 12070 18864
rect 12126 18808 12131 18864
rect 8753 18806 12131 18808
rect 12206 18866 12266 18942
rect 16849 18866 16915 18869
rect 12206 18864 16915 18866
rect 12206 18808 16854 18864
rect 16910 18808 16915 18864
rect 12206 18806 16915 18808
rect 8753 18803 8819 18806
rect 12065 18803 12131 18806
rect 16849 18803 16915 18806
rect 20161 18866 20227 18869
rect 22000 18866 22800 18896
rect 20161 18864 22800 18866
rect 20161 18808 20166 18864
rect 20222 18808 22800 18864
rect 20161 18806 22800 18808
rect 20161 18803 20227 18806
rect 22000 18776 22800 18806
rect 1945 18730 2011 18733
rect 17585 18730 17651 18733
rect 1945 18728 17651 18730
rect 1945 18672 1950 18728
rect 2006 18672 17590 18728
rect 17646 18672 17651 18728
rect 1945 18670 17651 18672
rect 1945 18667 2011 18670
rect 17585 18667 17651 18670
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 9673 18458 9739 18461
rect 10409 18458 10475 18461
rect 10961 18458 11027 18461
rect 9673 18456 11162 18458
rect 9673 18400 9678 18456
rect 9734 18400 10414 18456
rect 10470 18400 10966 18456
rect 11022 18400 11162 18456
rect 9673 18398 11162 18400
rect 9673 18395 9739 18398
rect 10409 18395 10475 18398
rect 10961 18395 11027 18398
rect 289 18322 355 18325
rect 10685 18322 10751 18325
rect 289 18320 10751 18322
rect 289 18264 294 18320
rect 350 18264 10690 18320
rect 10746 18264 10751 18320
rect 289 18262 10751 18264
rect 11102 18322 11162 18398
rect 12341 18322 12407 18325
rect 11102 18320 12407 18322
rect 11102 18264 12346 18320
rect 12402 18264 12407 18320
rect 11102 18262 12407 18264
rect 289 18259 355 18262
rect 10685 18259 10751 18262
rect 12341 18259 12407 18262
rect 20621 18322 20687 18325
rect 22000 18322 22800 18352
rect 20621 18320 22800 18322
rect 20621 18264 20626 18320
rect 20682 18264 22800 18320
rect 20621 18262 22800 18264
rect 20621 18259 20687 18262
rect 22000 18232 22800 18262
rect 8753 18186 8819 18189
rect 13905 18186 13971 18189
rect 18965 18186 19031 18189
rect 8753 18184 13971 18186
rect 8753 18128 8758 18184
rect 8814 18128 13910 18184
rect 13966 18128 13971 18184
rect 8753 18126 13971 18128
rect 8753 18123 8819 18126
rect 13905 18123 13971 18126
rect 14046 18184 19031 18186
rect 14046 18128 18970 18184
rect 19026 18128 19031 18184
rect 14046 18126 19031 18128
rect 10869 18050 10935 18053
rect 11237 18050 11303 18053
rect 10869 18048 11303 18050
rect 10869 17992 10874 18048
rect 10930 17992 11242 18048
rect 11298 17992 11303 18048
rect 10869 17990 11303 17992
rect 10869 17987 10935 17990
rect 11237 17987 11303 17990
rect 7808 17984 8128 17985
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 10317 17914 10383 17917
rect 14046 17914 14106 18126
rect 18965 18123 19031 18126
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 10317 17912 14106 17914
rect 10317 17856 10322 17912
rect 10378 17856 14106 17912
rect 10317 17854 14106 17856
rect 21725 17914 21791 17917
rect 22000 17914 22800 17944
rect 21725 17912 22800 17914
rect 21725 17856 21730 17912
rect 21786 17856 22800 17912
rect 21725 17854 22800 17856
rect 10317 17851 10383 17854
rect 21725 17851 21791 17854
rect 22000 17824 22800 17854
rect 10133 17778 10199 17781
rect 15745 17778 15811 17781
rect 10133 17776 15811 17778
rect 10133 17720 10138 17776
rect 10194 17720 15750 17776
rect 15806 17720 15811 17776
rect 10133 17718 15811 17720
rect 10133 17715 10199 17718
rect 15745 17715 15811 17718
rect 17033 17778 17099 17781
rect 18137 17778 18203 17781
rect 17033 17776 18203 17778
rect 17033 17720 17038 17776
rect 17094 17720 18142 17776
rect 18198 17720 18203 17776
rect 17033 17718 18203 17720
rect 17033 17715 17099 17718
rect 18137 17715 18203 17718
rect 17493 17642 17559 17645
rect 17861 17642 17927 17645
rect 17493 17640 17927 17642
rect 17493 17584 17498 17640
rect 17554 17584 17866 17640
rect 17922 17584 17927 17640
rect 17493 17582 17927 17584
rect 17493 17579 17559 17582
rect 17861 17579 17927 17582
rect 4376 17440 4696 17441
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 19241 17370 19307 17373
rect 22000 17370 22800 17400
rect 19241 17368 22800 17370
rect 19241 17312 19246 17368
rect 19302 17312 22800 17368
rect 19241 17310 22800 17312
rect 19241 17307 19307 17310
rect 22000 17280 22800 17310
rect 0 17234 800 17264
rect 3417 17234 3483 17237
rect 0 17232 3483 17234
rect 0 17176 3422 17232
rect 3478 17176 3483 17232
rect 0 17174 3483 17176
rect 0 17144 800 17174
rect 3417 17171 3483 17174
rect 14273 17234 14339 17237
rect 15510 17234 15516 17236
rect 14273 17232 15516 17234
rect 14273 17176 14278 17232
rect 14334 17176 15516 17232
rect 14273 17174 15516 17176
rect 14273 17171 14339 17174
rect 15510 17172 15516 17174
rect 15580 17172 15586 17236
rect 11973 17098 12039 17101
rect 15142 17098 15148 17100
rect 11973 17096 15148 17098
rect 11973 17040 11978 17096
rect 12034 17040 15148 17096
rect 11973 17038 15148 17040
rect 11973 17035 12039 17038
rect 15142 17036 15148 17038
rect 15212 17098 15218 17100
rect 18413 17098 18479 17101
rect 15212 17096 18479 17098
rect 15212 17040 18418 17096
rect 18474 17040 18479 17096
rect 15212 17038 18479 17040
rect 15212 17036 15218 17038
rect 18413 17035 18479 17038
rect 20161 16962 20227 16965
rect 22000 16962 22800 16992
rect 20161 16960 22800 16962
rect 20161 16904 20166 16960
rect 20222 16904 22800 16960
rect 20161 16902 22800 16904
rect 20161 16899 20227 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 22000 16872 22800 16902
rect 14672 16831 14992 16832
rect 10317 16690 10383 16693
rect 15101 16690 15167 16693
rect 10317 16688 15167 16690
rect 10317 16632 10322 16688
rect 10378 16632 15106 16688
rect 15162 16632 15167 16688
rect 10317 16630 15167 16632
rect 10317 16627 10383 16630
rect 15101 16627 15167 16630
rect 16389 16554 16455 16557
rect 18505 16554 18571 16557
rect 16389 16552 18571 16554
rect 16389 16496 16394 16552
rect 16450 16496 18510 16552
rect 18566 16496 18571 16552
rect 16389 16494 18571 16496
rect 16389 16491 16455 16494
rect 18505 16491 18571 16494
rect 19425 16554 19491 16557
rect 22000 16554 22800 16584
rect 19425 16552 22800 16554
rect 19425 16496 19430 16552
rect 19486 16496 22800 16552
rect 19425 16494 22800 16496
rect 19425 16491 19491 16494
rect 22000 16464 22800 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 13721 16282 13787 16285
rect 15837 16282 15903 16285
rect 13721 16280 15903 16282
rect 13721 16224 13726 16280
rect 13782 16224 15842 16280
rect 15898 16224 15903 16280
rect 13721 16222 15903 16224
rect 13721 16219 13787 16222
rect 15837 16219 15903 16222
rect 13445 16146 13511 16149
rect 16849 16146 16915 16149
rect 13445 16144 16915 16146
rect 13445 16088 13450 16144
rect 13506 16088 16854 16144
rect 16910 16088 16915 16144
rect 13445 16086 16915 16088
rect 13445 16083 13511 16086
rect 16849 16083 16915 16086
rect 13261 16010 13327 16013
rect 17309 16010 17375 16013
rect 13261 16008 17375 16010
rect 13261 15952 13266 16008
rect 13322 15952 17314 16008
rect 17370 15952 17375 16008
rect 13261 15950 17375 15952
rect 13261 15947 13327 15950
rect 17309 15947 17375 15950
rect 20713 16010 20779 16013
rect 22000 16010 22800 16040
rect 20713 16008 22800 16010
rect 20713 15952 20718 16008
rect 20774 15952 22800 16008
rect 20713 15950 22800 15952
rect 20713 15947 20779 15950
rect 22000 15920 22800 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 16849 15738 16915 15741
rect 16982 15738 16988 15740
rect 16849 15736 16988 15738
rect 16849 15680 16854 15736
rect 16910 15680 16988 15736
rect 16849 15678 16988 15680
rect 16849 15675 16915 15678
rect 16982 15676 16988 15678
rect 17052 15676 17058 15740
rect 10777 15602 10843 15605
rect 18045 15602 18111 15605
rect 10777 15600 18111 15602
rect 10777 15544 10782 15600
rect 10838 15544 18050 15600
rect 18106 15544 18111 15600
rect 10777 15542 18111 15544
rect 10777 15539 10843 15542
rect 18045 15539 18111 15542
rect 18229 15602 18295 15605
rect 22000 15602 22800 15632
rect 18229 15600 22800 15602
rect 18229 15544 18234 15600
rect 18290 15544 22800 15600
rect 18229 15542 22800 15544
rect 18229 15539 18295 15542
rect 22000 15512 22800 15542
rect 15377 15466 15443 15469
rect 17217 15466 17283 15469
rect 15377 15464 17283 15466
rect 15377 15408 15382 15464
rect 15438 15408 17222 15464
rect 17278 15408 17283 15464
rect 15377 15406 17283 15408
rect 15377 15403 15443 15406
rect 17217 15403 17283 15406
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 18597 15058 18663 15061
rect 22000 15058 22800 15088
rect 18597 15056 22800 15058
rect 18597 15000 18602 15056
rect 18658 15000 22800 15056
rect 18597 14998 22800 15000
rect 18597 14995 18663 14998
rect 22000 14968 22800 14998
rect 17309 14786 17375 14789
rect 19190 14786 19196 14788
rect 17309 14784 19196 14786
rect 17309 14728 17314 14784
rect 17370 14728 19196 14784
rect 17309 14726 19196 14728
rect 17309 14723 17375 14726
rect 19190 14724 19196 14726
rect 19260 14786 19266 14788
rect 20529 14786 20595 14789
rect 19260 14784 20595 14786
rect 19260 14728 20534 14784
rect 20590 14728 20595 14784
rect 19260 14726 20595 14728
rect 19260 14724 19266 14726
rect 20529 14723 20595 14726
rect 7808 14720 8128 14721
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 20437 14650 20503 14653
rect 22000 14650 22800 14680
rect 20437 14648 22800 14650
rect 20437 14592 20442 14648
rect 20498 14592 22800 14648
rect 20437 14590 22800 14592
rect 20437 14587 20503 14590
rect 22000 14560 22800 14590
rect 13537 14514 13603 14517
rect 19057 14514 19123 14517
rect 13537 14512 19123 14514
rect 13537 14456 13542 14512
rect 13598 14456 19062 14512
rect 19118 14456 19123 14512
rect 13537 14454 19123 14456
rect 13537 14451 13603 14454
rect 19057 14451 19123 14454
rect 4376 14176 4696 14177
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 20437 14106 20503 14109
rect 22000 14106 22800 14136
rect 20437 14104 22800 14106
rect 20437 14048 20442 14104
rect 20498 14048 22800 14104
rect 20437 14046 22800 14048
rect 20437 14043 20503 14046
rect 22000 14016 22800 14046
rect 10041 13698 10107 13701
rect 12801 13698 12867 13701
rect 10041 13696 12867 13698
rect 10041 13640 10046 13696
rect 10102 13640 12806 13696
rect 12862 13640 12867 13696
rect 10041 13638 12867 13640
rect 10041 13635 10107 13638
rect 12801 13635 12867 13638
rect 20621 13698 20687 13701
rect 22000 13698 22800 13728
rect 20621 13696 22800 13698
rect 20621 13640 20626 13696
rect 20682 13640 22800 13696
rect 20621 13638 22800 13640
rect 20621 13635 20687 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 22000 13608 22800 13638
rect 14672 13567 14992 13568
rect 13077 13426 13143 13429
rect 17861 13426 17927 13429
rect 18689 13428 18755 13429
rect 18638 13426 18644 13428
rect 13077 13424 17927 13426
rect 13077 13368 13082 13424
rect 13138 13368 17866 13424
rect 17922 13368 17927 13424
rect 13077 13366 17927 13368
rect 18598 13366 18644 13426
rect 18708 13424 18755 13428
rect 18750 13368 18755 13424
rect 13077 13363 13143 13366
rect 17861 13363 17927 13366
rect 18638 13364 18644 13366
rect 18708 13364 18755 13368
rect 18689 13363 18755 13364
rect 14273 13290 14339 13293
rect 14549 13290 14615 13293
rect 14273 13288 14615 13290
rect 14273 13232 14278 13288
rect 14334 13232 14554 13288
rect 14610 13232 14615 13288
rect 14273 13230 14615 13232
rect 14273 13227 14339 13230
rect 14549 13227 14615 13230
rect 20897 13290 20963 13293
rect 22000 13290 22800 13320
rect 20897 13288 22800 13290
rect 20897 13232 20902 13288
rect 20958 13232 22800 13288
rect 20897 13230 22800 13232
rect 20897 13227 20963 13230
rect 22000 13200 22800 13230
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 13261 13018 13327 13021
rect 14641 13018 14707 13021
rect 13261 13016 14707 13018
rect 13261 12960 13266 13016
rect 13322 12960 14646 13016
rect 14702 12960 14707 13016
rect 13261 12958 14707 12960
rect 13261 12955 13327 12958
rect 14641 12955 14707 12958
rect 15510 12956 15516 13020
rect 15580 13018 15586 13020
rect 15929 13018 15995 13021
rect 15580 13016 15995 13018
rect 15580 12960 15934 13016
rect 15990 12960 15995 13016
rect 15580 12958 15995 12960
rect 15580 12956 15586 12958
rect 15929 12955 15995 12958
rect 16297 13018 16363 13021
rect 16297 13016 18016 13018
rect 16297 12960 16302 13016
rect 16358 12960 18016 13016
rect 16297 12958 18016 12960
rect 16297 12955 16363 12958
rect 12801 12882 12867 12885
rect 16430 12882 16436 12884
rect 12801 12880 16436 12882
rect 12801 12824 12806 12880
rect 12862 12824 16436 12880
rect 12801 12822 16436 12824
rect 12801 12819 12867 12822
rect 16430 12820 16436 12822
rect 16500 12820 16506 12884
rect 17956 12882 18016 12958
rect 18321 12882 18387 12885
rect 17956 12880 18387 12882
rect 17956 12824 18326 12880
rect 18382 12824 18387 12880
rect 17956 12822 18387 12824
rect 18321 12819 18387 12822
rect 17861 12746 17927 12749
rect 22000 12746 22800 12776
rect 17861 12744 22800 12746
rect 17861 12688 17866 12744
rect 17922 12688 22800 12744
rect 17861 12686 22800 12688
rect 17861 12683 17927 12686
rect 22000 12656 22800 12686
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 16430 12412 16436 12476
rect 16500 12474 16506 12476
rect 18229 12474 18295 12477
rect 16500 12472 18295 12474
rect 16500 12416 18234 12472
rect 18290 12416 18295 12472
rect 16500 12414 18295 12416
rect 16500 12412 16506 12414
rect 18229 12411 18295 12414
rect 12065 12338 12131 12341
rect 15377 12338 15443 12341
rect 12065 12336 15443 12338
rect 12065 12280 12070 12336
rect 12126 12280 15382 12336
rect 15438 12280 15443 12336
rect 12065 12278 15443 12280
rect 12065 12275 12131 12278
rect 15377 12275 15443 12278
rect 16481 12338 16547 12341
rect 17401 12338 17467 12341
rect 22000 12338 22800 12368
rect 16481 12336 17234 12338
rect 16481 12280 16486 12336
rect 16542 12280 17234 12336
rect 16481 12278 17234 12280
rect 16481 12275 16547 12278
rect 16113 12202 16179 12205
rect 16389 12202 16455 12205
rect 16941 12204 17007 12205
rect 16941 12202 16988 12204
rect 16113 12200 16455 12202
rect 16113 12144 16118 12200
rect 16174 12144 16394 12200
rect 16450 12144 16455 12200
rect 16113 12142 16455 12144
rect 16896 12200 16988 12202
rect 16896 12144 16946 12200
rect 16896 12142 16988 12144
rect 16113 12139 16179 12142
rect 16389 12139 16455 12142
rect 16941 12140 16988 12142
rect 17052 12140 17058 12204
rect 17174 12202 17234 12278
rect 17401 12336 22800 12338
rect 17401 12280 17406 12336
rect 17462 12280 22800 12336
rect 17401 12278 22800 12280
rect 17401 12275 17467 12278
rect 22000 12248 22800 12278
rect 18045 12202 18111 12205
rect 17174 12200 18111 12202
rect 17174 12144 18050 12200
rect 18106 12144 18111 12200
rect 17174 12142 18111 12144
rect 16941 12139 17007 12140
rect 18045 12139 18111 12142
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 14549 11794 14615 11797
rect 22000 11794 22800 11824
rect 14549 11792 22800 11794
rect 14549 11736 14554 11792
rect 14610 11736 22800 11792
rect 14549 11734 22800 11736
rect 14549 11731 14615 11734
rect 22000 11704 22800 11734
rect 18965 11660 19031 11661
rect 18965 11658 19012 11660
rect 18920 11656 19012 11658
rect 18920 11600 18970 11656
rect 18920 11598 19012 11600
rect 18965 11596 19012 11598
rect 19076 11596 19082 11660
rect 18965 11595 19031 11596
rect 16481 11522 16547 11525
rect 19149 11522 19215 11525
rect 16481 11520 19215 11522
rect 16481 11464 16486 11520
rect 16542 11464 19154 11520
rect 19210 11464 19215 11520
rect 16481 11462 19215 11464
rect 16481 11459 16547 11462
rect 19149 11459 19215 11462
rect 7808 11456 8128 11457
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 15193 11386 15259 11389
rect 22000 11386 22800 11416
rect 15193 11384 22800 11386
rect 15193 11328 15198 11384
rect 15254 11328 22800 11384
rect 15193 11326 22800 11328
rect 15193 11323 15259 11326
rect 22000 11296 22800 11326
rect 10317 11114 10383 11117
rect 17309 11114 17375 11117
rect 17585 11114 17651 11117
rect 10317 11112 17651 11114
rect 10317 11056 10322 11112
rect 10378 11056 17314 11112
rect 17370 11056 17590 11112
rect 17646 11056 17651 11112
rect 10317 11054 17651 11056
rect 10317 11051 10383 11054
rect 17309 11051 17375 11054
rect 17585 11051 17651 11054
rect 4376 10912 4696 10913
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 22000 10842 22800 10872
rect 18646 10782 22800 10842
rect 18045 10706 18111 10709
rect 18646 10706 18706 10782
rect 22000 10752 22800 10782
rect 18045 10704 18706 10706
rect 18045 10648 18050 10704
rect 18106 10648 18706 10704
rect 18045 10646 18706 10648
rect 18045 10643 18111 10646
rect 12893 10570 12959 10573
rect 13445 10570 13511 10573
rect 12893 10568 13511 10570
rect 12893 10512 12898 10568
rect 12954 10512 13450 10568
rect 13506 10512 13511 10568
rect 12893 10510 13511 10512
rect 12893 10507 12959 10510
rect 13445 10507 13511 10510
rect 16389 10570 16455 10573
rect 18321 10570 18387 10573
rect 18638 10570 18644 10572
rect 16389 10568 18644 10570
rect 16389 10512 16394 10568
rect 16450 10512 18326 10568
rect 18382 10512 18644 10568
rect 16389 10510 18644 10512
rect 16389 10507 16455 10510
rect 18321 10507 18387 10510
rect 18638 10508 18644 10510
rect 18708 10508 18714 10572
rect 18965 10434 19031 10437
rect 19333 10434 19399 10437
rect 22000 10434 22800 10464
rect 18965 10432 22800 10434
rect 18965 10376 18970 10432
rect 19026 10376 19338 10432
rect 19394 10376 22800 10432
rect 18965 10374 22800 10376
rect 18965 10371 19031 10374
rect 19333 10371 19399 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 22000 10344 22800 10374
rect 14672 10303 14992 10304
rect 14917 10162 14983 10165
rect 15142 10162 15148 10164
rect 14917 10160 15148 10162
rect 14917 10104 14922 10160
rect 14978 10104 15148 10160
rect 14917 10102 15148 10104
rect 14917 10099 14983 10102
rect 15142 10100 15148 10102
rect 15212 10100 15218 10164
rect 20529 10026 20595 10029
rect 22000 10026 22800 10056
rect 20529 10024 22800 10026
rect 20529 9968 20534 10024
rect 20590 9968 22800 10024
rect 20529 9966 22800 9968
rect 20529 9963 20595 9966
rect 22000 9936 22800 9966
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 10225 9618 10291 9621
rect 10409 9618 10475 9621
rect 10225 9616 10475 9618
rect 10225 9560 10230 9616
rect 10286 9560 10414 9616
rect 10470 9560 10475 9616
rect 10225 9558 10475 9560
rect 10225 9555 10291 9558
rect 10409 9555 10475 9558
rect 14917 9482 14983 9485
rect 18413 9482 18479 9485
rect 22000 9482 22800 9512
rect 14917 9480 15210 9482
rect 14917 9424 14922 9480
rect 14978 9424 15210 9480
rect 14917 9422 15210 9424
rect 14917 9419 14983 9422
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 15150 9077 15210 9422
rect 18413 9480 22800 9482
rect 18413 9424 18418 9480
rect 18474 9424 22800 9480
rect 18413 9422 22800 9424
rect 18413 9419 18479 9422
rect 22000 9392 22800 9422
rect 18689 9346 18755 9349
rect 18822 9346 18828 9348
rect 18689 9344 18828 9346
rect 18689 9288 18694 9344
rect 18750 9288 18828 9344
rect 18689 9286 18828 9288
rect 18689 9283 18755 9286
rect 18822 9284 18828 9286
rect 18892 9284 18898 9348
rect 16389 9210 16455 9213
rect 16254 9208 16455 9210
rect 16254 9152 16394 9208
rect 16450 9152 16455 9208
rect 16254 9150 16455 9152
rect 13169 9074 13235 9077
rect 14733 9074 14799 9077
rect 13169 9072 14799 9074
rect 13169 9016 13174 9072
rect 13230 9016 14738 9072
rect 14794 9016 14799 9072
rect 13169 9014 14799 9016
rect 15150 9072 15259 9077
rect 15150 9016 15198 9072
rect 15254 9016 15259 9072
rect 15150 9014 15259 9016
rect 13169 9011 13235 9014
rect 14733 9011 14799 9014
rect 15193 9011 15259 9014
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 15929 8530 15995 8533
rect 16254 8530 16314 9150
rect 16389 9147 16455 9150
rect 18137 9074 18203 9077
rect 22000 9074 22800 9104
rect 18137 9072 22800 9074
rect 18137 9016 18142 9072
rect 18198 9016 22800 9072
rect 18137 9014 22800 9016
rect 18137 9011 18203 9014
rect 22000 8984 22800 9014
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 15929 8528 16314 8530
rect 15929 8472 15934 8528
rect 15990 8472 16314 8528
rect 15929 8470 16314 8472
rect 18045 8530 18111 8533
rect 22000 8530 22800 8560
rect 18045 8528 22800 8530
rect 18045 8472 18050 8528
rect 18106 8472 22800 8528
rect 18045 8470 22800 8472
rect 15929 8467 15995 8470
rect 18045 8467 18111 8470
rect 22000 8440 22800 8470
rect 16481 8258 16547 8261
rect 17125 8258 17191 8261
rect 16481 8256 17191 8258
rect 16481 8200 16486 8256
rect 16542 8200 17130 8256
rect 17186 8200 17191 8256
rect 16481 8198 17191 8200
rect 16481 8195 16547 8198
rect 17125 8195 17191 8198
rect 7808 8192 8128 8193
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 17861 8122 17927 8125
rect 22000 8122 22800 8152
rect 17861 8120 22800 8122
rect 17861 8064 17866 8120
rect 17922 8064 22800 8120
rect 17861 8062 22800 8064
rect 17861 8059 17927 8062
rect 22000 8032 22800 8062
rect 13261 7850 13327 7853
rect 19149 7850 19215 7853
rect 13261 7848 19215 7850
rect 13261 7792 13266 7848
rect 13322 7792 19154 7848
rect 19210 7792 19215 7848
rect 13261 7790 19215 7792
rect 13261 7787 13327 7790
rect 19149 7787 19215 7790
rect 19333 7714 19399 7717
rect 20253 7714 20319 7717
rect 19333 7712 20319 7714
rect 19333 7656 19338 7712
rect 19394 7656 20258 7712
rect 20314 7656 20319 7712
rect 19333 7654 20319 7656
rect 19333 7651 19399 7654
rect 20253 7651 20319 7654
rect 4376 7648 4696 7649
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 22000 7578 22800 7608
rect 18600 7518 22800 7578
rect 17585 7442 17651 7445
rect 18600 7442 18660 7518
rect 22000 7488 22800 7518
rect 17585 7440 18660 7442
rect 17585 7384 17590 7440
rect 17646 7384 18660 7440
rect 17585 7382 18660 7384
rect 17585 7379 17651 7382
rect 19149 7170 19215 7173
rect 22000 7170 22800 7200
rect 19149 7168 22800 7170
rect 19149 7112 19154 7168
rect 19210 7112 22800 7168
rect 19149 7110 22800 7112
rect 19149 7107 19215 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 22000 7080 22800 7110
rect 14672 7039 14992 7040
rect 19977 6762 20043 6765
rect 22000 6762 22800 6792
rect 19977 6760 22800 6762
rect 19977 6704 19982 6760
rect 20038 6704 22800 6760
rect 19977 6702 22800 6704
rect 19977 6699 20043 6702
rect 22000 6672 22800 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 10041 6354 10107 6357
rect 13997 6354 14063 6357
rect 10041 6352 14063 6354
rect 10041 6296 10046 6352
rect 10102 6296 14002 6352
rect 14058 6296 14063 6352
rect 10041 6294 14063 6296
rect 10041 6291 10107 6294
rect 13997 6291 14063 6294
rect 11789 6218 11855 6221
rect 17585 6218 17651 6221
rect 11789 6216 17651 6218
rect 11789 6160 11794 6216
rect 11850 6160 17590 6216
rect 17646 6160 17651 6216
rect 11789 6158 17651 6160
rect 11789 6155 11855 6158
rect 17585 6155 17651 6158
rect 18873 6218 18939 6221
rect 22000 6218 22800 6248
rect 18873 6216 22800 6218
rect 18873 6160 18878 6216
rect 18934 6160 22800 6216
rect 18873 6158 22800 6160
rect 18873 6155 18939 6158
rect 22000 6128 22800 6158
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 0 5810 800 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 800 5750
rect 4061 5747 4127 5750
rect 12065 5810 12131 5813
rect 15837 5810 15903 5813
rect 16757 5810 16823 5813
rect 12065 5808 16823 5810
rect 12065 5752 12070 5808
rect 12126 5752 15842 5808
rect 15898 5752 16762 5808
rect 16818 5752 16823 5808
rect 12065 5750 16823 5752
rect 12065 5747 12131 5750
rect 15837 5747 15903 5750
rect 16757 5747 16823 5750
rect 18045 5810 18111 5813
rect 22000 5810 22800 5840
rect 18045 5808 22800 5810
rect 18045 5752 18050 5808
rect 18106 5752 22800 5808
rect 18045 5750 22800 5752
rect 18045 5747 18111 5750
rect 22000 5720 22800 5750
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 18321 5266 18387 5269
rect 22000 5266 22800 5296
rect 18321 5264 22800 5266
rect 18321 5208 18326 5264
rect 18382 5208 22800 5264
rect 18321 5206 22800 5208
rect 18321 5203 18387 5206
rect 22000 5176 22800 5206
rect 7808 4928 8128 4929
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 22000 4858 22800 4888
rect 19014 4798 22800 4858
rect 18045 4586 18111 4589
rect 19014 4586 19074 4798
rect 22000 4768 22800 4798
rect 18045 4584 19074 4586
rect 18045 4528 18050 4584
rect 18106 4528 19074 4584
rect 18045 4526 19074 4528
rect 18045 4523 18111 4526
rect 4376 4384 4696 4385
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 18781 4314 18847 4317
rect 22000 4314 22800 4344
rect 18781 4312 22800 4314
rect 18781 4256 18786 4312
rect 18842 4256 22800 4312
rect 18781 4254 22800 4256
rect 18781 4251 18847 4254
rect 22000 4224 22800 4254
rect 20345 3906 20411 3909
rect 22000 3906 22800 3936
rect 20345 3904 22800 3906
rect 20345 3848 20350 3904
rect 20406 3848 22800 3904
rect 20345 3846 22800 3848
rect 20345 3843 20411 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 22000 3816 22800 3846
rect 14672 3775 14992 3776
rect 19190 3436 19196 3500
rect 19260 3498 19266 3500
rect 22000 3498 22800 3528
rect 19260 3438 22800 3498
rect 19260 3436 19266 3438
rect 22000 3408 22800 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 10225 2954 10291 2957
rect 15561 2954 15627 2957
rect 10225 2952 15627 2954
rect 10225 2896 10230 2952
rect 10286 2896 15566 2952
rect 15622 2896 15627 2952
rect 10225 2894 15627 2896
rect 10225 2891 10291 2894
rect 15561 2891 15627 2894
rect 18413 2954 18479 2957
rect 19006 2954 19012 2956
rect 18413 2952 19012 2954
rect 18413 2896 18418 2952
rect 18474 2896 19012 2952
rect 18413 2894 19012 2896
rect 18413 2891 18479 2894
rect 19006 2892 19012 2894
rect 19076 2954 19082 2956
rect 22000 2954 22800 2984
rect 19076 2894 22800 2954
rect 19076 2892 19082 2894
rect 22000 2864 22800 2894
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 17861 2546 17927 2549
rect 22000 2546 22800 2576
rect 17861 2544 22800 2546
rect 17861 2488 17866 2544
rect 17922 2488 22800 2544
rect 17861 2486 22800 2488
rect 17861 2483 17927 2486
rect 22000 2456 22800 2486
rect 16021 2410 16087 2413
rect 19149 2410 19215 2413
rect 16021 2408 19215 2410
rect 16021 2352 16026 2408
rect 16082 2352 19154 2408
rect 19210 2352 19215 2408
rect 16021 2350 19215 2352
rect 16021 2347 16087 2350
rect 19149 2347 19215 2350
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 18045 2002 18111 2005
rect 22000 2002 22800 2032
rect 18045 2000 22800 2002
rect 18045 1944 18050 2000
rect 18106 1944 22800 2000
rect 18045 1942 22800 1944
rect 18045 1939 18111 1942
rect 22000 1912 22800 1942
rect 10869 1594 10935 1597
rect 13353 1594 13419 1597
rect 22000 1594 22800 1624
rect 10869 1592 22800 1594
rect 10869 1536 10874 1592
rect 10930 1536 13358 1592
rect 13414 1536 22800 1592
rect 10869 1534 22800 1536
rect 10869 1531 10935 1534
rect 13353 1531 13419 1534
rect 22000 1504 22800 1534
rect 16430 988 16436 1052
rect 16500 1050 16506 1052
rect 22000 1050 22800 1080
rect 16500 990 22800 1050
rect 16500 988 16506 990
rect 22000 960 22800 990
rect 12157 642 12223 645
rect 22000 642 22800 672
rect 12157 640 22800 642
rect 12157 584 12162 640
rect 12218 584 22800 640
rect 12157 582 22800 584
rect 12157 579 12223 582
rect 22000 552 22800 582
rect 18822 172 18828 236
rect 18892 234 18898 236
rect 22000 234 22800 264
rect 18892 174 22800 234
rect 18892 172 18898 174
rect 22000 144 22800 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 15516 17172 15580 17236
rect 15148 17036 15212 17100
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 16988 15676 17052 15740
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 19196 14724 19260 14788
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 18644 13424 18708 13428
rect 18644 13368 18694 13424
rect 18694 13368 18708 13424
rect 18644 13364 18708 13368
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 15516 12956 15580 13020
rect 16436 12820 16500 12884
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 16436 12412 16500 12476
rect 16988 12200 17052 12204
rect 16988 12144 17002 12200
rect 17002 12144 17052 12200
rect 16988 12140 17052 12144
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 19012 11656 19076 11660
rect 19012 11600 19026 11656
rect 19026 11600 19076 11656
rect 19012 11596 19076 11600
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 18644 10508 18708 10572
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 15148 10100 15212 10164
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 18828 9284 18892 9348
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 19196 3436 19260 3500
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 19012 2892 19076 2956
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
rect 16436 988 16500 1052
rect 18828 172 18892 236
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 15515 17236 15581 17237
rect 15515 17172 15516 17236
rect 15580 17172 15581 17236
rect 15515 17171 15581 17172
rect 15147 17100 15213 17101
rect 15147 17036 15148 17100
rect 15212 17036 15213 17100
rect 15147 17035 15213 17036
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 15150 10165 15210 17035
rect 15518 13021 15578 17171
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 16987 15740 17053 15741
rect 16987 15676 16988 15740
rect 17052 15676 17053 15740
rect 16987 15675 17053 15676
rect 15515 13020 15581 13021
rect 15515 12956 15516 13020
rect 15580 12956 15581 13020
rect 15515 12955 15581 12956
rect 16435 12884 16501 12885
rect 16435 12820 16436 12884
rect 16500 12820 16501 12884
rect 16435 12819 16501 12820
rect 16438 12477 16498 12819
rect 16435 12476 16501 12477
rect 16435 12412 16436 12476
rect 16500 12412 16501 12476
rect 16435 12411 16501 12412
rect 15147 10164 15213 10165
rect 15147 10100 15148 10164
rect 15212 10100 15213 10164
rect 15147 10099 15213 10100
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 16438 1053 16498 12411
rect 16990 12205 17050 15675
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 19195 14788 19261 14789
rect 19195 14724 19196 14788
rect 19260 14724 19261 14788
rect 19195 14723 19261 14724
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18643 13428 18709 13429
rect 18643 13364 18644 13428
rect 18708 13364 18709 13428
rect 18643 13363 18709 13364
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 16987 12204 17053 12205
rect 16987 12140 16988 12204
rect 17052 12140 17053 12204
rect 16987 12139 17053 12140
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18646 10573 18706 13363
rect 19011 11660 19077 11661
rect 19011 11596 19012 11660
rect 19076 11596 19077 11660
rect 19011 11595 19077 11596
rect 18643 10572 18709 10573
rect 18643 10508 18644 10572
rect 18708 10508 18709 10572
rect 18643 10507 18709 10508
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18827 9348 18893 9349
rect 18827 9284 18828 9348
rect 18892 9284 18893 9348
rect 18827 9283 18893 9284
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
rect 16435 1052 16501 1053
rect 16435 988 16436 1052
rect 16500 988 16501 1052
rect 16435 987 16501 988
rect 18830 237 18890 9283
rect 19014 2957 19074 11595
rect 19198 3501 19258 14723
rect 19195 3500 19261 3501
rect 19195 3436 19196 3500
rect 19260 3436 19261 3500
rect 19195 3435 19261 3436
rect 19011 2956 19077 2957
rect 19011 2892 19012 2956
rect 19076 2892 19077 2956
rect 19011 2891 19077 2892
rect 18827 236 18893 237
rect 18827 172 18828 236
rect 18892 172 18893 236
rect 18827 171 18893 172
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1608761905
transform 1 0 20516 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1608761905
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1608761905
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1608761905
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1608761905
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1608761905
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1608761905
transform 1 0 19964 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1608761905
transform 1 0 19412 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1608761905
transform 1 0 18860 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_191
timestamp 1608761905
transform 1 0 18676 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1608761905
transform 1 0 19228 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_203
timestamp 1608761905
transform 1 0 19780 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1608761905
transform 1 0 17204 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1608761905
transform 1 0 18308 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1608761905
transform 1 0 16652 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1608761905
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_167
timestamp 1608761905
transform 1 0 16468 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_173
timestamp 1608761905
transform 1 0 17020 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_179
timestamp 1608761905
transform 1 0 17572 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_185
timestamp 1608761905
transform 1 0 18124 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1608761905
transform 1 0 14536 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1608761905
transform 1 0 15456 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1608761905
transform 1 0 16100 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1608761905
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_150
timestamp 1608761905
transform 1 0 14904 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_154
timestamp 1608761905
transform 1 0 15272 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_160
timestamp 1608761905
transform 1 0 15824 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1608761905
transform 1 0 13984 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1608761905
transform 1 0 13432 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_129
timestamp 1608761905
transform 1 0 12972 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_133
timestamp 1608761905
transform 1 0 13340 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1608761905
transform 1 0 13800 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_144
timestamp 1608761905
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1608761905
transform 1 0 12604 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1608761905
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1608761905
transform 1 0 10856 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1608761905
transform 1 0 11960 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1608761905
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1608761905
transform 1 0 9108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1608761905
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1608761905
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1608761905
transform 1 0 8004 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1608761905
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1608761905
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1608761905
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1608761905
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1608761905
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1608761905
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1608761905
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1608761905
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1608761905
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1608761905
transform 1 0 20792 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1608761905
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_212
timestamp 1608761905
transform 1 0 20608 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_218
timestamp 1608761905
transform 1 0 21160 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1608761905
transform 1 0 18952 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00
timestamp 1608761905
transform 1 0 19504 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_188
timestamp 1608761905
transform 1 0 18400 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_198
timestamp 1608761905
transform 1 0 19320 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1608761905
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1608761905
transform 1 0 16468 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1608761905
transform 1 0 17020 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1608761905
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_171
timestamp 1608761905
transform 1 0 16836 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_177
timestamp 1608761905
transform 1 0 17388 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1608761905
transform 1 0 15548 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 14628 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_153
timestamp 1608761905
transform 1 0 15180 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1608761905
transform 1 0 15916 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1608761905
transform 1 0 14076 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1608761905
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_145
timestamp 1608761905
transform 1 0 14444 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1608761905
transform 1 0 10948 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1608761905
transform 1 0 11776 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 12420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1608761905
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_106
timestamp 1608761905
transform 1 0 10856 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_111
timestamp 1608761905
transform 1 0 11316 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_115
timestamp 1608761905
transform 1 0 11684 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1608761905
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_98
timestamp 1608761905
transform 1 0 10120 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 8648 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_74
timestamp 1608761905
transform 1 0 7912 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1608761905
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1608761905
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1608761905
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1608761905
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1608761905
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1608761905
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1608761905
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1608761905
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1608761905
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1608761905
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1608761905
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_213
timestamp 1608761905
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1608761905
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1608761905
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1608761905
transform 1 0 19136 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 19596 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 18400 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1608761905
transform 1 0 18952 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_199
timestamp 1608761905
transform 1 0 19412 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_207
timestamp 1608761905
transform 1 0 20148 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1608761905
transform 1 0 17848 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 16928 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_170
timestamp 1608761905
transform 1 0 16744 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_178
timestamp 1608761905
transform 1 0 17480 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_186
timestamp 1608761905
transform 1 0 18216 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 15272 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1608761905
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1608761905
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1608761905
transform 1 0 13984 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1608761905
transform 1 0 14444 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1608761905
transform 1 0 12972 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_127
timestamp 1608761905
transform 1 0 12788 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1608761905
transform 1 0 13800 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_143
timestamp 1608761905
transform 1 0 14260 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 11316 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_109
timestamp 1608761905
transform 1 0 11132 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 9660 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1608761905
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1608761905
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1608761905
transform 1 0 8556 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1608761905
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_80
timestamp 1608761905
transform 1 0 8464 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1608761905
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1608761905
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1608761905
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1608761905
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1608761905
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1608761905
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1608761905
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1608761905
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1608761905
transform 1 0 20516 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1608761905
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_209
timestamp 1608761905
transform 1 0 20332 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1608761905
transform 1 0 20884 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_219
timestamp 1608761905
transform 1 0 21252 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1608761905
transform 1 0 19964 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1608761905
transform 1 0 19412 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_193
timestamp 1608761905
transform 1 0 18860 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_203
timestamp 1608761905
transform 1 0 19780 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1608761905
transform 1 0 17388 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_1_
timestamp 1608761905
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1608761905
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_172
timestamp 1608761905
transform 1 0 16928 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_176
timestamp 1608761905
transform 1 0 17296 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1608761905
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1608761905
transform 1 0 16100 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_161
timestamp 1608761905
transform 1 0 15916 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 12788 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 14444 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_143
timestamp 1608761905
transform 1 0 14260 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 11592 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1608761905
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_112
timestamp 1608761905
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1608761905
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_123
timestamp 1608761905
transform 1 0 12420 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1608761905
transform 1 0 9568 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_1_
timestamp 1608761905
transform 1 0 10580 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_29_89
timestamp 1608761905
transform 1 0 9292 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_101
timestamp 1608761905
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 7820 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 7084 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_71
timestamp 1608761905
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1608761905
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1608761905
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1608761905
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_62
timestamp 1608761905
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1608761905
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1608761905
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1608761905
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1608761905
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1608761905
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1608761905
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1608761905
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1608761905
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1608761905
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 19688 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_28_199
timestamp 1608761905
transform 1 0 19412 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_208
timestamp 1608761905
transform 1 0 20240 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 17940 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_181
timestamp 1608761905
transform 1 0 17756 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1608761905
transform 1 0 14720 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 16284 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1608761905
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1608761905
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_146
timestamp 1608761905
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1608761905
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_163
timestamp 1608761905
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1608761905
transform 1 0 12696 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_1_
timestamp 1608761905
transform 1 0 13708 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_135
timestamp 1608761905
transform 1 0 13524 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 11316 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_109
timestamp 1608761905
transform 1 0 11132 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_117
timestamp 1608761905
transform 1 0 11868 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_125
timestamp 1608761905
transform 1 0 12604 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1608761905
transform 1 0 9844 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l3_in_0_
timestamp 1608761905
transform 1 0 10304 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1608761905
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_86
timestamp 1608761905
transform 1 0 9016 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1608761905
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_98
timestamp 1608761905
transform 1 0 10120 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1608761905
transform 1 0 6992 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_1_
timestamp 1608761905
transform 1 0 8188 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_73
timestamp 1608761905
transform 1 0 7820 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1608761905
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_56
timestamp 1608761905
transform 1 0 6256 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1608761905
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1608761905
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1608761905
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1608761905
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1608761905
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1608761905
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 20516 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608761905
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608761905
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1608761905
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1608761905
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1608761905
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1608761905
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1608761905
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_217
timestamp 1608761905
transform 1 0 21068 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1608761905
transform 1 0 20240 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1608761905
transform 1 0 19228 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 19780 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_1_
timestamp 1608761905
transform 1 0 19136 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1608761905
transform 1 0 18952 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_205
timestamp 1608761905
transform 1 0 19964 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_193
timestamp 1608761905
transform 1 0 18860 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_201
timestamp 1608761905
transform 1 0 19596 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1608761905
transform 1 0 16928 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 17480 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1608761905
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1608761905
transform 1 0 16928 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1608761905
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_170
timestamp 1608761905
transform 1 0 16744 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_176
timestamp 1608761905
transform 1 0 17296 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_168
timestamp 1608761905
transform 1 0 16560 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1608761905
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1608761905
transform 1 0 16376 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1608761905
transform 1 0 15180 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1608761905
transform 1 0 15732 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1608761905
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1608761905
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_150
timestamp 1608761905
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_163
timestamp 1608761905
transform 1 0 16100 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_147
timestamp 1608761905
transform 1 0 14628 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_157
timestamp 1608761905
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l3_in_0_
timestamp 1608761905
transform 1 0 13064 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 14076 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1608761905
transform 1 0 14076 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1608761905
transform 1 0 13616 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_140
timestamp 1608761905
transform 1 0 13984 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_127
timestamp 1608761905
transform 1 0 12788 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_139
timestamp 1608761905
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1608761905
transform 1 0 12512 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 12144 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_3_
timestamp 1608761905
transform 1 0 11316 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1608761905
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_117
timestamp 1608761905
transform 1 0 11868 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_108
timestamp 1608761905
transform 1 0 11040 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1608761905
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1608761905
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 10396 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l3_in_0_
timestamp 1608761905
transform 1 0 9108 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1608761905
transform 1 0 10212 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 9660 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1608761905
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_88
timestamp 1608761905
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_99
timestamp 1608761905
transform 1 0 10212 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_85
timestamp 1608761905
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_96
timestamp 1608761905
transform 1 0 9936 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 6992 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 7452 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 8648 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_80
timestamp 1608761905
transform 1 0 8464 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_68
timestamp 1608761905
transform 1 0 7360 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1608761905
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1608761905
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_56
timestamp 1608761905
transform 1 0 6256 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1608761905
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1608761905
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_62
timestamp 1608761905
transform 1 0 6808 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1608761905
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1608761905
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1608761905
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1608761905
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1608761905
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608761905
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608761905
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1608761905
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1608761905
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1608761905
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1608761905
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 20608 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608761905
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_210
timestamp 1608761905
transform 1 0 20424 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_218
timestamp 1608761905
transform 1 0 21160 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1608761905
transform 1 0 18584 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1608761905
transform 1 0 19596 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_188
timestamp 1608761905
transform 1 0 18400 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_199
timestamp 1608761905
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1608761905
transform 1 0 18032 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1608761905
transform 1 0 16560 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1608761905
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1608761905
transform 1 0 17572 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_177
timestamp 1608761905
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1608761905
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1608761905
transform 1 0 15548 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_155
timestamp 1608761905
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1608761905
transform 1 0 16376 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 13892 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_2_
timestamp 1608761905
transform 1 0 12880 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_127
timestamp 1608761905
transform 1 0 12788 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_137
timestamp 1608761905
transform 1 0 13708 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1608761905
transform 1 0 11132 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1608761905
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_107
timestamp 1608761905
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1608761905
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_123
timestamp 1608761905
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 9476 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_89
timestamp 1608761905
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1608761905
transform 1 0 8464 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_78
timestamp 1608761905
transform 1 0 8280 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 6808 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1608761905
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1608761905
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1608761905
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1608761905
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1608761905
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608761905
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1608761905
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1608761905
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608761905
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1608761905
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_211
timestamp 1608761905
transform 1 0 20516 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1608761905
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1608761905
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1608761905
transform 1 0 19688 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_200
timestamp 1608761905
transform 1 0 19504 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 18032 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_182
timestamp 1608761905
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 16376 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1608761905
transform 1 0 15364 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1608761905
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1608761905
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_154
timestamp 1608761905
transform 1 0 15272 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_164
timestamp 1608761905
transform 1 0 16192 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 13524 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_131
timestamp 1608761905
transform 1 0 13156 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1608761905
transform 1 0 12328 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1608761905
transform 1 0 11316 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_109
timestamp 1608761905
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_120
timestamp 1608761905
transform 1 0 12144 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1608761905
transform 1 0 10304 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1608761905
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1608761905
transform 1 0 10028 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1608761905
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_93
timestamp 1608761905
transform 1 0 9660 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1608761905
transform 1 0 8096 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1608761905
transform 1 0 8556 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_24_73
timestamp 1608761905
transform 1 0 7820 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_79
timestamp 1608761905
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 6348 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1608761905
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_56
timestamp 1608761905
transform 1 0 6256 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1608761905
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1608761905
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1608761905
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608761905
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1608761905
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1608761905
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608761905
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_216
timestamp 1608761905
transform 1 0 20976 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 18492 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1608761905
transform 1 0 20148 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_205
timestamp 1608761905
transform 1 0 19964 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1608761905
transform 1 0 16560 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1608761905
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1608761905
transform 1 0 17388 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1608761905
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1608761905
transform 1 0 17020 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_171
timestamp 1608761905
transform 1 0 16836 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_176
timestamp 1608761905
transform 1 0 17296 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1608761905
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_187
timestamp 1608761905
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1608761905
transform 1 0 15548 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_155
timestamp 1608761905
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1608761905
transform 1 0 16376 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 13892 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1608761905
transform 1 0 12880 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_127
timestamp 1608761905
transform 1 0 12788 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_137
timestamp 1608761905
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1608761905
transform 1 0 11040 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1608761905
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_106
timestamp 1608761905
transform 1 0 10856 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_117
timestamp 1608761905
transform 1 0 11868 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1608761905
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_123
timestamp 1608761905
transform 1 0 12420 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1608761905
transform 1 0 9568 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1608761905
transform 1 0 10028 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_90
timestamp 1608761905
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_95
timestamp 1608761905
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 7912 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_23_71
timestamp 1608761905
transform 1 0 7636 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1608761905
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1608761905
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1608761905
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1608761905
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1608761905
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1608761905
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608761905
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1608761905
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1608761905
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1608761905
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608761905
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1608761905
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1608761905
transform 1 0 20424 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_218
timestamp 1608761905
transform 1 0 21160 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1608761905
transform 1 0 18400 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 18952 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_192
timestamp 1608761905
transform 1 0 18768 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1608761905
transform 1 0 17112 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_22_171
timestamp 1608761905
transform 1 0 16836 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_183
timestamp 1608761905
transform 1 0 17940 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_187
timestamp 1608761905
transform 1 0 18308 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1608761905
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 16284 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1608761905
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1608761905
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_163
timestamp 1608761905
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 12788 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 14444 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1608761905
transform 1 0 14260 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 11132 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1608761905
transform 1 0 10856 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_125
timestamp 1608761905
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1608761905
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 8832 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1608761905
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1608761905
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_102
timestamp 1608761905
transform 1 0 10488 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 6992 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1608761905
transform 1 0 8464 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1608761905
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_56
timestamp 1608761905
transform 1 0 6256 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1608761905
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1608761905
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1608761905
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608761905
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1608761905
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1608761905
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1608761905
transform 1 0 20792 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608761905
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_212
timestamp 1608761905
transform 1 0 20608 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_218
timestamp 1608761905
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 19044 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_1_
timestamp 1608761905
transform 1 0 19780 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_193
timestamp 1608761905
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_201
timestamp 1608761905
transform 1 0 19596 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1608761905
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1608761905
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_179
timestamp 1608761905
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 16100 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1608761905
transform 1 0 15088 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_150
timestamp 1608761905
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_161
timestamp 1608761905
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1608761905
transform 1 0 13616 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1608761905
transform 1 0 14076 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_132
timestamp 1608761905
transform 1 0 13248 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_139
timestamp 1608761905
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1608761905
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1608761905
transform 1 0 11316 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1608761905
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_110
timestamp 1608761905
transform 1 0 11224 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1608761905
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 9200 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_86
timestamp 1608761905
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_104
timestamp 1608761905
transform 1 0 10672 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1608761905
transform 1 0 8188 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_74
timestamp 1608761905
transform 1 0 7912 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1608761905
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1608761905
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1608761905
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1608761905
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1608761905
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1608761905
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608761905
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1608761905
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1608761905
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1608761905
transform 1 0 20700 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608761905
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608761905
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1608761905
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_211
timestamp 1608761905
transform 1 0 20516 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_217
timestamp 1608761905
transform 1 0 21068 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1608761905
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1608761905
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1608761905
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1608761905
transform 1 0 20240 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 19044 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1608761905
transform 1 0 19136 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_193
timestamp 1608761905
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1608761905
transform 1 0 18952 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_205
timestamp 1608761905
transform 1 0 19964 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 16468 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1608761905
transform 1 0 18124 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1608761905
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1608761905
transform 1 0 16744 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1608761905
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_168
timestamp 1608761905
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_179
timestamp 1608761905
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_183
timestamp 1608761905
transform 1 0 17940 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 15088 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1608761905
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1608761905
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_150
timestamp 1608761905
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1608761905
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1608761905
transform 1 0 16100 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 13432 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1608761905
transform 1 0 13432 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 14444 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1608761905
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_132
timestamp 1608761905
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_143
timestamp 1608761905
transform 1 0 14260 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1608761905
transform 1 0 10948 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 11684 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1608761905
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1608761905
transform 1 0 12420 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1608761905
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1608761905
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_105
timestamp 1608761905
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_116
timestamp 1608761905
transform 1 0 11776 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_121
timestamp 1608761905
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 9292 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1608761905
transform 1 0 9752 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1608761905
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1608761905
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_86
timestamp 1608761905
transform 1 0 9016 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_88
timestamp 1608761905
transform 1 0 9200 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1608761905
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_103
timestamp 1608761905
transform 1 0 10580 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1608761905
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1608761905
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_80
timestamp 1608761905
transform 1 0 8464 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1608761905
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1608761905
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1608761905
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1608761905
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1608761905
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1608761905
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1608761905
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1608761905
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1608761905
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1608761905
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1608761905
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608761905
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608761905
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1608761905
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1608761905
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1608761905
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1608761905
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608761905
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1608761905
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1608761905
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1608761905
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1608761905
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1608761905
transform 1 0 20240 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 18584 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_206
timestamp 1608761905
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1608761905
transform 1 0 16744 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 17756 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_168
timestamp 1608761905
transform 1 0 16560 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_179
timestamp 1608761905
transform 1 0 17572 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_187
timestamp 1608761905
transform 1 0 18308 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1608761905
transform 1 0 14720 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1608761905
transform 1 0 15732 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1608761905
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1608761905
transform 1 0 15456 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_146
timestamp 1608761905
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1608761905
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1608761905
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 13064 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_128
timestamp 1608761905
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 11408 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_18_106
timestamp 1608761905
transform 1 0 10856 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1608761905
transform 1 0 10028 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1608761905
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_93
timestamp 1608761905
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1608761905
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1608761905
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1608761905
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1608761905
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1608761905
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1608761905
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1608761905
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608761905
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1608761905
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1608761905
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 20608 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608761905
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_210
timestamp 1608761905
transform 1 0 20424 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_218
timestamp 1608761905
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1608761905
transform 1 0 19596 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1608761905
transform 1 0 18584 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_188
timestamp 1608761905
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_199
timestamp 1608761905
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1608761905
transform 1 0 18124 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1608761905
transform 1 0 17388 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1608761905
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1608761905
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_180
timestamp 1608761905
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_184
timestamp 1608761905
transform 1 0 18032 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 15732 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_17_153
timestamp 1608761905
transform 1 0 15180 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1608761905
transform 1 0 13524 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1608761905
transform 1 0 14352 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_133
timestamp 1608761905
transform 1 0 13340 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1608761905
transform 1 0 11408 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1608761905
transform 1 0 12512 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608761905
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1608761905
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_115
timestamp 1608761905
transform 1 0 11684 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1608761905
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_123
timestamp 1608761905
transform 1 0 12420 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1608761905
transform 1 0 10396 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_99
timestamp 1608761905
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 8740 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_17_74
timestamp 1608761905
transform 1 0 7912 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_82
timestamp 1608761905
transform 1 0 8648 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608761905
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1608761905
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1608761905
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1608761905
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1608761905
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1608761905
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608761905
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1608761905
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1608761905
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608761905
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608761905
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1608761905
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1608761905
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1608761905
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 19136 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 18400 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1608761905
transform 1 0 18952 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 16560 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_167
timestamp 1608761905
transform 1 0 16468 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_184
timestamp 1608761905
transform 1 0 18032 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1608761905
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608761905
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1608761905
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_163
timestamp 1608761905
transform 1 0 16100 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk
timestamp 1608761905
transform 1 0 12972 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_16_128
timestamp 1608761905
transform 1 0 12880 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 10856 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_105
timestamp 1608761905
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_122
timestamp 1608761905
transform 1 0 12328 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 9660 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608761905
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1608761905
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_99
timestamp 1608761905
transform 1 0 10212 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 7912 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_16_68
timestamp 1608761905
transform 1 0 7360 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1608761905
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1608761905
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608761905
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1608761905
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1608761905
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608761905
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1608761905
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1608761905
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608761905
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_218
timestamp 1608761905
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1608761905
transform 1 0 19044 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 19688 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_193
timestamp 1608761905
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1608761905
transform 1 0 19320 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1608761905
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608761905
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1608761905
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 16284 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1608761905
transform 1 0 15272 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_163
timestamp 1608761905
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1608761905
transform 1 0 13340 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1608761905
transform 1 0 14444 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_142
timestamp 1608761905
transform 1 0 14168 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1608761905
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1608761905
transform 1 0 10856 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1608761905
transform 1 0 12512 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608761905
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_115
timestamp 1608761905
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_123
timestamp 1608761905
transform 1 0 12420 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1608761905
transform 1 0 9844 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_93
timestamp 1608761905
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_104
timestamp 1608761905
transform 1 0 10672 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 8188 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_15_74
timestamp 1608761905
transform 1 0 7912 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608761905
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1608761905
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1608761905
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1608761905
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1608761905
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1608761905
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608761905
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1608761905
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1608761905
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1608761905
transform 1 0 20792 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608761905
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608761905
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608761905
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_212
timestamp 1608761905
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_217
timestamp 1608761905
transform 1 0 21068 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1608761905
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1608761905
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 19136 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1608761905
transform 1 0 19228 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_13_193
timestamp 1608761905
transform 1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_191
timestamp 1608761905
transform 1 0 18676 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_206
timestamp 1608761905
transform 1 0 20056 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1608761905
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1608761905
transform 1 0 16836 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1608761905
transform 1 0 17848 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608761905
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_174
timestamp 1608761905
transform 1 0 17112 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1608761905
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_180
timestamp 1608761905
transform 1 0 17664 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 14628 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1608761905
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1608761905
transform 1 0 16284 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608761905
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_163
timestamp 1608761905
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1608761905
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_163
timestamp 1608761905
transform 1 0 16100 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1608761905
transform 1 0 14168 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1608761905
transform 1 0 14168 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1608761905
transform 1 0 13156 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_140
timestamp 1608761905
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_145
timestamp 1608761905
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_140
timestamp 1608761905
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 12512 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 11592 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608761905
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_112
timestamp 1608761905
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1608761905
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_123
timestamp 1608761905
transform 1 0 12420 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_119
timestamp 1608761905
transform 1 0 12052 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 9936 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 10580 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_14_96
timestamp 1608761905
transform 1 0 9936 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_102
timestamp 1608761905
transform 1 0 10488 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1608761905
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608761905
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1608761905
transform 1 0 9660 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_88
timestamp 1608761905
transform 1 0 9200 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_92
timestamp 1608761905
transform 1 0 9568 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1608761905
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 7728 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1608761905
transform 1 0 8556 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_70
timestamp 1608761905
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1608761905
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_80
timestamp 1608761905
transform 1 0 8464 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608761905
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1608761905
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1608761905
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_62
timestamp 1608761905
transform 1 0 6808 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1608761905
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1608761905
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608761905
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1608761905
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1608761905
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1608761905
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1608761905
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608761905
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608761905
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1608761905
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1608761905
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1608761905
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1608761905
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608761905
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608761905
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1608761905
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1608761905
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1608761905
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 19136 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1608761905
transform 1 0 18952 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 17480 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1608761905
transform 1 0 16560 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_167
timestamp 1608761905
transform 1 0 16468 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_171
timestamp 1608761905
transform 1 0 16836 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_177
timestamp 1608761905
transform 1 0 17388 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1608761905
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608761905
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1608761905
transform 1 0 14536 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1608761905
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_163
timestamp 1608761905
transform 1 0 16100 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1608761905
transform 1 0 12880 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1608761905
transform 1 0 13524 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_126
timestamp 1608761905
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_131
timestamp 1608761905
transform 1 0 13156 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_144
timestamp 1608761905
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1608761905
transform 1 0 11868 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1608761905
transform 1 0 10856 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_115
timestamp 1608761905
transform 1 0 11684 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1608761905
transform 1 0 9844 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608761905
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1608761905
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1608761905
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_104
timestamp 1608761905
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1608761905
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1608761905
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_80
timestamp 1608761905
transform 1 0 8464 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1608761905
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1608761905
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608761905
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1608761905
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1608761905
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608761905
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1608761905
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1608761905
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608761905
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_215
timestamp 1608761905
transform 1 0 20884 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_219
timestamp 1608761905
transform 1 0 21252 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1608761905
transform 1 0 20056 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1608761905
transform 1 0 19044 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1608761905
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_204
timestamp 1608761905
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1608761905
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608761905
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_177
timestamp 1608761905
transform 1 0 17388 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 15916 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1608761905
transform 1 0 15088 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_146
timestamp 1608761905
transform 1 0 14536 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_155
timestamp 1608761905
transform 1 0 15364 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 13064 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_128
timestamp 1608761905
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 11500 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608761905
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1608761905
transform 1 0 12604 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_111
timestamp 1608761905
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_119
timestamp 1608761905
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1608761905
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 9844 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_91
timestamp 1608761905
transform 1 0 9476 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 8004 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_74
timestamp 1608761905
transform 1 0 7912 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608761905
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1608761905
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1608761905
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1608761905
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1608761905
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1608761905
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608761905
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1608761905
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1608761905
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1608761905
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608761905
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608761905
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_210
timestamp 1608761905
transform 1 0 20424 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_218
timestamp 1608761905
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1608761905
transform 1 0 19596 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_189
timestamp 1608761905
transform 1 0 18492 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1608761905
transform 1 0 17204 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1608761905
transform 1 0 17664 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_173
timestamp 1608761905
transform 1 0 17020 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_178
timestamp 1608761905
transform 1 0 17480 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 15548 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608761905
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_147
timestamp 1608761905
transform 1 0 14628 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_154
timestamp 1608761905
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1608761905
transform 1 0 13800 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1608761905
transform 1 0 12788 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_136
timestamp 1608761905
transform 1 0 13616 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 11132 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_107
timestamp 1608761905
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_125
timestamp 1608761905
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1608761905
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1608761905
transform 1 0 10120 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608761905
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1608761905
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_96
timestamp 1608761905
transform 1 0 9936 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1608761905
transform 1 0 8556 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1608761905
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_80
timestamp 1608761905
transform 1 0 8464 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1608761905
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1608761905
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608761905
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1608761905
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1608761905
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608761905
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1608761905
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1608761905
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1608761905
transform 1 0 20424 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608761905
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_214
timestamp 1608761905
transform 1 0 20792 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 18768 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_208
timestamp 1608761905
transform 1 0 20240 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608761905
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1608761905
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_184
timestamp 1608761905
transform 1 0 18032 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 16284 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1608761905
transform 1 0 15272 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_152
timestamp 1608761905
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_163
timestamp 1608761905
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 13616 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_134
timestamp 1608761905
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1608761905
transform 1 0 12604 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1608761905
transform 1 0 11316 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608761905
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_110
timestamp 1608761905
transform 1 0 11224 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1608761905
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1608761905
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 9200 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_86
timestamp 1608761905
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_104
timestamp 1608761905
transform 1 0 10672 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1608761905
transform 1 0 8188 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_74
timestamp 1608761905
transform 1 0 7912 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608761905
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1608761905
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1608761905
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1608761905
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1608761905
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1608761905
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608761905
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1608761905
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1608761905
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608761905
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608761905
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1608761905
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1608761905
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1608761905
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1608761905
transform 1 0 19780 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1608761905
transform 1 0 18768 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_190
timestamp 1608761905
transform 1 0 18584 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_201
timestamp 1608761905
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1608761905
transform 1 0 18216 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1608761905
transform 1 0 17204 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_173
timestamp 1608761905
transform 1 0 17020 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_184
timestamp 1608761905
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1608761905
transform 1 0 16192 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608761905
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_147
timestamp 1608761905
transform 1 0 14628 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_154
timestamp 1608761905
transform 1 0 15272 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_162
timestamp 1608761905
transform 1 0 16008 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1608761905
transform 1 0 13340 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1608761905
transform 1 0 13800 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_126
timestamp 1608761905
transform 1 0 12696 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_132
timestamp 1608761905
transform 1 0 13248 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_136
timestamp 1608761905
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 11224 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_8_107
timestamp 1608761905
transform 1 0 10948 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1608761905
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608761905
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1608761905
transform 1 0 10672 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1608761905
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1608761905
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 7912 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_8_68
timestamp 1608761905
transform 1 0 7360 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1608761905
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1608761905
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608761905
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1608761905
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1608761905
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608761905
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1608761905
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1608761905
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1608761905
transform 1 0 20792 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608761905
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608761905
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608761905
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_210
timestamp 1608761905
transform 1 0 20424 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1608761905
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1608761905
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_212
timestamp 1608761905
transform 1 0 20608 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_218
timestamp 1608761905
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 18952 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 19136 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_6_190
timestamp 1608761905
transform 1 0 18584 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_194
timestamp 1608761905
transform 1 0 18952 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1608761905
transform 1 0 16560 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 17112 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1608761905
transform 1 0 16836 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1608761905
transform 1 0 18124 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608761905
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_172
timestamp 1608761905
transform 1 0 16928 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1608761905
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_180
timestamp 1608761905
transform 1 0 17664 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_184
timestamp 1608761905
transform 1 0 18032 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1608761905
transform 1 0 14720 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1608761905
transform 1 0 15824 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1608761905
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1608761905
transform 1 0 14812 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608761905
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1608761905
transform 1 0 16284 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1608761905
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_163
timestamp 1608761905
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_158
timestamp 1608761905
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1608761905
transform 1 0 13248 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1608761905
transform 1 0 13524 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_133
timestamp 1608761905
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_144
timestamp 1608761905
transform 1 0 14352 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_126
timestamp 1608761905
transform 1 0 12696 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_141
timestamp 1608761905
transform 1 0 14076 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1608761905
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 10856 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1608761905
transform 1 0 12512 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1608761905
transform 1 0 11132 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608761905
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_122
timestamp 1608761905
transform 1 0 12328 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_107
timestamp 1608761905
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1608761905
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1608761905
transform 1 0 10120 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_6_102
timestamp 1608761905
transform 1 0 10488 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_96
timestamp 1608761905
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1608761905
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1608761905
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1608761905
transform 1 0 9108 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608761905
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_84
timestamp 1608761905
transform 1 0 8832 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1608761905
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_85
timestamp 1608761905
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 7452 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_6_72
timestamp 1608761905
transform 1 0 7728 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_68
timestamp 1608761905
transform 1 0 7360 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 6256 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608761905
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1608761905
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1608761905
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1608761905
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_62
timestamp 1608761905
transform 1 0 6808 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608761905
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608761905
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1608761905
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1608761905
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1608761905
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608761905
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608761905
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1608761905
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1608761905
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1608761905
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1608761905
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1608761905
transform 1 0 20884 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608761905
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_213
timestamp 1608761905
transform 1 0 20700 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_218
timestamp 1608761905
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1608761905
transform 1 0 19872 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_202
timestamp 1608761905
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 18216 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1608761905
transform 1 0 16744 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608761905
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_168
timestamp 1608761905
transform 1 0 16560 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_179
timestamp 1608761905
transform 1 0 17572 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_184
timestamp 1608761905
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 15088 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_150
timestamp 1608761905
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 13432 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_132
timestamp 1608761905
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1608761905
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1608761905
transform 1 0 11316 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608761905
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_110
timestamp 1608761905
transform 1 0 11224 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1608761905
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1608761905
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1608761905
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1608761905
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608761905
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1608761905
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1608761905
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1608761905
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1608761905
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1608761905
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608761905
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608761905
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1608761905
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1608761905
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608761905
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608761905
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1608761905
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_218
timestamp 1608761905
transform 1 0 21160 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1608761905
transform 1 0 18952 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1608761905
transform 1 0 19780 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_192
timestamp 1608761905
transform 1 0 18768 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_198
timestamp 1608761905
transform 1 0 19320 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_202
timestamp 1608761905
transform 1 0 19688 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 17296 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_174
timestamp 1608761905
transform 1 0 17112 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1608761905
transform 1 0 14628 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 15640 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608761905
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1608761905
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_154
timestamp 1608761905
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1608761905
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_134
timestamp 1608761905
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_145
timestamp 1608761905
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608761905
transform 1 0 11960 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1608761905
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_117
timestamp 1608761905
transform 1 0 11868 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608761905
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1608761905
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1608761905
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1608761905
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1608761905
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1608761905
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608761905
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1608761905
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1608761905
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608761905
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1608761905
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1608761905
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1608761905
transform 1 0 20608 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608761905
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_210
timestamp 1608761905
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_216
timestamp 1608761905
transform 1 0 20976 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1608761905
transform 1 0 19596 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1608761905
transform 1 0 18584 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_188
timestamp 1608761905
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_199
timestamp 1608761905
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1608761905
transform 1 0 17204 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1608761905
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608761905
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_173
timestamp 1608761905
transform 1 0 17020 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_179
timestamp 1608761905
transform 1 0 17572 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1608761905
transform 1 0 14720 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1608761905
transform 1 0 15180 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1608761905
transform 1 0 16192 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_146
timestamp 1608761905
transform 1 0 14536 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_151
timestamp 1608761905
transform 1 0 14996 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_162
timestamp 1608761905
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1608761905
transform 1 0 14168 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 13432 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1608761905
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_140
timestamp 1608761905
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 11592 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1608761905
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608761905
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1608761905
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 9016 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_3_102
timestamp 1608761905
transform 1 0 10488 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1608761905
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608761905
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1608761905
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1608761905
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1608761905
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1608761905
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1608761905
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608761905
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608761905
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1608761905
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1608761905
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608761905
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608761905
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_210
timestamp 1608761905
transform 1 0 20424 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_218
timestamp 1608761905
transform 1 0 21160 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1608761905
transform 1 0 20056 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 18400 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_204
timestamp 1608761905
transform 1 0 19872 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 16744 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_2_169
timestamp 1608761905
transform 1 0 16652 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_186
timestamp 1608761905
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1608761905
transform 1 0 15456 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608761905
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1608761905
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1608761905
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_165
timestamp 1608761905
transform 1 0 16284 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1608761905
transform 1 0 14444 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 12696 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1608761905
transform 1 0 13432 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_132
timestamp 1608761905
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_143
timestamp 1608761905
transform 1 0 14260 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 11040 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_106
timestamp 1608761905
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_124
timestamp 1608761905
transform 1 0 12512 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1608761905
transform 1 0 10580 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608761905
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_93
timestamp 1608761905
transform 1 0 9660 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101
timestamp 1608761905
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1608761905
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1608761905
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1608761905
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1608761905
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608761905
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1608761905
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608761905
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608761905
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1608761905
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1608761905
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608761905
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608761905
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_219
timestamp 1608761905
transform 1 0 21252 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608761905
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_214
timestamp 1608761905
transform 1 0 20792 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1608761905
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1608761905
transform 1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1608761905
transform 1 0 20424 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1608761905
transform 1 0 20516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1608761905
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1608761905
transform 1 0 19320 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1608761905
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 19044 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 19780 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1608761905
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_196
timestamp 1608761905
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_202
timestamp 1608761905
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_208
timestamp 1608761905
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_201
timestamp 1608761905
transform 1 0 19596 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1608761905
transform 1 0 17480 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1608761905
transform 1 0 16468 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1608761905
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1608761905
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608761905
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608761905
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_176
timestamp 1608761905
transform 1 0 17296 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1608761905
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1608761905
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608761905
transform 1 0 14628 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 16284 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 15732 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608761905
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1608761905
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_156
timestamp 1608761905
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1608761905
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_163
timestamp 1608761905
transform 1 0 16100 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 12972 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608761905
transform 1 0 12880 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1608761905
transform 1 0 13984 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134
timestamp 1608761905
transform 1 0 13432 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_127
timestamp 1608761905
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_145
timestamp 1608761905
transform 1 0 14444 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608761905
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125
timestamp 1608761905
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1608761905
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1608761905
transform 1 0 11776 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608761905
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1608761905
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1608761905
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1608761905
transform 1 0 11316 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_109
timestamp 1608761905
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 1608761905
transform 1 0 11500 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1608761905
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608761905
transform 1 0 10028 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1608761905
transform 1 0 10304 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608761905
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1608761905
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_98
timestamp 1608761905
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_86
timestamp 1608761905
transform 1 0 9016 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_94
timestamp 1608761905
transform 1 0 9752 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1608761905
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1608761905
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1608761905
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608761905
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608761905
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608761905
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56
timestamp 1608761905
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51
timestamp 1608761905
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1608761905
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1608761905
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608761905
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1608761905
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608761905
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1608761905
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1608761905
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608761905
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1608761905
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608761905
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608761905
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1608761905
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1608761905
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
<< labels >>
rlabel metal2 s 294 0 350 800 4 bottom_left_grid_pin_1_
port 1 nsew
rlabel metal3 s 0 5720 800 5840 4 ccff_head
port 2 nsew
rlabel metal3 s 0 17144 800 17264 4 ccff_tail
port 3 nsew
rlabel metal3 s 22000 3816 22800 3936 4 chanx_right_in[0]
port 4 nsew
rlabel metal3 s 22000 8440 22800 8560 4 chanx_right_in[10]
port 5 nsew
rlabel metal3 s 22000 8984 22800 9104 4 chanx_right_in[11]
port 6 nsew
rlabel metal3 s 22000 9392 22800 9512 4 chanx_right_in[12]
port 7 nsew
rlabel metal3 s 22000 9936 22800 10056 4 chanx_right_in[13]
port 8 nsew
rlabel metal3 s 22000 10344 22800 10464 4 chanx_right_in[14]
port 9 nsew
rlabel metal3 s 22000 10752 22800 10872 4 chanx_right_in[15]
port 10 nsew
rlabel metal3 s 22000 11296 22800 11416 4 chanx_right_in[16]
port 11 nsew
rlabel metal3 s 22000 11704 22800 11824 4 chanx_right_in[17]
port 12 nsew
rlabel metal3 s 22000 12248 22800 12368 4 chanx_right_in[18]
port 13 nsew
rlabel metal3 s 22000 12656 22800 12776 4 chanx_right_in[19]
port 14 nsew
rlabel metal3 s 22000 4224 22800 4344 4 chanx_right_in[1]
port 15 nsew
rlabel metal3 s 22000 4768 22800 4888 4 chanx_right_in[2]
port 16 nsew
rlabel metal3 s 22000 5176 22800 5296 4 chanx_right_in[3]
port 17 nsew
rlabel metal3 s 22000 5720 22800 5840 4 chanx_right_in[4]
port 18 nsew
rlabel metal3 s 22000 6128 22800 6248 4 chanx_right_in[5]
port 19 nsew
rlabel metal3 s 22000 6672 22800 6792 4 chanx_right_in[6]
port 20 nsew
rlabel metal3 s 22000 7080 22800 7200 4 chanx_right_in[7]
port 21 nsew
rlabel metal3 s 22000 7488 22800 7608 4 chanx_right_in[8]
port 22 nsew
rlabel metal3 s 22000 8032 22800 8152 4 chanx_right_in[9]
port 23 nsew
rlabel metal3 s 22000 13200 22800 13320 4 chanx_right_out[0]
port 24 nsew
rlabel metal3 s 22000 17824 22800 17944 4 chanx_right_out[10]
port 25 nsew
rlabel metal3 s 22000 18232 22800 18352 4 chanx_right_out[11]
port 26 nsew
rlabel metal3 s 22000 18776 22800 18896 4 chanx_right_out[12]
port 27 nsew
rlabel metal3 s 22000 19184 22800 19304 4 chanx_right_out[13]
port 28 nsew
rlabel metal3 s 22000 19728 22800 19848 4 chanx_right_out[14]
port 29 nsew
rlabel metal3 s 22000 20136 22800 20256 4 chanx_right_out[15]
port 30 nsew
rlabel metal3 s 22000 20544 22800 20664 4 chanx_right_out[16]
port 31 nsew
rlabel metal3 s 22000 21088 22800 21208 4 chanx_right_out[17]
port 32 nsew
rlabel metal3 s 22000 21496 22800 21616 4 chanx_right_out[18]
port 33 nsew
rlabel metal3 s 22000 22040 22800 22160 4 chanx_right_out[19]
port 34 nsew
rlabel metal3 s 22000 13608 22800 13728 4 chanx_right_out[1]
port 35 nsew
rlabel metal3 s 22000 14016 22800 14136 4 chanx_right_out[2]
port 36 nsew
rlabel metal3 s 22000 14560 22800 14680 4 chanx_right_out[3]
port 37 nsew
rlabel metal3 s 22000 14968 22800 15088 4 chanx_right_out[4]
port 38 nsew
rlabel metal3 s 22000 15512 22800 15632 4 chanx_right_out[5]
port 39 nsew
rlabel metal3 s 22000 15920 22800 16040 4 chanx_right_out[6]
port 40 nsew
rlabel metal3 s 22000 16464 22800 16584 4 chanx_right_out[7]
port 41 nsew
rlabel metal3 s 22000 16872 22800 16992 4 chanx_right_out[8]
port 42 nsew
rlabel metal3 s 22000 17280 22800 17400 4 chanx_right_out[9]
port 43 nsew
rlabel metal2 s 846 0 902 800 4 chany_bottom_in[0]
port 44 nsew
rlabel metal2 s 6366 0 6422 800 4 chany_bottom_in[10]
port 45 nsew
rlabel metal2 s 6918 0 6974 800 4 chany_bottom_in[11]
port 46 nsew
rlabel metal2 s 7470 0 7526 800 4 chany_bottom_in[12]
port 47 nsew
rlabel metal2 s 8022 0 8078 800 4 chany_bottom_in[13]
port 48 nsew
rlabel metal2 s 8574 0 8630 800 4 chany_bottom_in[14]
port 49 nsew
rlabel metal2 s 9126 0 9182 800 4 chany_bottom_in[15]
port 50 nsew
rlabel metal2 s 9678 0 9734 800 4 chany_bottom_in[16]
port 51 nsew
rlabel metal2 s 10230 0 10286 800 4 chany_bottom_in[17]
port 52 nsew
rlabel metal2 s 10782 0 10838 800 4 chany_bottom_in[18]
port 53 nsew
rlabel metal2 s 11334 0 11390 800 4 chany_bottom_in[19]
port 54 nsew
rlabel metal2 s 1398 0 1454 800 4 chany_bottom_in[1]
port 55 nsew
rlabel metal2 s 1950 0 2006 800 4 chany_bottom_in[2]
port 56 nsew
rlabel metal2 s 2502 0 2558 800 4 chany_bottom_in[3]
port 57 nsew
rlabel metal2 s 3054 0 3110 800 4 chany_bottom_in[4]
port 58 nsew
rlabel metal2 s 3606 0 3662 800 4 chany_bottom_in[5]
port 59 nsew
rlabel metal2 s 4158 0 4214 800 4 chany_bottom_in[6]
port 60 nsew
rlabel metal2 s 4710 0 4766 800 4 chany_bottom_in[7]
port 61 nsew
rlabel metal2 s 5262 0 5318 800 4 chany_bottom_in[8]
port 62 nsew
rlabel metal2 s 5814 0 5870 800 4 chany_bottom_in[9]
port 63 nsew
rlabel metal2 s 11978 0 12034 800 4 chany_bottom_out[0]
port 64 nsew
rlabel metal2 s 17498 0 17554 800 4 chany_bottom_out[10]
port 65 nsew
rlabel metal2 s 18050 0 18106 800 4 chany_bottom_out[11]
port 66 nsew
rlabel metal2 s 18602 0 18658 800 4 chany_bottom_out[12]
port 67 nsew
rlabel metal2 s 19154 0 19210 800 4 chany_bottom_out[13]
port 68 nsew
rlabel metal2 s 19706 0 19762 800 4 chany_bottom_out[14]
port 69 nsew
rlabel metal2 s 20258 0 20314 800 4 chany_bottom_out[15]
port 70 nsew
rlabel metal2 s 20810 0 20866 800 4 chany_bottom_out[16]
port 71 nsew
rlabel metal2 s 21362 0 21418 800 4 chany_bottom_out[17]
port 72 nsew
rlabel metal2 s 21914 0 21970 800 4 chany_bottom_out[18]
port 73 nsew
rlabel metal2 s 22466 0 22522 800 4 chany_bottom_out[19]
port 74 nsew
rlabel metal2 s 12530 0 12586 800 4 chany_bottom_out[1]
port 75 nsew
rlabel metal2 s 13082 0 13138 800 4 chany_bottom_out[2]
port 76 nsew
rlabel metal2 s 13634 0 13690 800 4 chany_bottom_out[3]
port 77 nsew
rlabel metal2 s 14186 0 14242 800 4 chany_bottom_out[4]
port 78 nsew
rlabel metal2 s 14738 0 14794 800 4 chany_bottom_out[5]
port 79 nsew
rlabel metal2 s 15290 0 15346 800 4 chany_bottom_out[6]
port 80 nsew
rlabel metal2 s 15842 0 15898 800 4 chany_bottom_out[7]
port 81 nsew
rlabel metal2 s 16394 0 16450 800 4 chany_bottom_out[8]
port 82 nsew
rlabel metal2 s 16946 0 17002 800 4 chany_bottom_out[9]
port 83 nsew
rlabel metal2 s 846 22000 902 22800 4 chany_top_in[0]
port 84 nsew
rlabel metal2 s 6366 22000 6422 22800 4 chany_top_in[10]
port 85 nsew
rlabel metal2 s 6918 22000 6974 22800 4 chany_top_in[11]
port 86 nsew
rlabel metal2 s 7470 22000 7526 22800 4 chany_top_in[12]
port 87 nsew
rlabel metal2 s 8022 22000 8078 22800 4 chany_top_in[13]
port 88 nsew
rlabel metal2 s 8574 22000 8630 22800 4 chany_top_in[14]
port 89 nsew
rlabel metal2 s 9126 22000 9182 22800 4 chany_top_in[15]
port 90 nsew
rlabel metal2 s 9678 22000 9734 22800 4 chany_top_in[16]
port 91 nsew
rlabel metal2 s 10230 22000 10286 22800 4 chany_top_in[17]
port 92 nsew
rlabel metal2 s 10782 22000 10838 22800 4 chany_top_in[18]
port 93 nsew
rlabel metal2 s 11334 22000 11390 22800 4 chany_top_in[19]
port 94 nsew
rlabel metal2 s 1398 22000 1454 22800 4 chany_top_in[1]
port 95 nsew
rlabel metal2 s 1950 22000 2006 22800 4 chany_top_in[2]
port 96 nsew
rlabel metal2 s 2502 22000 2558 22800 4 chany_top_in[3]
port 97 nsew
rlabel metal2 s 3054 22000 3110 22800 4 chany_top_in[4]
port 98 nsew
rlabel metal2 s 3606 22000 3662 22800 4 chany_top_in[5]
port 99 nsew
rlabel metal2 s 4158 22000 4214 22800 4 chany_top_in[6]
port 100 nsew
rlabel metal2 s 4710 22000 4766 22800 4 chany_top_in[7]
port 101 nsew
rlabel metal2 s 5262 22000 5318 22800 4 chany_top_in[8]
port 102 nsew
rlabel metal2 s 5814 22000 5870 22800 4 chany_top_in[9]
port 103 nsew
rlabel metal2 s 11978 22000 12034 22800 4 chany_top_out[0]
port 104 nsew
rlabel metal2 s 17498 22000 17554 22800 4 chany_top_out[10]
port 105 nsew
rlabel metal2 s 18050 22000 18106 22800 4 chany_top_out[11]
port 106 nsew
rlabel metal2 s 18602 22000 18658 22800 4 chany_top_out[12]
port 107 nsew
rlabel metal2 s 19154 22000 19210 22800 4 chany_top_out[13]
port 108 nsew
rlabel metal2 s 19706 22000 19762 22800 4 chany_top_out[14]
port 109 nsew
rlabel metal2 s 20258 22000 20314 22800 4 chany_top_out[15]
port 110 nsew
rlabel metal2 s 20810 22000 20866 22800 4 chany_top_out[16]
port 111 nsew
rlabel metal2 s 21362 22000 21418 22800 4 chany_top_out[17]
port 112 nsew
rlabel metal2 s 21914 22000 21970 22800 4 chany_top_out[18]
port 113 nsew
rlabel metal2 s 22466 22000 22522 22800 4 chany_top_out[19]
port 114 nsew
rlabel metal2 s 12530 22000 12586 22800 4 chany_top_out[1]
port 115 nsew
rlabel metal2 s 13082 22000 13138 22800 4 chany_top_out[2]
port 116 nsew
rlabel metal2 s 13634 22000 13690 22800 4 chany_top_out[3]
port 117 nsew
rlabel metal2 s 14186 22000 14242 22800 4 chany_top_out[4]
port 118 nsew
rlabel metal2 s 14738 22000 14794 22800 4 chany_top_out[5]
port 119 nsew
rlabel metal2 s 15290 22000 15346 22800 4 chany_top_out[6]
port 120 nsew
rlabel metal2 s 15842 22000 15898 22800 4 chany_top_out[7]
port 121 nsew
rlabel metal2 s 16394 22000 16450 22800 4 chany_top_out[8]
port 122 nsew
rlabel metal2 s 16946 22000 17002 22800 4 chany_top_out[9]
port 123 nsew
rlabel metal3 s 22000 22448 22800 22568 4 prog_clk_0_E_in
port 124 nsew
rlabel metal3 s 22000 144 22800 264 4 right_bottom_grid_pin_34_
port 125 nsew
rlabel metal3 s 22000 552 22800 672 4 right_bottom_grid_pin_35_
port 126 nsew
rlabel metal3 s 22000 960 22800 1080 4 right_bottom_grid_pin_36_
port 127 nsew
rlabel metal3 s 22000 1504 22800 1624 4 right_bottom_grid_pin_37_
port 128 nsew
rlabel metal3 s 22000 1912 22800 2032 4 right_bottom_grid_pin_38_
port 129 nsew
rlabel metal3 s 22000 2456 22800 2576 4 right_bottom_grid_pin_39_
port 130 nsew
rlabel metal3 s 22000 2864 22800 2984 4 right_bottom_grid_pin_40_
port 131 nsew
rlabel metal3 s 22000 3408 22800 3528 4 right_bottom_grid_pin_41_
port 132 nsew
rlabel metal2 s 294 22000 350 22800 4 top_left_grid_pin_1_
port 133 nsew
rlabel metal4 s 4376 2128 4696 20176 4 VPWR
port 134 nsew
rlabel metal4 s 7808 2128 8128 20176 4 VGND
port 135 nsew
<< properties >>
string FIXED_BBOX 0 0 22800 22800
string GDS_FILE /ef/openfpga/openlane/runs/sb_0__1_/results/magic/sb_0__1_.gds
string GDS_END 1098906
string GDS_START 81916
<< end >>
