* NGSPICE file created from cbx_1__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand3_4 abstract view
.subckt scs8hd_nand3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

.subckt cbx_1__0_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_grid_pin_0_ bottom_grid_pin_10_ bottom_grid_pin_12_ bottom_grid_pin_14_
+ bottom_grid_pin_2_ bottom_grid_pin_4_ bottom_grid_pin_6_ bottom_grid_pin_8_ chanx_left_in[0]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_right_in[0] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ data_in enable top_grid_pin_14_ top_grid_pin_2_ top_grid_pin_6_ vpwr vgnd
XFILLER_18_406 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_199 vpwr vgnd scs8hd_fill_2
XFILLER_13_177 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_0_.latch/Q mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_148 vpwr vgnd scs8hd_fill_2
XANTENNA__113__B _108_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_12 vpwr vgnd scs8hd_fill_2
XFILLER_3_34 vgnd vpwr scs8hd_decap_3
XFILLER_3_56 vgnd vpwr scs8hd_decap_3
XFILLER_5_332 vpwr vgnd scs8hd_fill_2
XFILLER_5_365 vgnd vpwr scs8hd_fill_1
XFILLER_5_376 vpwr vgnd scs8hd_fill_2
XFILLER_8_181 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_2.LATCH_1_.latch data_in mem_bottom_ipin_2.LATCH_1_.latch/Q _169_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_125 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_3.LATCH_3_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_269 vgnd vpwr scs8hd_decap_6
XANTENNA__124__A _124_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_4.LATCH_3_.latch/Q mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _154_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_200_ chanx_left_in[7] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
X_131_ _102_/X _126_/X _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_176 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_261 vgnd vpwr scs8hd_decap_4
XANTENNA__119__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_22 vpwr vgnd scs8hd_fill_2
XFILLER_9_77 vgnd vpwr scs8hd_decap_4
XFILLER_9_99 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_242 vgnd vpwr scs8hd_decap_6
XFILLER_18_86 vgnd vpwr scs8hd_decap_6
XFILLER_18_20 vgnd vpwr scs8hd_decap_8
XFILLER_11_253 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_5.LATCH_0_.latch data_in mem_top_ipin_5.LATCH_0_.latch/Q _132_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_235 vpwr vgnd scs8hd_fill_2
X_114_ _104_/X _108_/X _114_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_297 vpwr vgnd scs8hd_fill_2
XANTENNA__121__B _122_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_353 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _186_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XFILLER_4_205 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_87 vgnd vpwr scs8hd_decap_6
XFILLER_16_389 vgnd vpwr scs8hd_decap_8
Xmem_top_ipin_7.LATCH_3_.latch data_in mem_top_ipin_7.LATCH_3_.latch/Q _145_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__132__A _104_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_67 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _179_/HI mem_bottom_ipin_0.LATCH_5_.latch/Q
+ mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_1.LATCH_4_.latch_SLEEPB _078_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_348 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_4.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_319 vpwr vgnd scs8hd_fill_2
XFILLER_0_274 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_5.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_164 vgnd vpwr scs8hd_decap_4
XFILLER_16_120 vgnd vpwr scs8hd_decap_4
XANTENNA__127__A _068_/X vgnd vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_ipin_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_370 vgnd vpwr scs8hd_decap_8
XFILLER_13_156 vpwr vgnd scs8hd_fill_2
XFILLER_9_116 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_1_.latch/Q mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.INVTX1_0_.scs8hd_inv_1 chanx_left_in[3] mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_55 vgnd vpwr scs8hd_decap_6
XFILLER_2_325 vgnd vpwr scs8hd_decap_8
XFILLER_18_215 vgnd vpwr scs8hd_decap_12
XANTENNA__124__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_5_174 vpwr vgnd scs8hd_fill_2
XANTENNA__140__A _104_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_391 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_6.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_292 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_0_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_130_ _138_/A _126_/X _130_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_402 vgnd vpwr scs8hd_decap_4
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XANTENNA__119__B _122_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_284 vgnd vpwr scs8hd_decap_4
XANTENNA__135__A _068_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_45 vpwr vgnd scs8hd_fill_2
XFILLER_9_56 vgnd vpwr scs8hd_decap_3
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
X_113_ _102_/X _108_/X _113_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_203 vpwr vgnd scs8hd_fill_2
XFILLER_11_287 vpwr vgnd scs8hd_fill_2
XFILLER_7_258 vpwr vgnd scs8hd_fill_2
XFILLER_19_365 vgnd vpwr scs8hd_fill_1
XFILLER_6_291 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_0_.latch/Q mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_16_324 vgnd vpwr scs8hd_fill_1
XANTENNA__132__B _126_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_294 vpwr vgnd scs8hd_fill_2
XFILLER_19_195 vgnd vpwr scs8hd_decap_12
XFILLER_19_184 vgnd vpwr scs8hd_decap_3
XFILLER_13_316 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_77 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_3.LATCH_3_.latch/Q mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_0_242 vgnd vpwr scs8hd_decap_4
XFILLER_0_231 vpwr vgnd scs8hd_fill_2
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_187 vpwr vgnd scs8hd_fill_2
XFILLER_16_154 vgnd vpwr scs8hd_decap_3
XFILLER_12_360 vgnd vpwr scs8hd_fill_1
XFILLER_12_382 vgnd vpwr scs8hd_decap_12
XANTENNA__127__B _126_/X vgnd vpwr scs8hd_diode_2
XANTENNA__143__A _068_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_386 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_4_.latch data_in mem_top_ipin_0.LATCH_4_.latch/Q _174_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_301 vpwr vgnd scs8hd_fill_2
XFILLER_5_367 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__138__A _138_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_190 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_6.LATCH_4_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_304 vpwr vgnd scs8hd_fill_2
XFILLER_10_149 vpwr vgnd scs8hd_fill_2
XFILLER_12_23 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_6 vpwr vgnd scs8hd_fill_2
XFILLER_18_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_7.LATCH_4_.latch/Q mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_5_142 vpwr vgnd scs8hd_fill_2
XANTENNA__140__B _140_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_271 vgnd vpwr scs8hd_decap_12
XFILLER_17_260 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_3.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_219 vgnd vpwr scs8hd_decap_12
XFILLER_2_101 vgnd vpwr scs8hd_fill_1
XFILLER_14_274 vgnd vpwr scs8hd_fill_1
XFILLER_14_241 vgnd vpwr scs8hd_decap_4
XFILLER_0_37 vpwr vgnd scs8hd_fill_2
X_189_ _189_/HI _189_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__135__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA__151__A _073_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_211 vgnd vpwr scs8hd_decap_6
Xmux_top_ipin_4.INVTX1_4_.scs8hd_inv_1 chanx_left_in[7] mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_ipin_0.LATCH_4_.latch data_in mem_bottom_ipin_0.LATCH_4_.latch/Q _158_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_112_ _138_/A _108_/X _112_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_19_377 vpwr vgnd scs8hd_fill_2
XANTENNA__146__A _138_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _187_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_56 vgnd vpwr scs8hd_decap_6
Xmux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_1_.latch/Q mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_4.LATCH_5_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_303 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_3_240 vpwr vgnd scs8hd_fill_2
XFILLER_3_262 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_1.LATCH_0_.latch data_in mem_top_ipin_1.LATCH_0_.latch/Q _091_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_391 vgnd vpwr scs8hd_decap_12
XFILLER_15_12 vpwr vgnd scs8hd_fill_2
XFILLER_13_306 vgnd vpwr scs8hd_decap_3
XFILLER_0_287 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_332 vgnd vpwr scs8hd_fill_1
XFILLER_12_394 vgnd vpwr scs8hd_decap_3
XANTENNA__143__B _142_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_398 vgnd vpwr scs8hd_decap_8
Xmem_top_ipin_3.LATCH_3_.latch data_in mem_top_ipin_3.LATCH_3_.latch/Q _111_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_90 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_103 vpwr vgnd scs8hd_fill_2
XFILLER_9_129 vpwr vgnd scs8hd_fill_2
XFILLER_5_313 vpwr vgnd scs8hd_fill_2
XFILLER_5_357 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_2_.latch/Q mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_48 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__138__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _154_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_180 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_106 vgnd vpwr scs8hd_decap_4
XANTENNA__064__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_12_79 vgnd vpwr scs8hd_decap_4
XFILLER_18_206 vgnd vpwr scs8hd_decap_8
XFILLER_18_239 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_1.LATCH_0_.latch data_in _154_/A _152_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__149__A _141_/C vgnd vpwr scs8hd_diode_2
XFILLER_20_404 vgnd vpwr scs8hd_decap_3
XFILLER_17_283 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_0_.latch/Q mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_168 vpwr vgnd scs8hd_fill_2
XFILLER_2_146 vgnd vpwr scs8hd_decap_4
XFILLER_2_135 vpwr vgnd scs8hd_fill_2
XFILLER_0_16 vgnd vpwr scs8hd_decap_4
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_14_297 vpwr vgnd scs8hd_fill_2
X_188_ _188_/HI _188_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__151__B _152_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_2.LATCH_3_.latch/Q mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
Xmux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_56 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[3] mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_111_ _111_/A _108_/X _111_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_216 vgnd vpwr scs8hd_decap_3
XFILLER_11_234 vgnd vpwr scs8hd_fill_1
XFILLER_11_245 vgnd vpwr scs8hd_fill_1
XFILLER_19_367 vgnd vpwr scs8hd_decap_6
XFILLER_19_301 vgnd vpwr scs8hd_decap_4
XANTENNA__146__B _142_/X vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _104_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__072__A enable vgnd vpwr scs8hd_diode_2
XFILLER_16_348 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.INVTX1_4_.scs8hd_inv_1 chanx_left_in[5] mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__157__A _068_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_13_329 vpwr vgnd scs8hd_fill_2
XANTENNA__067__A _066_/X vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_6.LATCH_2_.latch data_in mem_top_ipin_6.LATCH_2_.latch/Q _138_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_6.LATCH_4_.latch/Q mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_0_200 vpwr vgnd scs8hd_fill_2
XFILLER_16_145 vgnd vpwr scs8hd_decap_8
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _153_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_16 vpwr vgnd scs8hd_fill_2
XFILLER_5_336 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_130 vpwr vgnd scs8hd_fill_2
XFILLER_8_163 vpwr vgnd scs8hd_fill_2
XFILLER_4_380 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__170__A _104_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_0_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_36 vpwr vgnd scs8hd_fill_2
XANTENNA__080__A _080_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_155 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_350 vgnd vpwr scs8hd_decap_12
XFILLER_5_199 vgnd vpwr scs8hd_decap_3
XFILLER_17_240 vgnd vpwr scs8hd_decap_4
XANTENNA__149__B address[6] vgnd vpwr scs8hd_diode_2
XANTENNA__165__A _068_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_1_.latch/Q mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__075__A _068_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_114 vpwr vgnd scs8hd_fill_2
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
XFILLER_14_265 vgnd vpwr scs8hd_fill_1
XFILLER_9_26 vpwr vgnd scs8hd_fill_2
X_187_ _187_/HI _187_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__151__C _163_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_110_ _096_/X _108_/X _110_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_213 vpwr vgnd scs8hd_fill_2
XFILLER_7_239 vgnd vpwr scs8hd_decap_3
XFILLER_11_268 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_6.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__162__B _156_/X vgnd vpwr scs8hd_diode_2
XFILLER_10_290 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _179_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _188_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__072__B _124_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_209 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_2_.latch/Q mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_404 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_231 vpwr vgnd scs8hd_fill_2
XFILLER_6_27 vpwr vgnd scs8hd_fill_2
XFILLER_19_121 vgnd vpwr scs8hd_fill_1
XFILLER_13_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__157__B _156_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _068_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__083__A _080_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_278 vgnd vpwr scs8hd_fill_1
XFILLER_16_179 vgnd vpwr scs8hd_fill_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_0_.latch/Q mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_356 vpwr vgnd scs8hd_fill_2
XANTENNA__168__A _168_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[7] mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_138 vgnd vpwr scs8hd_decap_4
XANTENNA__078__A _082_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_1.LATCH_3_.latch/Q mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__170__B _166_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_186 vgnd vpwr scs8hd_decap_3
XFILLER_4_392 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_6.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_119 vgnd vpwr scs8hd_decap_4
XFILLER_2_318 vgnd vpwr scs8hd_decap_4
XANTENNA__080__B address[2] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XFILLER_5_123 vpwr vgnd scs8hd_fill_2
XFILLER_5_178 vgnd vpwr scs8hd_decap_3
XFILLER_1_362 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__149__C address[5] vgnd vpwr scs8hd_diode_2
XANTENNA__165__B _166_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_60 vpwr vgnd scs8hd_fill_2
XFILLER_4_93 vpwr vgnd scs8hd_fill_2
XANTENNA__075__B _082_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_7.INVTX1_5_.scs8hd_inv_1 chanx_right_in[5] mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_406 vgnd vpwr scs8hd_fill_1
XFILLER_2_104 vgnd vpwr scs8hd_fill_1
XANTENNA__091__A _082_/A vgnd vpwr scs8hd_diode_2
XANTENNA__151__D _151_/D vgnd vpwr scs8hd_diode_2
X_186_ _186_/HI _186_/LO vgnd vpwr scs8hd_conb_1
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__176__A _168_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_5.LATCH_4_.latch/Q mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA__086__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_4
X_169_ _102_/A _166_/B _169_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_72 vgnd vpwr scs8hd_decap_3
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__072__C address[5] vgnd vpwr scs8hd_diode_2
XFILLER_16_328 vgnd vpwr scs8hd_decap_8
XFILLER_3_254 vpwr vgnd scs8hd_fill_2
XFILLER_3_298 vgnd vpwr scs8hd_decap_4
XFILLER_10_70 vgnd vpwr scs8hd_decap_4
XANTENNA__173__B _178_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_15_37 vgnd vpwr scs8hd_fill_1
XANTENNA__083__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_213 vpwr vgnd scs8hd_fill_2
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_1_.latch/Q mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_335 vgnd vpwr scs8hd_fill_1
XANTENNA__168__B _166_/B vgnd vpwr scs8hd_diode_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_7_82 vpwr vgnd scs8hd_fill_2
XANTENNA__078__B _166_/A vgnd vpwr scs8hd_diode_2
XANTENNA__094__A _094_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_349 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_6.LATCH_1_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_29 vgnd vpwr scs8hd_decap_3
Xmem_top_ipin_2.LATCH_2_.latch data_in mem_top_ipin_2.LATCH_2_.latch/Q _101_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_198 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_27 vpwr vgnd scs8hd_fill_2
XFILLER_2_308 vgnd vpwr scs8hd_fill_1
XANTENNA__080__C _151_/D vgnd vpwr scs8hd_diode_2
XANTENNA__089__A address[1] vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_4.LATCH_5_.latch data_in mem_top_ipin_4.LATCH_5_.latch/Q _117_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_341 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_2_.latch/Q mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_72 vgnd vpwr scs8hd_fill_1
XFILLER_4_190 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__091__B _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_245 vgnd vpwr scs8hd_fill_1
XFILLER_14_201 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_4.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_185_ _185_/HI _185_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_92 vpwr vgnd scs8hd_fill_2
XFILLER_1_182 vgnd vpwr scs8hd_fill_1
XANTENNA__176__B _178_/B vgnd vpwr scs8hd_diode_2
XANTENNA__192__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_9_271 vgnd vpwr scs8hd_decap_4
XFILLER_9_282 vgnd vpwr scs8hd_decap_4
XFILLER_18_15 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_0_.latch/Q mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__086__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_226 vpwr vgnd scs8hd_fill_2
XFILLER_11_237 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_2.LATCH_2_.latch data_in mem_bottom_ipin_2.LATCH_2_.latch/Q _168_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_337 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_4.LATCH_2_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
X_168_ _168_/A _166_/B _168_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_6_274 vgnd vpwr scs8hd_fill_1
X_099_ _111_/A _103_/B _099_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_40 vpwr vgnd scs8hd_fill_2
XFILLER_1_62 vgnd vpwr scs8hd_fill_1
XFILLER_1_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _189_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__097__A _096_/X vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_0.LATCH_3_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_3_277 vpwr vgnd scs8hd_fill_2
XFILLER_19_123 vgnd vpwr scs8hd_decap_12
XFILLER_15_351 vpwr vgnd scs8hd_fill_2
XFILLER_15_340 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_16 vpwr vgnd scs8hd_fill_2
XANTENNA__083__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_258 vpwr vgnd scs8hd_fill_2
XFILLER_16_126 vpwr vgnd scs8hd_fill_2
XFILLER_16_115 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_1_.latch/Q mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_369 vpwr vgnd scs8hd_fill_2
XFILLER_12_398 vgnd vpwr scs8hd_decap_8
XPHY_1 vgnd vpwr scs8hd_decap_3
Xmem_top_ipin_5.LATCH_1_.latch data_in mem_top_ipin_5.LATCH_1_.latch/Q _131_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_380 vpwr vgnd scs8hd_fill_2
XFILLER_7_391 vgnd vpwr scs8hd_decap_12
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_107 vpwr vgnd scs8hd_fill_2
XFILLER_5_317 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_4.LATCH_4_.latch/Q mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA_mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_350 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_7.LATCH_4_.latch data_in mem_top_ipin_7.LATCH_4_.latch/Q _144_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__195__A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_3_.latch_SLEEPB _099_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__089__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_5_114 vpwr vgnd scs8hd_fill_2
XFILLER_4_84 vpwr vgnd scs8hd_fill_2
XFILLER_14_268 vgnd vpwr scs8hd_decap_6
XFILLER_14_224 vgnd vpwr scs8hd_decap_8
XFILLER_14_213 vgnd vpwr scs8hd_fill_1
X_184_ _184_/HI _184_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_161 vgnd vpwr scs8hd_decap_3
XFILLER_20_249 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__086__C _151_/D vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_249 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
X_167_ _167_/A _166_/B _167_/Y vgnd vpwr scs8hd_nor2_4
X_098_ _167_/A _111_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_253 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_30 vgnd vpwr scs8hd_fill_1
XFILLER_16_308 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB _174_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XANTENNA__097__B _103_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_201 vpwr vgnd scs8hd_fill_2
XFILLER_19_135 vgnd vpwr scs8hd_decap_12
XFILLER_19_81 vpwr vgnd scs8hd_fill_2
XFILLER_19_70 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_3.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__198__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_ipin_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_348 vgnd vpwr scs8hd_decap_8
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_2_.latch/Q mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_311 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_182 vgnd vpwr scs8hd_fill_1
XFILLER_15_171 vpwr vgnd scs8hd_fill_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_7_62 vgnd vpwr scs8hd_decap_3
XFILLER_16_82 vpwr vgnd scs8hd_fill_2
XFILLER_8_145 vgnd vpwr scs8hd_decap_6
XFILLER_8_167 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_130 vgnd vpwr scs8hd_decap_4
XFILLER_12_163 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_0_.latch/Q mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__089__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_14_406 vgnd vpwr scs8hd_fill_1
XFILLER_5_159 vpwr vgnd scs8hd_fill_2
XFILLER_17_288 vpwr vgnd scs8hd_fill_2
XFILLER_4_41 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_118 vpwr vgnd scs8hd_fill_2
X_183_ _183_/HI _183_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_184 vpwr vgnd scs8hd_fill_2
XFILLER_1_140 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_0.LATCH_5_.latch data_in mem_top_ipin_0.LATCH_5_.latch/Q _173_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_28 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_7.LATCH_3_.latch_SLEEPB _145_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_1_.latch/Q mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_306 vgnd vpwr scs8hd_decap_12
XFILLER_10_250 vpwr vgnd scs8hd_fill_2
X_166_ _166_/A _166_/B _166_/Y vgnd vpwr scs8hd_nor2_4
X_097_ _096_/X _103_/B _097_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_232 vpwr vgnd scs8hd_fill_2
XFILLER_6_276 vgnd vpwr scs8hd_decap_6
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XFILLER_18_361 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _181_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB _160_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_3.LATCH_4_.latch/Q mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_3_213 vgnd vpwr scs8hd_fill_1
XFILLER_3_235 vgnd vpwr scs8hd_decap_3
XFILLER_10_40 vgnd vpwr scs8hd_decap_4
XFILLER_19_147 vgnd vpwr scs8hd_decap_12
XFILLER_10_84 vgnd vpwr scs8hd_decap_8
X_149_ _141_/C address[6] address[5] _149_/X vgnd vpwr scs8hd_or3_4
Xmux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_29 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_238 vpwr vgnd scs8hd_fill_2
XFILLER_0_227 vpwr vgnd scs8hd_fill_2
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_ipin_0.LATCH_5_.latch data_in mem_bottom_ipin_0.LATCH_5_.latch/Q _157_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_8 vpwr vgnd scs8hd_fill_2
XFILLER_15_150 vpwr vgnd scs8hd_fill_2
XPHY_3 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_1.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_5.LATCH_4_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_72 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _189_/HI mem_top_ipin_7.LATCH_5_.latch/Q
+ mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_186 vpwr vgnd scs8hd_fill_2
XFILLER_4_396 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_12_ vgnd vpwr scs8hd_inv_1
Xmem_top_ipin_1.LATCH_1_.latch data_in mem_top_ipin_1.LATCH_1_.latch/Q _088_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_138 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.INVTX1_2_.scs8hd_inv_1 chanx_left_in[1] mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_267 vpwr vgnd scs8hd_fill_2
XFILLER_17_256 vpwr vgnd scs8hd_fill_2
XFILLER_17_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_182 vpwr vgnd scs8hd_fill_2
XFILLER_4_64 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_3.LATCH_4_.latch data_in mem_top_ipin_3.LATCH_4_.latch/Q _110_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_248 vpwr vgnd scs8hd_fill_2
XFILLER_13_51 vpwr vgnd scs8hd_fill_2
X_182_ _182_/HI _182_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_62 vpwr vgnd scs8hd_fill_2
XANTENNA__100__A _168_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_218 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_2_.latch/Q mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_318 vgnd vpwr scs8hd_decap_12
XFILLER_1_7 vgnd vpwr scs8hd_fill_1
X_165_ _068_/A _166_/B _165_/Y vgnd vpwr scs8hd_nor2_4
X_096_ _166_/A _096_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mem_top_ipin_3.LATCH_5_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_266 vgnd vpwr scs8hd_decap_8
XFILLER_6_299 vgnd vpwr scs8hd_fill_1
XFILLER_18_373 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_1.LATCH_1_.latch data_in _153_/A _151_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_258 vpwr vgnd scs8hd_fill_2
XFILLER_10_74 vgnd vpwr scs8hd_fill_1
XFILLER_19_159 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_0_.latch/Q mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_365 vgnd vpwr scs8hd_fill_1
X_148_ _104_/X _142_/X _148_/Y vgnd vpwr scs8hd_nor2_4
X_079_ address[1] _080_/A vgnd vpwr scs8hd_inv_8
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_107 vgnd vpwr scs8hd_decap_8
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_328 vgnd vpwr scs8hd_decap_4
XFILLER_15_184 vgnd vpwr scs8hd_decap_3
XPHY_4 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_42 vpwr vgnd scs8hd_fill_2
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_7_86 vpwr vgnd scs8hd_fill_2
XFILLER_5_309 vpwr vgnd scs8hd_fill_2
XFILLER_17_405 vpwr vgnd scs8hd_fill_2
XFILLER_4_320 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_4.LATCH_0_.latch data_in mem_top_ipin_4.LATCH_0_.latch/Q _122_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__103__A _102_/X vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_1_.latch/Q mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_301 vpwr vgnd scs8hd_fill_2
XFILLER_1_367 vgnd vpwr scs8hd_decap_12
XFILLER_1_345 vgnd vpwr scs8hd_decap_3
XFILLER_17_213 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_6.LATCH_3_.latch data_in mem_top_ipin_6.LATCH_3_.latch/Q _137_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_161 vgnd vpwr scs8hd_decap_4
XFILLER_16_290 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_2.LATCH_4_.latch/Q mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_14_205 vpwr vgnd scs8hd_fill_2
X_181_ _181_/HI _181_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_96 vpwr vgnd scs8hd_fill_2
XFILLER_1_175 vgnd vpwr scs8hd_decap_4
XFILLER_1_153 vpwr vgnd scs8hd_fill_2
XFILLER_13_293 vpwr vgnd scs8hd_fill_2
XFILLER_13_271 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_5.INVTX1_2_.scs8hd_inv_1 chanx_left_in[7] mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_242 vpwr vgnd scs8hd_fill_2
XFILLER_9_275 vgnd vpwr scs8hd_fill_1
XFILLER_9_297 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__201__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_095_ _068_/X _103_/B _095_/Y vgnd vpwr scs8hd_nor2_4
X_164_ _163_/X _166_/B vgnd vpwr scs8hd_buf_1
XFILLER_10_263 vpwr vgnd scs8hd_fill_2
XFILLER_10_285 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_18_385 vgnd vpwr scs8hd_decap_12
XANTENNA__111__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_77 vpwr vgnd scs8hd_fill_2
XFILLER_1_88 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _188_/HI mem_top_ipin_6.LATCH_5_.latch/Q
+ mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_19_62 vgnd vpwr scs8hd_decap_4
XFILLER_15_355 vpwr vgnd scs8hd_fill_2
XFILLER_15_344 vgnd vpwr scs8hd_decap_4
XANTENNA__106__A address[4] vgnd vpwr scs8hd_diode_2
X_078_ _082_/A _166_/A _078_/Y vgnd vpwr scs8hd_nor2_4
X_147_ _102_/X _142_/X _147_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_292 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_207 vgnd vpwr scs8hd_decap_4
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_7_10 vpwr vgnd scs8hd_fill_2
XFILLER_11_380 vgnd vpwr scs8hd_decap_4
XFILLER_11_391 vgnd vpwr scs8hd_decap_4
XFILLER_7_362 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_41 vgnd vpwr scs8hd_decap_8
XFILLER_16_30 vgnd vpwr scs8hd_fill_1
XFILLER_16_96 vgnd vpwr scs8hd_decap_8
XFILLER_8_126 vpwr vgnd scs8hd_fill_2
XANTENNA__103__B _103_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_398 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_2_.latch/Q mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__204__A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_5_118 vpwr vgnd scs8hd_fill_2
XFILLER_1_379 vgnd vpwr scs8hd_decap_12
XFILLER_17_236 vpwr vgnd scs8hd_fill_2
XFILLER_17_225 vgnd vpwr scs8hd_decap_8
XFILLER_4_88 vgnd vpwr scs8hd_decap_4
XFILLER_4_140 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__114__A _104_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_75 vpwr vgnd scs8hd_fill_2
XFILLER_13_31 vpwr vgnd scs8hd_fill_2
X_180_ _180_/HI _180_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_1_132 vpwr vgnd scs8hd_fill_2
XANTENNA__109__A _068_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_254 vpwr vgnd scs8hd_fill_2
XFILLER_11_209 vpwr vgnd scs8hd_fill_2
X_163_ _163_/A _073_/B _163_/C _163_/X vgnd vpwr scs8hd_or3_4
X_094_ _094_/A _103_/B vgnd vpwr scs8hd_buf_1
XANTENNA__111__B _108_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB _177_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.INVTX1_2_.scs8hd_inv_1 chanx_left_in[5] mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_205 vpwr vgnd scs8hd_fill_2
XFILLER_3_227 vpwr vgnd scs8hd_fill_2
XFILLER_10_21 vgnd vpwr scs8hd_decap_8
XFILLER_19_85 vgnd vpwr scs8hd_decap_12
XFILLER_19_74 vgnd vpwr scs8hd_decap_4
XFILLER_15_323 vpwr vgnd scs8hd_fill_2
XFILLER_15_301 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_1_.latch/Q mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_367 vgnd vpwr scs8hd_decap_12
XANTENNA__122__A _104_/X vgnd vpwr scs8hd_diode_2
X_077_ _076_/X _166_/A vgnd vpwr scs8hd_buf_1
X_146_ _138_/A _142_/X _146_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_271 vpwr vgnd scs8hd_fill_2
XANTENNA__207__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_304 vgnd vpwr scs8hd_decap_4
XFILLER_12_348 vgnd vpwr scs8hd_decap_12
XFILLER_15_175 vgnd vpwr scs8hd_decap_4
XPHY_6 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_ipin_1.LATCH_4_.latch/Q mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_7_352 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__117__A _068_/X vgnd vpwr scs8hd_diode_2
X_129_ _111_/A _126_/X _129_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_86 vgnd vpwr scs8hd_decap_6
XFILLER_16_64 vpwr vgnd scs8hd_fill_2
XFILLER_16_20 vpwr vgnd scs8hd_fill_2
XFILLER_12_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_160 vpwr vgnd scs8hd_fill_2
XFILLER_7_193 vpwr vgnd scs8hd_fill_2
XFILLER_9_403 vgnd vpwr scs8hd_decap_4
XANTENNA__114__B _108_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_23 vgnd vpwr scs8hd_decap_6
XANTENNA__130__A _138_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _187_/HI mem_top_ipin_5.LATCH_5_.latch/Q
+ mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmem_top_ipin_0.LATCH_0_.latch data_in mem_top_ipin_0.LATCH_0_.latch/Q _178_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_0_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_406 vgnd vpwr scs8hd_fill_1
XFILLER_1_188 vpwr vgnd scs8hd_fill_2
XANTENNA__109__B _108_/X vgnd vpwr scs8hd_diode_2
XANTENNA__125__A _073_/A vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_2.LATCH_3_.latch data_in mem_top_ipin_2.LATCH_3_.latch/Q _099_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_162_ _104_/A _156_/X _162_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_232 vgnd vpwr scs8hd_fill_1
X_093_ _073_/A _152_/B _073_/C _094_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_236 vpwr vgnd scs8hd_fill_2
XFILLER_1_13 vpwr vgnd scs8hd_fill_2
XFILLER_1_24 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_398 vgnd vpwr scs8hd_decap_8
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_97 vgnd vpwr scs8hd_decap_12
XFILLER_15_379 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_145_ _111_/A _142_/X _145_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_2_.latch/Q mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__122__B _122_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_261 vgnd vpwr scs8hd_decap_3
X_076_ address[1] _076_/B address[0] _076_/X vgnd vpwr scs8hd_or3_4
XFILLER_18_151 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_0.LATCH_0_.latch data_in mem_bottom_ipin_0.LATCH_0_.latch/Q _162_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_195 vgnd vpwr scs8hd_decap_8
XFILLER_18_184 vgnd vpwr scs8hd_decap_8
XFILLER_18_173 vgnd vpwr scs8hd_decap_8
XFILLER_18_162 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_309 vgnd vpwr scs8hd_decap_6
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_ipin_1.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_198 vpwr vgnd scs8hd_fill_2
XFILLER_15_154 vpwr vgnd scs8hd_fill_2
XPHY_7 vgnd vpwr scs8hd_decap_3
X_128_ _096_/X _126_/X _128_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__133__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_7_23 vpwr vgnd scs8hd_fill_2
XFILLER_7_78 vpwr vgnd scs8hd_fill_2
XANTENNA__117__B _122_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_1_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_3_.latch data_in mem_bottom_ipin_2.LATCH_3_.latch/Q _167_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_6
XFILLER_12_102 vgnd vpwr scs8hd_decap_12
XFILLER_4_301 vgnd vpwr scs8hd_decap_4
XFILLER_12_168 vgnd vpwr scs8hd_decap_3
XANTENNA__128__A _096_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_190 vpwr vgnd scs8hd_fill_2
XFILLER_1_337 vpwr vgnd scs8hd_fill_2
XFILLER_1_326 vgnd vpwr scs8hd_decap_8
XFILLER_1_315 vpwr vgnd scs8hd_fill_2
XFILLER_17_249 vgnd vpwr scs8hd_decap_4
XFILLER_17_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_46 vgnd vpwr scs8hd_decap_3
XFILLER_4_68 vgnd vpwr scs8hd_decap_4
XFILLER_4_186 vpwr vgnd scs8hd_fill_2
XANTENNA__130__B _126_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_271 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_1_.latch/Q mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_11 vgnd vpwr scs8hd_decap_3
XFILLER_13_55 vgnd vpwr scs8hd_decap_4
XFILLER_13_44 vgnd vpwr scs8hd_decap_4
Xmem_top_ipin_5.LATCH_2_.latch data_in mem_top_ipin_5.LATCH_2_.latch/Q _130_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_101 vgnd vpwr scs8hd_decap_4
XFILLER_1_112 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__125__B _073_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_201 vgnd vpwr scs8hd_decap_3
XFILLER_9_234 vpwr vgnd scs8hd_fill_2
XFILLER_9_278 vpwr vgnd scs8hd_fill_2
XANTENNA__141__A _163_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_2_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_0.LATCH_4_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
Xmem_top_ipin_7.LATCH_5_.latch data_in mem_top_ipin_7.LATCH_5_.latch/Q _143_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_215 vgnd vpwr scs8hd_decap_4
X_161_ _102_/A _156_/X _161_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_211 vgnd vpwr scs8hd_fill_1
X_092_ address[3] _152_/B vgnd vpwr scs8hd_inv_8
XFILLER_18_300 vgnd vpwr scs8hd_decap_12
XFILLER_1_36 vpwr vgnd scs8hd_fill_2
XANTENNA__136__A _096_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_2_.latch/Q mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_075_ _068_/X _082_/A _075_/Y vgnd vpwr scs8hd_nor2_4
X_144_ _096_/X _142_/X _144_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_240 vpwr vgnd scs8hd_fill_2
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_328 vgnd vpwr scs8hd_decap_6
XFILLER_15_133 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _186_/HI mem_top_ipin_4.LATCH_5_.latch/Q
+ mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_127_ _068_/X _126_/X _127_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__133__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_46 vpwr vgnd scs8hd_fill_2
XFILLER_7_57 vgnd vpwr scs8hd_decap_4
XFILLER_7_376 vpwr vgnd scs8hd_fill_2
XFILLER_7_387 vpwr vgnd scs8hd_fill_2
XFILLER_16_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_1.LATCH_3_.latch_SLEEPB _082_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_114 vgnd vpwr scs8hd_decap_3
XFILLER_20_180 vgnd vpwr scs8hd_decap_6
XFILLER_4_324 vgnd vpwr scs8hd_decap_12
XFILLER_4_346 vpwr vgnd scs8hd_fill_2
XFILLER_4_357 vgnd vpwr scs8hd_decap_8
XFILLER_4_368 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__128__B _126_/X vgnd vpwr scs8hd_diode_2
XANTENNA__144__A _096_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_140 vgnd vpwr scs8hd_decap_3
XFILLER_4_121 vpwr vgnd scs8hd_fill_2
XFILLER_4_165 vgnd vpwr scs8hd_fill_1
XANTENNA__139__A _102_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_14_209 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_1_179 vgnd vpwr scs8hd_fill_1
XFILLER_1_157 vpwr vgnd scs8hd_fill_2
XFILLER_13_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_13_297 vpwr vgnd scs8hd_fill_2
XFILLER_13_275 vpwr vgnd scs8hd_fill_2
XANTENNA__125__C _141_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__141__B _073_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_091_ _082_/A _104_/A _091_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_249 vpwr vgnd scs8hd_fill_2
X_160_ _168_/A _156_/X _160_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_267 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_312 vgnd vpwr scs8hd_decap_12
XANTENNA__136__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _073_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_46 vgnd vpwr scs8hd_fill_1
XFILLER_19_109 vgnd vpwr scs8hd_decap_12
XFILLER_19_66 vgnd vpwr scs8hd_fill_1
XFILLER_19_11 vgnd vpwr scs8hd_decap_12
XFILLER_15_359 vgnd vpwr scs8hd_decap_6
XFILLER_15_315 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_074_ _073_/X _082_/A vgnd vpwr scs8hd_buf_1
X_143_ _068_/A _142_/X _143_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_296 vgnd vpwr scs8hd_decap_8
XFILLER_2_285 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_131 vgnd vpwr scs8hd_decap_12
XFILLER_18_7 vgnd vpwr scs8hd_decap_8
XANTENNA__147__A _102_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_373 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_123 vgnd vpwr scs8hd_fill_1
XFILLER_15_112 vgnd vpwr scs8hd_decap_4
XFILLER_15_101 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_167 vpwr vgnd scs8hd_fill_2
XFILLER_7_333 vpwr vgnd scs8hd_fill_2
XFILLER_11_351 vpwr vgnd scs8hd_fill_2
XFILLER_11_362 vpwr vgnd scs8hd_fill_2
X_126_ _125_/X _126_/X vgnd vpwr scs8hd_buf_1
XANTENNA__133__C _141_/C vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_1_.latch/Q mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_126 vpwr vgnd scs8hd_fill_2
XANTENNA__144__B _142_/X vgnd vpwr scs8hd_diode_2
X_109_ _068_/X _108_/X _109_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__160__A _168_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_281 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__070__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_4_100 vpwr vgnd scs8hd_fill_2
XANTENNA__155__A _073_/A vgnd vpwr scs8hd_diode_2
XANTENNA__139__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_2_.latch/Q mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_6.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_79 vpwr vgnd scs8hd_fill_2
XANTENNA__065__A address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_136 vpwr vgnd scs8hd_fill_2
XFILLER_8_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_6.LATCH_3_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_254 vpwr vgnd scs8hd_fill_2
XANTENNA__125__D _124_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_258 vpwr vgnd scs8hd_fill_2
XANTENNA__141__C _141_/C vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _185_/HI mem_top_ipin_3.LATCH_5_.latch/Q
+ mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_090_ _090_/A _104_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_206 vgnd vpwr scs8hd_decap_8
XFILLER_10_224 vpwr vgnd scs8hd_fill_2
XFILLER_10_246 vpwr vgnd scs8hd_fill_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_3
XFILLER_18_324 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_1.LATCH_2_.latch data_in mem_top_ipin_1.LATCH_2_.latch/Q _085_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__152__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_209 vgnd vpwr scs8hd_decap_4
XFILLER_10_36 vpwr vgnd scs8hd_fill_2
XFILLER_10_58 vgnd vpwr scs8hd_decap_12
XFILLER_19_23 vgnd vpwr scs8hd_decap_12
XFILLER_15_327 vpwr vgnd scs8hd_fill_2
X_142_ _142_/A _142_/X vgnd vpwr scs8hd_buf_1
X_073_ _073_/A _073_/B _073_/C _073_/X vgnd vpwr scs8hd_or3_4
Xmem_top_ipin_3.LATCH_5_.latch data_in mem_top_ipin_3.LATCH_5_.latch/Q _109_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.INVTX1_3_.scs8hd_inv_1 chanx_right_in[6] mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_154 vgnd vpwr scs8hd_decap_4
XFILLER_18_143 vgnd vpwr scs8hd_decap_8
XANTENNA__147__B _142_/X vgnd vpwr scs8hd_diode_2
XANTENNA__163__A _163_/A vgnd vpwr scs8hd_diode_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_308 vgnd vpwr scs8hd_fill_1
XFILLER_20_385 vgnd vpwr scs8hd_decap_12
XANTENNA__073__A _073_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_4_ vgnd vpwr scs8hd_inv_1
XFILLER_15_179 vgnd vpwr scs8hd_fill_1
X_125_ _073_/A _073_/B _141_/C _124_/X _125_/X vgnd vpwr scs8hd_or4_4
XFILLER_7_356 vgnd vpwr scs8hd_decap_4
XANTENNA__133__D _124_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_4_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__158__A _166_/A vgnd vpwr scs8hd_diode_2
XANTENNA__068__A _068_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_68 vgnd vpwr scs8hd_decap_4
XFILLER_16_24 vgnd vpwr scs8hd_decap_6
XFILLER_8_109 vgnd vpwr scs8hd_decap_8
XFILLER_12_149 vpwr vgnd scs8hd_fill_2
X_108_ _108_/A _108_/X vgnd vpwr scs8hd_buf_1
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
XFILLER_7_197 vgnd vpwr scs8hd_decap_4
XANTENNA__160__B _156_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_373 vgnd vpwr scs8hd_decap_12
XFILLER_4_178 vpwr vgnd scs8hd_fill_2
XANTENNA__155__B _073_/B vgnd vpwr scs8hd_diode_2
XANTENNA__171__A _163_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_406 vgnd vpwr scs8hd_fill_1
XANTENNA__081__A _080_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_215 vpwr vgnd scs8hd_fill_2
XANTENNA__141__D _124_/X vgnd vpwr scs8hd_diode_2
XANTENNA__166__A _166_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_2.LATCH_5_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_4.LATCH_1_.latch data_in mem_top_ipin_4.LATCH_1_.latch/Q _121_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__076__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_10_203 vpwr vgnd scs8hd_fill_2
XFILLER_1_17 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_1_.latch/Q mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__152__C _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_5_240 vpwr vgnd scs8hd_fill_2
XFILLER_5_284 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_6.LATCH_4_.latch data_in mem_top_ipin_6.LATCH_4_.latch/Q _136_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_35 vgnd vpwr scs8hd_decap_12
X_141_ _163_/A _073_/B _141_/C _124_/X _142_/A vgnd vpwr scs8hd_or4_4
X_072_ enable _124_/A address[5] _073_/C vgnd vpwr scs8hd_nand3_4
XFILLER_14_350 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_394 vgnd vpwr scs8hd_decap_3
XANTENNA__163__B _073_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_fill_1
XFILLER_20_342 vgnd vpwr scs8hd_decap_12
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_397 vgnd vpwr scs8hd_decap_6
XANTENNA__073__B _073_/B vgnd vpwr scs8hd_diode_2
X_124_ _124_/A address[5] _124_/X vgnd vpwr scs8hd_or2_4
XFILLER_7_27 vpwr vgnd scs8hd_fill_2
XFILLER_7_302 vgnd vpwr scs8hd_decap_3
XFILLER_7_313 vgnd vpwr scs8hd_decap_4
XFILLER_11_320 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_2_.latch/Q mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__158__B _156_/X vgnd vpwr scs8hd_diode_2
XANTENNA__174__A _166_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_58 vgnd vpwr scs8hd_decap_4
XANTENNA__084__A _083_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_305 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_107_ _163_/A _073_/B _073_/C _108_/A vgnd vpwr scs8hd_or3_4
XFILLER_7_132 vpwr vgnd scs8hd_fill_2
XFILLER_11_194 vpwr vgnd scs8hd_fill_2
XFILLER_3_371 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_3 vpwr vgnd scs8hd_fill_2
XANTENNA__169__A _102_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _184_/HI mem_top_ipin_2.LATCH_5_.latch/Q
+ mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_1_319 vgnd vpwr scs8hd_decap_4
XFILLER_17_209 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_0_385 vgnd vpwr scs8hd_decap_12
XFILLER_4_168 vgnd vpwr scs8hd_fill_1
XFILLER_16_231 vgnd vpwr scs8hd_decap_8
XANTENNA__155__C _163_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__171__B _152_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_13_48 vgnd vpwr scs8hd_fill_1
XFILLER_13_289 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_7.LATCH_0_.latch data_in mem_top_ipin_7.LATCH_0_.latch/Q _148_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_238 vpwr vgnd scs8hd_fill_2
XFILLER_0_182 vpwr vgnd scs8hd_fill_2
XFILLER_0_160 vgnd vpwr scs8hd_fill_1
XANTENNA__166__B _166_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB _167_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_60 vgnd vpwr scs8hd_fill_1
XANTENNA__076__B _076_/B vgnd vpwr scs8hd_diode_2
XANTENNA__092__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_18_337 vgnd vpwr scs8hd_decap_12
XFILLER_14_80 vpwr vgnd scs8hd_fill_2
XFILLER_5_230 vpwr vgnd scs8hd_fill_2
XANTENNA__152__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_5_263 vpwr vgnd scs8hd_fill_2
XANTENNA__177__A _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_381 vgnd vpwr scs8hd_decap_12
XFILLER_19_47 vgnd vpwr scs8hd_decap_12
XANTENNA__087__A _087_/A vgnd vpwr scs8hd_diode_2
X_140_ _104_/X _140_/B _140_/Y vgnd vpwr scs8hd_nor2_4
X_071_ address[6] _124_/A vgnd vpwr scs8hd_inv_8
XFILLER_2_244 vgnd vpwr scs8hd_decap_3
XFILLER_2_211 vgnd vpwr scs8hd_decap_3
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__163__C _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_2_83 vgnd vpwr scs8hd_decap_6
XFILLER_2_72 vgnd vpwr scs8hd_decap_8
XFILLER_20_354 vgnd vpwr scs8hd_decap_12
XANTENNA__073__C _073_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_5_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_137 vpwr vgnd scs8hd_fill_2
X_123_ enable _141_/C vgnd vpwr scs8hd_inv_8
XFILLER_11_343 vpwr vgnd scs8hd_fill_2
XFILLER_11_376 vpwr vgnd scs8hd_fill_2
XFILLER_11_387 vpwr vgnd scs8hd_fill_2
XFILLER_11_398 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB _091_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_92 vpwr vgnd scs8hd_fill_2
XFILLER_16_7 vgnd vpwr scs8hd_decap_4
XFILLER_14_181 vgnd vpwr scs8hd_fill_1
XANTENNA__174__B _178_/B vgnd vpwr scs8hd_diode_2
XANTENNA__190__A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
X_106_ address[4] _163_/A vgnd vpwr scs8hd_inv_8
XFILLER_11_184 vgnd vpwr scs8hd_decap_3
XFILLER_3_383 vgnd vpwr scs8hd_decap_12
XANTENNA__169__B _166_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_8_93 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_405 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__095__A _068_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_4_125 vpwr vgnd scs8hd_fill_2
XFILLER_4_136 vpwr vgnd scs8hd_fill_2
XFILLER_0_397 vgnd vpwr scs8hd_decap_6
XFILLER_0_342 vgnd vpwr scs8hd_decap_12
XFILLER_16_287 vgnd vpwr scs8hd_fill_1
XANTENNA__171__C _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_13_27 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_2_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_279 vgnd vpwr scs8hd_fill_1
XFILLER_13_235 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_6.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_94 vgnd vpwr scs8hd_decap_3
XANTENNA__076__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_18_349 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_2_.latch/Q mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_14_70 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_7.INVTX1_4_.scs8hd_inv_1 chanx_left_in[5] mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_297 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__177__B _178_/B vgnd vpwr scs8hd_diode_2
XANTENNA__193__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_17_393 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_ipin_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_0.LATCH_1_.latch data_in mem_top_ipin_0.LATCH_1_.latch/Q _177_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_070_ address[3] _073_/B vgnd vpwr scs8hd_buf_1
XFILLER_2_289 vgnd vpwr scs8hd_fill_1
XFILLER_2_267 vpwr vgnd scs8hd_fill_2
XFILLER_2_256 vgnd vpwr scs8hd_decap_3
XFILLER_2_201 vpwr vgnd scs8hd_fill_2
XFILLER_4_3 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _183_/HI mem_top_ipin_1.LATCH_5_.latch/Q
+ mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_14_374 vgnd vpwr scs8hd_decap_12
XFILLER_14_363 vgnd vpwr scs8hd_decap_8
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_199_ chanx_left_in[8] chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_366 vgnd vpwr scs8hd_decap_6
XFILLER_20_311 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_2.LATCH_4_.latch data_in mem_top_ipin_2.LATCH_4_.latch/Q _097_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_116 vgnd vpwr scs8hd_fill_1
XFILLER_15_105 vpwr vgnd scs8hd_fill_2
XANTENNA__098__A _167_/A vgnd vpwr scs8hd_diode_2
X_122_ _104_/X _122_/B _122_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_348 vpwr vgnd scs8hd_fill_2
XFILLER_14_193 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
X_105_ _104_/X _103_/B _105_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_156 vpwr vgnd scs8hd_fill_2
XFILLER_11_163 vgnd vpwr scs8hd_fill_1
XFILLER_3_362 vgnd vpwr scs8hd_decap_4
XFILLER_3_395 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_1_.latch data_in mem_bottom_ipin_0.LATCH_1_.latch/Q _161_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__095__B _103_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_104 vpwr vgnd scs8hd_fill_2
XFILLER_4_148 vgnd vpwr scs8hd_decap_3
XFILLER_0_354 vgnd vpwr scs8hd_decap_12
XFILLER_16_244 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_6.LATCH_0_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__196__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_4_.latch data_in mem_bottom_ipin_2.LATCH_4_.latch/Q _166_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_107 vpwr vgnd scs8hd_fill_2
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_258 vpwr vgnd scs8hd_fill_2
XFILLER_13_214 vpwr vgnd scs8hd_fill_2
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_40 vpwr vgnd scs8hd_fill_2
XFILLER_5_62 vpwr vgnd scs8hd_fill_2
XFILLER_8_295 vgnd vpwr scs8hd_fill_1
XFILLER_10_228 vgnd vpwr scs8hd_decap_4
XFILLER_5_254 vgnd vpwr scs8hd_decap_3
Xmem_top_ipin_3.LATCH_0_.latch data_in mem_top_ipin_3.LATCH_0_.latch/Q _114_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_158 vgnd vpwr scs8hd_fill_1
XFILLER_14_386 vgnd vpwr scs8hd_decap_8
XPHY_70 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_top_ipin_5.LATCH_3_.latch data_in mem_top_ipin_5.LATCH_3_.latch/Q _129_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_198_ chanx_right_in[0] chanx_left_out[0] vgnd vpwr scs8hd_buf_2
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_2.LATCH_3_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_10_ vgnd vpwr scs8hd_inv_1
XFILLER_2_30 vgnd vpwr scs8hd_fill_1
XFILLER_20_323 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_5.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_1_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
X_121_ _102_/X _122_/B _121_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_301 vgnd vpwr scs8hd_decap_4
XANTENNA__199__A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_4_308 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_104_ _104_/A _104_/X vgnd vpwr scs8hd_buf_1
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_175 vpwr vgnd scs8hd_fill_2
XFILLER_19_297 vpwr vgnd scs8hd_fill_2
XFILLER_19_231 vgnd vpwr scs8hd_decap_12
XFILLER_6_190 vpwr vgnd scs8hd_fill_2
XFILLER_8_84 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_2_.latch/Q mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_300 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_366 vgnd vpwr scs8hd_decap_6
XFILLER_17_93 vpwr vgnd scs8hd_fill_2
XFILLER_17_82 vpwr vgnd scs8hd_fill_2
XFILLER_17_71 vpwr vgnd scs8hd_fill_2
XFILLER_16_267 vpwr vgnd scs8hd_fill_2
XFILLER_16_256 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_3 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _182_/HI mem_top_ipin_0.LATCH_5_.latch/Q
+ mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_ipin_2.LATCH_2_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_219 vpwr vgnd scs8hd_fill_2
XFILLER_0_196 vpwr vgnd scs8hd_fill_2
XFILLER_8_241 vgnd vpwr scs8hd_decap_4
XFILLER_8_274 vgnd vpwr scs8hd_fill_1
XFILLER_8_285 vpwr vgnd scs8hd_fill_2
XFILLER_10_207 vgnd vpwr scs8hd_decap_4
XFILLER_2_406 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_8 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_211 vpwr vgnd scs8hd_fill_2
XFILLER_2_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_60 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_71 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_14_398 vgnd vpwr scs8hd_decap_8
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_197_ chanx_right_in[1] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_97 vgnd vpwr scs8hd_decap_4
XFILLER_2_20 vpwr vgnd scs8hd_fill_2
XFILLER_1_280 vpwr vgnd scs8hd_fill_2
XFILLER_20_335 vgnd vpwr scs8hd_decap_6
XFILLER_9_380 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_120_ _138_/A _122_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_324 vpwr vgnd scs8hd_fill_2
XFILLER_11_40 vgnd vpwr scs8hd_decap_4
XFILLER_11_51 vpwr vgnd scs8hd_fill_2
XFILLER_11_62 vpwr vgnd scs8hd_fill_2
XFILLER_11_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB _175_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_187 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_3.INVTX1_4_.scs8hd_inv_1 chanx_left_in[6] mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_103_ _102_/X _103_/B _103_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_136 vpwr vgnd scs8hd_fill_2
XFILLER_19_243 vgnd vpwr scs8hd_fill_1
XFILLER_14_7 vpwr vgnd scs8hd_fill_2
XFILLER_8_41 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_117 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_16_213 vgnd vpwr scs8hd_fill_1
XFILLER_16_279 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _153_/A mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_5_404 vgnd vpwr scs8hd_decap_3
XFILLER_0_120 vpwr vgnd scs8hd_fill_2
XFILLER_8_264 vpwr vgnd scs8hd_fill_2
XFILLER_12_271 vgnd vpwr scs8hd_decap_4
XFILLER_5_53 vgnd vpwr scs8hd_decap_4
XFILLER_14_84 vgnd vpwr scs8hd_decap_8
XFILLER_5_234 vgnd vpwr scs8hd_decap_4
XFILLER_5_278 vgnd vpwr scs8hd_decap_4
XFILLER_17_330 vgnd vpwr scs8hd_decap_12
XANTENNA__101__A _138_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_215 vpwr vgnd scs8hd_fill_2
XFILLER_14_333 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_ipin_7.LATCH_2_.latch_SLEEPB _146_/Y vgnd vpwr scs8hd_diode_2
X_196_ chanx_right_in[2] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_2_32 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_2_.latch/Q mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_171 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_392 vgnd vpwr scs8hd_decap_4
XFILLER_15_119 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_329 vpwr vgnd scs8hd_fill_2
XFILLER_11_347 vpwr vgnd scs8hd_fill_2
XFILLER_11_358 vpwr vgnd scs8hd_fill_2
XFILLER_2_3 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_163 vgnd vpwr scs8hd_decap_8
X_179_ _179_/HI _179_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_395 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_1.LATCH_3_.latch data_in mem_top_ipin_1.LATCH_3_.latch/Q _082_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_199 vgnd vpwr scs8hd_decap_12
XFILLER_16_406 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_155 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
X_102_ _102_/A _102_/X vgnd vpwr scs8hd_buf_1
XFILLER_3_332 vgnd vpwr scs8hd_decap_4
XFILLER_3_343 vpwr vgnd scs8hd_fill_2
XFILLER_3_354 vpwr vgnd scs8hd_fill_2
XFILLER_7_115 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_64 vgnd vpwr scs8hd_decap_3
XFILLER_8_97 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__104__A _104_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_162 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_3_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_239 vgnd vpwr scs8hd_decap_3
XFILLER_5_10 vpwr vgnd scs8hd_fill_2
XFILLER_8_298 vpwr vgnd scs8hd_fill_2
XFILLER_12_250 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_41 vgnd vpwr scs8hd_decap_3
XFILLER_14_30 vgnd vpwr scs8hd_fill_1
XFILLER_17_342 vgnd vpwr scs8hd_decap_12
XANTENNA__101__B _103_/B vgnd vpwr scs8hd_diode_2
XANTENNA__202__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_2_205 vgnd vpwr scs8hd_decap_4
XFILLER_4_7 vgnd vpwr scs8hd_decap_3
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_14_301 vgnd vpwr scs8hd_decap_4
XPHY_62 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_51 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_195_ chanx_right_in[3] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_2_55 vpwr vgnd scs8hd_fill_2
XFILLER_2_44 vgnd vpwr scs8hd_decap_8
XFILLER_1_293 vpwr vgnd scs8hd_fill_2
XANTENNA__112__A _138_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_194 vpwr vgnd scs8hd_fill_2
XFILLER_17_161 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_304 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_4_.latch_SLEEPB _110_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_319 vgnd vpwr scs8hd_fill_1
Xmem_top_ipin_4.LATCH_2_.latch data_in mem_top_ipin_4.LATCH_2_.latch/Q _120_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_175 vgnd vpwr scs8hd_decap_6
XANTENNA__107__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_370 vpwr vgnd scs8hd_fill_2
X_178_ _104_/A _178_/B _178_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_20_156 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_0.LATCH_3_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_top_ipin_6.LATCH_5_.latch data_in mem_top_ipin_6.LATCH_5_.latch/Q _135_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_101_ _138_/A _103_/B _101_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_105 vpwr vgnd scs8hd_fill_2
XFILLER_11_134 vpwr vgnd scs8hd_fill_2
XFILLER_19_245 vgnd vpwr scs8hd_decap_12
XFILLER_8_10 vpwr vgnd scs8hd_fill_2
XFILLER_0_325 vpwr vgnd scs8hd_fill_2
XFILLER_0_314 vpwr vgnd scs8hd_fill_2
XFILLER_16_248 vgnd vpwr scs8hd_decap_4
XFILLER_16_226 vpwr vgnd scs8hd_fill_2
XFILLER_3_141 vpwr vgnd scs8hd_fill_2
XANTENNA__120__A _138_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__205__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_5_.latch_SLEEPB _075_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_2_.latch/Q mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_177 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__115__A _163_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_222 vpwr vgnd scs8hd_fill_2
XFILLER_5_77 vpwr vgnd scs8hd_fill_2
XFILLER_5_99 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_3
XFILLER_14_20 vpwr vgnd scs8hd_fill_2
XFILLER_17_354 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_5.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_107 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_14_346 vpwr vgnd scs8hd_fill_2
XPHY_63 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_52 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_194_ chanx_right_in[4] chanx_left_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_2_89 vgnd vpwr scs8hd_fill_1
XANTENNA__112__B _108_/X vgnd vpwr scs8hd_diode_2
XFILLER_17_184 vgnd vpwr scs8hd_fill_1
Xmem_top_ipin_7.LATCH_1_.latch data_in mem_top_ipin_7.LATCH_1_.latch/Q _147_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_309 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_6.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_405 vpwr vgnd scs8hd_fill_2
XFILLER_14_132 vpwr vgnd scs8hd_fill_2
XANTENNA__107__B _073_/B vgnd vpwr scs8hd_diode_2
X_177_ _102_/A _178_/B _177_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_320 vpwr vgnd scs8hd_fill_2
XANTENNA__123__A enable vgnd vpwr scs8hd_diode_2
XFILLER_6_364 vpwr vgnd scs8hd_fill_2
XFILLER_6_375 vgnd vpwr scs8hd_decap_12
XFILLER_20_168 vgnd vpwr scs8hd_decap_12
X_100_ _168_/A _138_/A vgnd vpwr scs8hd_buf_1
XFILLER_11_179 vgnd vpwr scs8hd_decap_4
XFILLER_3_367 vpwr vgnd scs8hd_fill_2
XFILLER_19_257 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_183 vgnd vpwr scs8hd_fill_1
XFILLER_6_194 vgnd vpwr scs8hd_decap_3
XFILLER_8_88 vpwr vgnd scs8hd_fill_2
XFILLER_0_304 vpwr vgnd scs8hd_fill_2
XFILLER_16_205 vpwr vgnd scs8hd_fill_2
XFILLER_17_97 vpwr vgnd scs8hd_fill_2
XFILLER_17_86 vgnd vpwr scs8hd_decap_4
XFILLER_17_75 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_175 vpwr vgnd scs8hd_fill_2
XANTENNA__120__B _122_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_4
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__115__B _152_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_289 vgnd vpwr scs8hd_decap_6
XANTENNA__131__A _102_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_215 vpwr vgnd scs8hd_fill_2
XFILLER_5_259 vpwr vgnd scs8hd_fill_2
XFILLER_17_377 vpwr vgnd scs8hd_fill_2
XANTENNA__126__A _125_/X vgnd vpwr scs8hd_diode_2
XFILLER_18_119 vgnd vpwr scs8hd_decap_12
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_14_325 vgnd vpwr scs8hd_decap_6
XFILLER_14_314 vgnd vpwr scs8hd_decap_6
XPHY_64 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_53 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_42 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_20 vgnd vpwr scs8hd_decap_3
X_193_ chanx_right_in[5] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_top_ipin_6.LATCH_5_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_240 vpwr vgnd scs8hd_fill_2
XFILLER_2_24 vgnd vpwr scs8hd_decap_6
XFILLER_17_152 vgnd vpwr scs8hd_decap_6
XFILLER_17_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_362 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB _178_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_306 vgnd vpwr scs8hd_decap_3
XFILLER_11_328 vpwr vgnd scs8hd_fill_2
XFILLER_11_55 vgnd vpwr scs8hd_decap_4
XFILLER_11_88 vpwr vgnd scs8hd_fill_2
XFILLER_14_111 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_3.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_176_ _168_/A _178_/B _176_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__107__C _073_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_354 vgnd vpwr scs8hd_fill_1
XFILLER_6_387 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_398 vgnd vpwr scs8hd_decap_8
XFILLER_20_125 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_9_170 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_3_302 vgnd vpwr scs8hd_fill_1
XFILLER_0_3 vgnd vpwr scs8hd_decap_6
XFILLER_19_269 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_0.LATCH_2_.latch data_in mem_top_ipin_0.LATCH_2_.latch/Q _176_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
XANTENNA__118__B _122_/B vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_4.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_159_ _167_/A _156_/X _159_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__134__A _133_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_162 vgnd vpwr scs8hd_decap_4
XFILLER_16_239 vpwr vgnd scs8hd_fill_2
XFILLER_3_132 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_2.LATCH_5_.latch data_in mem_top_ipin_2.LATCH_5_.latch/Q _095_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_0_.latch/Q mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__129__A _111_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_202 vgnd vpwr scs8hd_decap_4
XFILLER_8_268 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__131__B _126_/X vgnd vpwr scs8hd_diode_2
XANTENNA__115__C _073_/C vgnd vpwr scs8hd_diode_2
XFILLER_5_57 vgnd vpwr scs8hd_fill_1
XFILLER_14_66 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_2_.latch data_in mem_bottom_ipin_0.LATCH_2_.latch/Q _160_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_367 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_ipin_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _142_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_219 vgnd vpwr scs8hd_decap_4
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_54 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_43 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_2.LATCH_5_.latch data_in mem_bottom_ipin_2.LATCH_5_.latch/Q _165_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_192_ chanx_right_in[6] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_1_263 vgnd vpwr scs8hd_fill_1
XFILLER_17_120 vpwr vgnd scs8hd_fill_2
XFILLER_2_36 vgnd vpwr scs8hd_decap_3
XFILLER_17_175 vgnd vpwr scs8hd_decap_6
XFILLER_13_381 vgnd vpwr scs8hd_decap_12
XANTENNA__137__A _111_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_352 vgnd vpwr scs8hd_fill_1
XFILLER_11_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_2_7 vpwr vgnd scs8hd_fill_2
XFILLER_14_145 vpwr vgnd scs8hd_fill_2
X_175_ _167_/A _178_/B _175_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_395 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_20_137 vgnd vpwr scs8hd_decap_12
XFILLER_9_193 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_3.LATCH_1_.latch data_in mem_top_ipin_3.LATCH_1_.latch/Q _113_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_ipin_5.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ _154_/A mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_3_336 vgnd vpwr scs8hd_fill_1
XFILLER_7_119 vgnd vpwr scs8hd_decap_3
XFILLER_11_159 vgnd vpwr scs8hd_decap_4
XFILLER_3_347 vgnd vpwr scs8hd_decap_4
XFILLER_3_358 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_6.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_158_ _166_/A _156_/X _158_/Y vgnd vpwr scs8hd_nor2_4
X_089_ address[1] address[2] address[0] _090_/A vgnd vpwr scs8hd_or3_4
XANTENNA__150__A _149_/X vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_5.LATCH_4_.latch data_in mem_top_ipin_5.LATCH_4_.latch/Q _128_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_5.LATCH_0_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_11 vgnd vpwr scs8hd_decap_4
XFILLER_16_218 vgnd vpwr scs8hd_decap_8
XFILLER_8_406 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_111 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_9 vgnd vpwr scs8hd_fill_1
XFILLER_15_240 vpwr vgnd scs8hd_fill_2
XANTENNA__129__B _126_/X vgnd vpwr scs8hd_diode_2
XANTENNA__145__A _111_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.INVTX1_5_.scs8hd_inv_1 chanx_right_in[5] mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_103 vpwr vgnd scs8hd_fill_2
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XFILLER_12_210 vpwr vgnd scs8hd_fill_2
XFILLER_8_247 vpwr vgnd scs8hd_fill_2
XFILLER_8_258 vgnd vpwr scs8hd_decap_4
XFILLER_12_254 vpwr vgnd scs8hd_fill_2
XFILLER_12_287 vgnd vpwr scs8hd_decap_8
XFILLER_5_25 vpwr vgnd scs8hd_fill_2
XFILLER_5_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_2_ vgnd vpwr scs8hd_inv_1
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_2.LATCH_4_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_283 vgnd vpwr scs8hd_fill_1
XPHY_33 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_66 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_55 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_44 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_3.LATCH_1_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
X_191_ chanx_right_in[7] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_2_59 vpwr vgnd scs8hd_fill_2
XFILLER_1_297 vpwr vgnd scs8hd_fill_2
XFILLER_17_198 vgnd vpwr scs8hd_decap_4
XFILLER_13_393 vgnd vpwr scs8hd_decap_12
XFILLER_13_360 vgnd vpwr scs8hd_decap_6
XANTENNA__137__B _140_/B vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _153_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_46 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_0_.latch/Q mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_102 vgnd vpwr scs8hd_decap_6
Xmem_top_ipin_6.LATCH_0_.latch data_in mem_top_ipin_6.LATCH_0_.latch/Q _140_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_174_ _166_/A _178_/B _174_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_374 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__148__A _104_/X vgnd vpwr scs8hd_diode_2
XFILLER_20_149 vgnd vpwr scs8hd_decap_6
XFILLER_7_109 vgnd vpwr scs8hd_decap_4
XFILLER_11_105 vpwr vgnd scs8hd_fill_2
XFILLER_11_138 vgnd vpwr scs8hd_decap_4
XFILLER_3_315 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_131 vpwr vgnd scs8hd_fill_2
XFILLER_8_58 vgnd vpwr scs8hd_decap_4
XFILLER_8_69 vgnd vpwr scs8hd_decap_4
XFILLER_10_182 vpwr vgnd scs8hd_fill_2
X_157_ _068_/A _156_/X _157_/Y vgnd vpwr scs8hd_nor2_4
X_088_ _082_/A _102_/A _088_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_186 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_329 vgnd vpwr scs8hd_decap_12
XFILLER_0_318 vgnd vpwr scs8hd_decap_4
XFILLER_17_23 vgnd vpwr scs8hd_decap_12
XFILLER_3_145 vpwr vgnd scs8hd_fill_2
XFILLER_15_285 vgnd vpwr scs8hd_fill_1
XFILLER_15_263 vgnd vpwr scs8hd_fill_1
XANTENNA__145__B _142_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_2_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__161__A _102_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__071__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_215 vpwr vgnd scs8hd_fill_2
XFILLER_8_226 vpwr vgnd scs8hd_fill_2
XANTENNA__156__A _156_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_24 vgnd vpwr scs8hd_decap_6
XANTENNA__066__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_14_46 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_251 vgnd vpwr scs8hd_decap_8
XFILLER_4_262 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
X_190_ chanx_right_in[8] chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XPHY_67 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_56 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_45 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XFILLER_1_276 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_6.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_376 vpwr vgnd scs8hd_fill_2
XFILLER_11_69 vpwr vgnd scs8hd_fill_2
X_173_ _068_/A _178_/B _173_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_302 vgnd vpwr scs8hd_decap_6
XFILLER_6_324 vpwr vgnd scs8hd_fill_2
XFILLER_6_346 vgnd vpwr scs8hd_decap_8
XFILLER_6_368 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_106 vgnd vpwr scs8hd_decap_12
XANTENNA__148__B _142_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__164__A _163_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_81 vpwr vgnd scs8hd_fill_2
XANTENNA__074__A _073_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
X_156_ _156_/A _156_/X vgnd vpwr scs8hd_buf_1
X_087_ _087_/A _102_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_110 vgnd vpwr scs8hd_decap_6
XFILLER_6_154 vgnd vpwr scs8hd_decap_3
XANTENNA__159__A _167_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_308 vpwr vgnd scs8hd_fill_2
XANTENNA__069__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
XFILLER_17_35 vgnd vpwr scs8hd_decap_12
XFILLER_16_209 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _180_/HI _153_/Y mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_297 vpwr vgnd scs8hd_fill_2
XFILLER_15_275 vpwr vgnd scs8hd_fill_2
XFILLER_15_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
X_139_ _102_/X _140_/B _139_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__161__B _156_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_1.LATCH_4_.latch data_in mem_top_ipin_1.LATCH_4_.latch/Q _078_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_267 vpwr vgnd scs8hd_fill_2
XFILLER_10_8 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _182_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__172__A _171_/X vgnd vpwr scs8hd_diode_2
XFILLER_7_271 vgnd vpwr scs8hd_decap_4
XFILLER_7_282 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_0_.latch/Q mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_58 vgnd vpwr scs8hd_decap_6
XANTENNA__066__B _076_/B vgnd vpwr scs8hd_diode_2
XANTENNA__082__A _082_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_403 vgnd vpwr scs8hd_decap_4
XFILLER_17_304 vgnd vpwr scs8hd_fill_1
XANTENNA__167__A _167_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_6.LATCH_2_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
XPHY_35 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A _076_/X vgnd vpwr scs8hd_diode_2
XPHY_46 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_13 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_68 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_222 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vgnd vpwr scs8hd_decap_4
XFILLER_17_112 vgnd vpwr scs8hd_decap_8
XFILLER_1_266 vgnd vpwr scs8hd_fill_1
XFILLER_17_167 vgnd vpwr scs8hd_fill_1
XFILLER_17_145 vgnd vpwr scs8hd_decap_4
XFILLER_17_123 vgnd vpwr scs8hd_decap_12
XFILLER_15_90 vgnd vpwr scs8hd_decap_3
XFILLER_9_344 vpwr vgnd scs8hd_fill_2
XFILLER_9_388 vpwr vgnd scs8hd_fill_2
XFILLER_9_399 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _180_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
X_172_ _171_/X _178_/B vgnd vpwr scs8hd_buf_1
XFILLER_10_387 vgnd vpwr scs8hd_decap_8
XFILLER_10_398 vgnd vpwr scs8hd_decap_8
XFILLER_20_118 vgnd vpwr scs8hd_decap_6
XFILLER_9_152 vpwr vgnd scs8hd_fill_2
XFILLER_5_380 vgnd vpwr scs8hd_decap_12
XFILLER_9_174 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_71 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_4.INVTX1_2_.scs8hd_inv_1 chanx_left_in[6] mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XANTENNA__090__A _090_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_339 vgnd vpwr scs8hd_fill_1
XFILLER_19_207 vgnd vpwr scs8hd_decap_12
XFILLER_8_27 vpwr vgnd scs8hd_fill_2
X_086_ address[1] address[2] _151_/D _087_/A vgnd vpwr scs8hd_or3_4
X_155_ _073_/A _073_/B _163_/C _156_/A vgnd vpwr scs8hd_or3_4
XFILLER_12_91 vgnd vpwr scs8hd_fill_1
XFILLER_18_284 vgnd vpwr scs8hd_fill_1
XANTENNA__159__B _156_/X vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_2.LATCH_0_.latch data_in mem_top_ipin_2.LATCH_0_.latch/Q _105_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__175__A _167_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_47 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_4.LATCH_3_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__085__A _082_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_136 vgnd vpwr scs8hd_decap_3
XFILLER_3_158 vpwr vgnd scs8hd_fill_2
X_207_ chanx_left_in[0] chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_top_ipin_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_138_ _138_/A _140_/B _138_/Y vgnd vpwr scs8hd_nor2_4
X_069_ address[4] _073_/A vgnd vpwr scs8hd_buf_1
Xmem_top_ipin_4.LATCH_3_.latch data_in mem_top_ipin_4.LATCH_3_.latch/Q _119_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_94 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_81 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_ipin_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_128 vgnd vpwr scs8hd_decap_4
XFILLER_12_224 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__066__C _151_/D vgnd vpwr scs8hd_diode_2
XANTENNA__082__B _167_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_0_.latch data_in mem_bottom_ipin_2.LATCH_0_.latch/Q _170_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_286 vpwr vgnd scs8hd_fill_2
XANTENNA__167__B _166_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_93 vpwr vgnd scs8hd_fill_2
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_47 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_69 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__093__A _073_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_245 vgnd vpwr scs8hd_decap_3
XFILLER_1_201 vpwr vgnd scs8hd_fill_2
XFILLER_17_135 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_ipin_6.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_4_.latch_SLEEPB _097_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_352 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _154_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_301 vpwr vgnd scs8hd_fill_2
XFILLER_9_323 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_7.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__178__A _104_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_0.LATCH_4_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_27 vpwr vgnd scs8hd_fill_2
XANTENNA__088__A _082_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_171_ _163_/A _152_/B _163_/C _171_/X vgnd vpwr scs8hd_or3_4
XFILLER_10_311 vpwr vgnd scs8hd_fill_2
XFILLER_13_160 vpwr vgnd scs8hd_fill_2
XFILLER_9_120 vpwr vgnd scs8hd_fill_2
XFILLER_5_392 vgnd vpwr scs8hd_decap_12
XFILLER_9_197 vpwr vgnd scs8hd_fill_2
XFILLER_3_94 vpwr vgnd scs8hd_fill_2
XFILLER_19_219 vgnd vpwr scs8hd_decap_12
XFILLER_15_403 vgnd vpwr scs8hd_decap_4
XFILLER_2_340 vgnd vpwr scs8hd_decap_8
X_085_ _082_/A _168_/A _085_/Y vgnd vpwr scs8hd_nor2_4
X_154_ _154_/A _154_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_145 vpwr vgnd scs8hd_fill_2
XFILLER_10_163 vgnd vpwr scs8hd_decap_3
XFILLER_2_395 vpwr vgnd scs8hd_fill_2
XFILLER_2_351 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_4.LATCH_0_.latch/Q mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__175__B _178_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__191__A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_7.LATCH_2_.latch data_in mem_top_ipin_7.LATCH_2_.latch/Q _146_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__085__B _168_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_406 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_2.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_115 vgnd vpwr scs8hd_fill_1
XFILLER_15_255 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_206_ chanx_left_in[1] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
X_137_ _111_/A _140_/B _137_/Y vgnd vpwr scs8hd_nor2_4
X_068_ _068_/A _068_/X vgnd vpwr scs8hd_buf_1
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB _173_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_71 vgnd vpwr scs8hd_decap_4
XANTENNA__096__A _166_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_280 vgnd vpwr scs8hd_decap_12
XFILLER_12_236 vgnd vpwr scs8hd_decap_3
XFILLER_5_29 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_8_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _183_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_291 vgnd vpwr scs8hd_decap_4
XFILLER_17_306 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_59 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_48 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_15 vgnd vpwr scs8hd_decap_3
XANTENNA__093__B _152_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_158 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_191 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__194__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA__178__B _178_/B vgnd vpwr scs8hd_diode_2
XANTENNA__088__B _102_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_128 vpwr vgnd scs8hd_fill_2
X_170_ _104_/A _166_/B _170_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_334 vpwr vgnd scs8hd_fill_2
XFILLER_10_356 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_109 vgnd vpwr scs8hd_decap_3
XFILLER_3_319 vpwr vgnd scs8hd_fill_2
XANTENNA__099__A _111_/A vgnd vpwr scs8hd_diode_2
X_153_ _153_/A _153_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_135 vgnd vpwr scs8hd_fill_1
XFILLER_10_186 vgnd vpwr scs8hd_decap_6
XFILLER_2_363 vgnd vpwr scs8hd_decap_12
X_084_ _083_/X _168_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_168 vpwr vgnd scs8hd_fill_2
XFILLER_6_179 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_7.LATCH_4_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_7 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_245 vgnd vpwr scs8hd_fill_1
X_205_ chanx_left_in[2] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
X_136_ _096_/X _140_/B _136_/Y vgnd vpwr scs8hd_nor2_4
X_067_ _066_/X _068_/A vgnd vpwr scs8hd_buf_1
Xmux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_7.LATCH_3_.latch/Q mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_41 vpwr vgnd scs8hd_fill_2
XFILLER_0_63 vpwr vgnd scs8hd_fill_2
XFILLER_0_74 vpwr vgnd scs8hd_fill_2
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XFILLER_20_292 vgnd vpwr scs8hd_decap_12
XFILLER_8_208 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[3] mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_119_ _111_/A _122_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_296 vgnd vpwr scs8hd_decap_4
XFILLER_19_381 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_0.LATCH_3_.latch data_in mem_top_ipin_0.LATCH_3_.latch/Q _175_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__197__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_17_318 vgnd vpwr scs8hd_decap_12
XFILLER_4_266 vgnd vpwr scs8hd_fill_1
XFILLER_16_340 vgnd vpwr scs8hd_decap_8
XFILLER_6_51 vgnd vpwr scs8hd_decap_4
XFILLER_6_84 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_5.LATCH_5_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_16 vgnd vpwr scs8hd_decap_3
XANTENNA__093__C _073_/C vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_3.LATCH_0_.latch/Q mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_236 vpwr vgnd scs8hd_fill_2
XFILLER_17_104 vpwr vgnd scs8hd_fill_2
XFILLER_9_358 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_7.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_324 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_328 vgnd vpwr scs8hd_decap_8
XFILLER_13_195 vpwr vgnd scs8hd_fill_2
XFILLER_13_173 vpwr vgnd scs8hd_fill_2
XFILLER_9_144 vpwr vgnd scs8hd_fill_2
XFILLER_3_52 vpwr vgnd scs8hd_fill_2
XFILLER_5_361 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_0.LATCH_3_.latch data_in mem_bottom_ipin_0.LATCH_3_.latch/Q _159_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__099__B _103_/B vgnd vpwr scs8hd_diode_2
X_083_ _080_/A address[2] address[0] _083_/X vgnd vpwr scs8hd_or3_4
X_152_ _073_/A _152_/B _163_/C address[0] _152_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_2_375 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_7.LATCH_1_.latch/Q mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_276 vgnd vpwr scs8hd_decap_8
XFILLER_15_202 vpwr vgnd scs8hd_fill_2
X_204_ chanx_left_in[3] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_15_279 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_066_ address[1] _076_/B _151_/D _066_/X vgnd vpwr scs8hd_or3_4
X_135_ _068_/X _140_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_172 vpwr vgnd scs8hd_fill_2
XFILLER_2_150 vgnd vpwr scs8hd_fill_1
XFILLER_9_95 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_3.LATCH_2_.latch data_in mem_top_ipin_3.LATCH_2_.latch/Q _112_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _184_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_275 vgnd vpwr scs8hd_fill_1
X_118_ _096_/X _122_/B _118_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_19_393 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_5.LATCH_5_.latch data_in mem_top_ipin_5.LATCH_5_.latch/Q _127_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_94 vgnd vpwr scs8hd_decap_12
XFILLER_4_201 vpwr vgnd scs8hd_fill_2
XFILLER_4_234 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_41 vgnd vpwr scs8hd_decap_8
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_1_259 vgnd vpwr scs8hd_decap_4
XFILLER_13_333 vgnd vpwr scs8hd_decap_4
XFILLER_13_377 vpwr vgnd scs8hd_fill_2
XFILLER_9_315 vpwr vgnd scs8hd_fill_2
XFILLER_9_348 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_0_270 vpwr vgnd scs8hd_fill_2
XFILLER_16_171 vgnd vpwr scs8hd_decap_8
XFILLER_16_160 vpwr vgnd scs8hd_fill_2
XFILLER_14_108 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ _154_/Y mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_14_ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_ipin_6.LATCH_3_.latch/Q mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_9_112 vpwr vgnd scs8hd_fill_2
XFILLER_9_123 vgnd vpwr scs8hd_decap_4
XFILLER_9_156 vgnd vpwr scs8hd_decap_3
XFILLER_9_178 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_4.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_5.INVTX1_3_.scs8hd_inv_1 chanx_right_in[7] mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_151_ _073_/A _152_/B _163_/C _151_/D _151_/Y vgnd vpwr scs8hd_nor4_4
X_082_ _082_/A _167_/A _082_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_133 vgnd vpwr scs8hd_fill_1
XFILLER_12_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_398 vgnd vpwr scs8hd_decap_8
XFILLER_2_387 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_4.LATCH_0_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_288 vgnd vpwr scs8hd_decap_12
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
X_203_ chanx_left_in[4] chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_15_236 vpwr vgnd scs8hd_fill_2
X_065_ address[0] _151_/D vgnd vpwr scs8hd_inv_8
X_134_ _133_/X _140_/B vgnd vpwr scs8hd_buf_1
XFILLER_0_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XFILLER_14_280 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_6.LATCH_1_.latch data_in mem_top_ipin_6.LATCH_1_.latch/Q _139_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_9_41 vpwr vgnd scs8hd_fill_2
XFILLER_9_52 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_2.LATCH_0_.latch/Q mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_206 vpwr vgnd scs8hd_fill_2
XFILLER_12_228 vgnd vpwr scs8hd_decap_8
XFILLER_20_261 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _153_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _181_/HI mem_bottom_ipin_2.LATCH_5_.latch/Q
+ mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_7_221 vgnd vpwr scs8hd_decap_3
XFILLER_7_254 vpwr vgnd scs8hd_fill_2
X_117_ _068_/X _122_/B _117_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_272 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_213 vgnd vpwr scs8hd_fill_1
XFILLER_4_279 vgnd vpwr scs8hd_decap_4
XFILLER_16_353 vgnd vpwr scs8hd_decap_12
XFILLER_16_320 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB _103_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_97 vpwr vgnd scs8hd_fill_2
XFILLER_19_191 vpwr vgnd scs8hd_fill_2
XPHY_29 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
XFILLER_1_205 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_6.LATCH_1_.latch/Q mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_73 vpwr vgnd scs8hd_fill_2
XFILLER_15_62 vpwr vgnd scs8hd_fill_2
XFILLER_15_40 vpwr vgnd scs8hd_fill_2
XFILLER_13_367 vgnd vpwr scs8hd_decap_4
XFILLER_13_356 vpwr vgnd scs8hd_fill_2
XFILLER_13_312 vpwr vgnd scs8hd_fill_2
XFILLER_13_301 vpwr vgnd scs8hd_fill_2
XFILLER_15_95 vgnd vpwr scs8hd_decap_3
XANTENNA__102__A _102_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_183 vpwr vgnd scs8hd_fill_2
XFILLER_6_308 vgnd vpwr scs8hd_fill_1
XFILLER_10_348 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_142 vgnd vpwr scs8hd_fill_1
XFILLER_3_98 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_150_ _149_/X _163_/C vgnd vpwr scs8hd_buf_1
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_322 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_081_ _080_/X _167_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_127 vpwr vgnd scs8hd_fill_2
XFILLER_6_149 vpwr vgnd scs8hd_fill_2
XFILLER_10_145 vpwr vgnd scs8hd_fill_2
XFILLER_12_74 vgnd vpwr scs8hd_decap_3
XFILLER_12_85 vgnd vpwr scs8hd_decap_6
XFILLER_2_333 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_193 vgnd vpwr scs8hd_decap_4
XFILLER_17_19 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB _176_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__200__A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_15_259 vgnd vpwr scs8hd_decap_4
XFILLER_15_215 vpwr vgnd scs8hd_fill_2
X_202_ chanx_left_in[5] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
X_133_ address[4] _152_/B _141_/C _124_/X _133_/X vgnd vpwr scs8hd_or4_4
XFILLER_7_403 vgnd vpwr scs8hd_decap_4
XFILLER_2_163 vgnd vpwr scs8hd_decap_3
X_064_ address[2] _076_/B vgnd vpwr scs8hd_inv_8
XFILLER_17_7 vpwr vgnd scs8hd_fill_2
XANTENNA__110__A _096_/X vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_3.INVTX1_3_.scs8hd_inv_1 chanx_right_in[5] mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_99 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_14_ vgnd vpwr scs8hd_inv_1
XFILLER_20_273 vgnd vpwr scs8hd_decap_6
XFILLER_4_406 vgnd vpwr scs8hd_fill_1
XANTENNA__105__A _104_/X vgnd vpwr scs8hd_diode_2
X_116_ _116_/A _122_/B vgnd vpwr scs8hd_buf_1
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _185_/HI vgnd vpwr
+ scs8hd_diode_2
Xmux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_5.LATCH_3_.latch/Q mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_20_63 vgnd vpwr scs8hd_decap_12
XFILLER_4_269 vgnd vpwr scs8hd_decap_6
XFILLER_16_398 vgnd vpwr scs8hd_decap_8
XFILLER_16_365 vgnd vpwr scs8hd_decap_12
XPHY_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_9 vpwr vgnd scs8hd_fill_2
XFILLER_0_283 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_1.LATCH_5_.latch data_in mem_top_ipin_1.LATCH_5_.latch/Q _075_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_195 vgnd vpwr scs8hd_fill_1
XFILLER_8_394 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_10_305 vgnd vpwr scs8hd_decap_4
XANTENNA__203__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_7_6 vpwr vgnd scs8hd_fill_2
XFILLER_13_132 vgnd vpwr scs8hd_decap_4
XANTENNA__113__A _102_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_353 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_1.LATCH_0_.latch/Q mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_77 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_7.LATCH_1_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_080_ _080_/A address[2] _151_/D _080_/X vgnd vpwr scs8hd_or3_4
XFILLER_10_102 vpwr vgnd scs8hd_fill_2
XFILLER_10_168 vgnd vpwr scs8hd_decap_3
XFILLER_18_257 vgnd vpwr scs8hd_decap_12
XFILLER_18_246 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__108__A _108_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
X_201_ chanx_left_in[6] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
X_132_ _104_/X _126_/X _132_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_197 vpwr vgnd scs8hd_fill_2
XFILLER_2_142 vpwr vgnd scs8hd_fill_2
XFILLER_2_131 vpwr vgnd scs8hd_fill_2
XANTENNA__110__B _108_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_12 vpwr vgnd scs8hd_fill_2
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_78 vgnd vpwr scs8hd_decap_4
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_5.LATCH_1_.latch/Q mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_230 vgnd vpwr scs8hd_decap_12
XFILLER_18_74 vgnd vpwr scs8hd_decap_12
XFILLER_18_63 vgnd vpwr scs8hd_decap_8
XFILLER_18_96 vgnd vpwr scs8hd_decap_8
XFILLER_11_230 vgnd vpwr scs8hd_decap_4
XFILLER_11_241 vgnd vpwr scs8hd_decap_3
XANTENNA__105__B _103_/B vgnd vpwr scs8hd_diode_2
X_115_ _163_/A _152_/B _073_/C _116_/A vgnd vpwr scs8hd_or3_4
XFILLER_7_278 vpwr vgnd scs8hd_fill_2
XANTENNA__121__A _102_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_341 vgnd vpwr scs8hd_decap_12
XFILLER_19_330 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_top_ipin_2.LATCH_1_.latch data_in mem_top_ipin_2.LATCH_1_.latch/Q _103_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_top_ipin_5.LATCH_2_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__206__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_6
XFILLER_20_75 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_377 vgnd vpwr scs8hd_decap_12
XANTENNA__116__A _116_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_3_281 vpwr vgnd scs8hd_fill_2
XFILLER_6_55 vgnd vpwr scs8hd_fill_1
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_19_171 vgnd vpwr scs8hd_decap_12
Xmem_top_ipin_4.LATCH_4_.latch data_in mem_top_ipin_4.LATCH_4_.latch/Q _118_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_1_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_17_108 vpwr vgnd scs8hd_fill_2
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_9_329 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_7.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_262 vpwr vgnd scs8hd_fill_2
XFILLER_16_130 vgnd vpwr scs8hd_decap_12
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_373 vgnd vpwr scs8hd_decap_4
.ends

