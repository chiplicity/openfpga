magic
tech sky130A
magscale 1 2
timestamp 1605200248
<< locali >>
rect 2881 18275 2915 18377
rect 17785 18071 17819 18377
rect 9965 12767 9999 12937
rect 12909 12087 12943 12393
rect 14013 8483 14047 8585
rect 9137 8279 9171 8449
rect 4905 7803 4939 8041
rect 11989 7803 12023 8041
rect 3801 7191 3835 7293
rect 10057 7191 10091 7361
rect 1961 6239 1995 6409
rect 10149 6103 10183 6409
rect 9413 5559 9447 5661
rect 7665 5083 7699 5185
rect 7757 4607 7791 4709
rect 9781 4063 9815 4165
rect 8125 1411 8159 1717
rect 10425 1411 10459 1649
<< viali >>
rect 4261 20553 4295 20587
rect 5273 20553 5307 20587
rect 12633 20553 12667 20587
rect 15761 20553 15795 20587
rect 18797 20553 18831 20587
rect 20177 20553 20211 20587
rect 6929 20485 6963 20519
rect 9781 20485 9815 20519
rect 5825 20417 5859 20451
rect 7481 20417 7515 20451
rect 10333 20417 10367 20451
rect 13185 20417 13219 20451
rect 16865 20417 16899 20451
rect 1777 20349 1811 20383
rect 4077 20349 4111 20383
rect 8493 20349 8527 20383
rect 11345 20349 11379 20383
rect 14197 20349 14231 20383
rect 15577 20349 15611 20383
rect 16681 20349 16715 20383
rect 18613 20349 18647 20383
rect 19993 20349 20027 20383
rect 2044 20281 2078 20315
rect 5733 20281 5767 20315
rect 7389 20281 7423 20315
rect 3157 20213 3191 20247
rect 5641 20213 5675 20247
rect 7297 20213 7331 20247
rect 8677 20213 8711 20247
rect 10149 20213 10183 20247
rect 10241 20213 10275 20247
rect 11529 20213 11563 20247
rect 13001 20213 13035 20247
rect 13093 20213 13127 20247
rect 14381 20213 14415 20247
rect 1961 20009 1995 20043
rect 3065 20009 3099 20043
rect 10609 20009 10643 20043
rect 11069 20009 11103 20043
rect 14289 20009 14323 20043
rect 15761 20009 15795 20043
rect 17693 20009 17727 20043
rect 18797 20009 18831 20043
rect 19901 20009 19935 20043
rect 1777 19873 1811 19907
rect 2881 19873 2915 19907
rect 4445 19873 4479 19907
rect 4537 19873 4571 19907
rect 6633 19873 6667 19907
rect 10977 19873 11011 19907
rect 12541 19873 12575 19907
rect 14105 19873 14139 19907
rect 15577 19873 15611 19907
rect 17509 19873 17543 19907
rect 18613 19873 18647 19907
rect 19717 19873 19751 19907
rect 4629 19805 4663 19839
rect 6377 19805 6411 19839
rect 8585 19805 8619 19839
rect 11253 19805 11287 19839
rect 12633 19805 12667 19839
rect 12817 19805 12851 19839
rect 4077 19737 4111 19771
rect 7757 19669 7791 19703
rect 12173 19669 12207 19703
rect 5549 19465 5583 19499
rect 11529 19465 11563 19499
rect 3157 19329 3191 19363
rect 15025 19329 15059 19363
rect 1501 19261 1535 19295
rect 4169 19261 4203 19295
rect 7113 19261 7147 19295
rect 10149 19261 10183 19295
rect 12449 19261 12483 19295
rect 13737 19261 13771 19295
rect 14841 19261 14875 19295
rect 16129 19261 16163 19295
rect 19533 19261 19567 19295
rect 3065 19193 3099 19227
rect 4436 19193 4470 19227
rect 7380 19193 7414 19227
rect 10416 19193 10450 19227
rect 12725 19193 12759 19227
rect 16405 19193 16439 19227
rect 20637 19193 20671 19227
rect 1685 19125 1719 19159
rect 2605 19125 2639 19159
rect 2973 19125 3007 19159
rect 8493 19125 8527 19159
rect 13921 19125 13955 19159
rect 18061 19125 18095 19159
rect 19717 19125 19751 19159
rect 3065 18921 3099 18955
rect 4077 18921 4111 18955
rect 6101 18921 6135 18955
rect 10149 18921 10183 18955
rect 15669 18921 15703 18955
rect 17325 18921 17359 18955
rect 19901 18921 19935 18955
rect 4537 18853 4571 18887
rect 15761 18853 15795 18887
rect 1777 18785 1811 18819
rect 2881 18785 2915 18819
rect 4445 18785 4479 18819
rect 6009 18785 6043 18819
rect 7461 18785 7495 18819
rect 10057 18785 10091 18819
rect 13001 18785 13035 18819
rect 14105 18785 14139 18819
rect 17233 18785 17267 18819
rect 19717 18785 19751 18819
rect 4629 18717 4663 18751
rect 6193 18717 6227 18751
rect 7205 18717 7239 18751
rect 10241 18717 10275 18751
rect 11253 18717 11287 18751
rect 15945 18717 15979 18751
rect 17509 18717 17543 18751
rect 18429 18717 18463 18751
rect 1961 18581 1995 18615
rect 5641 18581 5675 18615
rect 8585 18581 8619 18615
rect 9689 18581 9723 18615
rect 13185 18581 13219 18615
rect 14289 18581 14323 18615
rect 15301 18581 15335 18615
rect 16865 18581 16899 18615
rect 2881 18377 2915 18411
rect 16957 18377 16991 18411
rect 17785 18377 17819 18411
rect 20729 18377 20763 18411
rect 5917 18309 5951 18343
rect 14013 18309 14047 18343
rect 2881 18241 2915 18275
rect 3617 18241 3651 18275
rect 8217 18241 8251 18275
rect 13001 18241 13035 18275
rect 14657 18241 14691 18275
rect 15577 18241 15611 18275
rect 1777 18173 1811 18207
rect 4537 18173 4571 18207
rect 14473 18173 14507 18207
rect 3433 18105 3467 18139
rect 4804 18105 4838 18139
rect 8484 18105 8518 18139
rect 12909 18105 12943 18139
rect 15822 18105 15856 18139
rect 18521 18241 18555 18275
rect 18705 18241 18739 18275
rect 20545 18173 20579 18207
rect 18429 18105 18463 18139
rect 18889 18105 18923 18139
rect 1961 18037 1995 18071
rect 2973 18037 3007 18071
rect 3341 18037 3375 18071
rect 6837 18037 6871 18071
rect 9597 18037 9631 18071
rect 10425 18037 10459 18071
rect 12449 18037 12483 18071
rect 12817 18037 12851 18071
rect 14381 18037 14415 18071
rect 17785 18037 17819 18071
rect 18061 18037 18095 18071
rect 12081 17833 12115 17867
rect 14289 17833 14323 17867
rect 15301 17833 15335 17867
rect 18797 17833 18831 17867
rect 2053 17697 2087 17731
rect 4344 17697 4378 17731
rect 7389 17697 7423 17731
rect 7656 17697 7690 17731
rect 11989 17697 12023 17731
rect 14105 17697 14139 17731
rect 15669 17697 15703 17731
rect 15761 17697 15795 17731
rect 17233 17697 17267 17731
rect 18889 17697 18923 17731
rect 2329 17629 2363 17663
rect 4077 17629 4111 17663
rect 6285 17629 6319 17663
rect 10609 17629 10643 17663
rect 12173 17629 12207 17663
rect 15853 17629 15887 17663
rect 17325 17629 17359 17663
rect 17509 17629 17543 17663
rect 19073 17629 19107 17663
rect 18429 17561 18463 17595
rect 5457 17493 5491 17527
rect 8769 17493 8803 17527
rect 11621 17493 11655 17527
rect 16865 17493 16899 17527
rect 18245 17493 18279 17527
rect 19257 17493 19291 17527
rect 4445 17289 4479 17323
rect 3617 17221 3651 17255
rect 7665 17221 7699 17255
rect 10241 17221 10275 17255
rect 18061 17221 18095 17255
rect 5089 17153 5123 17187
rect 8217 17153 8251 17187
rect 10885 17153 10919 17187
rect 14289 17153 14323 17187
rect 18521 17153 18555 17187
rect 18613 17153 18647 17187
rect 20177 17153 20211 17187
rect 2237 17085 2271 17119
rect 2504 17085 2538 17119
rect 4905 17085 4939 17119
rect 10609 17085 10643 17119
rect 14105 17085 14139 17119
rect 14197 17085 14231 17119
rect 15301 17085 15335 17119
rect 19993 17085 20027 17119
rect 8033 17017 8067 17051
rect 15557 17017 15591 17051
rect 4813 16949 4847 16983
rect 8125 16949 8159 16983
rect 9229 16949 9263 16983
rect 10701 16949 10735 16983
rect 12449 16949 12483 16983
rect 13737 16949 13771 16983
rect 16681 16949 16715 16983
rect 18429 16949 18463 16983
rect 19625 16949 19659 16983
rect 20085 16949 20119 16983
rect 4537 16745 4571 16779
rect 10149 16745 10183 16779
rect 12265 16745 12299 16779
rect 2329 16677 2363 16711
rect 4445 16677 4479 16711
rect 6377 16677 6411 16711
rect 13645 16677 13679 16711
rect 13829 16677 13863 16711
rect 16120 16677 16154 16711
rect 18429 16677 18463 16711
rect 18521 16677 18555 16711
rect 2053 16609 2087 16643
rect 7389 16609 7423 16643
rect 7656 16609 7690 16643
rect 10517 16609 10551 16643
rect 12633 16609 12667 16643
rect 19625 16609 19659 16643
rect 4721 16541 4755 16575
rect 10609 16541 10643 16575
rect 10701 16541 10735 16575
rect 12725 16541 12759 16575
rect 12909 16541 12943 16575
rect 15853 16541 15887 16575
rect 18613 16541 18647 16575
rect 18061 16473 18095 16507
rect 19809 16473 19843 16507
rect 4077 16405 4111 16439
rect 8769 16405 8803 16439
rect 17233 16405 17267 16439
rect 4721 16201 4755 16235
rect 10793 16133 10827 16167
rect 18061 16133 18095 16167
rect 2421 16065 2455 16099
rect 5365 16065 5399 16099
rect 7665 16065 7699 16099
rect 8585 16065 8619 16099
rect 11345 16065 11379 16099
rect 15669 16065 15703 16099
rect 16773 16065 16807 16099
rect 18613 16065 18647 16099
rect 20177 16065 20211 16099
rect 2145 15997 2179 16031
rect 3433 15997 3467 16031
rect 7481 15997 7515 16031
rect 12817 15997 12851 16031
rect 16589 15997 16623 16031
rect 19993 15997 20027 16031
rect 20085 15997 20119 16031
rect 3709 15929 3743 15963
rect 5089 15929 5123 15963
rect 5181 15929 5215 15963
rect 8830 15929 8864 15963
rect 11161 15929 11195 15963
rect 11253 15929 11287 15963
rect 13084 15929 13118 15963
rect 15485 15929 15519 15963
rect 18429 15929 18463 15963
rect 7021 15861 7055 15895
rect 7389 15861 7423 15895
rect 9965 15861 9999 15895
rect 14197 15861 14231 15895
rect 15025 15861 15059 15895
rect 15393 15861 15427 15895
rect 18521 15861 18555 15895
rect 19625 15861 19659 15895
rect 1409 15657 1443 15691
rect 4261 15657 4295 15691
rect 4721 15657 4755 15691
rect 8033 15657 8067 15691
rect 8401 15657 8435 15691
rect 11253 15657 11287 15691
rect 13645 15657 13679 15691
rect 14013 15657 14047 15691
rect 14105 15657 14139 15691
rect 2881 15589 2915 15623
rect 4629 15589 4663 15623
rect 19257 15589 19291 15623
rect 2789 15521 2823 15555
rect 6092 15521 6126 15555
rect 10057 15521 10091 15555
rect 10149 15521 10183 15555
rect 11621 15521 11655 15555
rect 15301 15521 15335 15555
rect 16856 15521 16890 15555
rect 19165 15521 19199 15555
rect 3065 15453 3099 15487
rect 4813 15453 4847 15487
rect 5825 15453 5859 15487
rect 8493 15453 8527 15487
rect 8585 15453 8619 15487
rect 10241 15453 10275 15487
rect 11713 15453 11747 15487
rect 11805 15453 11839 15487
rect 14197 15453 14231 15487
rect 15577 15453 15611 15487
rect 16589 15453 16623 15487
rect 19349 15453 19383 15487
rect 18797 15385 18831 15419
rect 2421 15317 2455 15351
rect 7205 15317 7239 15351
rect 9689 15317 9723 15351
rect 17969 15317 18003 15351
rect 6837 15113 6871 15147
rect 19625 15113 19659 15147
rect 6469 15045 6503 15079
rect 14933 15045 14967 15079
rect 2881 14977 2915 15011
rect 7389 14977 7423 15011
rect 8585 14977 8619 15011
rect 11345 14977 11379 15011
rect 13185 14977 13219 15011
rect 13369 14977 13403 15011
rect 15393 14977 15427 15011
rect 15485 14977 15519 15011
rect 18613 14977 18647 15011
rect 20177 14977 20211 15011
rect 3801 14909 3835 14943
rect 6653 14909 6687 14943
rect 14841 14909 14875 14943
rect 16681 14909 16715 14943
rect 16957 14909 16991 14943
rect 20085 14909 20119 14943
rect 2605 14841 2639 14875
rect 4068 14841 4102 14875
rect 7205 14841 7239 14875
rect 8852 14841 8886 14875
rect 11161 14841 11195 14875
rect 19993 14841 20027 14875
rect 2237 14773 2271 14807
rect 2697 14773 2731 14807
rect 5181 14773 5215 14807
rect 7297 14773 7331 14807
rect 9965 14773 9999 14807
rect 10793 14773 10827 14807
rect 11253 14773 11287 14807
rect 12725 14773 12759 14807
rect 13093 14773 13127 14807
rect 14657 14773 14691 14807
rect 15301 14773 15335 14807
rect 18061 14773 18095 14807
rect 18429 14773 18463 14807
rect 18521 14773 18555 14807
rect 6469 14569 6503 14603
rect 6837 14569 6871 14603
rect 8033 14569 8067 14603
rect 8401 14569 8435 14603
rect 14289 14569 14323 14603
rect 17141 14569 17175 14603
rect 18245 14569 18279 14603
rect 18705 14569 18739 14603
rect 2044 14501 2078 14535
rect 6929 14501 6963 14535
rect 8493 14501 8527 14535
rect 12164 14501 12198 14535
rect 17049 14501 17083 14535
rect 4813 14433 4847 14467
rect 4905 14433 4939 14467
rect 10057 14433 10091 14467
rect 11437 14433 11471 14467
rect 14105 14433 14139 14467
rect 15301 14433 15335 14467
rect 18613 14433 18647 14467
rect 1777 14365 1811 14399
rect 4997 14365 5031 14399
rect 7113 14365 7147 14399
rect 8677 14365 8711 14399
rect 10149 14365 10183 14399
rect 10241 14365 10275 14399
rect 11897 14365 11931 14399
rect 15485 14365 15519 14399
rect 17325 14365 17359 14399
rect 18889 14365 18923 14399
rect 19809 14365 19843 14399
rect 3157 14297 3191 14331
rect 13277 14297 13311 14331
rect 4445 14229 4479 14263
rect 9689 14229 9723 14263
rect 10609 14229 10643 14263
rect 11253 14229 11287 14263
rect 16681 14229 16715 14263
rect 9689 14025 9723 14059
rect 11437 14025 11471 14059
rect 17049 14025 17083 14059
rect 20821 14025 20855 14059
rect 5457 13957 5491 13991
rect 8861 13957 8895 13991
rect 4169 13889 4203 13923
rect 4353 13889 4387 13923
rect 10241 13889 10275 13923
rect 13553 13889 13587 13923
rect 13737 13889 13771 13923
rect 14657 13889 14691 13923
rect 1501 13821 1535 13855
rect 1768 13821 1802 13855
rect 5273 13821 5307 13855
rect 7481 13821 7515 13855
rect 11253 13821 11287 13855
rect 14924 13821 14958 13855
rect 16865 13821 16899 13855
rect 18061 13821 18095 13855
rect 19441 13821 19475 13855
rect 19697 13821 19731 13855
rect 4077 13753 4111 13787
rect 7748 13753 7782 13787
rect 10149 13753 10183 13787
rect 18337 13753 18371 13787
rect 2881 13685 2915 13719
rect 3709 13685 3743 13719
rect 10057 13685 10091 13719
rect 13093 13685 13127 13719
rect 13461 13685 13495 13719
rect 16037 13685 16071 13719
rect 7757 13481 7791 13515
rect 8585 13481 8619 13515
rect 11897 13481 11931 13515
rect 12357 13481 12391 13515
rect 18153 13481 18187 13515
rect 18981 13481 19015 13515
rect 19349 13481 19383 13515
rect 2329 13413 2363 13447
rect 4445 13413 4479 13447
rect 6622 13413 6656 13447
rect 9934 13413 9968 13447
rect 14105 13413 14139 13447
rect 15577 13413 15611 13447
rect 2053 13345 2087 13379
rect 4537 13345 4571 13379
rect 6009 13345 6043 13379
rect 12265 13345 12299 13379
rect 14013 13345 14047 13379
rect 15301 13345 15335 13379
rect 16773 13345 16807 13379
rect 17040 13345 17074 13379
rect 4721 13277 4755 13311
rect 6377 13277 6411 13311
rect 9689 13277 9723 13311
rect 12541 13277 12575 13311
rect 14289 13277 14323 13311
rect 19441 13277 19475 13311
rect 19625 13277 19659 13311
rect 5825 13209 5859 13243
rect 4077 13141 4111 13175
rect 11069 13141 11103 13175
rect 13645 13141 13679 13175
rect 2789 12937 2823 12971
rect 4353 12937 4387 12971
rect 6469 12937 6503 12971
rect 6837 12937 6871 12971
rect 9965 12937 9999 12971
rect 11529 12937 11563 12971
rect 3249 12801 3283 12835
rect 3341 12801 3375 12835
rect 4905 12801 4939 12835
rect 7297 12801 7331 12835
rect 7481 12801 7515 12835
rect 8953 12801 8987 12835
rect 13829 12869 13863 12903
rect 16037 12869 16071 12903
rect 17049 12869 17083 12903
rect 18061 12869 18095 12903
rect 10149 12801 10183 12835
rect 18613 12801 18647 12835
rect 20177 12801 20211 12835
rect 1691 12733 1725 12767
rect 3157 12733 3191 12767
rect 6653 12733 6687 12767
rect 8769 12733 8803 12767
rect 9965 12733 9999 12767
rect 10405 12733 10439 12767
rect 12449 12733 12483 12767
rect 12705 12733 12739 12767
rect 14657 12733 14691 12767
rect 16865 12733 16899 12767
rect 18521 12733 18555 12767
rect 20085 12733 20119 12767
rect 7205 12665 7239 12699
rect 14902 12665 14936 12699
rect 18429 12665 18463 12699
rect 1869 12597 1903 12631
rect 4721 12597 4755 12631
rect 4813 12597 4847 12631
rect 8401 12597 8435 12631
rect 8861 12597 8895 12631
rect 19625 12597 19659 12631
rect 19993 12597 20027 12631
rect 2605 12393 2639 12427
rect 6377 12393 6411 12427
rect 8309 12393 8343 12427
rect 11713 12393 11747 12427
rect 12909 12393 12943 12427
rect 15301 12393 15335 12427
rect 19717 12393 19751 12427
rect 2513 12257 2547 12291
rect 4169 12257 4203 12291
rect 4436 12257 4470 12291
rect 6745 12257 6779 12291
rect 8401 12257 8435 12291
rect 10057 12257 10091 12291
rect 11621 12257 11655 12291
rect 2697 12189 2731 12223
rect 6837 12189 6871 12223
rect 6929 12189 6963 12223
rect 8493 12189 8527 12223
rect 10149 12189 10183 12223
rect 10333 12189 10367 12223
rect 11805 12189 11839 12223
rect 13268 12325 13302 12359
rect 17316 12325 17350 12359
rect 19625 12325 19659 12359
rect 15669 12257 15703 12291
rect 17049 12257 17083 12291
rect 13001 12189 13035 12223
rect 15761 12189 15795 12223
rect 15945 12189 15979 12223
rect 19809 12189 19843 12223
rect 2145 12053 2179 12087
rect 5549 12053 5583 12087
rect 7941 12053 7975 12087
rect 9689 12053 9723 12087
rect 11253 12053 11287 12087
rect 12909 12053 12943 12087
rect 14381 12053 14415 12087
rect 18429 12053 18463 12087
rect 19257 12053 19291 12087
rect 3801 11849 3835 11883
rect 7021 11849 7055 11883
rect 8585 11849 8619 11883
rect 12449 11849 12483 11883
rect 14013 11849 14047 11883
rect 1409 11713 1443 11747
rect 5181 11713 5215 11747
rect 7481 11713 7515 11747
rect 7665 11713 7699 11747
rect 9229 11713 9263 11747
rect 11713 11713 11747 11747
rect 13001 11713 13035 11747
rect 15577 11713 15611 11747
rect 18705 11713 18739 11747
rect 20177 11713 20211 11747
rect 2421 11645 2455 11679
rect 9045 11645 9079 11679
rect 9689 11645 9723 11679
rect 9956 11645 9990 11679
rect 11621 11645 11655 11679
rect 12909 11645 12943 11679
rect 14197 11645 14231 11679
rect 16497 11645 16531 11679
rect 18521 11645 18555 11679
rect 19993 11645 20027 11679
rect 2688 11577 2722 11611
rect 4997 11577 5031 11611
rect 7389 11577 7423 11611
rect 11529 11577 11563 11611
rect 15301 11577 15335 11611
rect 16773 11577 16807 11611
rect 20085 11577 20119 11611
rect 4629 11509 4663 11543
rect 5089 11509 5123 11543
rect 8953 11509 8987 11543
rect 11069 11509 11103 11543
rect 11161 11509 11195 11543
rect 12817 11509 12851 11543
rect 14933 11509 14967 11543
rect 15393 11509 15427 11543
rect 18061 11509 18095 11543
rect 18429 11509 18463 11543
rect 19625 11509 19659 11543
rect 2421 11305 2455 11339
rect 2881 11305 2915 11339
rect 5917 11305 5951 11339
rect 12725 11305 12759 11339
rect 13645 11305 13679 11339
rect 14105 11305 14139 11339
rect 18153 11305 18187 11339
rect 18981 11305 19015 11339
rect 19349 11305 19383 11339
rect 4804 11237 4838 11271
rect 7656 11237 7690 11271
rect 12633 11237 12667 11271
rect 14013 11237 14047 11271
rect 15577 11237 15611 11271
rect 2789 11169 2823 11203
rect 7389 11169 7423 11203
rect 10425 11169 10459 11203
rect 15301 11169 15335 11203
rect 16773 11169 16807 11203
rect 17040 11169 17074 11203
rect 1409 11101 1443 11135
rect 3065 11101 3099 11135
rect 4537 11101 4571 11135
rect 12817 11101 12851 11135
rect 14289 11101 14323 11135
rect 19441 11101 19475 11135
rect 19533 11101 19567 11135
rect 8769 11033 8803 11067
rect 12265 11033 12299 11067
rect 11713 10965 11747 10999
rect 9045 10761 9079 10795
rect 10977 10761 11011 10795
rect 15853 10761 15887 10795
rect 18061 10761 18095 10795
rect 19625 10761 19659 10795
rect 3433 10693 3467 10727
rect 12081 10693 12115 10727
rect 4813 10625 4847 10659
rect 13001 10625 13035 10659
rect 18613 10625 18647 10659
rect 20177 10625 20211 10659
rect 2053 10557 2087 10591
rect 2320 10557 2354 10591
rect 4629 10557 4663 10591
rect 6837 10557 6871 10591
rect 9229 10557 9263 10591
rect 9597 10557 9631 10591
rect 12265 10557 12299 10591
rect 14473 10557 14507 10591
rect 16681 10557 16715 10591
rect 19441 10557 19475 10591
rect 19993 10557 20027 10591
rect 20085 10557 20119 10591
rect 20453 10557 20487 10591
rect 4721 10489 4755 10523
rect 7104 10489 7138 10523
rect 9864 10489 9898 10523
rect 12909 10489 12943 10523
rect 14740 10489 14774 10523
rect 16957 10489 16991 10523
rect 18429 10489 18463 10523
rect 4261 10421 4295 10455
rect 8217 10421 8251 10455
rect 12449 10421 12483 10455
rect 12817 10421 12851 10455
rect 18521 10421 18555 10455
rect 18889 10421 18923 10455
rect 7941 10217 7975 10251
rect 15301 10217 15335 10251
rect 15761 10217 15795 10251
rect 18429 10217 18463 10251
rect 18797 10217 18831 10251
rect 1768 10149 1802 10183
rect 4353 10149 4387 10183
rect 8033 10149 8067 10183
rect 10508 10149 10542 10183
rect 15669 10149 15703 10183
rect 18889 10149 18923 10183
rect 1501 10081 1535 10115
rect 4077 10081 4111 10115
rect 5632 10081 5666 10115
rect 12705 10081 12739 10115
rect 17233 10081 17267 10115
rect 5365 10013 5399 10047
rect 8125 10013 8159 10047
rect 10241 10013 10275 10047
rect 12449 10013 12483 10047
rect 15945 10013 15979 10047
rect 17325 10013 17359 10047
rect 17417 10013 17451 10047
rect 18981 10013 19015 10047
rect 6745 9945 6779 9979
rect 11621 9945 11655 9979
rect 2881 9877 2915 9911
rect 7573 9877 7607 9911
rect 13829 9877 13863 9911
rect 16865 9877 16899 9911
rect 1961 9673 1995 9707
rect 16129 9673 16163 9707
rect 7021 9605 7055 9639
rect 12541 9605 12575 9639
rect 2789 9537 2823 9571
rect 4261 9537 4295 9571
rect 5457 9537 5491 9571
rect 8585 9537 8619 9571
rect 10333 9537 10367 9571
rect 10517 9537 10551 9571
rect 13185 9537 13219 9571
rect 14749 9537 14783 9571
rect 16957 9537 16991 9571
rect 1409 9469 1443 9503
rect 1777 9469 1811 9503
rect 2513 9469 2547 9503
rect 5304 9469 5338 9503
rect 6837 9469 6871 9503
rect 8309 9469 8343 9503
rect 9689 9469 9723 9503
rect 14289 9469 14323 9503
rect 18061 9469 18095 9503
rect 20269 9469 20303 9503
rect 4169 9401 4203 9435
rect 8401 9401 8435 9435
rect 12909 9401 12943 9435
rect 15016 9401 15050 9435
rect 18306 9401 18340 9435
rect 1593 9333 1627 9367
rect 2145 9333 2179 9367
rect 2605 9333 2639 9367
rect 3709 9333 3743 9367
rect 4077 9333 4111 9367
rect 7941 9333 7975 9367
rect 9505 9333 9539 9367
rect 9873 9333 9907 9367
rect 10241 9333 10275 9367
rect 13001 9333 13035 9367
rect 14105 9333 14139 9367
rect 19441 9333 19475 9367
rect 1409 9129 1443 9163
rect 3249 9129 3283 9163
rect 4445 9129 4479 9163
rect 5457 9129 5491 9163
rect 5825 9129 5859 9163
rect 9873 9129 9907 9163
rect 12357 9129 12391 9163
rect 12817 9129 12851 9163
rect 13921 9129 13955 9163
rect 14197 9129 14231 9163
rect 18889 9129 18923 9163
rect 2881 9061 2915 9095
rect 7481 9061 7515 9095
rect 8585 9061 8619 9095
rect 1777 8993 1811 9027
rect 1869 8993 1903 9027
rect 2789 8993 2823 9027
rect 4905 8993 4939 9027
rect 7389 8993 7423 9027
rect 10241 8993 10275 9027
rect 10333 8993 10367 9027
rect 11897 8993 11931 9027
rect 12725 8993 12759 9027
rect 14097 8993 14131 9027
rect 15669 8993 15703 9027
rect 17417 8993 17451 9027
rect 18797 8993 18831 9027
rect 2053 8925 2087 8959
rect 3065 8925 3099 8959
rect 4537 8925 4571 8959
rect 4721 8925 4755 8959
rect 5089 8925 5123 8959
rect 5917 8925 5951 8959
rect 6009 8925 6043 8959
rect 7573 8925 7607 8959
rect 10517 8925 10551 8959
rect 12909 8925 12943 8959
rect 15761 8925 15795 8959
rect 15945 8925 15979 8959
rect 18981 8925 19015 8959
rect 4077 8857 4111 8891
rect 7021 8857 7055 8891
rect 15301 8857 15335 8891
rect 2421 8789 2455 8823
rect 11713 8789 11747 8823
rect 18429 8789 18463 8823
rect 5089 8585 5123 8619
rect 5733 8585 5767 8619
rect 14013 8585 14047 8619
rect 15485 8585 15519 8619
rect 19441 8585 19475 8619
rect 2881 8517 2915 8551
rect 5457 8517 5491 8551
rect 7573 8517 7607 8551
rect 16405 8517 16439 8551
rect 3157 8449 3191 8483
rect 6377 8449 6411 8483
rect 8033 8449 8067 8483
rect 8217 8449 8251 8483
rect 9137 8449 9171 8483
rect 9229 8449 9263 8483
rect 10241 8449 10275 8483
rect 14013 8449 14047 8483
rect 14105 8449 14139 8483
rect 16957 8449 16991 8483
rect 1501 8381 1535 8415
rect 1768 8381 1802 8415
rect 2973 8381 3007 8415
rect 3709 8381 3743 8415
rect 5641 8381 5675 8415
rect 6101 8381 6135 8415
rect 7941 8381 7975 8415
rect 3976 8313 4010 8347
rect 12909 8381 12943 8415
rect 16773 8381 16807 8415
rect 18061 8381 18095 8415
rect 11345 8313 11379 8347
rect 14350 8313 14384 8347
rect 16865 8313 16899 8347
rect 18306 8313 18340 8347
rect 20269 8313 20303 8347
rect 6193 8245 6227 8279
rect 9137 8245 9171 8279
rect 2421 8041 2455 8075
rect 2881 8041 2915 8075
rect 4537 8041 4571 8075
rect 4905 8041 4939 8075
rect 6653 8041 6687 8075
rect 7205 8041 7239 8075
rect 11069 8041 11103 8075
rect 11989 8041 12023 8075
rect 12541 8041 12575 8075
rect 13645 8041 13679 8075
rect 15761 8041 15795 8075
rect 2789 7973 2823 8007
rect 1777 7905 1811 7939
rect 4445 7905 4479 7939
rect 1869 7837 1903 7871
rect 2053 7837 2087 7871
rect 2973 7837 3007 7871
rect 4721 7837 4755 7871
rect 5253 7905 5287 7939
rect 6469 7905 6503 7939
rect 7573 7905 7607 7939
rect 7665 7905 7699 7939
rect 8953 7905 8987 7939
rect 9689 7905 9723 7939
rect 9956 7905 9990 7939
rect 4997 7837 5031 7871
rect 7757 7837 7791 7871
rect 14013 7973 14047 8007
rect 12449 7905 12483 7939
rect 15669 7905 15703 7939
rect 17509 7905 17543 7939
rect 17776 7905 17810 7939
rect 19717 7905 19751 7939
rect 12725 7837 12759 7871
rect 14105 7837 14139 7871
rect 14289 7837 14323 7871
rect 15853 7837 15887 7871
rect 2329 7769 2363 7803
rect 4905 7769 4939 7803
rect 8769 7769 8803 7803
rect 11989 7769 12023 7803
rect 12081 7769 12115 7803
rect 1409 7701 1443 7735
rect 4077 7701 4111 7735
rect 6377 7701 6411 7735
rect 15301 7701 15335 7735
rect 18889 7701 18923 7735
rect 19901 7701 19935 7735
rect 2237 7497 2271 7531
rect 4077 7497 4111 7531
rect 5733 7497 5767 7531
rect 19441 7497 19475 7531
rect 8217 7429 8251 7463
rect 11529 7429 11563 7463
rect 15025 7429 15059 7463
rect 19625 7429 19659 7463
rect 2053 7361 2087 7395
rect 2697 7361 2731 7395
rect 2881 7361 2915 7395
rect 4629 7361 4663 7395
rect 5457 7361 5491 7395
rect 6193 7361 6227 7395
rect 6377 7361 6411 7395
rect 9045 7361 9079 7395
rect 10057 7361 10091 7395
rect 15669 7361 15703 7395
rect 18613 7361 18647 7395
rect 20085 7361 20119 7395
rect 20177 7361 20211 7395
rect 1777 7293 1811 7327
rect 3801 7293 3835 7327
rect 3985 7293 4019 7327
rect 4445 7293 4479 7327
rect 6837 7293 6871 7327
rect 7104 7293 7138 7327
rect 4537 7225 4571 7259
rect 5273 7225 5307 7259
rect 5365 7225 5399 7259
rect 6101 7225 6135 7259
rect 10149 7293 10183 7327
rect 10416 7293 10450 7327
rect 12449 7293 12483 7327
rect 15393 7293 15427 7327
rect 16589 7293 16623 7327
rect 18337 7293 18371 7327
rect 19993 7293 20027 7327
rect 12694 7225 12728 7259
rect 16865 7225 16899 7259
rect 1409 7157 1443 7191
rect 1869 7157 1903 7191
rect 2605 7157 2639 7191
rect 3801 7157 3835 7191
rect 4905 7157 4939 7191
rect 10057 7157 10091 7191
rect 13829 7157 13863 7191
rect 15485 7157 15519 7191
rect 3341 6953 3375 6987
rect 4445 6953 4479 6987
rect 5273 6953 5307 6987
rect 5365 6953 5399 6987
rect 5733 6953 5767 6987
rect 6101 6953 6135 6987
rect 12081 6953 12115 6987
rect 3249 6885 3283 6919
rect 7665 6885 7699 6919
rect 7757 6885 7791 6919
rect 11989 6885 12023 6919
rect 16466 6885 16500 6919
rect 1676 6817 1710 6851
rect 6193 6817 6227 6851
rect 10425 6817 10459 6851
rect 14013 6817 14047 6851
rect 14105 6817 14139 6851
rect 16221 6817 16255 6851
rect 18685 6817 18719 6851
rect 1409 6749 1443 6783
rect 3525 6749 3559 6783
rect 4537 6749 4571 6783
rect 4721 6749 4755 6783
rect 5457 6749 5491 6783
rect 6285 6749 6319 6783
rect 6561 6749 6595 6783
rect 7849 6749 7883 6783
rect 10517 6749 10551 6783
rect 10701 6749 10735 6783
rect 12265 6749 12299 6783
rect 14197 6749 14231 6783
rect 18429 6749 18463 6783
rect 4905 6681 4939 6715
rect 10057 6681 10091 6715
rect 2789 6613 2823 6647
rect 2881 6613 2915 6647
rect 4077 6613 4111 6647
rect 7297 6613 7331 6647
rect 11621 6613 11655 6647
rect 13645 6613 13679 6647
rect 17601 6613 17635 6647
rect 19809 6613 19843 6647
rect 1961 6409 1995 6443
rect 3433 6409 3467 6443
rect 5917 6409 5951 6443
rect 6193 6409 6227 6443
rect 6561 6409 6595 6443
rect 8309 6409 8343 6443
rect 8401 6409 8435 6443
rect 9413 6409 9447 6443
rect 10149 6409 10183 6443
rect 14657 6409 14691 6443
rect 19625 6409 19659 6443
rect 4169 6273 4203 6307
rect 4537 6273 4571 6307
rect 6929 6273 6963 6307
rect 8861 6273 8895 6307
rect 9045 6273 9079 6307
rect 1409 6205 1443 6239
rect 1961 6205 1995 6239
rect 2053 6205 2087 6239
rect 6009 6205 6043 6239
rect 6377 6205 6411 6239
rect 8769 6205 8803 6239
rect 9229 6205 9263 6239
rect 1685 6137 1719 6171
rect 2320 6137 2354 6171
rect 3985 6137 4019 6171
rect 4804 6137 4838 6171
rect 7196 6137 7230 6171
rect 10241 6341 10275 6375
rect 10885 6273 10919 6307
rect 12449 6273 12483 6307
rect 15301 6273 15335 6307
rect 16865 6273 16899 6307
rect 18613 6273 18647 6307
rect 20177 6273 20211 6307
rect 10701 6205 10735 6239
rect 12716 6205 12750 6239
rect 15025 6205 15059 6239
rect 16589 6205 16623 6239
rect 16681 6205 16715 6239
rect 18429 6205 18463 6239
rect 18521 6205 18555 6239
rect 19993 6205 20027 6239
rect 3525 6069 3559 6103
rect 3893 6069 3927 6103
rect 10149 6069 10183 6103
rect 10609 6069 10643 6103
rect 13829 6069 13863 6103
rect 15117 6069 15151 6103
rect 16221 6069 16255 6103
rect 18061 6069 18095 6103
rect 20085 6069 20119 6103
rect 2881 5865 2915 5899
rect 5733 5865 5767 5899
rect 6193 5865 6227 5899
rect 7021 5865 7055 5899
rect 7481 5865 7515 5899
rect 8953 5865 8987 5899
rect 13921 5865 13955 5899
rect 1676 5797 1710 5831
rect 12265 5797 12299 5831
rect 3249 5729 3283 5763
rect 4261 5729 4295 5763
rect 4528 5729 4562 5763
rect 6101 5729 6135 5763
rect 6929 5729 6963 5763
rect 7849 5729 7883 5763
rect 9956 5729 9990 5763
rect 13829 5729 13863 5763
rect 15853 5729 15887 5763
rect 16120 5729 16154 5763
rect 18337 5729 18371 5763
rect 18604 5729 18638 5763
rect 3341 5661 3375 5695
rect 3525 5661 3559 5695
rect 6377 5661 6411 5695
rect 7205 5661 7239 5695
rect 7941 5661 7975 5695
rect 8125 5661 8159 5695
rect 9045 5661 9079 5695
rect 9229 5661 9263 5695
rect 9413 5661 9447 5695
rect 9689 5661 9723 5695
rect 12357 5661 12391 5695
rect 12449 5661 12483 5695
rect 14013 5661 14047 5695
rect 2789 5593 2823 5627
rect 6561 5593 6595 5627
rect 8585 5593 8619 5627
rect 11069 5593 11103 5627
rect 19717 5593 19751 5627
rect 5641 5525 5675 5559
rect 9413 5525 9447 5559
rect 11897 5525 11931 5559
rect 13461 5525 13495 5559
rect 17233 5525 17267 5559
rect 7757 5321 7791 5355
rect 4261 5253 4295 5287
rect 8677 5253 8711 5287
rect 16037 5253 16071 5287
rect 17049 5253 17083 5287
rect 6377 5185 6411 5219
rect 7297 5185 7331 5219
rect 7481 5185 7515 5219
rect 7665 5185 7699 5219
rect 8401 5185 8435 5219
rect 9137 5185 9171 5219
rect 9321 5185 9355 5219
rect 10333 5185 10367 5219
rect 10425 5185 10459 5219
rect 12449 5185 12483 5219
rect 18613 5185 18647 5219
rect 20177 5185 20211 5219
rect 2881 5117 2915 5151
rect 3137 5117 3171 5151
rect 4353 5117 4387 5151
rect 4620 5117 4654 5151
rect 6193 5117 6227 5151
rect 8125 5117 8159 5151
rect 8217 5117 8251 5151
rect 9045 5117 9079 5151
rect 10241 5117 10275 5151
rect 12705 5117 12739 5151
rect 14657 5117 14691 5151
rect 16865 5117 16899 5151
rect 18429 5117 18463 5151
rect 18521 5117 18555 5151
rect 1676 5049 1710 5083
rect 7205 5049 7239 5083
rect 7665 5049 7699 5083
rect 14902 5049 14936 5083
rect 20085 5049 20119 5083
rect 2789 4981 2823 5015
rect 5733 4981 5767 5015
rect 5825 4981 5859 5015
rect 6285 4981 6319 5015
rect 6837 4981 6871 5015
rect 9873 4981 9907 5015
rect 13829 4981 13863 5015
rect 18061 4981 18095 5015
rect 19625 4981 19659 5015
rect 19993 4981 20027 5015
rect 3341 4777 3375 4811
rect 5457 4777 5491 4811
rect 6745 4777 6779 4811
rect 8309 4777 8343 4811
rect 8677 4777 8711 4811
rect 9965 4777 9999 4811
rect 10333 4777 10367 4811
rect 13185 4777 13219 4811
rect 3249 4709 3283 4743
rect 7757 4709 7791 4743
rect 8217 4709 8251 4743
rect 9045 4709 9079 4743
rect 10425 4709 10459 4743
rect 11069 4709 11103 4743
rect 11989 4709 12023 4743
rect 13645 4709 13679 4743
rect 16221 4709 16255 4743
rect 17662 4709 17696 4743
rect 1676 4641 1710 4675
rect 4077 4641 4111 4675
rect 4344 4641 4378 4675
rect 5917 4641 5951 4675
rect 6009 4641 6043 4675
rect 7205 4641 7239 4675
rect 10793 4641 10827 4675
rect 13553 4641 13587 4675
rect 19717 4641 19751 4675
rect 3525 4573 3559 4607
rect 6101 4573 6135 4607
rect 6837 4573 6871 4607
rect 6929 4573 6963 4607
rect 7481 4573 7515 4607
rect 7757 4573 7791 4607
rect 8493 4573 8527 4607
rect 9137 4573 9171 4607
rect 9321 4573 9355 4607
rect 10609 4573 10643 4607
rect 12081 4573 12115 4607
rect 12265 4573 12299 4607
rect 13737 4573 13771 4607
rect 16313 4573 16347 4607
rect 16497 4573 16531 4607
rect 17417 4573 17451 4607
rect 2789 4505 2823 4539
rect 15853 4505 15887 4539
rect 2881 4437 2915 4471
rect 5549 4437 5583 4471
rect 6377 4437 6411 4471
rect 7849 4437 7883 4471
rect 11621 4437 11655 4471
rect 18797 4437 18831 4471
rect 19901 4437 19935 4471
rect 5733 4233 5767 4267
rect 15853 4233 15887 4267
rect 9137 4165 9171 4199
rect 9781 4165 9815 4199
rect 6377 4097 6411 4131
rect 7297 4097 7331 4131
rect 7481 4097 7515 4131
rect 7757 4097 7791 4131
rect 10517 4097 10551 4131
rect 11345 4097 11379 4131
rect 14473 4097 14507 4131
rect 18521 4097 18555 4131
rect 18705 4097 18739 4131
rect 20085 4097 20119 4131
rect 20177 4097 20211 4131
rect 1665 4029 1699 4063
rect 3137 4029 3171 4063
rect 4353 4029 4387 4063
rect 4620 4029 4654 4063
rect 8013 4029 8047 4063
rect 9229 4029 9263 4063
rect 9781 4029 9815 4063
rect 11652 4029 11686 4063
rect 11897 4029 11931 4063
rect 12541 4029 12575 4063
rect 14740 4029 14774 4063
rect 16681 4029 16715 4063
rect 19993 4029 20027 4063
rect 6285 3961 6319 3995
rect 7205 3961 7239 3995
rect 9505 3961 9539 3995
rect 10425 3961 10459 3995
rect 11253 3961 11287 3995
rect 2789 3893 2823 3927
rect 4261 3893 4295 3927
rect 5825 3893 5859 3927
rect 6193 3893 6227 3927
rect 6837 3893 6871 3927
rect 9965 3893 9999 3927
rect 10333 3893 10367 3927
rect 10793 3893 10827 3927
rect 11161 3893 11195 3927
rect 12725 3893 12759 3927
rect 16865 3893 16899 3927
rect 18061 3893 18095 3927
rect 18429 3893 18463 3927
rect 19625 3893 19659 3927
rect 7205 3689 7239 3723
rect 7481 3689 7515 3723
rect 7665 3689 7699 3723
rect 8125 3689 8159 3723
rect 9229 3689 9263 3723
rect 9321 3689 9355 3723
rect 10057 3689 10091 3723
rect 11713 3689 11747 3723
rect 17601 3689 17635 3723
rect 1654 3621 1688 3655
rect 4344 3621 4378 3655
rect 6092 3621 6126 3655
rect 10885 3621 10919 3655
rect 11805 3621 11839 3655
rect 17969 3621 18003 3655
rect 1409 3553 1443 3587
rect 3249 3553 3283 3587
rect 8033 3553 8067 3587
rect 12173 3553 12207 3587
rect 12541 3553 12575 3587
rect 12817 3553 12851 3587
rect 14105 3553 14139 3587
rect 15301 3553 15335 3587
rect 16497 3553 16531 3587
rect 19625 3553 19659 3587
rect 3341 3485 3375 3519
rect 3433 3485 3467 3519
rect 5825 3485 5859 3519
rect 8217 3485 8251 3519
rect 10149 3485 10183 3519
rect 10333 3485 10367 3519
rect 10977 3485 11011 3519
rect 11069 3485 11103 3519
rect 11897 3485 11931 3519
rect 18061 3485 18095 3519
rect 18153 3485 18187 3519
rect 2789 3417 2823 3451
rect 9689 3417 9723 3451
rect 11345 3417 11379 3451
rect 2881 3349 2915 3383
rect 5457 3349 5491 3383
rect 10517 3349 10551 3383
rect 12357 3349 12391 3383
rect 14289 3349 14323 3383
rect 15485 3349 15519 3383
rect 16681 3349 16715 3383
rect 19809 3349 19843 3383
rect 5917 3145 5951 3179
rect 8125 3145 8159 3179
rect 11345 3145 11379 3179
rect 12449 3145 12483 3179
rect 2789 3077 2823 3111
rect 4261 3077 4295 3111
rect 7113 3077 7147 3111
rect 19349 3077 19383 3111
rect 7665 3009 7699 3043
rect 11115 3009 11149 3043
rect 11897 3009 11931 3043
rect 13093 3009 13127 3043
rect 14565 3009 14599 3043
rect 20453 3009 20487 3043
rect 1676 2941 1710 2975
rect 3148 2941 3182 2975
rect 4537 2941 4571 2975
rect 6193 2941 6227 2975
rect 7573 2941 7607 2975
rect 7941 2941 7975 2975
rect 8309 2941 8343 2975
rect 9781 2941 9815 2975
rect 14381 2941 14415 2975
rect 15577 2941 15611 2975
rect 16681 2941 16715 2975
rect 18049 2941 18083 2975
rect 19165 2941 19199 2975
rect 20269 2941 20303 2975
rect 4782 2873 4816 2907
rect 6469 2873 6503 2907
rect 8576 2873 8610 2907
rect 10057 2873 10091 2907
rect 11713 2873 11747 2907
rect 11805 2873 11839 2907
rect 12817 2873 12851 2907
rect 7481 2805 7515 2839
rect 9689 2805 9723 2839
rect 10517 2805 10551 2839
rect 10885 2805 10919 2839
rect 10977 2805 11011 2839
rect 12909 2805 12943 2839
rect 14013 2805 14047 2839
rect 14473 2805 14507 2839
rect 15761 2805 15795 2839
rect 16865 2805 16899 2839
rect 18245 2805 18279 2839
rect 5457 2601 5491 2635
rect 5549 2601 5583 2635
rect 5917 2601 5951 2635
rect 6009 2601 6043 2635
rect 8861 2601 8895 2635
rect 9413 2601 9447 2635
rect 10609 2601 10643 2635
rect 11069 2601 11103 2635
rect 11437 2601 11471 2635
rect 12633 2601 12667 2635
rect 13001 2601 13035 2635
rect 15945 2601 15979 2635
rect 20177 2601 20211 2635
rect 1676 2533 1710 2567
rect 4344 2533 4378 2567
rect 8769 2533 8803 2567
rect 13093 2533 13127 2567
rect 15853 2533 15887 2567
rect 1409 2465 1443 2499
rect 3249 2465 3283 2499
rect 6377 2465 6411 2499
rect 7196 2465 7230 2499
rect 9229 2465 9263 2499
rect 10149 2465 10183 2499
rect 10241 2465 10275 2499
rect 10977 2465 11011 2499
rect 11805 2465 11839 2499
rect 11897 2465 11931 2499
rect 14197 2465 14231 2499
rect 17049 2465 17083 2499
rect 18889 2465 18923 2499
rect 19993 2465 20027 2499
rect 3341 2397 3375 2431
rect 3433 2397 3467 2431
rect 3709 2397 3743 2431
rect 6101 2397 6135 2431
rect 8953 2397 8987 2431
rect 10333 2397 10367 2431
rect 11161 2397 11195 2431
rect 11989 2397 12023 2431
rect 13185 2397 13219 2431
rect 16037 2397 16071 2431
rect 8401 2329 8435 2363
rect 15485 2329 15519 2363
rect 2789 2261 2823 2295
rect 2881 2261 2915 2295
rect 6561 2261 6595 2295
rect 8309 2261 8343 2295
rect 9781 2261 9815 2295
rect 14381 2261 14415 2295
rect 17233 2261 17267 2295
rect 19073 2261 19107 2295
rect 8125 1717 8159 1751
rect 8125 1377 8159 1411
rect 10425 1649 10459 1683
rect 10425 1377 10459 1411
<< metal1 >>
rect 7006 20748 7012 20800
rect 7064 20788 7070 20800
rect 8110 20788 8116 20800
rect 7064 20760 8116 20788
rect 7064 20748 7070 20760
rect 8110 20748 8116 20760
rect 8168 20748 8174 20800
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 4154 20544 4160 20596
rect 4212 20584 4218 20596
rect 4249 20587 4307 20593
rect 4249 20584 4261 20587
rect 4212 20556 4261 20584
rect 4212 20544 4218 20556
rect 4249 20553 4261 20556
rect 4295 20553 4307 20587
rect 4249 20547 4307 20553
rect 5261 20587 5319 20593
rect 5261 20553 5273 20587
rect 5307 20584 5319 20587
rect 12526 20584 12532 20596
rect 5307 20556 12532 20584
rect 5307 20553 5319 20556
rect 5261 20547 5319 20553
rect 12526 20544 12532 20556
rect 12584 20544 12590 20596
rect 12621 20587 12679 20593
rect 12621 20553 12633 20587
rect 12667 20584 12679 20587
rect 14090 20584 14096 20596
rect 12667 20556 14096 20584
rect 12667 20553 12679 20556
rect 12621 20547 12679 20553
rect 14090 20544 14096 20556
rect 14148 20544 14154 20596
rect 15194 20544 15200 20596
rect 15252 20584 15258 20596
rect 15749 20587 15807 20593
rect 15749 20584 15761 20587
rect 15252 20556 15761 20584
rect 15252 20544 15258 20556
rect 15749 20553 15761 20556
rect 15795 20553 15807 20587
rect 15749 20547 15807 20553
rect 18785 20587 18843 20593
rect 18785 20553 18797 20587
rect 18831 20584 18843 20587
rect 19426 20584 19432 20596
rect 18831 20556 19432 20584
rect 18831 20553 18843 20556
rect 18785 20547 18843 20553
rect 19426 20544 19432 20556
rect 19484 20544 19490 20596
rect 20165 20587 20223 20593
rect 20165 20553 20177 20587
rect 20211 20584 20223 20587
rect 21266 20584 21272 20596
rect 20211 20556 21272 20584
rect 20211 20553 20223 20556
rect 20165 20547 20223 20553
rect 21266 20544 21272 20556
rect 21324 20544 21330 20596
rect 6917 20519 6975 20525
rect 6917 20485 6929 20519
rect 6963 20516 6975 20519
rect 9674 20516 9680 20528
rect 6963 20488 9680 20516
rect 6963 20485 6975 20488
rect 6917 20479 6975 20485
rect 9674 20476 9680 20488
rect 9732 20476 9738 20528
rect 9769 20519 9827 20525
rect 9769 20485 9781 20519
rect 9815 20516 9827 20519
rect 9815 20488 11100 20516
rect 9815 20485 9827 20488
rect 9769 20479 9827 20485
rect 5718 20408 5724 20460
rect 5776 20448 5782 20460
rect 5813 20451 5871 20457
rect 5813 20448 5825 20451
rect 5776 20420 5825 20448
rect 5776 20408 5782 20420
rect 5813 20417 5825 20420
rect 5859 20417 5871 20451
rect 5813 20411 5871 20417
rect 7098 20408 7104 20460
rect 7156 20448 7162 20460
rect 7469 20451 7527 20457
rect 7469 20448 7481 20451
rect 7156 20420 7481 20448
rect 7156 20408 7162 20420
rect 7469 20417 7481 20420
rect 7515 20417 7527 20451
rect 7469 20411 7527 20417
rect 8312 20420 10272 20448
rect 1765 20383 1823 20389
rect 1765 20349 1777 20383
rect 1811 20380 1823 20383
rect 3970 20380 3976 20392
rect 1811 20352 3976 20380
rect 1811 20349 1823 20352
rect 1765 20343 1823 20349
rect 3970 20340 3976 20352
rect 4028 20340 4034 20392
rect 4065 20383 4123 20389
rect 4065 20349 4077 20383
rect 4111 20380 4123 20383
rect 4154 20380 4160 20392
rect 4111 20352 4160 20380
rect 4111 20349 4123 20352
rect 4065 20343 4123 20349
rect 4154 20340 4160 20352
rect 4212 20340 4218 20392
rect 8312 20380 8340 20420
rect 8478 20380 8484 20392
rect 5736 20352 8340 20380
rect 8439 20352 8484 20380
rect 2032 20315 2090 20321
rect 2032 20281 2044 20315
rect 2078 20312 2090 20315
rect 4614 20312 4620 20324
rect 2078 20284 4620 20312
rect 2078 20281 2090 20284
rect 2032 20275 2090 20281
rect 4614 20272 4620 20284
rect 4672 20272 4678 20324
rect 5736 20321 5764 20352
rect 8478 20340 8484 20352
rect 8536 20340 8542 20392
rect 10244 20380 10272 20420
rect 10318 20408 10324 20460
rect 10376 20448 10382 20460
rect 11072 20448 11100 20488
rect 12894 20448 12900 20460
rect 10376 20420 10421 20448
rect 11072 20420 12900 20448
rect 10376 20408 10382 20420
rect 12894 20408 12900 20420
rect 12952 20408 12958 20460
rect 13173 20451 13231 20457
rect 13173 20417 13185 20451
rect 13219 20417 13231 20451
rect 16853 20451 16911 20457
rect 16853 20448 16865 20451
rect 13173 20411 13231 20417
rect 15580 20420 16865 20448
rect 10410 20380 10416 20392
rect 10244 20352 10416 20380
rect 10410 20340 10416 20352
rect 10468 20340 10474 20392
rect 11330 20380 11336 20392
rect 11291 20352 11336 20380
rect 11330 20340 11336 20352
rect 11388 20340 11394 20392
rect 12986 20340 12992 20392
rect 13044 20380 13050 20392
rect 13188 20380 13216 20411
rect 15580 20389 15608 20420
rect 16853 20417 16865 20420
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 14185 20383 14243 20389
rect 14185 20380 14197 20383
rect 13044 20352 13216 20380
rect 13280 20352 14197 20380
rect 13044 20340 13050 20352
rect 5721 20315 5779 20321
rect 5721 20281 5733 20315
rect 5767 20281 5779 20315
rect 5721 20275 5779 20281
rect 7377 20315 7435 20321
rect 7377 20281 7389 20315
rect 7423 20312 7435 20315
rect 10962 20312 10968 20324
rect 7423 20284 10968 20312
rect 7423 20281 7435 20284
rect 7377 20275 7435 20281
rect 10962 20272 10968 20284
rect 11020 20272 11026 20324
rect 11238 20272 11244 20324
rect 11296 20312 11302 20324
rect 13280 20312 13308 20352
rect 14185 20349 14197 20352
rect 14231 20349 14243 20383
rect 14185 20343 14243 20349
rect 15565 20383 15623 20389
rect 15565 20349 15577 20383
rect 15611 20349 15623 20383
rect 15565 20343 15623 20349
rect 16669 20383 16727 20389
rect 16669 20349 16681 20383
rect 16715 20380 16727 20383
rect 17770 20380 17776 20392
rect 16715 20352 17776 20380
rect 16715 20349 16727 20352
rect 16669 20343 16727 20349
rect 17770 20340 17776 20352
rect 17828 20340 17834 20392
rect 18601 20383 18659 20389
rect 18601 20349 18613 20383
rect 18647 20349 18659 20383
rect 19978 20380 19984 20392
rect 19939 20352 19984 20380
rect 18601 20343 18659 20349
rect 11296 20284 13308 20312
rect 11296 20272 11302 20284
rect 13538 20272 13544 20324
rect 13596 20312 13602 20324
rect 18616 20312 18644 20343
rect 19978 20340 19984 20352
rect 20036 20340 20042 20392
rect 13596 20284 18644 20312
rect 13596 20272 13602 20284
rect 2682 20204 2688 20256
rect 2740 20244 2746 20256
rect 3145 20247 3203 20253
rect 3145 20244 3157 20247
rect 2740 20216 3157 20244
rect 2740 20204 2746 20216
rect 3145 20213 3157 20216
rect 3191 20213 3203 20247
rect 5626 20244 5632 20256
rect 5587 20216 5632 20244
rect 3145 20207 3203 20213
rect 5626 20204 5632 20216
rect 5684 20204 5690 20256
rect 6638 20204 6644 20256
rect 6696 20244 6702 20256
rect 7285 20247 7343 20253
rect 7285 20244 7297 20247
rect 6696 20216 7297 20244
rect 6696 20204 6702 20216
rect 7285 20213 7297 20216
rect 7331 20213 7343 20247
rect 8662 20244 8668 20256
rect 8623 20216 8668 20244
rect 7285 20207 7343 20213
rect 8662 20204 8668 20216
rect 8720 20204 8726 20256
rect 10134 20244 10140 20256
rect 10095 20216 10140 20244
rect 10134 20204 10140 20216
rect 10192 20204 10198 20256
rect 10229 20247 10287 20253
rect 10229 20213 10241 20247
rect 10275 20244 10287 20247
rect 10594 20244 10600 20256
rect 10275 20216 10600 20244
rect 10275 20213 10287 20216
rect 10229 20207 10287 20213
rect 10594 20204 10600 20216
rect 10652 20204 10658 20256
rect 11517 20247 11575 20253
rect 11517 20213 11529 20247
rect 11563 20244 11575 20247
rect 11698 20244 11704 20256
rect 11563 20216 11704 20244
rect 11563 20213 11575 20216
rect 11517 20207 11575 20213
rect 11698 20204 11704 20216
rect 11756 20204 11762 20256
rect 11790 20204 11796 20256
rect 11848 20244 11854 20256
rect 12989 20247 13047 20253
rect 12989 20244 13001 20247
rect 11848 20216 13001 20244
rect 11848 20204 11854 20216
rect 12989 20213 13001 20216
rect 13035 20213 13047 20247
rect 12989 20207 13047 20213
rect 13078 20204 13084 20256
rect 13136 20244 13142 20256
rect 13136 20216 13181 20244
rect 13136 20204 13142 20216
rect 13354 20204 13360 20256
rect 13412 20244 13418 20256
rect 14369 20247 14427 20253
rect 14369 20244 14381 20247
rect 13412 20216 14381 20244
rect 13412 20204 13418 20216
rect 14369 20213 14381 20216
rect 14415 20213 14427 20247
rect 14369 20207 14427 20213
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 1946 20040 1952 20052
rect 1907 20012 1952 20040
rect 1946 20000 1952 20012
rect 2004 20000 2010 20052
rect 3050 20040 3056 20052
rect 3011 20012 3056 20040
rect 3050 20000 3056 20012
rect 3108 20000 3114 20052
rect 3786 20000 3792 20052
rect 3844 20040 3850 20052
rect 7282 20040 7288 20052
rect 3844 20012 7288 20040
rect 3844 20000 3850 20012
rect 7282 20000 7288 20012
rect 7340 20000 7346 20052
rect 7374 20000 7380 20052
rect 7432 20040 7438 20052
rect 7432 20012 9168 20040
rect 7432 20000 7438 20012
rect 5626 19932 5632 19984
rect 5684 19972 5690 19984
rect 7834 19972 7840 19984
rect 5684 19944 7840 19972
rect 5684 19932 5690 19944
rect 7834 19932 7840 19944
rect 7892 19932 7898 19984
rect 9140 19972 9168 20012
rect 9214 20000 9220 20052
rect 9272 20040 9278 20052
rect 10318 20040 10324 20052
rect 9272 20012 10324 20040
rect 9272 20000 9278 20012
rect 10318 20000 10324 20012
rect 10376 20000 10382 20052
rect 10594 20040 10600 20052
rect 10555 20012 10600 20040
rect 10594 20000 10600 20012
rect 10652 20000 10658 20052
rect 11057 20043 11115 20049
rect 11057 20009 11069 20043
rect 11103 20040 11115 20043
rect 12802 20040 12808 20052
rect 11103 20012 12808 20040
rect 11103 20009 11115 20012
rect 11057 20003 11115 20009
rect 12802 20000 12808 20012
rect 12860 20000 12866 20052
rect 14277 20043 14335 20049
rect 14277 20009 14289 20043
rect 14323 20040 14335 20043
rect 14734 20040 14740 20052
rect 14323 20012 14740 20040
rect 14323 20009 14335 20012
rect 14277 20003 14335 20009
rect 14734 20000 14740 20012
rect 14792 20000 14798 20052
rect 15749 20043 15807 20049
rect 15749 20009 15761 20043
rect 15795 20040 15807 20043
rect 16114 20040 16120 20052
rect 15795 20012 16120 20040
rect 15795 20009 15807 20012
rect 15749 20003 15807 20009
rect 16114 20000 16120 20012
rect 16172 20000 16178 20052
rect 17681 20043 17739 20049
rect 17681 20009 17693 20043
rect 17727 20040 17739 20043
rect 18138 20040 18144 20052
rect 17727 20012 18144 20040
rect 17727 20009 17739 20012
rect 17681 20003 17739 20009
rect 18138 20000 18144 20012
rect 18196 20000 18202 20052
rect 18785 20043 18843 20049
rect 18785 20009 18797 20043
rect 18831 20040 18843 20043
rect 19794 20040 19800 20052
rect 18831 20012 19800 20040
rect 18831 20009 18843 20012
rect 18785 20003 18843 20009
rect 19794 20000 19800 20012
rect 19852 20000 19858 20052
rect 19889 20043 19947 20049
rect 19889 20009 19901 20043
rect 19935 20040 19947 20043
rect 20806 20040 20812 20052
rect 19935 20012 20812 20040
rect 19935 20009 19947 20012
rect 19889 20003 19947 20009
rect 20806 20000 20812 20012
rect 20864 20000 20870 20052
rect 11238 19972 11244 19984
rect 9140 19944 11244 19972
rect 11238 19932 11244 19944
rect 11296 19932 11302 19984
rect 11330 19932 11336 19984
rect 11388 19972 11394 19984
rect 16942 19972 16948 19984
rect 11388 19944 16948 19972
rect 11388 19932 11394 19944
rect 16942 19932 16948 19944
rect 17000 19932 17006 19984
rect 1765 19907 1823 19913
rect 1765 19873 1777 19907
rect 1811 19904 1823 19907
rect 1854 19904 1860 19916
rect 1811 19876 1860 19904
rect 1811 19873 1823 19876
rect 1765 19867 1823 19873
rect 1854 19864 1860 19876
rect 1912 19864 1918 19916
rect 2869 19907 2927 19913
rect 2869 19873 2881 19907
rect 2915 19904 2927 19907
rect 3510 19904 3516 19916
rect 2915 19876 3516 19904
rect 2915 19873 2927 19876
rect 2869 19867 2927 19873
rect 3510 19864 3516 19876
rect 3568 19864 3574 19916
rect 3602 19864 3608 19916
rect 3660 19904 3666 19916
rect 4433 19907 4491 19913
rect 4433 19904 4445 19907
rect 3660 19876 4445 19904
rect 3660 19864 3666 19876
rect 4433 19873 4445 19876
rect 4479 19873 4491 19907
rect 4433 19867 4491 19873
rect 4522 19864 4528 19916
rect 4580 19904 4586 19916
rect 6621 19907 6679 19913
rect 6621 19904 6633 19907
rect 4580 19876 4625 19904
rect 5644 19876 6633 19904
rect 4580 19864 4586 19876
rect 5644 19848 5672 19876
rect 6621 19873 6633 19876
rect 6667 19904 6679 19907
rect 7098 19904 7104 19916
rect 6667 19876 7104 19904
rect 6667 19873 6679 19876
rect 6621 19867 6679 19873
rect 7098 19864 7104 19876
rect 7156 19864 7162 19916
rect 9858 19864 9864 19916
rect 9916 19904 9922 19916
rect 10965 19907 11023 19913
rect 10965 19904 10977 19907
rect 9916 19876 10977 19904
rect 9916 19864 9922 19876
rect 10965 19873 10977 19876
rect 11011 19873 11023 19907
rect 10965 19867 11023 19873
rect 12526 19864 12532 19916
rect 12584 19904 12590 19916
rect 12584 19876 12629 19904
rect 12584 19864 12590 19876
rect 12710 19864 12716 19916
rect 12768 19904 12774 19916
rect 12768 19876 13124 19904
rect 12768 19864 12774 19876
rect 4614 19836 4620 19848
rect 4575 19808 4620 19836
rect 4614 19796 4620 19808
rect 4672 19836 4678 19848
rect 5534 19836 5540 19848
rect 4672 19808 5540 19836
rect 4672 19796 4678 19808
rect 5534 19796 5540 19808
rect 5592 19796 5598 19848
rect 5626 19796 5632 19848
rect 5684 19796 5690 19848
rect 6365 19839 6423 19845
rect 6365 19805 6377 19839
rect 6411 19805 6423 19839
rect 6365 19799 6423 19805
rect 8573 19839 8631 19845
rect 8573 19805 8585 19839
rect 8619 19836 8631 19839
rect 8754 19836 8760 19848
rect 8619 19808 8760 19836
rect 8619 19805 8631 19808
rect 8573 19799 8631 19805
rect 4062 19768 4068 19780
rect 4023 19740 4068 19768
rect 4062 19728 4068 19740
rect 4120 19728 4126 19780
rect 6380 19700 6408 19799
rect 8754 19796 8760 19808
rect 8812 19796 8818 19848
rect 8846 19796 8852 19848
rect 8904 19836 8910 19848
rect 10226 19836 10232 19848
rect 8904 19808 10232 19836
rect 8904 19796 8910 19808
rect 10226 19796 10232 19808
rect 10284 19796 10290 19848
rect 11238 19836 11244 19848
rect 11199 19808 11244 19836
rect 11238 19796 11244 19808
rect 11296 19796 11302 19848
rect 11330 19796 11336 19848
rect 11388 19836 11394 19848
rect 12621 19839 12679 19845
rect 12621 19836 12633 19839
rect 11388 19808 12633 19836
rect 11388 19796 11394 19808
rect 12621 19805 12633 19808
rect 12667 19805 12679 19839
rect 12802 19836 12808 19848
rect 12763 19808 12808 19836
rect 12621 19799 12679 19805
rect 12802 19796 12808 19808
rect 12860 19796 12866 19848
rect 13096 19836 13124 19876
rect 13906 19864 13912 19916
rect 13964 19904 13970 19916
rect 14093 19907 14151 19913
rect 14093 19904 14105 19907
rect 13964 19876 14105 19904
rect 13964 19864 13970 19876
rect 14093 19873 14105 19876
rect 14139 19873 14151 19907
rect 14093 19867 14151 19873
rect 15565 19907 15623 19913
rect 15565 19873 15577 19907
rect 15611 19904 15623 19907
rect 17402 19904 17408 19916
rect 15611 19876 17408 19904
rect 15611 19873 15623 19876
rect 15565 19867 15623 19873
rect 17402 19864 17408 19876
rect 17460 19864 17466 19916
rect 17497 19907 17555 19913
rect 17497 19873 17509 19907
rect 17543 19873 17555 19907
rect 17497 19867 17555 19873
rect 18601 19907 18659 19913
rect 18601 19873 18613 19907
rect 18647 19904 18659 19907
rect 18874 19904 18880 19916
rect 18647 19876 18880 19904
rect 18647 19873 18659 19876
rect 18601 19867 18659 19873
rect 13096 19808 15332 19836
rect 7834 19728 7840 19780
rect 7892 19768 7898 19780
rect 15194 19768 15200 19780
rect 7892 19740 15200 19768
rect 7892 19728 7898 19740
rect 15194 19728 15200 19740
rect 15252 19728 15258 19780
rect 15304 19768 15332 19808
rect 16298 19768 16304 19780
rect 15304 19740 16304 19768
rect 16298 19728 16304 19740
rect 16356 19728 16362 19780
rect 7098 19700 7104 19712
rect 6380 19672 7104 19700
rect 7098 19660 7104 19672
rect 7156 19660 7162 19712
rect 7558 19660 7564 19712
rect 7616 19700 7622 19712
rect 7745 19703 7803 19709
rect 7745 19700 7757 19703
rect 7616 19672 7757 19700
rect 7616 19660 7622 19672
rect 7745 19669 7757 19672
rect 7791 19669 7803 19703
rect 7745 19663 7803 19669
rect 9766 19660 9772 19712
rect 9824 19700 9830 19712
rect 12161 19703 12219 19709
rect 12161 19700 12173 19703
rect 9824 19672 12173 19700
rect 9824 19660 9830 19672
rect 12161 19669 12173 19672
rect 12207 19669 12219 19703
rect 12161 19663 12219 19669
rect 12434 19660 12440 19712
rect 12492 19700 12498 19712
rect 17512 19700 17540 19867
rect 18874 19864 18880 19876
rect 18932 19864 18938 19916
rect 19705 19907 19763 19913
rect 19705 19873 19717 19907
rect 19751 19873 19763 19907
rect 19705 19867 19763 19873
rect 17862 19796 17868 19848
rect 17920 19836 17926 19848
rect 19720 19836 19748 19867
rect 17920 19808 19748 19836
rect 17920 19796 17926 19808
rect 12492 19672 17540 19700
rect 12492 19660 12498 19672
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 5534 19496 5540 19508
rect 5495 19468 5540 19496
rect 5534 19456 5540 19468
rect 5592 19456 5598 19508
rect 5902 19456 5908 19508
rect 5960 19496 5966 19508
rect 9214 19496 9220 19508
rect 5960 19468 9220 19496
rect 5960 19456 5966 19468
rect 9214 19456 9220 19468
rect 9272 19456 9278 19508
rect 11517 19499 11575 19505
rect 11517 19465 11529 19499
rect 11563 19496 11575 19499
rect 11974 19496 11980 19508
rect 11563 19468 11980 19496
rect 11563 19465 11575 19468
rect 11517 19459 11575 19465
rect 11974 19456 11980 19468
rect 12032 19456 12038 19508
rect 12894 19456 12900 19508
rect 12952 19496 12958 19508
rect 14550 19496 14556 19508
rect 12952 19468 14556 19496
rect 12952 19456 12958 19468
rect 14550 19456 14556 19468
rect 14608 19456 14614 19508
rect 13998 19388 14004 19440
rect 14056 19428 14062 19440
rect 14056 19400 18000 19428
rect 14056 19388 14062 19400
rect 2130 19320 2136 19372
rect 2188 19360 2194 19372
rect 2682 19360 2688 19372
rect 2188 19332 2688 19360
rect 2188 19320 2194 19332
rect 2682 19320 2688 19332
rect 2740 19360 2746 19372
rect 3145 19363 3203 19369
rect 3145 19360 3157 19363
rect 2740 19332 3157 19360
rect 2740 19320 2746 19332
rect 3145 19329 3157 19332
rect 3191 19329 3203 19363
rect 3145 19323 3203 19329
rect 3896 19332 4292 19360
rect 1486 19292 1492 19304
rect 1447 19264 1492 19292
rect 1486 19252 1492 19264
rect 1544 19252 1550 19304
rect 3418 19252 3424 19304
rect 3476 19292 3482 19304
rect 3896 19292 3924 19332
rect 3476 19264 3924 19292
rect 3476 19252 3482 19264
rect 3970 19252 3976 19304
rect 4028 19292 4034 19304
rect 4157 19295 4215 19301
rect 4157 19292 4169 19295
rect 4028 19264 4169 19292
rect 4028 19252 4034 19264
rect 4157 19261 4169 19264
rect 4203 19261 4215 19295
rect 4264 19292 4292 19332
rect 8846 19320 8852 19372
rect 8904 19360 8910 19372
rect 12250 19360 12256 19372
rect 8904 19332 10272 19360
rect 8904 19320 8910 19332
rect 6914 19292 6920 19304
rect 4264 19264 6920 19292
rect 4157 19255 4215 19261
rect 6914 19252 6920 19264
rect 6972 19252 6978 19304
rect 7098 19292 7104 19304
rect 7011 19264 7104 19292
rect 7098 19252 7104 19264
rect 7156 19292 7162 19304
rect 8202 19292 8208 19304
rect 7156 19264 8208 19292
rect 7156 19252 7162 19264
rect 8202 19252 8208 19264
rect 8260 19292 8266 19304
rect 10137 19295 10195 19301
rect 10137 19292 10149 19295
rect 8260 19264 10149 19292
rect 8260 19252 8266 19264
rect 10137 19261 10149 19264
rect 10183 19261 10195 19295
rect 10244 19292 10272 19332
rect 11164 19332 12256 19360
rect 11164 19292 11192 19332
rect 12250 19320 12256 19332
rect 12308 19320 12314 19372
rect 15010 19320 15016 19372
rect 15068 19360 15074 19372
rect 15068 19332 15113 19360
rect 15068 19320 15074 19332
rect 12434 19292 12440 19304
rect 10244 19264 11192 19292
rect 12395 19264 12440 19292
rect 10137 19255 10195 19261
rect 12434 19252 12440 19264
rect 12492 19252 12498 19304
rect 13078 19252 13084 19304
rect 13136 19292 13142 19304
rect 13725 19295 13783 19301
rect 13725 19292 13737 19295
rect 13136 19264 13737 19292
rect 13136 19252 13142 19264
rect 13725 19261 13737 19264
rect 13771 19261 13783 19295
rect 13725 19255 13783 19261
rect 14458 19252 14464 19304
rect 14516 19292 14522 19304
rect 14829 19295 14887 19301
rect 14829 19292 14841 19295
rect 14516 19264 14841 19292
rect 14516 19252 14522 19264
rect 14829 19261 14841 19264
rect 14875 19261 14887 19295
rect 14829 19255 14887 19261
rect 15286 19252 15292 19304
rect 15344 19292 15350 19304
rect 16117 19295 16175 19301
rect 16117 19292 16129 19295
rect 15344 19264 16129 19292
rect 15344 19252 15350 19264
rect 16117 19261 16129 19264
rect 16163 19261 16175 19295
rect 17034 19292 17040 19304
rect 16117 19255 16175 19261
rect 16224 19264 17040 19292
rect 2774 19224 2780 19236
rect 1688 19196 2780 19224
rect 1688 19165 1716 19196
rect 2774 19184 2780 19196
rect 2832 19184 2838 19236
rect 3053 19227 3111 19233
rect 3053 19193 3065 19227
rect 3099 19224 3111 19227
rect 4246 19224 4252 19236
rect 3099 19196 4252 19224
rect 3099 19193 3111 19196
rect 3053 19187 3111 19193
rect 4246 19184 4252 19196
rect 4304 19184 4310 19236
rect 4424 19227 4482 19233
rect 4424 19193 4436 19227
rect 4470 19224 4482 19227
rect 5442 19224 5448 19236
rect 4470 19196 5448 19224
rect 4470 19193 4482 19196
rect 4424 19187 4482 19193
rect 5442 19184 5448 19196
rect 5500 19184 5506 19236
rect 7368 19227 7426 19233
rect 7368 19193 7380 19227
rect 7414 19224 7426 19227
rect 7558 19224 7564 19236
rect 7414 19196 7564 19224
rect 7414 19193 7426 19196
rect 7368 19187 7426 19193
rect 7558 19184 7564 19196
rect 7616 19184 7622 19236
rect 7668 19196 8616 19224
rect 1673 19159 1731 19165
rect 1673 19125 1685 19159
rect 1719 19125 1731 19159
rect 1673 19119 1731 19125
rect 2593 19159 2651 19165
rect 2593 19125 2605 19159
rect 2639 19156 2651 19159
rect 2682 19156 2688 19168
rect 2639 19128 2688 19156
rect 2639 19125 2651 19128
rect 2593 19119 2651 19125
rect 2682 19116 2688 19128
rect 2740 19116 2746 19168
rect 2958 19156 2964 19168
rect 2919 19128 2964 19156
rect 2958 19116 2964 19128
rect 3016 19116 3022 19168
rect 4062 19116 4068 19168
rect 4120 19156 4126 19168
rect 7668 19156 7696 19196
rect 8478 19156 8484 19168
rect 4120 19128 7696 19156
rect 8439 19128 8484 19156
rect 4120 19116 4126 19128
rect 8478 19116 8484 19128
rect 8536 19116 8542 19168
rect 8588 19156 8616 19196
rect 9122 19184 9128 19236
rect 9180 19224 9186 19236
rect 10226 19224 10232 19236
rect 9180 19196 10232 19224
rect 9180 19184 9186 19196
rect 10226 19184 10232 19196
rect 10284 19184 10290 19236
rect 10404 19227 10462 19233
rect 10404 19193 10416 19227
rect 10450 19224 10462 19227
rect 10962 19224 10968 19236
rect 10450 19196 10968 19224
rect 10450 19193 10462 19196
rect 10404 19187 10462 19193
rect 10962 19184 10968 19196
rect 11020 19184 11026 19236
rect 12713 19227 12771 19233
rect 12713 19193 12725 19227
rect 12759 19224 12771 19227
rect 13446 19224 13452 19236
rect 12759 19196 13452 19224
rect 12759 19193 12771 19196
rect 12713 19187 12771 19193
rect 13446 19184 13452 19196
rect 13504 19184 13510 19236
rect 16224 19224 16252 19264
rect 17034 19252 17040 19264
rect 17092 19252 17098 19304
rect 16390 19224 16396 19236
rect 15120 19196 16252 19224
rect 16351 19196 16396 19224
rect 13909 19159 13967 19165
rect 13909 19156 13921 19159
rect 8588 19128 13921 19156
rect 13909 19125 13921 19128
rect 13955 19125 13967 19159
rect 13909 19119 13967 19125
rect 13998 19116 14004 19168
rect 14056 19156 14062 19168
rect 15120 19156 15148 19196
rect 16390 19184 16396 19196
rect 16448 19184 16454 19236
rect 17972 19224 18000 19400
rect 19521 19295 19579 19301
rect 19521 19261 19533 19295
rect 19567 19292 19579 19295
rect 19610 19292 19616 19304
rect 19567 19264 19616 19292
rect 19567 19261 19579 19264
rect 19521 19255 19579 19261
rect 19610 19252 19616 19264
rect 19668 19252 19674 19304
rect 20625 19227 20683 19233
rect 20625 19224 20637 19227
rect 17972 19196 20637 19224
rect 20625 19193 20637 19196
rect 20671 19193 20683 19227
rect 20625 19187 20683 19193
rect 14056 19128 15148 19156
rect 14056 19116 14062 19128
rect 15194 19116 15200 19168
rect 15252 19156 15258 19168
rect 18049 19159 18107 19165
rect 18049 19156 18061 19159
rect 15252 19128 18061 19156
rect 15252 19116 15258 19128
rect 18049 19125 18061 19128
rect 18095 19125 18107 19159
rect 18049 19119 18107 19125
rect 19705 19159 19763 19165
rect 19705 19125 19717 19159
rect 19751 19156 19763 19159
rect 20346 19156 20352 19168
rect 19751 19128 20352 19156
rect 19751 19125 19763 19128
rect 19705 19119 19763 19125
rect 20346 19116 20352 19128
rect 20404 19116 20410 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 2866 18912 2872 18964
rect 2924 18952 2930 18964
rect 3053 18955 3111 18961
rect 3053 18952 3065 18955
rect 2924 18924 3065 18952
rect 2924 18912 2930 18924
rect 3053 18921 3065 18924
rect 3099 18921 3111 18955
rect 3053 18915 3111 18921
rect 4065 18955 4123 18961
rect 4065 18921 4077 18955
rect 4111 18952 4123 18955
rect 6089 18955 6147 18961
rect 6089 18952 6101 18955
rect 4111 18924 6101 18952
rect 4111 18921 4123 18924
rect 4065 18915 4123 18921
rect 6089 18921 6101 18924
rect 6135 18921 6147 18955
rect 6089 18915 6147 18921
rect 6914 18912 6920 18964
rect 6972 18952 6978 18964
rect 6972 18924 7604 18952
rect 6972 18912 6978 18924
rect 198 18844 204 18896
rect 256 18884 262 18896
rect 4525 18887 4583 18893
rect 256 18856 4384 18884
rect 256 18844 262 18856
rect 1762 18816 1768 18828
rect 1723 18788 1768 18816
rect 1762 18776 1768 18788
rect 1820 18776 1826 18828
rect 2869 18819 2927 18825
rect 2869 18785 2881 18819
rect 2915 18816 2927 18819
rect 4246 18816 4252 18828
rect 2915 18788 4252 18816
rect 2915 18785 2927 18788
rect 2869 18779 2927 18785
rect 4246 18776 4252 18788
rect 4304 18776 4310 18828
rect 658 18708 664 18760
rect 716 18748 722 18760
rect 3786 18748 3792 18760
rect 716 18720 3792 18748
rect 716 18708 722 18720
rect 3786 18708 3792 18720
rect 3844 18708 3850 18760
rect 1118 18640 1124 18692
rect 1176 18680 1182 18692
rect 3694 18680 3700 18692
rect 1176 18652 3700 18680
rect 1176 18640 1182 18652
rect 3694 18640 3700 18652
rect 3752 18640 3758 18692
rect 4356 18680 4384 18856
rect 4525 18853 4537 18887
rect 4571 18884 4583 18887
rect 7190 18884 7196 18896
rect 4571 18856 7196 18884
rect 4571 18853 4583 18856
rect 4525 18847 4583 18853
rect 7190 18844 7196 18856
rect 7248 18844 7254 18896
rect 4433 18819 4491 18825
rect 4433 18785 4445 18819
rect 4479 18816 4491 18819
rect 4706 18816 4712 18828
rect 4479 18788 4712 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 4706 18776 4712 18788
rect 4764 18776 4770 18828
rect 4890 18776 4896 18828
rect 4948 18816 4954 18828
rect 5997 18819 6055 18825
rect 5997 18816 6009 18819
rect 4948 18788 6009 18816
rect 4948 18776 4954 18788
rect 5997 18785 6009 18788
rect 6043 18785 6055 18819
rect 5997 18779 6055 18785
rect 7282 18776 7288 18828
rect 7340 18816 7346 18828
rect 7449 18819 7507 18825
rect 7449 18816 7461 18819
rect 7340 18788 7461 18816
rect 7340 18776 7346 18788
rect 7449 18785 7461 18788
rect 7495 18785 7507 18819
rect 7576 18816 7604 18924
rect 7650 18912 7656 18964
rect 7708 18952 7714 18964
rect 8202 18952 8208 18964
rect 7708 18924 8208 18952
rect 7708 18912 7714 18924
rect 8202 18912 8208 18924
rect 8260 18912 8266 18964
rect 9674 18912 9680 18964
rect 9732 18952 9738 18964
rect 10137 18955 10195 18961
rect 10137 18952 10149 18955
rect 9732 18924 10149 18952
rect 9732 18912 9738 18924
rect 10137 18921 10149 18924
rect 10183 18921 10195 18955
rect 10137 18915 10195 18921
rect 12250 18912 12256 18964
rect 12308 18952 12314 18964
rect 15657 18955 15715 18961
rect 15657 18952 15669 18955
rect 12308 18924 15669 18952
rect 12308 18912 12314 18924
rect 15657 18921 15669 18924
rect 15703 18952 15715 18955
rect 17313 18955 17371 18961
rect 17313 18952 17325 18955
rect 15703 18924 17325 18952
rect 15703 18921 15715 18924
rect 15657 18915 15715 18921
rect 17313 18921 17325 18924
rect 17359 18921 17371 18955
rect 17313 18915 17371 18921
rect 19889 18955 19947 18961
rect 19889 18921 19901 18955
rect 19935 18952 19947 18955
rect 22186 18952 22192 18964
rect 19935 18924 22192 18952
rect 19935 18921 19947 18924
rect 19889 18915 19947 18921
rect 22186 18912 22192 18924
rect 22244 18912 22250 18964
rect 7834 18844 7840 18896
rect 7892 18884 7898 18896
rect 15194 18884 15200 18896
rect 7892 18856 10272 18884
rect 7892 18844 7898 18856
rect 9950 18816 9956 18828
rect 7576 18788 9956 18816
rect 7449 18779 7507 18785
rect 9950 18776 9956 18788
rect 10008 18776 10014 18828
rect 10045 18819 10103 18825
rect 10045 18785 10057 18819
rect 10091 18785 10103 18819
rect 10045 18779 10103 18785
rect 4614 18748 4620 18760
rect 4575 18720 4620 18748
rect 4614 18708 4620 18720
rect 4672 18708 4678 18760
rect 4798 18708 4804 18760
rect 4856 18748 4862 18760
rect 6181 18751 6239 18757
rect 6181 18748 6193 18751
rect 4856 18720 6193 18748
rect 4856 18708 4862 18720
rect 6181 18717 6193 18720
rect 6227 18717 6239 18751
rect 6181 18711 6239 18717
rect 7098 18708 7104 18760
rect 7156 18748 7162 18760
rect 7193 18751 7251 18757
rect 7193 18748 7205 18751
rect 7156 18720 7205 18748
rect 7156 18708 7162 18720
rect 7193 18717 7205 18720
rect 7239 18717 7251 18751
rect 7193 18711 7251 18717
rect 8202 18708 8208 18760
rect 8260 18748 8266 18760
rect 8260 18720 9996 18748
rect 8260 18708 8266 18720
rect 9214 18680 9220 18692
rect 4356 18652 5764 18680
rect 1949 18615 2007 18621
rect 1949 18581 1961 18615
rect 1995 18612 2007 18615
rect 2866 18612 2872 18624
rect 1995 18584 2872 18612
rect 1995 18581 2007 18584
rect 1949 18575 2007 18581
rect 2866 18572 2872 18584
rect 2924 18572 2930 18624
rect 4246 18572 4252 18624
rect 4304 18612 4310 18624
rect 5258 18612 5264 18624
rect 4304 18584 5264 18612
rect 4304 18572 4310 18584
rect 5258 18572 5264 18584
rect 5316 18572 5322 18624
rect 5626 18612 5632 18624
rect 5587 18584 5632 18612
rect 5626 18572 5632 18584
rect 5684 18572 5690 18624
rect 5736 18612 5764 18652
rect 8128 18652 9220 18680
rect 8128 18612 8156 18652
rect 9214 18640 9220 18652
rect 9272 18640 9278 18692
rect 8570 18612 8576 18624
rect 5736 18584 8156 18612
rect 8531 18584 8576 18612
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 9306 18572 9312 18624
rect 9364 18612 9370 18624
rect 9677 18615 9735 18621
rect 9677 18612 9689 18615
rect 9364 18584 9689 18612
rect 9364 18572 9370 18584
rect 9677 18581 9689 18584
rect 9723 18581 9735 18615
rect 9968 18612 9996 18720
rect 10060 18680 10088 18779
rect 10244 18757 10272 18856
rect 13004 18856 15200 18884
rect 10778 18776 10784 18828
rect 10836 18816 10842 18828
rect 11698 18816 11704 18828
rect 10836 18788 11704 18816
rect 10836 18776 10842 18788
rect 11698 18776 11704 18788
rect 11756 18776 11762 18828
rect 13004 18825 13032 18856
rect 15194 18844 15200 18856
rect 15252 18844 15258 18896
rect 15470 18844 15476 18896
rect 15528 18884 15534 18896
rect 15749 18887 15807 18893
rect 15749 18884 15761 18887
rect 15528 18856 15761 18884
rect 15528 18844 15534 18856
rect 15749 18853 15761 18856
rect 15795 18853 15807 18887
rect 17954 18884 17960 18896
rect 15749 18847 15807 18853
rect 16500 18856 17960 18884
rect 12989 18819 13047 18825
rect 12989 18785 13001 18819
rect 13035 18785 13047 18819
rect 12989 18779 13047 18785
rect 13538 18776 13544 18828
rect 13596 18816 13602 18828
rect 14093 18819 14151 18825
rect 14093 18816 14105 18819
rect 13596 18788 14105 18816
rect 13596 18776 13602 18788
rect 14093 18785 14105 18788
rect 14139 18785 14151 18819
rect 14093 18779 14151 18785
rect 16022 18776 16028 18828
rect 16080 18816 16086 18828
rect 16500 18816 16528 18856
rect 17954 18844 17960 18856
rect 18012 18844 18018 18896
rect 17218 18816 17224 18828
rect 16080 18788 16528 18816
rect 17179 18788 17224 18816
rect 16080 18776 16086 18788
rect 17218 18776 17224 18788
rect 17276 18776 17282 18828
rect 18690 18776 18696 18828
rect 18748 18816 18754 18828
rect 19705 18819 19763 18825
rect 19705 18816 19717 18819
rect 18748 18788 19717 18816
rect 18748 18776 18754 18788
rect 19705 18785 19717 18788
rect 19751 18785 19763 18819
rect 19705 18779 19763 18785
rect 10229 18751 10287 18757
rect 10229 18717 10241 18751
rect 10275 18717 10287 18751
rect 10229 18711 10287 18717
rect 11241 18751 11299 18757
rect 11241 18717 11253 18751
rect 11287 18748 11299 18751
rect 11974 18748 11980 18760
rect 11287 18720 11980 18748
rect 11287 18717 11299 18720
rect 11241 18711 11299 18717
rect 11974 18708 11980 18720
rect 12032 18708 12038 18760
rect 12434 18708 12440 18760
rect 12492 18748 12498 18760
rect 12618 18748 12624 18760
rect 12492 18720 12624 18748
rect 12492 18708 12498 18720
rect 12618 18708 12624 18720
rect 12676 18708 12682 18760
rect 12802 18708 12808 18760
rect 12860 18748 12866 18760
rect 13262 18748 13268 18760
rect 12860 18720 13268 18748
rect 12860 18708 12866 18720
rect 13262 18708 13268 18720
rect 13320 18708 13326 18760
rect 13630 18708 13636 18760
rect 13688 18748 13694 18760
rect 15286 18748 15292 18760
rect 13688 18720 15292 18748
rect 13688 18708 13694 18720
rect 15286 18708 15292 18720
rect 15344 18708 15350 18760
rect 15933 18751 15991 18757
rect 15933 18717 15945 18751
rect 15979 18748 15991 18751
rect 16114 18748 16120 18760
rect 15979 18720 16120 18748
rect 15979 18717 15991 18720
rect 15933 18711 15991 18717
rect 16114 18708 16120 18720
rect 16172 18708 16178 18760
rect 17497 18751 17555 18757
rect 17497 18717 17509 18751
rect 17543 18748 17555 18751
rect 17678 18748 17684 18760
rect 17543 18720 17684 18748
rect 17543 18717 17555 18720
rect 17497 18711 17555 18717
rect 17678 18708 17684 18720
rect 17736 18708 17742 18760
rect 18417 18751 18475 18757
rect 18417 18717 18429 18751
rect 18463 18717 18475 18751
rect 18417 18711 18475 18717
rect 18432 18680 18460 18711
rect 10060 18652 15700 18680
rect 12894 18612 12900 18624
rect 9968 18584 12900 18612
rect 9677 18575 9735 18581
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 13173 18615 13231 18621
rect 13173 18581 13185 18615
rect 13219 18612 13231 18615
rect 13998 18612 14004 18624
rect 13219 18584 14004 18612
rect 13219 18581 13231 18584
rect 13173 18575 13231 18581
rect 13998 18572 14004 18584
rect 14056 18572 14062 18624
rect 14277 18615 14335 18621
rect 14277 18581 14289 18615
rect 14323 18612 14335 18615
rect 15194 18612 15200 18624
rect 14323 18584 15200 18612
rect 14323 18581 14335 18584
rect 14277 18575 14335 18581
rect 15194 18572 15200 18584
rect 15252 18572 15258 18624
rect 15289 18615 15347 18621
rect 15289 18581 15301 18615
rect 15335 18612 15347 18615
rect 15562 18612 15568 18624
rect 15335 18584 15568 18612
rect 15335 18581 15347 18584
rect 15289 18575 15347 18581
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 15672 18612 15700 18652
rect 15948 18652 18460 18680
rect 15948 18612 15976 18652
rect 15672 18584 15976 18612
rect 16853 18615 16911 18621
rect 16853 18581 16865 18615
rect 16899 18612 16911 18615
rect 18138 18612 18144 18624
rect 16899 18584 18144 18612
rect 16899 18581 16911 18584
rect 16853 18575 16911 18581
rect 18138 18572 18144 18584
rect 18196 18572 18202 18624
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 1670 18368 1676 18420
rect 1728 18408 1734 18420
rect 2590 18408 2596 18420
rect 1728 18380 2596 18408
rect 1728 18368 1734 18380
rect 2590 18368 2596 18380
rect 2648 18368 2654 18420
rect 2869 18411 2927 18417
rect 2869 18377 2881 18411
rect 2915 18408 2927 18411
rect 12710 18408 12716 18420
rect 2915 18380 12716 18408
rect 2915 18377 2927 18380
rect 2869 18371 2927 18377
rect 12710 18368 12716 18380
rect 12768 18368 12774 18420
rect 16945 18411 17003 18417
rect 16945 18408 16957 18411
rect 12820 18380 16957 18408
rect 2498 18300 2504 18352
rect 2556 18340 2562 18352
rect 5905 18343 5963 18349
rect 2556 18312 4375 18340
rect 2556 18300 2562 18312
rect 2038 18232 2044 18284
rect 2096 18272 2102 18284
rect 2869 18275 2927 18281
rect 2869 18272 2881 18275
rect 2096 18244 2881 18272
rect 2096 18232 2102 18244
rect 2869 18241 2881 18244
rect 2915 18241 2927 18275
rect 2869 18235 2927 18241
rect 3605 18275 3663 18281
rect 3605 18241 3617 18275
rect 3651 18272 3663 18275
rect 4246 18272 4252 18284
rect 3651 18244 4252 18272
rect 3651 18241 3663 18244
rect 3605 18235 3663 18241
rect 4246 18232 4252 18244
rect 4304 18232 4310 18284
rect 4347 18272 4375 18312
rect 5905 18309 5917 18343
rect 5951 18340 5963 18343
rect 7282 18340 7288 18352
rect 5951 18312 7288 18340
rect 5951 18309 5963 18312
rect 5905 18303 5963 18309
rect 7282 18300 7288 18312
rect 7340 18300 7346 18352
rect 9214 18300 9220 18352
rect 9272 18340 9278 18352
rect 12342 18340 12348 18352
rect 9272 18312 12348 18340
rect 9272 18300 9278 18312
rect 12342 18300 12348 18312
rect 12400 18300 12406 18352
rect 4347 18244 4660 18272
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18204 1823 18207
rect 2314 18204 2320 18216
rect 1811 18176 2320 18204
rect 1811 18173 1823 18176
rect 1765 18167 1823 18173
rect 2314 18164 2320 18176
rect 2372 18164 2378 18216
rect 3142 18164 3148 18216
rect 3200 18204 3206 18216
rect 3200 18176 3556 18204
rect 3200 18164 3206 18176
rect 2590 18096 2596 18148
rect 2648 18136 2654 18148
rect 3421 18139 3479 18145
rect 3421 18136 3433 18139
rect 2648 18108 3433 18136
rect 2648 18096 2654 18108
rect 3421 18105 3433 18108
rect 3467 18105 3479 18139
rect 3528 18136 3556 18176
rect 3970 18164 3976 18216
rect 4028 18204 4034 18216
rect 4525 18207 4583 18213
rect 4525 18204 4537 18207
rect 4028 18176 4537 18204
rect 4028 18164 4034 18176
rect 4525 18173 4537 18176
rect 4571 18173 4583 18207
rect 4632 18204 4660 18244
rect 5626 18232 5632 18284
rect 5684 18272 5690 18284
rect 7466 18272 7472 18284
rect 5684 18244 7472 18272
rect 5684 18232 5690 18244
rect 7466 18232 7472 18244
rect 7524 18232 7530 18284
rect 8202 18272 8208 18284
rect 8163 18244 8208 18272
rect 8202 18232 8208 18244
rect 8260 18232 8266 18284
rect 9674 18232 9680 18284
rect 9732 18272 9738 18284
rect 9858 18272 9864 18284
rect 9732 18244 9864 18272
rect 9732 18232 9738 18244
rect 9858 18232 9864 18244
rect 9916 18232 9922 18284
rect 10686 18232 10692 18284
rect 10744 18272 10750 18284
rect 12820 18272 12848 18380
rect 10744 18244 12848 18272
rect 10744 18232 10750 18244
rect 12894 18232 12900 18284
rect 12952 18232 12958 18284
rect 13004 18281 13032 18380
rect 16945 18377 16957 18380
rect 16991 18377 17003 18411
rect 16945 18371 17003 18377
rect 17678 18368 17684 18420
rect 17736 18408 17742 18420
rect 17773 18411 17831 18417
rect 17773 18408 17785 18411
rect 17736 18380 17785 18408
rect 17736 18368 17742 18380
rect 17773 18377 17785 18380
rect 17819 18377 17831 18411
rect 17773 18371 17831 18377
rect 20717 18411 20775 18417
rect 20717 18377 20729 18411
rect 20763 18408 20775 18411
rect 21726 18408 21732 18420
rect 20763 18380 21732 18408
rect 20763 18377 20775 18380
rect 20717 18371 20775 18377
rect 21726 18368 21732 18380
rect 21784 18368 21790 18420
rect 14001 18343 14059 18349
rect 14001 18309 14013 18343
rect 14047 18340 14059 18343
rect 15194 18340 15200 18352
rect 14047 18312 15200 18340
rect 14047 18309 14059 18312
rect 14001 18303 14059 18309
rect 15194 18300 15200 18312
rect 15252 18300 15258 18352
rect 12989 18275 13047 18281
rect 12989 18241 13001 18275
rect 13035 18241 13047 18275
rect 12989 18235 13047 18241
rect 14645 18275 14703 18281
rect 14645 18241 14657 18275
rect 14691 18272 14703 18275
rect 14734 18272 14740 18284
rect 14691 18244 14740 18272
rect 14691 18241 14703 18244
rect 14645 18235 14703 18241
rect 14734 18232 14740 18244
rect 14792 18232 14798 18284
rect 15286 18232 15292 18284
rect 15344 18272 15350 18284
rect 15565 18275 15623 18281
rect 15565 18272 15577 18275
rect 15344 18244 15577 18272
rect 15344 18232 15350 18244
rect 15565 18241 15577 18244
rect 15611 18241 15623 18275
rect 15565 18235 15623 18241
rect 16850 18232 16856 18284
rect 16908 18272 16914 18284
rect 17034 18272 17040 18284
rect 16908 18244 17040 18272
rect 16908 18232 16914 18244
rect 17034 18232 17040 18244
rect 17092 18272 17098 18284
rect 18509 18275 18567 18281
rect 18509 18272 18521 18275
rect 17092 18244 18521 18272
rect 17092 18232 17098 18244
rect 18509 18241 18521 18244
rect 18555 18241 18567 18275
rect 18509 18235 18567 18241
rect 18693 18275 18751 18281
rect 18693 18241 18705 18275
rect 18739 18272 18751 18275
rect 18966 18272 18972 18284
rect 18739 18244 18972 18272
rect 18739 18241 18751 18244
rect 18693 18235 18751 18241
rect 18966 18232 18972 18244
rect 19024 18232 19030 18284
rect 4632 18176 8616 18204
rect 4525 18167 4583 18173
rect 4792 18139 4850 18145
rect 3528 18108 4375 18136
rect 3421 18099 3479 18105
rect 1949 18071 2007 18077
rect 1949 18037 1961 18071
rect 1995 18068 2007 18071
rect 2774 18068 2780 18080
rect 1995 18040 2780 18068
rect 1995 18037 2007 18040
rect 1949 18031 2007 18037
rect 2774 18028 2780 18040
rect 2832 18028 2838 18080
rect 2961 18071 3019 18077
rect 2961 18037 2973 18071
rect 3007 18068 3019 18071
rect 3142 18068 3148 18080
rect 3007 18040 3148 18068
rect 3007 18037 3019 18040
rect 2961 18031 3019 18037
rect 3142 18028 3148 18040
rect 3200 18028 3206 18080
rect 3326 18068 3332 18080
rect 3287 18040 3332 18068
rect 3326 18028 3332 18040
rect 3384 18028 3390 18080
rect 3878 18028 3884 18080
rect 3936 18068 3942 18080
rect 4246 18068 4252 18080
rect 3936 18040 4252 18068
rect 3936 18028 3942 18040
rect 4246 18028 4252 18040
rect 4304 18028 4310 18080
rect 4347 18068 4375 18108
rect 4792 18105 4804 18139
rect 4838 18136 4850 18139
rect 5994 18136 6000 18148
rect 4838 18108 6000 18136
rect 4838 18105 4850 18108
rect 4792 18099 4850 18105
rect 5994 18096 6000 18108
rect 6052 18096 6058 18148
rect 8478 18145 8484 18148
rect 8472 18136 8484 18145
rect 8439 18108 8484 18136
rect 8472 18099 8484 18108
rect 8478 18096 8484 18099
rect 8536 18096 8542 18148
rect 8588 18136 8616 18176
rect 8938 18164 8944 18216
rect 8996 18204 9002 18216
rect 10870 18204 10876 18216
rect 8996 18176 10876 18204
rect 8996 18164 9002 18176
rect 10870 18164 10876 18176
rect 10928 18164 10934 18216
rect 12912 18204 12940 18232
rect 12636 18176 12940 18204
rect 12636 18136 12664 18176
rect 14182 18164 14188 18216
rect 14240 18204 14246 18216
rect 14461 18207 14519 18213
rect 14461 18204 14473 18207
rect 14240 18176 14473 18204
rect 14240 18164 14246 18176
rect 14461 18173 14473 18176
rect 14507 18173 14519 18207
rect 20533 18207 20591 18213
rect 20533 18204 20545 18207
rect 14461 18167 14519 18173
rect 14568 18176 20545 18204
rect 12897 18139 12955 18145
rect 12897 18136 12909 18139
rect 8588 18108 12664 18136
rect 12728 18108 12909 18136
rect 12728 18080 12756 18108
rect 12897 18105 12909 18108
rect 12943 18105 12955 18139
rect 12897 18099 12955 18105
rect 13814 18096 13820 18148
rect 13872 18136 13878 18148
rect 14568 18136 14596 18176
rect 20533 18173 20545 18176
rect 20579 18173 20591 18207
rect 20533 18167 20591 18173
rect 13872 18108 14596 18136
rect 13872 18096 13878 18108
rect 15378 18096 15384 18148
rect 15436 18136 15442 18148
rect 15810 18139 15868 18145
rect 15810 18136 15822 18139
rect 15436 18108 15822 18136
rect 15436 18096 15442 18108
rect 15810 18105 15822 18108
rect 15856 18105 15868 18139
rect 15810 18099 15868 18105
rect 17678 18096 17684 18148
rect 17736 18136 17742 18148
rect 18417 18139 18475 18145
rect 18417 18136 18429 18139
rect 17736 18108 18429 18136
rect 17736 18096 17742 18108
rect 18417 18105 18429 18108
rect 18463 18136 18475 18139
rect 18877 18139 18935 18145
rect 18877 18136 18889 18139
rect 18463 18108 18889 18136
rect 18463 18105 18475 18108
rect 18417 18099 18475 18105
rect 18877 18105 18889 18108
rect 18923 18105 18935 18139
rect 18877 18099 18935 18105
rect 6178 18068 6184 18080
rect 4347 18040 6184 18068
rect 6178 18028 6184 18040
rect 6236 18028 6242 18080
rect 6822 18068 6828 18080
rect 6783 18040 6828 18068
rect 6822 18028 6828 18040
rect 6880 18028 6886 18080
rect 9582 18068 9588 18080
rect 9543 18040 9588 18068
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 10413 18071 10471 18077
rect 10413 18037 10425 18071
rect 10459 18068 10471 18071
rect 11146 18068 11152 18080
rect 10459 18040 11152 18068
rect 10459 18037 10471 18040
rect 10413 18031 10471 18037
rect 11146 18028 11152 18040
rect 11204 18028 11210 18080
rect 12158 18028 12164 18080
rect 12216 18068 12222 18080
rect 12437 18071 12495 18077
rect 12437 18068 12449 18071
rect 12216 18040 12449 18068
rect 12216 18028 12222 18040
rect 12437 18037 12449 18040
rect 12483 18037 12495 18071
rect 12437 18031 12495 18037
rect 12710 18028 12716 18080
rect 12768 18028 12774 18080
rect 12805 18071 12863 18077
rect 12805 18037 12817 18071
rect 12851 18068 12863 18071
rect 13998 18068 14004 18080
rect 12851 18040 14004 18068
rect 12851 18037 12863 18040
rect 12805 18031 12863 18037
rect 13998 18028 14004 18040
rect 14056 18028 14062 18080
rect 14366 18068 14372 18080
rect 14327 18040 14372 18068
rect 14366 18028 14372 18040
rect 14424 18028 14430 18080
rect 14734 18028 14740 18080
rect 14792 18068 14798 18080
rect 16114 18068 16120 18080
rect 14792 18040 16120 18068
rect 14792 18028 14798 18040
rect 16114 18028 16120 18040
rect 16172 18028 16178 18080
rect 16390 18028 16396 18080
rect 16448 18068 16454 18080
rect 17773 18071 17831 18077
rect 17773 18068 17785 18071
rect 16448 18040 17785 18068
rect 16448 18028 16454 18040
rect 17773 18037 17785 18040
rect 17819 18037 17831 18071
rect 18046 18068 18052 18080
rect 18007 18040 18052 18068
rect 17773 18031 17831 18037
rect 18046 18028 18052 18040
rect 18104 18028 18110 18080
rect 20254 18028 20260 18080
rect 20312 18068 20318 18080
rect 22646 18068 22652 18080
rect 20312 18040 22652 18068
rect 20312 18028 20318 18040
rect 22646 18028 22652 18040
rect 22704 18028 22710 18080
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 7650 17864 7656 17876
rect 2056 17836 7656 17864
rect 2056 17737 2084 17836
rect 7650 17824 7656 17836
rect 7708 17824 7714 17876
rect 9030 17824 9036 17876
rect 9088 17864 9094 17876
rect 9490 17864 9496 17876
rect 9088 17836 9496 17864
rect 9088 17824 9094 17836
rect 9490 17824 9496 17836
rect 9548 17824 9554 17876
rect 9582 17824 9588 17876
rect 9640 17864 9646 17876
rect 11698 17864 11704 17876
rect 9640 17836 11704 17864
rect 9640 17824 9646 17836
rect 11698 17824 11704 17836
rect 11756 17824 11762 17876
rect 11882 17824 11888 17876
rect 11940 17864 11946 17876
rect 12069 17867 12127 17873
rect 12069 17864 12081 17867
rect 11940 17836 12081 17864
rect 11940 17824 11946 17836
rect 12069 17833 12081 17836
rect 12115 17864 12127 17867
rect 12250 17864 12256 17876
rect 12115 17836 12256 17864
rect 12115 17833 12127 17836
rect 12069 17827 12127 17833
rect 12250 17824 12256 17836
rect 12308 17824 12314 17876
rect 14277 17867 14335 17873
rect 14277 17833 14289 17867
rect 14323 17833 14335 17867
rect 14277 17827 14335 17833
rect 15289 17867 15347 17873
rect 15289 17833 15301 17867
rect 15335 17864 15347 17867
rect 18598 17864 18604 17876
rect 15335 17836 18604 17864
rect 15335 17833 15347 17836
rect 15289 17827 15347 17833
rect 4062 17756 4068 17808
rect 4120 17796 4126 17808
rect 13354 17796 13360 17808
rect 4120 17768 13360 17796
rect 4120 17756 4126 17768
rect 13354 17756 13360 17768
rect 13412 17756 13418 17808
rect 14292 17796 14320 17827
rect 18598 17824 18604 17836
rect 18656 17824 18662 17876
rect 18785 17867 18843 17873
rect 18785 17833 18797 17867
rect 18831 17864 18843 17867
rect 19058 17864 19064 17876
rect 18831 17836 19064 17864
rect 18831 17833 18843 17836
rect 18785 17827 18843 17833
rect 19058 17824 19064 17836
rect 19116 17824 19122 17876
rect 16482 17796 16488 17808
rect 13464 17768 14228 17796
rect 14292 17768 16488 17796
rect 2041 17731 2099 17737
rect 2041 17697 2053 17731
rect 2087 17697 2099 17731
rect 2041 17691 2099 17697
rect 4332 17731 4390 17737
rect 4332 17697 4344 17731
rect 4378 17728 4390 17731
rect 4798 17728 4804 17740
rect 4378 17700 4804 17728
rect 4378 17697 4390 17700
rect 4332 17691 4390 17697
rect 4798 17688 4804 17700
rect 4856 17688 4862 17740
rect 7190 17688 7196 17740
rect 7248 17728 7254 17740
rect 7377 17731 7435 17737
rect 7377 17728 7389 17731
rect 7248 17700 7389 17728
rect 7248 17688 7254 17700
rect 7377 17697 7389 17700
rect 7423 17697 7435 17731
rect 7377 17691 7435 17697
rect 7644 17731 7702 17737
rect 7644 17697 7656 17731
rect 7690 17728 7702 17731
rect 8570 17728 8576 17740
rect 7690 17700 8576 17728
rect 7690 17697 7702 17700
rect 7644 17691 7702 17697
rect 8570 17688 8576 17700
rect 8628 17688 8634 17740
rect 8938 17688 8944 17740
rect 8996 17728 9002 17740
rect 11606 17728 11612 17740
rect 8996 17700 11612 17728
rect 8996 17688 9002 17700
rect 11606 17688 11612 17700
rect 11664 17688 11670 17740
rect 11977 17731 12035 17737
rect 11977 17697 11989 17731
rect 12023 17728 12035 17731
rect 12342 17728 12348 17740
rect 12023 17700 12348 17728
rect 12023 17697 12035 17700
rect 11977 17691 12035 17697
rect 12342 17688 12348 17700
rect 12400 17688 12406 17740
rect 12894 17688 12900 17740
rect 12952 17728 12958 17740
rect 13464 17728 13492 17768
rect 14093 17731 14151 17737
rect 14093 17728 14105 17731
rect 12952 17700 13492 17728
rect 14016 17700 14105 17728
rect 12952 17688 12958 17700
rect 2317 17663 2375 17669
rect 2317 17629 2329 17663
rect 2363 17660 2375 17663
rect 2406 17660 2412 17672
rect 2363 17632 2412 17660
rect 2363 17629 2375 17632
rect 2317 17623 2375 17629
rect 2406 17620 2412 17632
rect 2464 17620 2470 17672
rect 4065 17663 4123 17669
rect 4065 17629 4077 17663
rect 4111 17629 4123 17663
rect 4065 17623 4123 17629
rect 2038 17552 2044 17604
rect 2096 17592 2102 17604
rect 3970 17592 3976 17604
rect 2096 17564 3976 17592
rect 2096 17552 2102 17564
rect 3970 17552 3976 17564
rect 4028 17592 4034 17604
rect 4080 17592 4108 17623
rect 5534 17620 5540 17672
rect 5592 17660 5598 17672
rect 6273 17663 6331 17669
rect 6273 17660 6285 17663
rect 5592 17632 6285 17660
rect 5592 17620 5598 17632
rect 6273 17629 6285 17632
rect 6319 17629 6331 17663
rect 10594 17660 10600 17672
rect 10555 17632 10600 17660
rect 6273 17623 6331 17629
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 10962 17620 10968 17672
rect 11020 17660 11026 17672
rect 12161 17663 12219 17669
rect 12161 17660 12173 17663
rect 11020 17632 12173 17660
rect 11020 17620 11026 17632
rect 12161 17629 12173 17632
rect 12207 17629 12219 17663
rect 12360 17660 12388 17688
rect 14016 17672 14044 17700
rect 14093 17697 14105 17700
rect 14139 17697 14151 17731
rect 14200 17728 14228 17768
rect 16482 17756 16488 17768
rect 16540 17756 16546 17808
rect 16666 17756 16672 17808
rect 16724 17796 16730 17808
rect 20254 17796 20260 17808
rect 16724 17768 20260 17796
rect 16724 17756 16730 17768
rect 20254 17756 20260 17768
rect 20312 17756 20318 17808
rect 15378 17728 15384 17740
rect 14200 17700 15384 17728
rect 14093 17691 14151 17697
rect 15378 17688 15384 17700
rect 15436 17728 15442 17740
rect 15657 17731 15715 17737
rect 15657 17728 15669 17731
rect 15436 17700 15669 17728
rect 15436 17688 15442 17700
rect 15657 17697 15669 17700
rect 15703 17697 15715 17731
rect 15657 17691 15715 17697
rect 15746 17688 15752 17740
rect 15804 17728 15810 17740
rect 15804 17700 15849 17728
rect 15804 17688 15810 17700
rect 16022 17688 16028 17740
rect 16080 17728 16086 17740
rect 17221 17731 17279 17737
rect 17221 17728 17233 17731
rect 16080 17700 17233 17728
rect 16080 17688 16086 17700
rect 17221 17697 17233 17700
rect 17267 17697 17279 17731
rect 17221 17691 17279 17697
rect 18506 17688 18512 17740
rect 18564 17728 18570 17740
rect 18877 17731 18935 17737
rect 18877 17728 18889 17731
rect 18564 17700 18889 17728
rect 18564 17688 18570 17700
rect 18877 17697 18889 17700
rect 18923 17728 18935 17731
rect 19886 17728 19892 17740
rect 18923 17700 19892 17728
rect 18923 17697 18935 17700
rect 18877 17691 18935 17697
rect 19886 17688 19892 17700
rect 19944 17688 19950 17740
rect 13814 17660 13820 17672
rect 12360 17632 13820 17660
rect 12161 17623 12219 17629
rect 13814 17620 13820 17632
rect 13872 17620 13878 17672
rect 13998 17620 14004 17672
rect 14056 17620 14062 17672
rect 14274 17620 14280 17672
rect 14332 17660 14338 17672
rect 14332 17632 15516 17660
rect 14332 17620 14338 17632
rect 15488 17592 15516 17632
rect 15838 17620 15844 17672
rect 15896 17660 15902 17672
rect 16390 17660 16396 17672
rect 15896 17632 16396 17660
rect 15896 17620 15902 17632
rect 16390 17620 16396 17632
rect 16448 17620 16454 17672
rect 17310 17660 17316 17672
rect 17271 17632 17316 17660
rect 17310 17620 17316 17632
rect 17368 17620 17374 17672
rect 17497 17663 17555 17669
rect 17497 17629 17509 17663
rect 17543 17660 17555 17663
rect 18230 17660 18236 17672
rect 17543 17632 18236 17660
rect 17543 17629 17555 17632
rect 17497 17623 17555 17629
rect 18230 17620 18236 17632
rect 18288 17660 18294 17672
rect 19061 17663 19119 17669
rect 18288 17632 18552 17660
rect 18288 17620 18294 17632
rect 18417 17595 18475 17601
rect 18417 17592 18429 17595
rect 4028 17564 4108 17592
rect 5368 17564 5672 17592
rect 4028 17552 4034 17564
rect 2406 17484 2412 17536
rect 2464 17524 2470 17536
rect 5368 17524 5396 17564
rect 2464 17496 5396 17524
rect 2464 17484 2470 17496
rect 5442 17484 5448 17536
rect 5500 17524 5506 17536
rect 5644 17524 5672 17564
rect 8312 17564 15240 17592
rect 15488 17564 18429 17592
rect 8312 17524 8340 17564
rect 5500 17496 5545 17524
rect 5644 17496 8340 17524
rect 8757 17527 8815 17533
rect 5500 17484 5506 17496
rect 8757 17493 8769 17527
rect 8803 17524 8815 17527
rect 10962 17524 10968 17536
rect 8803 17496 10968 17524
rect 8803 17493 8815 17496
rect 8757 17487 8815 17493
rect 10962 17484 10968 17496
rect 11020 17484 11026 17536
rect 11238 17484 11244 17536
rect 11296 17524 11302 17536
rect 11609 17527 11667 17533
rect 11609 17524 11621 17527
rect 11296 17496 11621 17524
rect 11296 17484 11302 17496
rect 11609 17493 11621 17496
rect 11655 17493 11667 17527
rect 11609 17487 11667 17493
rect 11698 17484 11704 17536
rect 11756 17524 11762 17536
rect 13078 17524 13084 17536
rect 11756 17496 13084 17524
rect 11756 17484 11762 17496
rect 13078 17484 13084 17496
rect 13136 17484 13142 17536
rect 15212 17524 15240 17564
rect 18417 17561 18429 17564
rect 18463 17561 18475 17595
rect 18524 17592 18552 17632
rect 19061 17629 19073 17663
rect 19107 17660 19119 17663
rect 19242 17660 19248 17672
rect 19107 17632 19248 17660
rect 19107 17629 19119 17632
rect 19061 17623 19119 17629
rect 19242 17620 19248 17632
rect 19300 17620 19306 17672
rect 20806 17592 20812 17604
rect 18524 17564 20812 17592
rect 18417 17555 18475 17561
rect 20806 17552 20812 17564
rect 20864 17552 20870 17604
rect 16206 17524 16212 17536
rect 15212 17496 16212 17524
rect 16206 17484 16212 17496
rect 16264 17484 16270 17536
rect 16853 17527 16911 17533
rect 16853 17493 16865 17527
rect 16899 17524 16911 17527
rect 17126 17524 17132 17536
rect 16899 17496 17132 17524
rect 16899 17493 16911 17496
rect 16853 17487 16911 17493
rect 17126 17484 17132 17496
rect 17184 17484 17190 17536
rect 17218 17484 17224 17536
rect 17276 17524 17282 17536
rect 18233 17527 18291 17533
rect 18233 17524 18245 17527
rect 17276 17496 18245 17524
rect 17276 17484 17282 17496
rect 18233 17493 18245 17496
rect 18279 17524 18291 17527
rect 19058 17524 19064 17536
rect 18279 17496 19064 17524
rect 18279 17493 18291 17496
rect 18233 17487 18291 17493
rect 19058 17484 19064 17496
rect 19116 17524 19122 17536
rect 19245 17527 19303 17533
rect 19245 17524 19257 17527
rect 19116 17496 19257 17524
rect 19116 17484 19122 17496
rect 19245 17493 19257 17496
rect 19291 17493 19303 17527
rect 19245 17487 19303 17493
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 3326 17280 3332 17332
rect 3384 17320 3390 17332
rect 3384 17292 4292 17320
rect 3384 17280 3390 17292
rect 3605 17255 3663 17261
rect 3605 17221 3617 17255
rect 3651 17221 3663 17255
rect 4264 17252 4292 17292
rect 4338 17280 4344 17332
rect 4396 17320 4402 17332
rect 4433 17323 4491 17329
rect 4433 17320 4445 17323
rect 4396 17292 4445 17320
rect 4396 17280 4402 17292
rect 4433 17289 4445 17292
rect 4479 17289 4491 17323
rect 4433 17283 4491 17289
rect 4982 17280 4988 17332
rect 5040 17320 5046 17332
rect 5166 17320 5172 17332
rect 5040 17292 5172 17320
rect 5040 17280 5046 17292
rect 5166 17280 5172 17292
rect 5224 17280 5230 17332
rect 14274 17320 14280 17332
rect 6472 17292 14280 17320
rect 6472 17252 6500 17292
rect 14274 17280 14280 17292
rect 14332 17280 14338 17332
rect 15304 17292 20024 17320
rect 7650 17252 7656 17264
rect 4264 17224 6500 17252
rect 7611 17224 7656 17252
rect 3605 17215 3663 17221
rect 3620 17184 3648 17215
rect 7650 17212 7656 17224
rect 7708 17212 7714 17264
rect 10134 17252 10140 17264
rect 7760 17224 10140 17252
rect 4798 17184 4804 17196
rect 3620 17156 4804 17184
rect 4798 17144 4804 17156
rect 4856 17144 4862 17196
rect 5077 17187 5135 17193
rect 5077 17153 5089 17187
rect 5123 17184 5135 17187
rect 5442 17184 5448 17196
rect 5123 17156 5448 17184
rect 5123 17153 5135 17156
rect 5077 17147 5135 17153
rect 5442 17144 5448 17156
rect 5500 17144 5506 17196
rect 5718 17144 5724 17196
rect 5776 17184 5782 17196
rect 7760 17184 7788 17224
rect 10134 17212 10140 17224
rect 10192 17212 10198 17264
rect 10229 17255 10287 17261
rect 10229 17221 10241 17255
rect 10275 17252 10287 17255
rect 12434 17252 12440 17264
rect 10275 17224 12440 17252
rect 10275 17221 10287 17224
rect 10229 17215 10287 17221
rect 12434 17212 12440 17224
rect 12492 17212 12498 17264
rect 12526 17212 12532 17264
rect 12584 17252 12590 17264
rect 15304 17252 15332 17292
rect 12584 17224 15332 17252
rect 12584 17212 12590 17224
rect 17586 17212 17592 17264
rect 17644 17252 17650 17264
rect 18049 17255 18107 17261
rect 18049 17252 18061 17255
rect 17644 17224 18061 17252
rect 17644 17212 17650 17224
rect 18049 17221 18061 17224
rect 18095 17221 18107 17255
rect 18049 17215 18107 17221
rect 18414 17212 18420 17264
rect 18472 17252 18478 17264
rect 18472 17224 18644 17252
rect 18472 17212 18478 17224
rect 5776 17156 7788 17184
rect 8205 17187 8263 17193
rect 5776 17144 5782 17156
rect 8205 17153 8217 17187
rect 8251 17184 8263 17187
rect 8570 17184 8576 17196
rect 8251 17156 8576 17184
rect 8251 17153 8263 17156
rect 8205 17147 8263 17153
rect 8570 17144 8576 17156
rect 8628 17144 8634 17196
rect 10778 17184 10784 17196
rect 8680 17156 10784 17184
rect 2038 17076 2044 17128
rect 2096 17116 2102 17128
rect 2498 17125 2504 17128
rect 2225 17119 2283 17125
rect 2225 17116 2237 17119
rect 2096 17088 2237 17116
rect 2096 17076 2102 17088
rect 2225 17085 2237 17088
rect 2271 17085 2283 17119
rect 2492 17116 2504 17125
rect 2459 17088 2504 17116
rect 2225 17079 2283 17085
rect 2492 17079 2504 17088
rect 2498 17076 2504 17079
rect 2556 17076 2562 17128
rect 4893 17119 4951 17125
rect 4893 17085 4905 17119
rect 4939 17116 4951 17119
rect 5350 17116 5356 17128
rect 4939 17088 5356 17116
rect 4939 17085 4951 17088
rect 4893 17079 4951 17085
rect 5350 17076 5356 17088
rect 5408 17076 5414 17128
rect 6546 17116 6552 17128
rect 6288 17088 6552 17116
rect 6288 17048 6316 17088
rect 6546 17076 6552 17088
rect 6604 17076 6610 17128
rect 7006 17076 7012 17128
rect 7064 17116 7070 17128
rect 7374 17116 7380 17128
rect 7064 17088 7380 17116
rect 7064 17076 7070 17088
rect 7374 17076 7380 17088
rect 7432 17076 7438 17128
rect 8680 17116 8708 17156
rect 10778 17144 10784 17156
rect 10836 17144 10842 17196
rect 10873 17187 10931 17193
rect 10873 17153 10885 17187
rect 10919 17184 10931 17187
rect 10962 17184 10968 17196
rect 10919 17156 10968 17184
rect 10919 17153 10931 17156
rect 10873 17147 10931 17153
rect 10962 17144 10968 17156
rect 11020 17144 11026 17196
rect 12986 17144 12992 17196
rect 13044 17184 13050 17196
rect 14277 17187 14335 17193
rect 14277 17184 14289 17187
rect 13044 17156 14289 17184
rect 13044 17144 13050 17156
rect 14277 17153 14289 17156
rect 14323 17184 14335 17187
rect 14734 17184 14740 17196
rect 14323 17156 14740 17184
rect 14323 17153 14335 17156
rect 14277 17147 14335 17153
rect 14734 17144 14740 17156
rect 14792 17144 14798 17196
rect 17310 17144 17316 17196
rect 17368 17184 17374 17196
rect 18506 17184 18512 17196
rect 17368 17156 18512 17184
rect 17368 17144 17374 17156
rect 18506 17144 18512 17156
rect 18564 17144 18570 17196
rect 18616 17193 18644 17224
rect 18601 17187 18659 17193
rect 18601 17153 18613 17187
rect 18647 17153 18659 17187
rect 18601 17147 18659 17153
rect 10594 17116 10600 17128
rect 7944 17088 8708 17116
rect 10555 17088 10600 17116
rect 4816 17020 6316 17048
rect 2498 16940 2504 16992
rect 2556 16980 2562 16992
rect 4816 16989 4844 17020
rect 4801 16983 4859 16989
rect 4801 16980 4813 16983
rect 2556 16952 4813 16980
rect 2556 16940 2562 16952
rect 4801 16949 4813 16952
rect 4847 16949 4859 16983
rect 4801 16943 4859 16949
rect 4982 16940 4988 16992
rect 5040 16980 5046 16992
rect 7944 16980 7972 17088
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 11698 17076 11704 17128
rect 11756 17116 11762 17128
rect 13906 17116 13912 17128
rect 11756 17088 13912 17116
rect 11756 17076 11762 17088
rect 13906 17076 13912 17088
rect 13964 17116 13970 17128
rect 14093 17119 14151 17125
rect 14093 17116 14105 17119
rect 13964 17088 14105 17116
rect 13964 17076 13970 17088
rect 14093 17085 14105 17088
rect 14139 17085 14151 17119
rect 14093 17079 14151 17085
rect 14185 17119 14243 17125
rect 14185 17085 14197 17119
rect 14231 17116 14243 17119
rect 15102 17116 15108 17128
rect 14231 17088 15108 17116
rect 14231 17085 14243 17088
rect 14185 17079 14243 17085
rect 15102 17076 15108 17088
rect 15160 17076 15166 17128
rect 15286 17116 15292 17128
rect 15247 17088 15292 17116
rect 15286 17076 15292 17088
rect 15344 17076 15350 17128
rect 19702 17116 19708 17128
rect 15396 17088 19708 17116
rect 8021 17051 8079 17057
rect 8021 17017 8033 17051
rect 8067 17048 8079 17051
rect 8202 17048 8208 17060
rect 8067 17020 8208 17048
rect 8067 17017 8079 17020
rect 8021 17011 8079 17017
rect 8202 17008 8208 17020
rect 8260 17008 8266 17060
rect 9030 17008 9036 17060
rect 9088 17048 9094 17060
rect 9088 17020 10824 17048
rect 9088 17008 9094 17020
rect 5040 16952 7972 16980
rect 8113 16983 8171 16989
rect 5040 16940 5046 16952
rect 8113 16949 8125 16983
rect 8159 16980 8171 16983
rect 8570 16980 8576 16992
rect 8159 16952 8576 16980
rect 8159 16949 8171 16952
rect 8113 16943 8171 16949
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 9122 16940 9128 16992
rect 9180 16980 9186 16992
rect 9217 16983 9275 16989
rect 9217 16980 9229 16983
rect 9180 16952 9229 16980
rect 9180 16940 9186 16952
rect 9217 16949 9229 16952
rect 9263 16949 9275 16983
rect 9217 16943 9275 16949
rect 9950 16940 9956 16992
rect 10008 16980 10014 16992
rect 10689 16983 10747 16989
rect 10689 16980 10701 16983
rect 10008 16952 10701 16980
rect 10008 16940 10014 16952
rect 10689 16949 10701 16952
rect 10735 16949 10747 16983
rect 10796 16980 10824 17020
rect 12526 17008 12532 17060
rect 12584 17048 12590 17060
rect 15396 17048 15424 17088
rect 19702 17076 19708 17088
rect 19760 17076 19766 17128
rect 19996 17125 20024 17292
rect 20165 17187 20223 17193
rect 20165 17153 20177 17187
rect 20211 17153 20223 17187
rect 20165 17147 20223 17153
rect 19981 17119 20039 17125
rect 19981 17085 19993 17119
rect 20027 17085 20039 17119
rect 19981 17079 20039 17085
rect 12584 17020 15424 17048
rect 15545 17051 15603 17057
rect 12584 17008 12590 17020
rect 15545 17017 15557 17051
rect 15591 17017 15603 17051
rect 15545 17011 15603 17017
rect 12342 16980 12348 16992
rect 10796 16952 12348 16980
rect 10689 16943 10747 16949
rect 12342 16940 12348 16952
rect 12400 16940 12406 16992
rect 12437 16983 12495 16989
rect 12437 16949 12449 16983
rect 12483 16980 12495 16983
rect 12618 16980 12624 16992
rect 12483 16952 12624 16980
rect 12483 16949 12495 16952
rect 12437 16943 12495 16949
rect 12618 16940 12624 16952
rect 12676 16940 12682 16992
rect 12894 16940 12900 16992
rect 12952 16980 12958 16992
rect 13725 16983 13783 16989
rect 13725 16980 13737 16983
rect 12952 16952 13737 16980
rect 12952 16940 12958 16952
rect 13725 16949 13737 16952
rect 13771 16949 13783 16983
rect 13725 16943 13783 16949
rect 14734 16940 14740 16992
rect 14792 16980 14798 16992
rect 15549 16980 15577 17011
rect 15654 17008 15660 17060
rect 15712 17048 15718 17060
rect 20180 17048 20208 17147
rect 15712 17020 20208 17048
rect 15712 17008 15718 17020
rect 14792 16952 15577 16980
rect 14792 16940 14798 16952
rect 16114 16940 16120 16992
rect 16172 16980 16178 16992
rect 16669 16983 16727 16989
rect 16669 16980 16681 16983
rect 16172 16952 16681 16980
rect 16172 16940 16178 16952
rect 16669 16949 16681 16952
rect 16715 16949 16727 16983
rect 16669 16943 16727 16949
rect 18417 16983 18475 16989
rect 18417 16949 18429 16983
rect 18463 16980 18475 16983
rect 19058 16980 19064 16992
rect 18463 16952 19064 16980
rect 18463 16949 18475 16952
rect 18417 16943 18475 16949
rect 19058 16940 19064 16952
rect 19116 16940 19122 16992
rect 19613 16983 19671 16989
rect 19613 16949 19625 16983
rect 19659 16980 19671 16983
rect 19794 16980 19800 16992
rect 19659 16952 19800 16980
rect 19659 16949 19671 16952
rect 19613 16943 19671 16949
rect 19794 16940 19800 16952
rect 19852 16940 19858 16992
rect 20070 16940 20076 16992
rect 20128 16980 20134 16992
rect 20128 16952 20173 16980
rect 20128 16940 20134 16952
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 4338 16736 4344 16788
rect 4396 16776 4402 16788
rect 4525 16779 4583 16785
rect 4525 16776 4537 16779
rect 4396 16748 4537 16776
rect 4396 16736 4402 16748
rect 4525 16745 4537 16748
rect 4571 16745 4583 16779
rect 4525 16739 4583 16745
rect 5074 16736 5080 16788
rect 5132 16776 5138 16788
rect 5718 16776 5724 16788
rect 5132 16748 5724 16776
rect 5132 16736 5138 16748
rect 2317 16711 2375 16717
rect 2317 16677 2329 16711
rect 2363 16708 2375 16711
rect 4433 16711 4491 16717
rect 2363 16680 4384 16708
rect 2363 16677 2375 16680
rect 2317 16671 2375 16677
rect 2041 16643 2099 16649
rect 2041 16609 2053 16643
rect 2087 16640 2099 16643
rect 4154 16640 4160 16652
rect 2087 16612 4160 16640
rect 2087 16609 2099 16612
rect 2041 16603 2099 16609
rect 4154 16600 4160 16612
rect 4212 16600 4218 16652
rect 4356 16640 4384 16680
rect 4433 16677 4445 16711
rect 4479 16708 4491 16711
rect 5276 16708 5304 16748
rect 5718 16736 5724 16748
rect 5776 16736 5782 16788
rect 7650 16736 7656 16788
rect 7708 16776 7714 16788
rect 7708 16748 7779 16776
rect 7708 16736 7714 16748
rect 4479 16680 5304 16708
rect 6365 16711 6423 16717
rect 4479 16677 4491 16680
rect 4433 16671 4491 16677
rect 6365 16677 6377 16711
rect 6411 16708 6423 16711
rect 7558 16708 7564 16720
rect 6411 16680 7564 16708
rect 6411 16677 6423 16680
rect 6365 16671 6423 16677
rect 7558 16668 7564 16680
rect 7616 16668 7622 16720
rect 7006 16640 7012 16652
rect 4356 16612 7012 16640
rect 7006 16600 7012 16612
rect 7064 16600 7070 16652
rect 7190 16600 7196 16652
rect 7248 16640 7254 16652
rect 7377 16643 7435 16649
rect 7377 16640 7389 16643
rect 7248 16612 7389 16640
rect 7248 16600 7254 16612
rect 7377 16609 7389 16612
rect 7423 16609 7435 16643
rect 7377 16603 7435 16609
rect 7644 16643 7702 16649
rect 7644 16609 7656 16643
rect 7690 16640 7702 16643
rect 7751 16640 7779 16748
rect 8570 16736 8576 16788
rect 8628 16776 8634 16788
rect 10137 16779 10195 16785
rect 10137 16776 10149 16779
rect 8628 16748 10149 16776
rect 8628 16736 8634 16748
rect 10137 16745 10149 16748
rect 10183 16745 10195 16779
rect 10137 16739 10195 16745
rect 11790 16736 11796 16788
rect 11848 16776 11854 16788
rect 12253 16779 12311 16785
rect 12253 16776 12265 16779
rect 11848 16748 12265 16776
rect 11848 16736 11854 16748
rect 12253 16745 12265 16748
rect 12299 16745 12311 16779
rect 12253 16739 12311 16745
rect 12342 16736 12348 16788
rect 12400 16776 12406 16788
rect 20070 16776 20076 16788
rect 12400 16748 20076 16776
rect 12400 16736 12406 16748
rect 20070 16736 20076 16748
rect 20128 16736 20134 16788
rect 7926 16668 7932 16720
rect 7984 16708 7990 16720
rect 12434 16708 12440 16720
rect 7984 16680 12440 16708
rect 7984 16668 7990 16680
rect 12434 16668 12440 16680
rect 12492 16668 12498 16720
rect 16114 16717 16120 16720
rect 13633 16711 13691 16717
rect 13633 16708 13645 16711
rect 12544 16680 13645 16708
rect 7690 16612 7779 16640
rect 7690 16609 7702 16612
rect 7644 16603 7702 16609
rect 8018 16600 8024 16652
rect 8076 16640 8082 16652
rect 8076 16612 8432 16640
rect 8076 16600 8082 16612
rect 3510 16532 3516 16584
rect 3568 16532 3574 16584
rect 4709 16575 4767 16581
rect 4709 16541 4721 16575
rect 4755 16572 4767 16575
rect 4982 16572 4988 16584
rect 4755 16544 4988 16572
rect 4755 16541 4767 16544
rect 4709 16535 4767 16541
rect 4982 16532 4988 16544
rect 5040 16532 5046 16584
rect 8404 16572 8432 16612
rect 8570 16600 8576 16652
rect 8628 16640 8634 16652
rect 9858 16640 9864 16652
rect 8628 16612 9864 16640
rect 8628 16600 8634 16612
rect 9858 16600 9864 16612
rect 9916 16600 9922 16652
rect 10505 16643 10563 16649
rect 10505 16609 10517 16643
rect 10551 16640 10563 16643
rect 10778 16640 10784 16652
rect 10551 16612 10784 16640
rect 10551 16609 10563 16612
rect 10505 16603 10563 16609
rect 10778 16600 10784 16612
rect 10836 16640 10842 16652
rect 11054 16640 11060 16652
rect 10836 16612 11060 16640
rect 10836 16600 10842 16612
rect 11054 16600 11060 16612
rect 11112 16600 11118 16652
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 12544 16640 12572 16680
rect 13633 16677 13645 16680
rect 13679 16708 13691 16711
rect 13817 16711 13875 16717
rect 13817 16708 13829 16711
rect 13679 16680 13829 16708
rect 13679 16677 13691 16680
rect 13633 16671 13691 16677
rect 13817 16677 13829 16680
rect 13863 16677 13875 16711
rect 16108 16708 16120 16717
rect 16075 16680 16120 16708
rect 13817 16671 13875 16677
rect 16108 16671 16120 16680
rect 16114 16668 16120 16671
rect 16172 16668 16178 16720
rect 16206 16668 16212 16720
rect 16264 16708 16270 16720
rect 16264 16680 18092 16708
rect 16264 16668 16270 16680
rect 11756 16612 12572 16640
rect 12621 16643 12679 16649
rect 11756 16600 11762 16612
rect 12621 16609 12633 16643
rect 12667 16640 12679 16643
rect 13078 16640 13084 16652
rect 12667 16612 13084 16640
rect 12667 16609 12679 16612
rect 12621 16603 12679 16609
rect 9766 16572 9772 16584
rect 8404 16544 9772 16572
rect 9766 16532 9772 16544
rect 9824 16532 9830 16584
rect 10594 16572 10600 16584
rect 10555 16544 10600 16572
rect 10594 16532 10600 16544
rect 10652 16532 10658 16584
rect 10689 16575 10747 16581
rect 10689 16541 10701 16575
rect 10735 16541 10747 16575
rect 10689 16535 10747 16541
rect 3528 16504 3556 16532
rect 7374 16504 7380 16516
rect 3528 16476 4752 16504
rect 2958 16396 2964 16448
rect 3016 16436 3022 16448
rect 3510 16436 3516 16448
rect 3016 16408 3516 16436
rect 3016 16396 3022 16408
rect 3510 16396 3516 16408
rect 3568 16396 3574 16448
rect 4062 16436 4068 16448
rect 4023 16408 4068 16436
rect 4062 16396 4068 16408
rect 4120 16396 4126 16448
rect 4724 16436 4752 16476
rect 7208 16476 7380 16504
rect 7208 16436 7236 16476
rect 7374 16464 7380 16476
rect 7432 16464 7438 16516
rect 10704 16504 10732 16535
rect 10870 16532 10876 16584
rect 10928 16572 10934 16584
rect 12636 16572 12664 16603
rect 13078 16600 13084 16612
rect 13136 16600 13142 16652
rect 13998 16600 14004 16652
rect 14056 16640 14062 16652
rect 18064 16640 18092 16680
rect 18138 16668 18144 16720
rect 18196 16708 18202 16720
rect 18417 16711 18475 16717
rect 18417 16708 18429 16711
rect 18196 16680 18429 16708
rect 18196 16668 18202 16680
rect 18417 16677 18429 16680
rect 18463 16677 18475 16711
rect 18417 16671 18475 16677
rect 18509 16711 18567 16717
rect 18509 16677 18521 16711
rect 18555 16708 18567 16711
rect 18598 16708 18604 16720
rect 18555 16680 18604 16708
rect 18555 16677 18567 16680
rect 18509 16671 18567 16677
rect 18598 16668 18604 16680
rect 18656 16668 18662 16720
rect 19613 16643 19671 16649
rect 19613 16640 19625 16643
rect 14056 16612 18000 16640
rect 18064 16612 19625 16640
rect 14056 16600 14062 16612
rect 10928 16544 12664 16572
rect 12713 16575 12771 16581
rect 10928 16532 10934 16544
rect 12713 16541 12725 16575
rect 12759 16541 12771 16575
rect 12713 16535 12771 16541
rect 12897 16575 12955 16581
rect 12897 16541 12909 16575
rect 12943 16572 12955 16575
rect 13170 16572 13176 16584
rect 12943 16544 13176 16572
rect 12943 16541 12955 16544
rect 12897 16535 12955 16541
rect 8588 16476 10732 16504
rect 4724 16408 7236 16436
rect 7282 16396 7288 16448
rect 7340 16436 7346 16448
rect 8588 16436 8616 16476
rect 12342 16464 12348 16516
rect 12400 16504 12406 16516
rect 12728 16504 12756 16535
rect 13170 16532 13176 16544
rect 13228 16532 13234 16584
rect 13262 16532 13268 16584
rect 13320 16572 13326 16584
rect 13630 16572 13636 16584
rect 13320 16544 13636 16572
rect 13320 16532 13326 16544
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 15286 16532 15292 16584
rect 15344 16572 15350 16584
rect 15470 16572 15476 16584
rect 15344 16544 15476 16572
rect 15344 16532 15350 16544
rect 15470 16532 15476 16544
rect 15528 16572 15534 16584
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 15528 16544 15853 16572
rect 15528 16532 15534 16544
rect 15841 16541 15853 16544
rect 15887 16541 15899 16575
rect 17972 16572 18000 16612
rect 19613 16609 19625 16612
rect 19659 16609 19671 16643
rect 19613 16603 19671 16609
rect 17972 16544 18092 16572
rect 15841 16535 15899 16541
rect 13354 16504 13360 16516
rect 12400 16476 13360 16504
rect 12400 16464 12406 16476
rect 13354 16464 13360 16476
rect 13412 16464 13418 16516
rect 18064 16513 18092 16544
rect 18138 16532 18144 16584
rect 18196 16572 18202 16584
rect 18601 16575 18659 16581
rect 18601 16572 18613 16575
rect 18196 16544 18613 16572
rect 18196 16532 18202 16544
rect 18601 16541 18613 16544
rect 18647 16541 18659 16575
rect 18601 16535 18659 16541
rect 18049 16507 18107 16513
rect 17144 16476 18000 16504
rect 7340 16408 8616 16436
rect 7340 16396 7346 16408
rect 8662 16396 8668 16448
rect 8720 16436 8726 16448
rect 8757 16439 8815 16445
rect 8757 16436 8769 16439
rect 8720 16408 8769 16436
rect 8720 16396 8726 16408
rect 8757 16405 8769 16408
rect 8803 16405 8815 16439
rect 8757 16399 8815 16405
rect 8846 16396 8852 16448
rect 8904 16436 8910 16448
rect 12526 16436 12532 16448
rect 8904 16408 12532 16436
rect 8904 16396 8910 16408
rect 12526 16396 12532 16408
rect 12584 16396 12590 16448
rect 13170 16396 13176 16448
rect 13228 16436 13234 16448
rect 15838 16436 15844 16448
rect 13228 16408 15844 16436
rect 13228 16396 13234 16408
rect 15838 16396 15844 16408
rect 15896 16436 15902 16448
rect 16022 16436 16028 16448
rect 15896 16408 16028 16436
rect 15896 16396 15902 16408
rect 16022 16396 16028 16408
rect 16080 16436 16086 16448
rect 17144 16436 17172 16476
rect 16080 16408 17172 16436
rect 17221 16439 17279 16445
rect 16080 16396 16086 16408
rect 17221 16405 17233 16439
rect 17267 16436 17279 16439
rect 17310 16436 17316 16448
rect 17267 16408 17316 16436
rect 17267 16405 17279 16408
rect 17221 16399 17279 16405
rect 17310 16396 17316 16408
rect 17368 16396 17374 16448
rect 17972 16436 18000 16476
rect 18049 16473 18061 16507
rect 18095 16473 18107 16507
rect 18049 16467 18107 16473
rect 18414 16464 18420 16516
rect 18472 16464 18478 16516
rect 19702 16464 19708 16516
rect 19760 16504 19766 16516
rect 19797 16507 19855 16513
rect 19797 16504 19809 16507
rect 19760 16476 19809 16504
rect 19760 16464 19766 16476
rect 19797 16473 19809 16476
rect 19843 16473 19855 16507
rect 19797 16467 19855 16473
rect 18432 16436 18460 16464
rect 19334 16436 19340 16448
rect 17972 16408 19340 16436
rect 19334 16396 19340 16408
rect 19392 16396 19398 16448
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 4154 16192 4160 16244
rect 4212 16232 4218 16244
rect 4709 16235 4767 16241
rect 4709 16232 4721 16235
rect 4212 16204 4721 16232
rect 4212 16192 4218 16204
rect 4709 16201 4721 16204
rect 4755 16201 4767 16235
rect 9766 16232 9772 16244
rect 4709 16195 4767 16201
rect 4816 16204 9772 16232
rect 3436 16136 3924 16164
rect 2406 16096 2412 16108
rect 2367 16068 2412 16096
rect 2406 16056 2412 16068
rect 2464 16056 2470 16108
rect 2133 16031 2191 16037
rect 2133 15997 2145 16031
rect 2179 16028 2191 16031
rect 3050 16028 3056 16040
rect 2179 16000 3056 16028
rect 2179 15997 2191 16000
rect 2133 15991 2191 15997
rect 3050 15988 3056 16000
rect 3108 15988 3114 16040
rect 3436 16037 3464 16136
rect 3421 16031 3479 16037
rect 3421 15997 3433 16031
rect 3467 15997 3479 16031
rect 3896 16028 3924 16136
rect 3970 16124 3976 16176
rect 4028 16164 4034 16176
rect 4816 16164 4844 16204
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 9858 16192 9864 16244
rect 9916 16232 9922 16244
rect 9916 16204 16804 16232
rect 9916 16192 9922 16204
rect 4028 16136 4844 16164
rect 4028 16124 4034 16136
rect 7190 16124 7196 16176
rect 7248 16164 7254 16176
rect 7742 16164 7748 16176
rect 7248 16136 7748 16164
rect 7248 16124 7254 16136
rect 7742 16124 7748 16136
rect 7800 16164 7806 16176
rect 10781 16167 10839 16173
rect 7800 16136 8616 16164
rect 7800 16124 7806 16136
rect 5350 16096 5356 16108
rect 5311 16068 5356 16096
rect 5350 16056 5356 16068
rect 5408 16096 5414 16108
rect 5994 16096 6000 16108
rect 5408 16068 6000 16096
rect 5408 16056 5414 16068
rect 5994 16056 6000 16068
rect 6052 16056 6058 16108
rect 7653 16099 7711 16105
rect 7300 16068 7604 16096
rect 7300 16028 7328 16068
rect 3896 16000 7328 16028
rect 3421 15991 3479 15997
rect 7374 15988 7380 16040
rect 7432 16028 7438 16040
rect 7469 16031 7527 16037
rect 7469 16028 7481 16031
rect 7432 16000 7481 16028
rect 7432 15988 7438 16000
rect 7469 15997 7481 16000
rect 7515 15997 7527 16031
rect 7576 16028 7604 16068
rect 7653 16065 7665 16099
rect 7699 16096 7711 16099
rect 8294 16096 8300 16108
rect 7699 16068 8300 16096
rect 7699 16065 7711 16068
rect 7653 16059 7711 16065
rect 8294 16056 8300 16068
rect 8352 16056 8358 16108
rect 8588 16105 8616 16136
rect 10781 16133 10793 16167
rect 10827 16164 10839 16167
rect 12710 16164 12716 16176
rect 10827 16136 12716 16164
rect 10827 16133 10839 16136
rect 10781 16127 10839 16133
rect 12710 16124 12716 16136
rect 12768 16124 12774 16176
rect 16574 16164 16580 16176
rect 13832 16136 16580 16164
rect 8573 16099 8631 16105
rect 8573 16065 8585 16099
rect 8619 16065 8631 16099
rect 11330 16096 11336 16108
rect 11291 16068 11336 16096
rect 8573 16059 8631 16065
rect 11330 16056 11336 16068
rect 11388 16056 11394 16108
rect 8018 16028 8024 16040
rect 7576 16000 8024 16028
rect 7469 15991 7527 15997
rect 8018 15988 8024 16000
rect 8076 15988 8082 16040
rect 10410 15988 10416 16040
rect 10468 16028 10474 16040
rect 10594 16028 10600 16040
rect 10468 16000 10600 16028
rect 10468 15988 10474 16000
rect 10594 15988 10600 16000
rect 10652 15988 10658 16040
rect 12710 15988 12716 16040
rect 12768 16028 12774 16040
rect 12805 16031 12863 16037
rect 12805 16028 12817 16031
rect 12768 16000 12817 16028
rect 12768 15988 12774 16000
rect 12805 15997 12817 16000
rect 12851 15997 12863 16031
rect 13832 16028 13860 16136
rect 16574 16124 16580 16136
rect 16632 16124 16638 16176
rect 15470 16056 15476 16108
rect 15528 16096 15534 16108
rect 15657 16099 15715 16105
rect 15528 16068 15599 16096
rect 15528 16056 15534 16068
rect 12805 15991 12863 15997
rect 13004 16000 13860 16028
rect 3694 15960 3700 15972
rect 3655 15932 3700 15960
rect 3694 15920 3700 15932
rect 3752 15920 3758 15972
rect 4430 15920 4436 15972
rect 4488 15960 4494 15972
rect 5077 15963 5135 15969
rect 5077 15960 5089 15963
rect 4488 15932 5089 15960
rect 4488 15920 4494 15932
rect 5077 15929 5089 15932
rect 5123 15929 5135 15963
rect 5077 15923 5135 15929
rect 5169 15963 5227 15969
rect 5169 15929 5181 15963
rect 5215 15960 5227 15963
rect 5215 15932 7779 15960
rect 5215 15929 5227 15932
rect 5169 15923 5227 15929
rect 5994 15852 6000 15904
rect 6052 15892 6058 15904
rect 7009 15895 7067 15901
rect 7009 15892 7021 15895
rect 6052 15864 7021 15892
rect 6052 15852 6058 15864
rect 7009 15861 7021 15864
rect 7055 15861 7067 15895
rect 7009 15855 7067 15861
rect 7377 15895 7435 15901
rect 7377 15861 7389 15895
rect 7423 15892 7435 15895
rect 7650 15892 7656 15904
rect 7423 15864 7656 15892
rect 7423 15861 7435 15864
rect 7377 15855 7435 15861
rect 7650 15852 7656 15864
rect 7708 15852 7714 15904
rect 7751 15892 7779 15932
rect 8662 15920 8668 15972
rect 8720 15960 8726 15972
rect 8818 15963 8876 15969
rect 8818 15960 8830 15963
rect 8720 15932 8830 15960
rect 8720 15920 8726 15932
rect 8818 15929 8830 15932
rect 8864 15929 8876 15963
rect 8818 15923 8876 15929
rect 9122 15920 9128 15972
rect 9180 15960 9186 15972
rect 11149 15963 11207 15969
rect 11149 15960 11161 15963
rect 9180 15932 11161 15960
rect 9180 15920 9186 15932
rect 11149 15929 11161 15932
rect 11195 15929 11207 15963
rect 11149 15923 11207 15929
rect 11241 15963 11299 15969
rect 11241 15929 11253 15963
rect 11287 15960 11299 15963
rect 13004 15960 13032 16000
rect 11287 15932 13032 15960
rect 13072 15963 13130 15969
rect 11287 15929 11299 15932
rect 11241 15923 11299 15929
rect 13072 15929 13084 15963
rect 13118 15960 13130 15963
rect 13170 15960 13176 15972
rect 13118 15932 13176 15960
rect 13118 15929 13130 15932
rect 13072 15923 13130 15929
rect 13170 15920 13176 15932
rect 13228 15920 13234 15972
rect 13630 15920 13636 15972
rect 13688 15960 13694 15972
rect 15473 15963 15531 15969
rect 15473 15960 15485 15963
rect 13688 15932 15485 15960
rect 13688 15920 13694 15932
rect 15473 15929 15485 15932
rect 15519 15929 15531 15963
rect 15571 15960 15599 16068
rect 15657 16065 15669 16099
rect 15703 16096 15715 16099
rect 16114 16096 16120 16108
rect 15703 16068 16120 16096
rect 15703 16065 15715 16068
rect 15657 16059 15715 16065
rect 16114 16056 16120 16068
rect 16172 16056 16178 16108
rect 16776 16105 16804 16204
rect 18049 16167 18107 16173
rect 18049 16133 18061 16167
rect 18095 16164 18107 16167
rect 19058 16164 19064 16176
rect 18095 16136 19064 16164
rect 18095 16133 18107 16136
rect 18049 16127 18107 16133
rect 19058 16124 19064 16136
rect 19116 16124 19122 16176
rect 16761 16099 16819 16105
rect 16761 16065 16773 16099
rect 16807 16065 16819 16099
rect 18138 16096 18144 16108
rect 16761 16059 16819 16065
rect 16859 16068 18144 16096
rect 16298 15988 16304 16040
rect 16356 16028 16362 16040
rect 16577 16031 16635 16037
rect 16577 16028 16589 16031
rect 16356 16000 16589 16028
rect 16356 15988 16362 16000
rect 16577 15997 16589 16000
rect 16623 15997 16635 16031
rect 16577 15991 16635 15997
rect 16482 15960 16488 15972
rect 15571 15932 16488 15960
rect 15473 15923 15531 15929
rect 16482 15920 16488 15932
rect 16540 15920 16546 15972
rect 9858 15892 9864 15904
rect 7751 15864 9864 15892
rect 9858 15852 9864 15864
rect 9916 15852 9922 15904
rect 9950 15852 9956 15904
rect 10008 15892 10014 15904
rect 10410 15892 10416 15904
rect 10008 15864 10416 15892
rect 10008 15852 10014 15864
rect 10410 15852 10416 15864
rect 10468 15852 10474 15904
rect 13906 15852 13912 15904
rect 13964 15892 13970 15904
rect 14185 15895 14243 15901
rect 14185 15892 14197 15895
rect 13964 15864 14197 15892
rect 13964 15852 13970 15864
rect 14185 15861 14197 15864
rect 14231 15861 14243 15895
rect 14185 15855 14243 15861
rect 15013 15895 15071 15901
rect 15013 15861 15025 15895
rect 15059 15892 15071 15895
rect 15286 15892 15292 15904
rect 15059 15864 15292 15892
rect 15059 15861 15071 15864
rect 15013 15855 15071 15861
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 15378 15852 15384 15904
rect 15436 15892 15442 15904
rect 15436 15864 15481 15892
rect 15436 15852 15442 15864
rect 16390 15852 16396 15904
rect 16448 15892 16454 15904
rect 16859 15892 16887 16068
rect 18138 16056 18144 16068
rect 18196 16096 18202 16108
rect 18601 16099 18659 16105
rect 18601 16096 18613 16099
rect 18196 16068 18613 16096
rect 18196 16056 18202 16068
rect 18601 16065 18613 16068
rect 18647 16065 18659 16099
rect 18601 16059 18659 16065
rect 19334 16056 19340 16108
rect 19392 16096 19398 16108
rect 20165 16099 20223 16105
rect 20165 16096 20177 16099
rect 19392 16068 20177 16096
rect 19392 16056 19398 16068
rect 20165 16065 20177 16068
rect 20211 16065 20223 16099
rect 20165 16059 20223 16065
rect 17402 15988 17408 16040
rect 17460 16028 17466 16040
rect 17586 16028 17592 16040
rect 17460 16000 17592 16028
rect 17460 15988 17466 16000
rect 17586 15988 17592 16000
rect 17644 16028 17650 16040
rect 19981 16031 20039 16037
rect 19981 16028 19993 16031
rect 17644 16000 19993 16028
rect 17644 15988 17650 16000
rect 19981 15997 19993 16000
rect 20027 15997 20039 16031
rect 19981 15991 20039 15997
rect 20073 16031 20131 16037
rect 20073 15997 20085 16031
rect 20119 16028 20131 16031
rect 20254 16028 20260 16040
rect 20119 16000 20260 16028
rect 20119 15997 20131 16000
rect 20073 15991 20131 15997
rect 20254 15988 20260 16000
rect 20312 15988 20318 16040
rect 18417 15963 18475 15969
rect 18417 15929 18429 15963
rect 18463 15960 18475 15963
rect 19518 15960 19524 15972
rect 18463 15932 19524 15960
rect 18463 15929 18475 15932
rect 18417 15923 18475 15929
rect 19518 15920 19524 15932
rect 19576 15920 19582 15972
rect 16448 15864 16887 15892
rect 16448 15852 16454 15864
rect 17034 15852 17040 15904
rect 17092 15892 17098 15904
rect 17402 15892 17408 15904
rect 17092 15864 17408 15892
rect 17092 15852 17098 15864
rect 17402 15852 17408 15864
rect 17460 15852 17466 15904
rect 18509 15895 18567 15901
rect 18509 15861 18521 15895
rect 18555 15892 18567 15895
rect 19613 15895 19671 15901
rect 19613 15892 19625 15895
rect 18555 15864 19625 15892
rect 18555 15861 18567 15864
rect 18509 15855 18567 15861
rect 19613 15861 19625 15864
rect 19659 15861 19671 15895
rect 19613 15855 19671 15861
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 1397 15691 1455 15697
rect 1397 15657 1409 15691
rect 1443 15688 1455 15691
rect 3602 15688 3608 15700
rect 1443 15660 3608 15688
rect 1443 15657 1455 15660
rect 1397 15651 1455 15657
rect 3602 15648 3608 15660
rect 3660 15648 3666 15700
rect 4249 15691 4307 15697
rect 4249 15657 4261 15691
rect 4295 15688 4307 15691
rect 4430 15688 4436 15700
rect 4295 15660 4436 15688
rect 4295 15657 4307 15660
rect 4249 15651 4307 15657
rect 4430 15648 4436 15660
rect 4488 15648 4494 15700
rect 4709 15691 4767 15697
rect 4709 15657 4721 15691
rect 4755 15688 4767 15691
rect 5166 15688 5172 15700
rect 4755 15660 5172 15688
rect 4755 15657 4767 15660
rect 4709 15651 4767 15657
rect 5166 15648 5172 15660
rect 5224 15688 5230 15700
rect 5442 15688 5448 15700
rect 5224 15660 5448 15688
rect 5224 15648 5230 15660
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 5534 15648 5540 15700
rect 5592 15648 5598 15700
rect 7190 15648 7196 15700
rect 7248 15688 7254 15700
rect 7466 15688 7472 15700
rect 7248 15660 7472 15688
rect 7248 15648 7254 15660
rect 7466 15648 7472 15660
rect 7524 15648 7530 15700
rect 8021 15691 8079 15697
rect 8021 15657 8033 15691
rect 8067 15688 8079 15691
rect 8202 15688 8208 15700
rect 8067 15660 8208 15688
rect 8067 15657 8079 15660
rect 8021 15651 8079 15657
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 8389 15691 8447 15697
rect 8389 15657 8401 15691
rect 8435 15688 8447 15691
rect 9214 15688 9220 15700
rect 8435 15660 9220 15688
rect 8435 15657 8447 15660
rect 8389 15651 8447 15657
rect 9214 15648 9220 15660
rect 9272 15648 9278 15700
rect 10134 15648 10140 15700
rect 10192 15648 10198 15700
rect 10410 15648 10416 15700
rect 10468 15648 10474 15700
rect 10962 15648 10968 15700
rect 11020 15688 11026 15700
rect 11241 15691 11299 15697
rect 11241 15688 11253 15691
rect 11020 15660 11253 15688
rect 11020 15648 11026 15660
rect 11241 15657 11253 15660
rect 11287 15657 11299 15691
rect 13630 15688 13636 15700
rect 13591 15660 13636 15688
rect 11241 15651 11299 15657
rect 13630 15648 13636 15660
rect 13688 15648 13694 15700
rect 13998 15688 14004 15700
rect 13959 15660 14004 15688
rect 13998 15648 14004 15660
rect 14056 15648 14062 15700
rect 14090 15648 14096 15700
rect 14148 15688 14154 15700
rect 14148 15660 14193 15688
rect 14148 15648 14154 15660
rect 16666 15648 16672 15700
rect 16724 15688 16730 15700
rect 17586 15688 17592 15700
rect 16724 15660 17592 15688
rect 16724 15648 16730 15660
rect 17586 15648 17592 15660
rect 17644 15648 17650 15700
rect 2590 15580 2596 15632
rect 2648 15620 2654 15632
rect 2869 15623 2927 15629
rect 2869 15620 2881 15623
rect 2648 15592 2881 15620
rect 2648 15580 2654 15592
rect 2869 15589 2881 15592
rect 2915 15589 2927 15623
rect 2869 15583 2927 15589
rect 4617 15623 4675 15629
rect 4617 15589 4629 15623
rect 4663 15620 4675 15623
rect 5552 15620 5580 15648
rect 9950 15620 9956 15632
rect 4663 15592 5580 15620
rect 6012 15592 9956 15620
rect 4663 15589 4675 15592
rect 4617 15583 4675 15589
rect 2777 15555 2835 15561
rect 2777 15521 2789 15555
rect 2823 15552 2835 15555
rect 3878 15552 3884 15564
rect 2823 15524 3884 15552
rect 2823 15521 2835 15524
rect 2777 15515 2835 15521
rect 3878 15512 3884 15524
rect 3936 15512 3942 15564
rect 6012 15552 6040 15592
rect 9950 15580 9956 15592
rect 10008 15580 10014 15632
rect 4816 15524 6040 15552
rect 6080 15555 6138 15561
rect 3050 15484 3056 15496
rect 3011 15456 3056 15484
rect 3050 15444 3056 15456
rect 3108 15444 3114 15496
rect 4816 15493 4844 15524
rect 6080 15521 6092 15555
rect 6126 15552 6138 15555
rect 6454 15552 6460 15564
rect 6126 15524 6460 15552
rect 6126 15521 6138 15524
rect 6080 15515 6138 15521
rect 6454 15512 6460 15524
rect 6512 15512 6518 15564
rect 6546 15512 6552 15564
rect 6604 15552 6610 15564
rect 6604 15524 6868 15552
rect 6604 15512 6610 15524
rect 4801 15487 4859 15493
rect 4801 15453 4813 15487
rect 4847 15453 4859 15487
rect 4801 15447 4859 15453
rect 1394 15376 1400 15428
rect 1452 15416 1458 15428
rect 4816 15416 4844 15447
rect 5626 15444 5632 15496
rect 5684 15484 5690 15496
rect 5813 15487 5871 15493
rect 5813 15484 5825 15487
rect 5684 15456 5825 15484
rect 5684 15444 5690 15456
rect 5813 15453 5825 15456
rect 5859 15453 5871 15487
rect 6840 15484 6868 15524
rect 7282 15512 7288 15564
rect 7340 15552 7346 15564
rect 10042 15552 10048 15564
rect 7340 15524 8616 15552
rect 10003 15524 10048 15552
rect 7340 15512 7346 15524
rect 8588 15493 8616 15524
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 10152 15561 10180 15648
rect 10428 15620 10456 15648
rect 10428 15592 11836 15620
rect 10137 15555 10195 15561
rect 10137 15521 10149 15555
rect 10183 15552 10195 15555
rect 10183 15524 10364 15552
rect 10183 15521 10195 15524
rect 10137 15515 10195 15521
rect 8481 15487 8539 15493
rect 8481 15484 8493 15487
rect 6840 15456 8493 15484
rect 5813 15447 5871 15453
rect 8481 15453 8493 15456
rect 8527 15453 8539 15487
rect 8481 15447 8539 15453
rect 8573 15487 8631 15493
rect 8573 15453 8585 15487
rect 8619 15453 8631 15487
rect 8573 15447 8631 15453
rect 9674 15444 9680 15496
rect 9732 15484 9738 15496
rect 10229 15487 10287 15493
rect 9732 15456 9996 15484
rect 9732 15444 9738 15456
rect 1452 15388 4844 15416
rect 1452 15376 1458 15388
rect 8294 15376 8300 15428
rect 8352 15416 8358 15428
rect 9858 15416 9864 15428
rect 8352 15388 9864 15416
rect 8352 15376 8358 15388
rect 9858 15376 9864 15388
rect 9916 15376 9922 15428
rect 2222 15308 2228 15360
rect 2280 15348 2286 15360
rect 2409 15351 2467 15357
rect 2409 15348 2421 15351
rect 2280 15320 2421 15348
rect 2280 15308 2286 15320
rect 2409 15317 2421 15320
rect 2455 15317 2467 15351
rect 2409 15311 2467 15317
rect 7193 15351 7251 15357
rect 7193 15317 7205 15351
rect 7239 15348 7251 15351
rect 7282 15348 7288 15360
rect 7239 15320 7288 15348
rect 7239 15317 7251 15320
rect 7193 15311 7251 15317
rect 7282 15308 7288 15320
rect 7340 15308 7346 15360
rect 8202 15308 8208 15360
rect 8260 15348 8266 15360
rect 9122 15348 9128 15360
rect 8260 15320 9128 15348
rect 8260 15308 8266 15320
rect 9122 15308 9128 15320
rect 9180 15308 9186 15360
rect 9674 15348 9680 15360
rect 9635 15320 9680 15348
rect 9674 15308 9680 15320
rect 9732 15308 9738 15360
rect 9968 15348 9996 15456
rect 10229 15453 10241 15487
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 10244 15360 10272 15447
rect 10336 15416 10364 15524
rect 10410 15512 10416 15564
rect 10468 15552 10474 15564
rect 11606 15552 11612 15564
rect 10468 15524 11612 15552
rect 10468 15512 10474 15524
rect 11606 15512 11612 15524
rect 11664 15512 11670 15564
rect 10502 15444 10508 15496
rect 10560 15484 10566 15496
rect 10962 15484 10968 15496
rect 10560 15456 10968 15484
rect 10560 15444 10566 15456
rect 10962 15444 10968 15456
rect 11020 15484 11026 15496
rect 11808 15493 11836 15592
rect 14550 15580 14556 15632
rect 14608 15620 14614 15632
rect 14918 15620 14924 15632
rect 14608 15592 14924 15620
rect 14608 15580 14614 15592
rect 14918 15580 14924 15592
rect 14976 15580 14982 15632
rect 16206 15580 16212 15632
rect 16264 15620 16270 15632
rect 19245 15623 19303 15629
rect 19245 15620 19257 15623
rect 16264 15592 19257 15620
rect 16264 15580 16270 15592
rect 19245 15589 19257 15592
rect 19291 15589 19303 15623
rect 19245 15583 19303 15589
rect 15286 15552 15292 15564
rect 15247 15524 15292 15552
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 16844 15555 16902 15561
rect 16844 15521 16856 15555
rect 16890 15552 16902 15555
rect 17310 15552 17316 15564
rect 16890 15524 17316 15552
rect 16890 15521 16902 15524
rect 16844 15515 16902 15521
rect 17310 15512 17316 15524
rect 17368 15512 17374 15564
rect 19150 15552 19156 15564
rect 19111 15524 19156 15552
rect 19150 15512 19156 15524
rect 19208 15512 19214 15564
rect 11701 15487 11759 15493
rect 11701 15484 11713 15487
rect 11020 15456 11713 15484
rect 11020 15444 11026 15456
rect 11701 15453 11713 15456
rect 11747 15453 11759 15487
rect 11701 15447 11759 15453
rect 11793 15487 11851 15493
rect 11793 15453 11805 15487
rect 11839 15453 11851 15487
rect 11793 15447 11851 15453
rect 13998 15444 14004 15496
rect 14056 15484 14062 15496
rect 14185 15487 14243 15493
rect 14185 15484 14197 15487
rect 14056 15456 14197 15484
rect 14056 15444 14062 15456
rect 14185 15453 14197 15456
rect 14231 15484 14243 15487
rect 14734 15484 14740 15496
rect 14231 15456 14740 15484
rect 14231 15453 14243 15456
rect 14185 15447 14243 15453
rect 14734 15444 14740 15456
rect 14792 15444 14798 15496
rect 15565 15487 15623 15493
rect 15565 15453 15577 15487
rect 15611 15484 15623 15487
rect 15838 15484 15844 15496
rect 15611 15456 15844 15484
rect 15611 15453 15623 15456
rect 15565 15447 15623 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 16482 15444 16488 15496
rect 16540 15484 16546 15496
rect 16577 15487 16635 15493
rect 16577 15484 16589 15487
rect 16540 15456 16589 15484
rect 16540 15444 16546 15456
rect 16577 15453 16589 15456
rect 16623 15453 16635 15487
rect 16577 15447 16635 15453
rect 18138 15444 18144 15496
rect 18196 15484 18202 15496
rect 19334 15484 19340 15496
rect 18196 15456 18920 15484
rect 19295 15456 19340 15484
rect 18196 15444 18202 15456
rect 12158 15416 12164 15428
rect 10336 15388 12164 15416
rect 12158 15376 12164 15388
rect 12216 15376 12222 15428
rect 17586 15376 17592 15428
rect 17644 15416 17650 15428
rect 18785 15419 18843 15425
rect 18785 15416 18797 15419
rect 17644 15388 18797 15416
rect 17644 15376 17650 15388
rect 18785 15385 18797 15388
rect 18831 15385 18843 15419
rect 18892 15416 18920 15456
rect 19334 15444 19340 15456
rect 19392 15444 19398 15496
rect 19610 15416 19616 15428
rect 18892 15388 19616 15416
rect 18785 15379 18843 15385
rect 19610 15376 19616 15388
rect 19668 15416 19674 15428
rect 20070 15416 20076 15428
rect 19668 15388 20076 15416
rect 19668 15376 19674 15388
rect 20070 15376 20076 15388
rect 20128 15376 20134 15428
rect 10226 15348 10232 15360
rect 9968 15320 10232 15348
rect 10226 15308 10232 15320
rect 10284 15308 10290 15360
rect 12710 15308 12716 15360
rect 12768 15348 12774 15360
rect 14090 15348 14096 15360
rect 12768 15320 14096 15348
rect 12768 15308 12774 15320
rect 14090 15308 14096 15320
rect 14148 15308 14154 15360
rect 17957 15351 18015 15357
rect 17957 15317 17969 15351
rect 18003 15348 18015 15351
rect 18874 15348 18880 15360
rect 18003 15320 18880 15348
rect 18003 15317 18015 15320
rect 17957 15311 18015 15317
rect 18874 15308 18880 15320
rect 18932 15308 18938 15360
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 1946 15104 1952 15156
rect 2004 15144 2010 15156
rect 3234 15144 3240 15156
rect 2004 15116 3240 15144
rect 2004 15104 2010 15116
rect 3234 15104 3240 15116
rect 3292 15104 3298 15156
rect 6825 15147 6883 15153
rect 6825 15113 6837 15147
rect 6871 15144 6883 15147
rect 10870 15144 10876 15156
rect 6871 15116 10876 15144
rect 6871 15113 6883 15116
rect 6825 15107 6883 15113
rect 10870 15104 10876 15116
rect 10928 15104 10934 15156
rect 15746 15104 15752 15156
rect 15804 15144 15810 15156
rect 15804 15116 18460 15144
rect 15804 15104 15810 15116
rect 18432 15088 18460 15116
rect 19518 15104 19524 15156
rect 19576 15144 19582 15156
rect 19613 15147 19671 15153
rect 19613 15144 19625 15147
rect 19576 15116 19625 15144
rect 19576 15104 19582 15116
rect 19613 15113 19625 15116
rect 19659 15113 19671 15147
rect 19613 15107 19671 15113
rect 1670 15036 1676 15088
rect 1728 15076 1734 15088
rect 2130 15076 2136 15088
rect 1728 15048 2136 15076
rect 1728 15036 1734 15048
rect 2130 15036 2136 15048
rect 2188 15036 2194 15088
rect 5626 15036 5632 15088
rect 5684 15076 5690 15088
rect 6457 15079 6515 15085
rect 6457 15076 6469 15079
rect 5684 15048 6469 15076
rect 5684 15036 5690 15048
rect 6457 15045 6469 15048
rect 6503 15076 6515 15079
rect 7466 15076 7472 15088
rect 6503 15048 7472 15076
rect 6503 15045 6515 15048
rect 6457 15039 6515 15045
rect 7466 15036 7472 15048
rect 7524 15076 7530 15088
rect 7524 15048 7788 15076
rect 7524 15036 7530 15048
rect 7760 15020 7788 15048
rect 9766 15036 9772 15088
rect 9824 15076 9830 15088
rect 14274 15076 14280 15088
rect 9824 15048 14280 15076
rect 9824 15036 9830 15048
rect 14274 15036 14280 15048
rect 14332 15036 14338 15088
rect 14550 15036 14556 15088
rect 14608 15076 14614 15088
rect 14921 15079 14979 15085
rect 14921 15076 14933 15079
rect 14608 15048 14933 15076
rect 14608 15036 14614 15048
rect 14921 15045 14933 15048
rect 14967 15045 14979 15079
rect 17586 15076 17592 15088
rect 14921 15039 14979 15045
rect 15396 15048 17592 15076
rect 2869 15011 2927 15017
rect 2869 14977 2881 15011
rect 2915 15008 2927 15011
rect 3510 15008 3516 15020
rect 2915 14980 3516 15008
rect 2915 14977 2927 14980
rect 2869 14971 2927 14977
rect 3510 14968 3516 14980
rect 3568 14968 3574 15020
rect 5460 14980 6776 15008
rect 1486 14900 1492 14952
rect 1544 14940 1550 14952
rect 2038 14940 2044 14952
rect 1544 14912 2044 14940
rect 1544 14900 1550 14912
rect 2038 14900 2044 14912
rect 2096 14940 2102 14952
rect 3789 14943 3847 14949
rect 3789 14940 3801 14943
rect 2096 14912 3801 14940
rect 2096 14900 2102 14912
rect 3789 14909 3801 14912
rect 3835 14909 3847 14943
rect 3789 14903 3847 14909
rect 2593 14875 2651 14881
rect 2593 14841 2605 14875
rect 2639 14872 2651 14875
rect 3326 14872 3332 14884
rect 2639 14844 3332 14872
rect 2639 14841 2651 14844
rect 2593 14835 2651 14841
rect 3326 14832 3332 14844
rect 3384 14832 3390 14884
rect 4056 14875 4114 14881
rect 4056 14841 4068 14875
rect 4102 14872 4114 14875
rect 4982 14872 4988 14884
rect 4102 14844 4988 14872
rect 4102 14841 4114 14844
rect 4056 14835 4114 14841
rect 4982 14832 4988 14844
rect 5040 14832 5046 14884
rect 2130 14764 2136 14816
rect 2188 14804 2194 14816
rect 2225 14807 2283 14813
rect 2225 14804 2237 14807
rect 2188 14776 2237 14804
rect 2188 14764 2194 14776
rect 2225 14773 2237 14776
rect 2271 14773 2283 14807
rect 2225 14767 2283 14773
rect 2498 14764 2504 14816
rect 2556 14804 2562 14816
rect 2685 14807 2743 14813
rect 2685 14804 2697 14807
rect 2556 14776 2697 14804
rect 2556 14764 2562 14776
rect 2685 14773 2697 14776
rect 2731 14773 2743 14807
rect 5166 14804 5172 14816
rect 5127 14776 5172 14804
rect 2685 14767 2743 14773
rect 5166 14764 5172 14776
rect 5224 14764 5230 14816
rect 5350 14764 5356 14816
rect 5408 14804 5414 14816
rect 5460 14804 5488 14980
rect 6638 14940 6644 14952
rect 6599 14912 6644 14940
rect 6638 14900 6644 14912
rect 6696 14900 6702 14952
rect 6748 14940 6776 14980
rect 7282 14968 7288 15020
rect 7340 15008 7346 15020
rect 7377 15011 7435 15017
rect 7377 15008 7389 15011
rect 7340 14980 7389 15008
rect 7340 14968 7346 14980
rect 7377 14977 7389 14980
rect 7423 14977 7435 15011
rect 7377 14971 7435 14977
rect 7742 14968 7748 15020
rect 7800 15008 7806 15020
rect 8573 15011 8631 15017
rect 8573 15008 8585 15011
rect 7800 14980 8585 15008
rect 7800 14968 7806 14980
rect 8573 14977 8585 14980
rect 8619 14977 8631 15011
rect 8573 14971 8631 14977
rect 10226 14968 10232 15020
rect 10284 15008 10290 15020
rect 11333 15011 11391 15017
rect 11333 15008 11345 15011
rect 10284 14980 11345 15008
rect 10284 14968 10290 14980
rect 11333 14977 11345 14980
rect 11379 14977 11391 15011
rect 11882 15008 11888 15020
rect 11333 14971 11391 14977
rect 11440 14980 11888 15008
rect 6748 14912 8984 14940
rect 6546 14832 6552 14884
rect 6604 14872 6610 14884
rect 8846 14881 8852 14884
rect 7193 14875 7251 14881
rect 7193 14872 7205 14875
rect 6604 14844 7205 14872
rect 6604 14832 6610 14844
rect 7193 14841 7205 14844
rect 7239 14841 7251 14875
rect 8840 14872 8852 14881
rect 8807 14844 8852 14872
rect 7193 14835 7251 14841
rect 8840 14835 8852 14844
rect 8846 14832 8852 14835
rect 8904 14832 8910 14884
rect 8956 14872 8984 14912
rect 9306 14900 9312 14952
rect 9364 14940 9370 14952
rect 11440 14940 11468 14980
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 12526 14968 12532 15020
rect 12584 15008 12590 15020
rect 13170 15008 13176 15020
rect 12584 14980 13176 15008
rect 12584 14968 12590 14980
rect 13170 14968 13176 14980
rect 13228 14968 13234 15020
rect 13357 15011 13415 15017
rect 13357 14977 13369 15011
rect 13403 15008 13415 15011
rect 13630 15008 13636 15020
rect 13403 14980 13636 15008
rect 13403 14977 13415 14980
rect 13357 14971 13415 14977
rect 13630 14968 13636 14980
rect 13688 14968 13694 15020
rect 15396 15017 15424 15048
rect 17586 15036 17592 15048
rect 17644 15036 17650 15088
rect 18414 15036 18420 15088
rect 18472 15036 18478 15088
rect 15381 15011 15439 15017
rect 15381 14977 15393 15011
rect 15427 14977 15439 15011
rect 15381 14971 15439 14977
rect 15473 15011 15531 15017
rect 15473 14977 15485 15011
rect 15519 15008 15531 15011
rect 16390 15008 16396 15020
rect 15519 14980 16396 15008
rect 15519 14977 15531 14980
rect 15473 14971 15531 14977
rect 9364 14912 11468 14940
rect 9364 14900 9370 14912
rect 14734 14900 14740 14952
rect 14792 14940 14798 14952
rect 14829 14943 14887 14949
rect 14829 14940 14841 14943
rect 14792 14912 14841 14940
rect 14792 14900 14798 14912
rect 14829 14909 14841 14912
rect 14875 14909 14887 14943
rect 14829 14903 14887 14909
rect 15102 14900 15108 14952
rect 15160 14940 15166 14952
rect 15488 14940 15516 14971
rect 16390 14968 16396 14980
rect 16448 14968 16454 15020
rect 17310 14968 17316 15020
rect 17368 15008 17374 15020
rect 18601 15011 18659 15017
rect 18601 15008 18613 15011
rect 17368 14980 18613 15008
rect 17368 14968 17374 14980
rect 18601 14977 18613 14980
rect 18647 14977 18659 15011
rect 18601 14971 18659 14977
rect 19334 14968 19340 15020
rect 19392 15008 19398 15020
rect 20165 15011 20223 15017
rect 20165 15008 20177 15011
rect 19392 14980 20177 15008
rect 19392 14968 19398 14980
rect 20165 14977 20177 14980
rect 20211 14977 20223 15011
rect 20165 14971 20223 14977
rect 15160 14912 15516 14940
rect 16669 14943 16727 14949
rect 15160 14900 15166 14912
rect 16669 14909 16681 14943
rect 16715 14940 16727 14943
rect 16850 14940 16856 14952
rect 16715 14912 16856 14940
rect 16715 14909 16727 14912
rect 16669 14903 16727 14909
rect 16850 14900 16856 14912
rect 16908 14900 16914 14952
rect 16945 14943 17003 14949
rect 16945 14909 16957 14943
rect 16991 14940 17003 14943
rect 17862 14940 17868 14952
rect 16991 14912 17868 14940
rect 16991 14909 17003 14912
rect 16945 14903 17003 14909
rect 17862 14900 17868 14912
rect 17920 14900 17926 14952
rect 18138 14900 18144 14952
rect 18196 14940 18202 14952
rect 18966 14940 18972 14952
rect 18196 14912 18972 14940
rect 18196 14900 18202 14912
rect 18966 14900 18972 14912
rect 19024 14900 19030 14952
rect 20070 14940 20076 14952
rect 20031 14912 20076 14940
rect 20070 14900 20076 14912
rect 20128 14900 20134 14952
rect 11146 14872 11152 14884
rect 8956 14844 10916 14872
rect 11107 14844 11152 14872
rect 5408 14776 5488 14804
rect 5408 14764 5414 14776
rect 5626 14764 5632 14816
rect 5684 14804 5690 14816
rect 5902 14804 5908 14816
rect 5684 14776 5908 14804
rect 5684 14764 5690 14776
rect 5902 14764 5908 14776
rect 5960 14764 5966 14816
rect 7285 14807 7343 14813
rect 7285 14773 7297 14807
rect 7331 14804 7343 14807
rect 9582 14804 9588 14816
rect 7331 14776 9588 14804
rect 7331 14773 7343 14776
rect 7285 14767 7343 14773
rect 9582 14764 9588 14776
rect 9640 14764 9646 14816
rect 9950 14804 9956 14816
rect 9911 14776 9956 14804
rect 9950 14764 9956 14776
rect 10008 14764 10014 14816
rect 10778 14804 10784 14816
rect 10739 14776 10784 14804
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 10888 14804 10916 14844
rect 11146 14832 11152 14844
rect 11204 14832 11210 14884
rect 12434 14832 12440 14884
rect 12492 14872 12498 14884
rect 13354 14872 13360 14884
rect 12492 14844 13360 14872
rect 12492 14832 12498 14844
rect 13354 14832 13360 14844
rect 13412 14832 13418 14884
rect 14918 14832 14924 14884
rect 14976 14872 14982 14884
rect 14976 14844 15424 14872
rect 14976 14832 14982 14844
rect 11241 14807 11299 14813
rect 11241 14804 11253 14807
rect 10888 14776 11253 14804
rect 11241 14773 11253 14776
rect 11287 14773 11299 14807
rect 12710 14804 12716 14816
rect 12671 14776 12716 14804
rect 11241 14767 11299 14773
rect 12710 14764 12716 14776
rect 12768 14764 12774 14816
rect 13078 14804 13084 14816
rect 13039 14776 13084 14804
rect 13078 14764 13084 14776
rect 13136 14764 13142 14816
rect 14090 14764 14096 14816
rect 14148 14804 14154 14816
rect 14645 14807 14703 14813
rect 14645 14804 14657 14807
rect 14148 14776 14657 14804
rect 14148 14764 14154 14776
rect 14645 14773 14657 14776
rect 14691 14773 14703 14807
rect 14645 14767 14703 14773
rect 14734 14764 14740 14816
rect 14792 14804 14798 14816
rect 15289 14807 15347 14813
rect 15289 14804 15301 14807
rect 14792 14776 15301 14804
rect 14792 14764 14798 14776
rect 15289 14773 15301 14776
rect 15335 14773 15347 14807
rect 15396 14804 15424 14844
rect 16390 14832 16396 14884
rect 16448 14872 16454 14884
rect 19981 14875 20039 14881
rect 19981 14872 19993 14875
rect 16448 14844 19993 14872
rect 16448 14832 16454 14844
rect 19981 14841 19993 14844
rect 20027 14841 20039 14875
rect 19981 14835 20039 14841
rect 17034 14804 17040 14816
rect 15396 14776 17040 14804
rect 15289 14767 15347 14773
rect 17034 14764 17040 14776
rect 17092 14764 17098 14816
rect 18049 14807 18107 14813
rect 18049 14773 18061 14807
rect 18095 14804 18107 14807
rect 18230 14804 18236 14816
rect 18095 14776 18236 14804
rect 18095 14773 18107 14776
rect 18049 14767 18107 14773
rect 18230 14764 18236 14776
rect 18288 14764 18294 14816
rect 18414 14804 18420 14816
rect 18375 14776 18420 14804
rect 18414 14764 18420 14776
rect 18472 14764 18478 14816
rect 18509 14807 18567 14813
rect 18509 14773 18521 14807
rect 18555 14804 18567 14807
rect 18598 14804 18604 14816
rect 18555 14776 18604 14804
rect 18555 14773 18567 14776
rect 18509 14767 18567 14773
rect 18598 14764 18604 14776
rect 18656 14764 18662 14816
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 6457 14603 6515 14609
rect 6457 14569 6469 14603
rect 6503 14600 6515 14603
rect 6546 14600 6552 14612
rect 6503 14572 6552 14600
rect 6503 14569 6515 14572
rect 6457 14563 6515 14569
rect 6546 14560 6552 14572
rect 6604 14560 6610 14612
rect 6822 14600 6828 14612
rect 6783 14572 6828 14600
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 7006 14560 7012 14612
rect 7064 14600 7070 14612
rect 8021 14603 8079 14609
rect 8021 14600 8033 14603
rect 7064 14572 8033 14600
rect 7064 14560 7070 14572
rect 8021 14569 8033 14572
rect 8067 14569 8079 14603
rect 8021 14563 8079 14569
rect 8389 14603 8447 14609
rect 8389 14569 8401 14603
rect 8435 14600 8447 14603
rect 10778 14600 10784 14612
rect 8435 14572 10784 14600
rect 8435 14569 8447 14572
rect 8389 14563 8447 14569
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 10870 14560 10876 14612
rect 10928 14600 10934 14612
rect 12434 14600 12440 14612
rect 10928 14572 12440 14600
rect 10928 14560 10934 14572
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 12526 14560 12532 14612
rect 12584 14600 12590 14612
rect 14274 14600 14280 14612
rect 12584 14572 13952 14600
rect 14235 14572 14280 14600
rect 12584 14560 12590 14572
rect 2032 14535 2090 14541
rect 2032 14501 2044 14535
rect 2078 14532 2090 14535
rect 5902 14532 5908 14544
rect 2078 14504 5908 14532
rect 2078 14501 2090 14504
rect 2032 14495 2090 14501
rect 5902 14492 5908 14504
rect 5960 14492 5966 14544
rect 6730 14492 6736 14544
rect 6788 14532 6794 14544
rect 6917 14535 6975 14541
rect 6917 14532 6929 14535
rect 6788 14504 6929 14532
rect 6788 14492 6794 14504
rect 6917 14501 6929 14504
rect 6963 14532 6975 14535
rect 8481 14535 8539 14541
rect 6963 14504 7052 14532
rect 6963 14501 6975 14504
rect 6917 14495 6975 14501
rect 7024 14476 7052 14504
rect 8481 14501 8493 14535
rect 8527 14532 8539 14535
rect 9674 14532 9680 14544
rect 8527 14504 9680 14532
rect 8527 14501 8539 14504
rect 8481 14495 8539 14501
rect 9674 14492 9680 14504
rect 9732 14492 9738 14544
rect 11330 14532 11336 14544
rect 9784 14504 11336 14532
rect 3970 14424 3976 14476
rect 4028 14464 4034 14476
rect 4706 14464 4712 14476
rect 4028 14436 4712 14464
rect 4028 14424 4034 14436
rect 4706 14424 4712 14436
rect 4764 14464 4770 14476
rect 4801 14467 4859 14473
rect 4801 14464 4813 14467
rect 4764 14436 4813 14464
rect 4764 14424 4770 14436
rect 4801 14433 4813 14436
rect 4847 14433 4859 14467
rect 4801 14427 4859 14433
rect 4893 14467 4951 14473
rect 4893 14433 4905 14467
rect 4939 14464 4951 14467
rect 5074 14464 5080 14476
rect 4939 14436 5080 14464
rect 4939 14433 4951 14436
rect 4893 14427 4951 14433
rect 5074 14424 5080 14436
rect 5132 14464 5138 14476
rect 6362 14464 6368 14476
rect 5132 14436 6368 14464
rect 5132 14424 5138 14436
rect 6362 14424 6368 14436
rect 6420 14424 6426 14476
rect 7006 14424 7012 14476
rect 7064 14424 7070 14476
rect 9214 14424 9220 14476
rect 9272 14464 9278 14476
rect 9784 14464 9812 14504
rect 11330 14492 11336 14504
rect 11388 14492 11394 14544
rect 12152 14535 12210 14541
rect 12152 14501 12164 14535
rect 12198 14532 12210 14535
rect 12986 14532 12992 14544
rect 12198 14504 12992 14532
rect 12198 14501 12210 14504
rect 12152 14495 12210 14501
rect 12986 14492 12992 14504
rect 13044 14492 13050 14544
rect 13924 14532 13952 14572
rect 14274 14560 14280 14572
rect 14332 14560 14338 14612
rect 17129 14603 17187 14609
rect 17129 14569 17141 14603
rect 17175 14600 17187 14603
rect 18233 14603 18291 14609
rect 18233 14600 18245 14603
rect 17175 14572 18245 14600
rect 17175 14569 17187 14572
rect 17129 14563 17187 14569
rect 18233 14569 18245 14572
rect 18279 14569 18291 14603
rect 18233 14563 18291 14569
rect 18322 14560 18328 14612
rect 18380 14600 18386 14612
rect 18693 14603 18751 14609
rect 18693 14600 18705 14603
rect 18380 14572 18705 14600
rect 18380 14560 18386 14572
rect 18693 14569 18705 14572
rect 18739 14569 18751 14603
rect 18693 14563 18751 14569
rect 17037 14535 17095 14541
rect 13924 14504 15424 14532
rect 9272 14436 9812 14464
rect 10045 14467 10103 14473
rect 9272 14424 9278 14436
rect 10045 14433 10057 14467
rect 10091 14464 10103 14467
rect 11422 14464 11428 14476
rect 10091 14436 10640 14464
rect 11383 14436 11428 14464
rect 10091 14433 10103 14436
rect 10045 14427 10103 14433
rect 1486 14356 1492 14408
rect 1544 14396 1550 14408
rect 1765 14399 1823 14405
rect 1765 14396 1777 14399
rect 1544 14368 1777 14396
rect 1544 14356 1550 14368
rect 1765 14365 1777 14368
rect 1811 14365 1823 14399
rect 4982 14396 4988 14408
rect 4943 14368 4988 14396
rect 1765 14359 1823 14365
rect 4982 14356 4988 14368
rect 5040 14356 5046 14408
rect 6454 14356 6460 14408
rect 6512 14396 6518 14408
rect 7101 14399 7159 14405
rect 7101 14396 7113 14399
rect 6512 14368 7113 14396
rect 6512 14356 6518 14368
rect 7101 14365 7113 14368
rect 7147 14365 7159 14399
rect 8662 14396 8668 14408
rect 8623 14368 8668 14396
rect 7101 14359 7159 14365
rect 3145 14331 3203 14337
rect 3145 14297 3157 14331
rect 3191 14328 3203 14331
rect 6362 14328 6368 14340
rect 3191 14300 6368 14328
rect 3191 14297 3203 14300
rect 3145 14291 3203 14297
rect 6362 14288 6368 14300
rect 6420 14288 6426 14340
rect 7116 14328 7144 14359
rect 8662 14356 8668 14368
rect 8720 14356 8726 14408
rect 9674 14356 9680 14408
rect 9732 14396 9738 14408
rect 10137 14399 10195 14405
rect 10137 14396 10149 14399
rect 9732 14368 10149 14396
rect 9732 14356 9738 14368
rect 10137 14365 10149 14368
rect 10183 14365 10195 14399
rect 10137 14359 10195 14365
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14365 10287 14399
rect 10229 14359 10287 14365
rect 9950 14328 9956 14340
rect 7116 14300 9956 14328
rect 9950 14288 9956 14300
rect 10008 14328 10014 14340
rect 10244 14328 10272 14359
rect 10008 14300 10272 14328
rect 10008 14288 10014 14300
rect 4154 14220 4160 14272
rect 4212 14260 4218 14272
rect 4433 14263 4491 14269
rect 4433 14260 4445 14263
rect 4212 14232 4445 14260
rect 4212 14220 4218 14232
rect 4433 14229 4445 14232
rect 4479 14229 4491 14263
rect 4433 14223 4491 14229
rect 6178 14220 6184 14272
rect 6236 14260 6242 14272
rect 9306 14260 9312 14272
rect 6236 14232 9312 14260
rect 6236 14220 6242 14232
rect 9306 14220 9312 14232
rect 9364 14220 9370 14272
rect 9582 14220 9588 14272
rect 9640 14260 9646 14272
rect 10612 14269 10640 14436
rect 11422 14424 11428 14436
rect 11480 14424 11486 14476
rect 12434 14424 12440 14476
rect 12492 14464 12498 14476
rect 14093 14467 14151 14473
rect 14093 14464 14105 14467
rect 12492 14436 14105 14464
rect 12492 14424 12498 14436
rect 14093 14433 14105 14436
rect 14139 14433 14151 14467
rect 14093 14427 14151 14433
rect 14274 14424 14280 14476
rect 14332 14464 14338 14476
rect 14458 14464 14464 14476
rect 14332 14436 14464 14464
rect 14332 14424 14338 14436
rect 14458 14424 14464 14436
rect 14516 14424 14522 14476
rect 15194 14424 15200 14476
rect 15252 14464 15258 14476
rect 15289 14467 15347 14473
rect 15289 14464 15301 14467
rect 15252 14436 15301 14464
rect 15252 14424 15258 14436
rect 15289 14433 15301 14436
rect 15335 14433 15347 14467
rect 15396 14464 15424 14504
rect 17037 14501 17049 14535
rect 17083 14532 17095 14535
rect 18966 14532 18972 14544
rect 17083 14504 18972 14532
rect 17083 14501 17095 14504
rect 17037 14495 17095 14501
rect 18966 14492 18972 14504
rect 19024 14492 19030 14544
rect 18138 14464 18144 14476
rect 15396 14436 18144 14464
rect 15289 14427 15347 14433
rect 18138 14424 18144 14436
rect 18196 14424 18202 14476
rect 18601 14467 18659 14473
rect 18601 14433 18613 14467
rect 18647 14464 18659 14467
rect 20254 14464 20260 14476
rect 18647 14436 20260 14464
rect 18647 14433 18659 14436
rect 18601 14427 18659 14433
rect 20254 14424 20260 14436
rect 20312 14424 20318 14476
rect 11882 14396 11888 14408
rect 11843 14368 11888 14396
rect 11882 14356 11888 14368
rect 11940 14356 11946 14408
rect 13906 14356 13912 14408
rect 13964 14396 13970 14408
rect 15473 14399 15531 14405
rect 15473 14396 15485 14399
rect 13964 14368 15485 14396
rect 13964 14356 13970 14368
rect 15473 14365 15485 14368
rect 15519 14365 15531 14399
rect 17310 14396 17316 14408
rect 17271 14368 17316 14396
rect 15473 14359 15531 14365
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 18874 14396 18880 14408
rect 18835 14368 18880 14396
rect 18874 14356 18880 14368
rect 18932 14356 18938 14408
rect 19797 14399 19855 14405
rect 19797 14365 19809 14399
rect 19843 14365 19855 14399
rect 19797 14359 19855 14365
rect 13170 14288 13176 14340
rect 13228 14328 13234 14340
rect 13265 14331 13323 14337
rect 13265 14328 13277 14331
rect 13228 14300 13277 14328
rect 13228 14288 13234 14300
rect 13265 14297 13277 14300
rect 13311 14328 13323 14331
rect 15654 14328 15660 14340
rect 13311 14300 15660 14328
rect 13311 14297 13323 14300
rect 13265 14291 13323 14297
rect 15654 14288 15660 14300
rect 15712 14288 15718 14340
rect 17954 14288 17960 14340
rect 18012 14328 18018 14340
rect 19812 14328 19840 14359
rect 18012 14300 19840 14328
rect 18012 14288 18018 14300
rect 9677 14263 9735 14269
rect 9677 14260 9689 14263
rect 9640 14232 9689 14260
rect 9640 14220 9646 14232
rect 9677 14229 9689 14232
rect 9723 14229 9735 14263
rect 9677 14223 9735 14229
rect 10597 14263 10655 14269
rect 10597 14229 10609 14263
rect 10643 14260 10655 14263
rect 11146 14260 11152 14272
rect 10643 14232 11152 14260
rect 10643 14229 10655 14232
rect 10597 14223 10655 14229
rect 11146 14220 11152 14232
rect 11204 14220 11210 14272
rect 11241 14263 11299 14269
rect 11241 14229 11253 14263
rect 11287 14260 11299 14263
rect 11882 14260 11888 14272
rect 11287 14232 11888 14260
rect 11287 14229 11299 14232
rect 11241 14223 11299 14229
rect 11882 14220 11888 14232
rect 11940 14220 11946 14272
rect 13354 14220 13360 14272
rect 13412 14260 13418 14272
rect 15930 14260 15936 14272
rect 13412 14232 15936 14260
rect 13412 14220 13418 14232
rect 15930 14220 15936 14232
rect 15988 14220 15994 14272
rect 16669 14263 16727 14269
rect 16669 14229 16681 14263
rect 16715 14260 16727 14263
rect 18138 14260 18144 14272
rect 16715 14232 18144 14260
rect 16715 14229 16727 14232
rect 16669 14223 16727 14229
rect 18138 14220 18144 14232
rect 18196 14220 18202 14272
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 3142 14016 3148 14068
rect 3200 14056 3206 14068
rect 9674 14056 9680 14068
rect 3200 14028 8984 14056
rect 9635 14028 9680 14056
rect 3200 14016 3206 14028
rect 3786 13948 3792 14000
rect 3844 13988 3850 14000
rect 5445 13991 5503 13997
rect 5445 13988 5457 13991
rect 3844 13960 5457 13988
rect 3844 13948 3850 13960
rect 5445 13957 5457 13960
rect 5491 13957 5503 13991
rect 8846 13988 8852 14000
rect 8759 13960 8852 13988
rect 5445 13951 5503 13957
rect 8846 13948 8852 13960
rect 8904 13948 8910 14000
rect 8956 13988 8984 14028
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 11425 14059 11483 14065
rect 11425 14056 11437 14059
rect 9784 14028 11437 14056
rect 9784 13988 9812 14028
rect 11425 14025 11437 14028
rect 11471 14025 11483 14059
rect 11425 14019 11483 14025
rect 11790 14016 11796 14068
rect 11848 14056 11854 14068
rect 17037 14059 17095 14065
rect 17037 14056 17049 14059
rect 11848 14028 17049 14056
rect 11848 14016 11854 14028
rect 17037 14025 17049 14028
rect 17083 14025 17095 14059
rect 20806 14056 20812 14068
rect 20767 14028 20812 14056
rect 17037 14019 17095 14025
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 13906 13988 13912 14000
rect 8956 13960 9812 13988
rect 12636 13960 13912 13988
rect 4062 13880 4068 13932
rect 4120 13920 4126 13932
rect 4157 13923 4215 13929
rect 4157 13920 4169 13923
rect 4120 13892 4169 13920
rect 4120 13880 4126 13892
rect 4157 13889 4169 13892
rect 4203 13889 4215 13923
rect 4157 13883 4215 13889
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13920 4399 13923
rect 5166 13920 5172 13932
rect 4387 13892 5172 13920
rect 4387 13889 4399 13892
rect 4341 13883 4399 13889
rect 1486 13852 1492 13864
rect 1447 13824 1492 13852
rect 1486 13812 1492 13824
rect 1544 13812 1550 13864
rect 1756 13855 1814 13861
rect 1756 13821 1768 13855
rect 1802 13852 1814 13855
rect 4356 13852 4384 13883
rect 5166 13880 5172 13892
rect 5224 13880 5230 13932
rect 8864 13920 8892 13948
rect 10229 13923 10287 13929
rect 10229 13920 10241 13923
rect 8864 13892 10241 13920
rect 10229 13889 10241 13892
rect 10275 13889 10287 13923
rect 12636 13920 12664 13960
rect 13906 13948 13912 13960
rect 13964 13948 13970 14000
rect 14090 13948 14096 14000
rect 14148 13988 14154 14000
rect 14148 13960 14688 13988
rect 14148 13948 14154 13960
rect 10229 13883 10287 13889
rect 10336 13892 12664 13920
rect 1802 13824 4384 13852
rect 5261 13855 5319 13861
rect 1802 13821 1814 13824
rect 1756 13815 1814 13821
rect 5261 13821 5273 13855
rect 5307 13821 5319 13855
rect 7466 13852 7472 13864
rect 7427 13824 7472 13852
rect 5261 13815 5319 13821
rect 4065 13787 4123 13793
rect 4065 13753 4077 13787
rect 4111 13784 4123 13787
rect 4154 13784 4160 13796
rect 4111 13756 4160 13784
rect 4111 13753 4123 13756
rect 4065 13747 4123 13753
rect 4154 13744 4160 13756
rect 4212 13744 4218 13796
rect 2866 13716 2872 13728
rect 2827 13688 2872 13716
rect 2866 13676 2872 13688
rect 2924 13676 2930 13728
rect 3234 13676 3240 13728
rect 3292 13716 3298 13728
rect 3697 13719 3755 13725
rect 3697 13716 3709 13719
rect 3292 13688 3709 13716
rect 3292 13676 3298 13688
rect 3697 13685 3709 13688
rect 3743 13685 3755 13719
rect 5276 13716 5304 13815
rect 7466 13812 7472 13824
rect 7524 13812 7530 13864
rect 10336 13852 10364 13892
rect 12710 13880 12716 13932
rect 12768 13920 12774 13932
rect 13541 13923 13599 13929
rect 13541 13920 13553 13923
rect 12768 13892 13553 13920
rect 12768 13880 12774 13892
rect 13541 13889 13553 13892
rect 13587 13889 13599 13923
rect 13541 13883 13599 13889
rect 13725 13923 13783 13929
rect 13725 13889 13737 13923
rect 13771 13920 13783 13923
rect 14458 13920 14464 13932
rect 13771 13892 14464 13920
rect 13771 13889 13783 13892
rect 13725 13883 13783 13889
rect 14458 13880 14464 13892
rect 14516 13880 14522 13932
rect 14660 13929 14688 13960
rect 15930 13948 15936 14000
rect 15988 13988 15994 14000
rect 19334 13988 19340 14000
rect 15988 13960 19340 13988
rect 15988 13948 15994 13960
rect 19334 13948 19340 13960
rect 19392 13948 19398 14000
rect 14645 13923 14703 13929
rect 14645 13889 14657 13923
rect 14691 13889 14703 13923
rect 14645 13883 14703 13889
rect 19150 13880 19156 13932
rect 19208 13920 19214 13932
rect 19208 13892 19564 13920
rect 19208 13880 19214 13892
rect 7944 13824 10364 13852
rect 11241 13855 11299 13861
rect 7742 13793 7748 13796
rect 7736 13747 7748 13793
rect 7800 13784 7806 13796
rect 7800 13756 7836 13784
rect 7742 13744 7748 13747
rect 7800 13744 7806 13756
rect 7944 13716 7972 13824
rect 11241 13821 11253 13855
rect 11287 13852 11299 13855
rect 11287 13824 12388 13852
rect 11287 13821 11299 13824
rect 11241 13815 11299 13821
rect 9398 13744 9404 13796
rect 9456 13784 9462 13796
rect 10137 13787 10195 13793
rect 10137 13784 10149 13787
rect 9456 13756 10149 13784
rect 9456 13744 9462 13756
rect 10137 13753 10149 13756
rect 10183 13753 10195 13787
rect 12360 13784 12388 13824
rect 13354 13812 13360 13864
rect 13412 13852 13418 13864
rect 14090 13852 14096 13864
rect 13412 13824 14096 13852
rect 13412 13812 13418 13824
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 14912 13855 14970 13861
rect 14912 13821 14924 13855
rect 14958 13852 14970 13855
rect 16022 13852 16028 13864
rect 14958 13824 16028 13852
rect 14958 13821 14970 13824
rect 14912 13815 14970 13821
rect 16022 13812 16028 13824
rect 16080 13812 16086 13864
rect 16114 13812 16120 13864
rect 16172 13812 16178 13864
rect 16850 13852 16856 13864
rect 16811 13824 16856 13852
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 17034 13812 17040 13864
rect 17092 13852 17098 13864
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 17092 13824 18061 13852
rect 17092 13812 17098 13824
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 18230 13812 18236 13864
rect 18288 13852 18294 13864
rect 19429 13855 19487 13861
rect 18288 13824 19380 13852
rect 18288 13812 18294 13824
rect 15194 13784 15200 13796
rect 12360 13756 15200 13784
rect 10137 13747 10195 13753
rect 15194 13744 15200 13756
rect 15252 13744 15258 13796
rect 5276 13688 7972 13716
rect 3697 13679 3755 13685
rect 8662 13676 8668 13728
rect 8720 13716 8726 13728
rect 9766 13716 9772 13728
rect 8720 13688 9772 13716
rect 8720 13676 8726 13688
rect 9766 13676 9772 13688
rect 9824 13676 9830 13728
rect 10042 13716 10048 13728
rect 10003 13688 10048 13716
rect 10042 13676 10048 13688
rect 10100 13716 10106 13728
rect 10318 13716 10324 13728
rect 10100 13688 10324 13716
rect 10100 13676 10106 13688
rect 10318 13676 10324 13688
rect 10376 13676 10382 13728
rect 10778 13676 10784 13728
rect 10836 13716 10842 13728
rect 12618 13716 12624 13728
rect 10836 13688 12624 13716
rect 10836 13676 10842 13688
rect 12618 13676 12624 13688
rect 12676 13676 12682 13728
rect 13081 13719 13139 13725
rect 13081 13685 13093 13719
rect 13127 13716 13139 13719
rect 13354 13716 13360 13728
rect 13127 13688 13360 13716
rect 13127 13685 13139 13688
rect 13081 13679 13139 13685
rect 13354 13676 13360 13688
rect 13412 13676 13418 13728
rect 13449 13719 13507 13725
rect 13449 13685 13461 13719
rect 13495 13716 13507 13719
rect 15470 13716 15476 13728
rect 13495 13688 15476 13716
rect 13495 13685 13507 13688
rect 13449 13679 13507 13685
rect 15470 13676 15476 13688
rect 15528 13676 15534 13728
rect 16025 13719 16083 13725
rect 16025 13685 16037 13719
rect 16071 13716 16083 13719
rect 16132 13716 16160 13812
rect 17954 13744 17960 13796
rect 18012 13784 18018 13796
rect 18325 13787 18383 13793
rect 18325 13784 18337 13787
rect 18012 13756 18337 13784
rect 18012 13744 18018 13756
rect 18325 13753 18337 13756
rect 18371 13753 18383 13787
rect 19352 13784 19380 13824
rect 19429 13821 19441 13855
rect 19475 13821 19487 13855
rect 19536 13852 19564 13892
rect 19685 13855 19743 13861
rect 19685 13852 19697 13855
rect 19536 13824 19697 13852
rect 19429 13815 19487 13821
rect 19685 13821 19697 13824
rect 19731 13821 19743 13855
rect 19685 13815 19743 13821
rect 19444 13784 19472 13815
rect 19352 13756 19472 13784
rect 18325 13747 18383 13753
rect 16071 13688 16160 13716
rect 16071 13685 16083 13688
rect 16025 13679 16083 13685
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 3970 13472 3976 13524
rect 4028 13512 4034 13524
rect 7742 13512 7748 13524
rect 4028 13484 6776 13512
rect 7703 13484 7748 13512
rect 4028 13472 4034 13484
rect 2314 13444 2320 13456
rect 2275 13416 2320 13444
rect 2314 13404 2320 13416
rect 2372 13404 2378 13456
rect 2406 13404 2412 13456
rect 2464 13444 2470 13456
rect 4433 13447 4491 13453
rect 4433 13444 4445 13447
rect 2464 13416 4445 13444
rect 2464 13404 2470 13416
rect 4433 13413 4445 13416
rect 4479 13413 4491 13447
rect 4433 13407 4491 13413
rect 6362 13404 6368 13456
rect 6420 13444 6426 13456
rect 6610 13447 6668 13453
rect 6610 13444 6622 13447
rect 6420 13416 6622 13444
rect 6420 13404 6426 13416
rect 6610 13413 6622 13416
rect 6656 13413 6668 13447
rect 6610 13407 6668 13413
rect 2041 13379 2099 13385
rect 2041 13345 2053 13379
rect 2087 13376 2099 13379
rect 2774 13376 2780 13388
rect 2087 13348 2780 13376
rect 2087 13345 2099 13348
rect 2041 13339 2099 13345
rect 2774 13336 2780 13348
rect 2832 13336 2838 13388
rect 4338 13336 4344 13388
rect 4396 13376 4402 13388
rect 4525 13379 4583 13385
rect 4525 13376 4537 13379
rect 4396 13348 4537 13376
rect 4396 13336 4402 13348
rect 4525 13345 4537 13348
rect 4571 13345 4583 13379
rect 4525 13339 4583 13345
rect 5997 13379 6055 13385
rect 5997 13345 6009 13379
rect 6043 13376 6055 13379
rect 6454 13376 6460 13388
rect 6043 13348 6460 13376
rect 6043 13345 6055 13348
rect 5997 13339 6055 13345
rect 6454 13336 6460 13348
rect 6512 13336 6518 13388
rect 6748 13376 6776 13484
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 8573 13515 8631 13521
rect 8573 13481 8585 13515
rect 8619 13512 8631 13515
rect 8938 13512 8944 13524
rect 8619 13484 8944 13512
rect 8619 13481 8631 13484
rect 8573 13475 8631 13481
rect 8938 13472 8944 13484
rect 8996 13472 9002 13524
rect 9306 13472 9312 13524
rect 9364 13512 9370 13524
rect 11790 13512 11796 13524
rect 9364 13484 11796 13512
rect 9364 13472 9370 13484
rect 11790 13472 11796 13484
rect 11848 13472 11854 13524
rect 11885 13515 11943 13521
rect 11885 13481 11897 13515
rect 11931 13481 11943 13515
rect 12342 13512 12348 13524
rect 12303 13484 12348 13512
rect 11885 13475 11943 13481
rect 6822 13404 6828 13456
rect 6880 13444 6886 13456
rect 9766 13444 9772 13456
rect 6880 13416 9772 13444
rect 6880 13404 6886 13416
rect 9766 13404 9772 13416
rect 9824 13404 9830 13456
rect 9858 13404 9864 13456
rect 9916 13453 9922 13456
rect 9916 13447 9980 13453
rect 9916 13413 9934 13447
rect 9968 13413 9980 13447
rect 11900 13444 11928 13475
rect 12342 13472 12348 13484
rect 12400 13472 12406 13524
rect 17310 13472 17316 13524
rect 17368 13512 17374 13524
rect 17862 13512 17868 13524
rect 17368 13484 17868 13512
rect 17368 13472 17374 13484
rect 17862 13472 17868 13484
rect 17920 13512 17926 13524
rect 18141 13515 18199 13521
rect 18141 13512 18153 13515
rect 17920 13484 18153 13512
rect 17920 13472 17926 13484
rect 18141 13481 18153 13484
rect 18187 13481 18199 13515
rect 18966 13512 18972 13524
rect 18927 13484 18972 13512
rect 18141 13475 18199 13481
rect 18966 13472 18972 13484
rect 19024 13472 19030 13524
rect 19337 13515 19395 13521
rect 19337 13481 19349 13515
rect 19383 13512 19395 13515
rect 19978 13512 19984 13524
rect 19383 13484 19984 13512
rect 19383 13481 19395 13484
rect 19337 13475 19395 13481
rect 19978 13472 19984 13484
rect 20036 13472 20042 13524
rect 9916 13407 9980 13413
rect 11808 13416 11928 13444
rect 9916 13404 9922 13407
rect 6748 13348 10732 13376
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13308 4767 13311
rect 5166 13308 5172 13320
rect 4755 13280 5172 13308
rect 4755 13277 4767 13280
rect 4709 13271 4767 13277
rect 5166 13268 5172 13280
rect 5224 13268 5230 13320
rect 6365 13311 6423 13317
rect 6365 13277 6377 13311
rect 6411 13277 6423 13311
rect 6365 13271 6423 13277
rect 5813 13243 5871 13249
rect 5813 13209 5825 13243
rect 5859 13240 5871 13243
rect 6178 13240 6184 13252
rect 5859 13212 6184 13240
rect 5859 13209 5871 13212
rect 5813 13203 5871 13209
rect 6178 13200 6184 13212
rect 6236 13240 6242 13252
rect 6380 13240 6408 13271
rect 8662 13268 8668 13320
rect 8720 13308 8726 13320
rect 9214 13308 9220 13320
rect 8720 13280 9220 13308
rect 8720 13268 8726 13280
rect 9214 13268 9220 13280
rect 9272 13268 9278 13320
rect 9306 13268 9312 13320
rect 9364 13308 9370 13320
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 9364 13280 9689 13308
rect 9364 13268 9370 13280
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 9677 13271 9735 13277
rect 6236 13212 6408 13240
rect 10704 13240 10732 13348
rect 11808 13320 11836 13416
rect 12618 13404 12624 13456
rect 12676 13444 12682 13456
rect 12894 13444 12900 13456
rect 12676 13416 12900 13444
rect 12676 13404 12682 13416
rect 12894 13404 12900 13416
rect 12952 13404 12958 13456
rect 13538 13404 13544 13456
rect 13596 13444 13602 13456
rect 14093 13447 14151 13453
rect 14093 13444 14105 13447
rect 13596 13416 14105 13444
rect 13596 13404 13602 13416
rect 14093 13413 14105 13416
rect 14139 13413 14151 13447
rect 14093 13407 14151 13413
rect 15565 13447 15623 13453
rect 15565 13413 15577 13447
rect 15611 13444 15623 13447
rect 16850 13444 16856 13456
rect 15611 13416 16856 13444
rect 15611 13413 15623 13416
rect 15565 13407 15623 13413
rect 16850 13404 16856 13416
rect 16908 13404 16914 13456
rect 18230 13444 18236 13456
rect 16960 13416 18236 13444
rect 12253 13379 12311 13385
rect 12253 13345 12265 13379
rect 12299 13376 12311 13379
rect 12342 13376 12348 13388
rect 12299 13348 12348 13376
rect 12299 13345 12311 13348
rect 12253 13339 12311 13345
rect 12342 13336 12348 13348
rect 12400 13336 12406 13388
rect 14001 13379 14059 13385
rect 14001 13376 14013 13379
rect 12452 13348 14013 13376
rect 11790 13268 11796 13320
rect 11848 13268 11854 13320
rect 12452 13240 12480 13348
rect 14001 13345 14013 13348
rect 14047 13345 14059 13379
rect 14001 13339 14059 13345
rect 15289 13379 15347 13385
rect 15289 13345 15301 13379
rect 15335 13376 15347 13379
rect 15930 13376 15936 13388
rect 15335 13348 15936 13376
rect 15335 13345 15347 13348
rect 15289 13339 15347 13345
rect 15930 13336 15936 13348
rect 15988 13336 15994 13388
rect 16482 13336 16488 13388
rect 16540 13376 16546 13388
rect 16758 13376 16764 13388
rect 16540 13348 16764 13376
rect 16540 13336 16546 13348
rect 16758 13336 16764 13348
rect 16816 13376 16822 13388
rect 16960 13376 16988 13416
rect 18230 13404 18236 13416
rect 18288 13404 18294 13456
rect 18874 13404 18880 13456
rect 18932 13444 18938 13456
rect 18932 13416 19656 13444
rect 18932 13404 18938 13416
rect 16816 13348 16988 13376
rect 17028 13379 17086 13385
rect 16816 13336 16822 13348
rect 17028 13345 17040 13379
rect 17074 13376 17086 13379
rect 18892 13376 18920 13404
rect 17074 13348 18920 13376
rect 17074 13345 17086 13348
rect 17028 13339 17086 13345
rect 12529 13311 12587 13317
rect 12529 13277 12541 13311
rect 12575 13308 12587 13311
rect 12802 13308 12808 13320
rect 12575 13280 12808 13308
rect 12575 13277 12587 13280
rect 12529 13271 12587 13277
rect 12802 13268 12808 13280
rect 12860 13268 12866 13320
rect 14277 13311 14335 13317
rect 14277 13277 14289 13311
rect 14323 13308 14335 13311
rect 14458 13308 14464 13320
rect 14323 13280 14464 13308
rect 14323 13277 14335 13280
rect 14277 13271 14335 13277
rect 14458 13268 14464 13280
rect 14516 13308 14522 13320
rect 15654 13308 15660 13320
rect 14516 13280 15660 13308
rect 14516 13268 14522 13280
rect 15654 13268 15660 13280
rect 15712 13268 15718 13320
rect 19628 13317 19656 13416
rect 19429 13311 19487 13317
rect 19429 13277 19441 13311
rect 19475 13277 19487 13311
rect 19429 13271 19487 13277
rect 19613 13311 19671 13317
rect 19613 13277 19625 13311
rect 19659 13308 19671 13311
rect 20162 13308 20168 13320
rect 19659 13280 20168 13308
rect 19659 13277 19671 13280
rect 19613 13271 19671 13277
rect 10704 13212 12480 13240
rect 6236 13200 6242 13212
rect 12894 13200 12900 13252
rect 12952 13240 12958 13252
rect 13262 13240 13268 13252
rect 12952 13212 13268 13240
rect 12952 13200 12958 13212
rect 13262 13200 13268 13212
rect 13320 13200 13326 13252
rect 3142 13132 3148 13184
rect 3200 13172 3206 13184
rect 4065 13175 4123 13181
rect 4065 13172 4077 13175
rect 3200 13144 4077 13172
rect 3200 13132 3206 13144
rect 4065 13141 4077 13144
rect 4111 13141 4123 13175
rect 4065 13135 4123 13141
rect 4154 13132 4160 13184
rect 4212 13172 4218 13184
rect 5350 13172 5356 13184
rect 4212 13144 5356 13172
rect 4212 13132 4218 13144
rect 5350 13132 5356 13144
rect 5408 13132 5414 13184
rect 5718 13132 5724 13184
rect 5776 13172 5782 13184
rect 8202 13172 8208 13184
rect 5776 13144 8208 13172
rect 5776 13132 5782 13144
rect 8202 13132 8208 13144
rect 8260 13132 8266 13184
rect 10042 13132 10048 13184
rect 10100 13172 10106 13184
rect 11057 13175 11115 13181
rect 11057 13172 11069 13175
rect 10100 13144 11069 13172
rect 10100 13132 10106 13144
rect 11057 13141 11069 13144
rect 11103 13172 11115 13175
rect 11882 13172 11888 13184
rect 11103 13144 11888 13172
rect 11103 13141 11115 13144
rect 11057 13135 11115 13141
rect 11882 13132 11888 13144
rect 11940 13132 11946 13184
rect 13633 13175 13691 13181
rect 13633 13141 13645 13175
rect 13679 13172 13691 13175
rect 13998 13172 14004 13184
rect 13679 13144 14004 13172
rect 13679 13141 13691 13144
rect 13633 13135 13691 13141
rect 13998 13132 14004 13144
rect 14056 13132 14062 13184
rect 14458 13132 14464 13184
rect 14516 13172 14522 13184
rect 19444 13172 19472 13271
rect 20162 13268 20168 13280
rect 20220 13268 20226 13320
rect 14516 13144 19472 13172
rect 14516 13132 14522 13144
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 2774 12928 2780 12980
rect 2832 12968 2838 12980
rect 4338 12968 4344 12980
rect 2832 12940 2877 12968
rect 4299 12940 4344 12968
rect 2832 12928 2838 12940
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 6457 12971 6515 12977
rect 6457 12937 6469 12971
rect 6503 12968 6515 12971
rect 6638 12968 6644 12980
rect 6503 12940 6644 12968
rect 6503 12937 6515 12940
rect 6457 12931 6515 12937
rect 6638 12928 6644 12940
rect 6696 12928 6702 12980
rect 6822 12968 6828 12980
rect 6783 12940 6828 12968
rect 6822 12928 6828 12940
rect 6880 12928 6886 12980
rect 7190 12928 7196 12980
rect 7248 12968 7254 12980
rect 9214 12968 9220 12980
rect 7248 12940 9220 12968
rect 7248 12928 7254 12940
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 9953 12971 10011 12977
rect 9953 12937 9965 12971
rect 9999 12968 10011 12971
rect 10778 12968 10784 12980
rect 9999 12940 10784 12968
rect 9999 12937 10011 12940
rect 9953 12931 10011 12937
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 11238 12928 11244 12980
rect 11296 12968 11302 12980
rect 11517 12971 11575 12977
rect 11517 12968 11529 12971
rect 11296 12940 11529 12968
rect 11296 12928 11302 12940
rect 11517 12937 11529 12940
rect 11563 12937 11575 12971
rect 11517 12931 11575 12937
rect 2866 12860 2872 12912
rect 2924 12900 2930 12912
rect 2924 12872 3372 12900
rect 2924 12860 2930 12872
rect 2590 12792 2596 12844
rect 2648 12832 2654 12844
rect 2774 12832 2780 12844
rect 2648 12804 2780 12832
rect 2648 12792 2654 12804
rect 2774 12792 2780 12804
rect 2832 12792 2838 12844
rect 3234 12832 3240 12844
rect 3195 12804 3240 12832
rect 3234 12792 3240 12804
rect 3292 12792 3298 12844
rect 3344 12841 3372 12872
rect 4430 12860 4436 12912
rect 4488 12900 4494 12912
rect 9858 12900 9864 12912
rect 4488 12872 9864 12900
rect 4488 12860 4494 12872
rect 9858 12860 9864 12872
rect 9916 12860 9922 12912
rect 3329 12835 3387 12841
rect 3329 12801 3341 12835
rect 3375 12801 3387 12835
rect 3329 12795 3387 12801
rect 4522 12792 4528 12844
rect 4580 12832 4586 12844
rect 4893 12835 4951 12841
rect 4893 12832 4905 12835
rect 4580 12804 4905 12832
rect 4580 12792 4586 12804
rect 4893 12801 4905 12804
rect 4939 12832 4951 12835
rect 4982 12832 4988 12844
rect 4939 12804 4988 12832
rect 4939 12801 4951 12804
rect 4893 12795 4951 12801
rect 4982 12792 4988 12804
rect 5040 12792 5046 12844
rect 7282 12832 7288 12844
rect 7243 12804 7288 12832
rect 7282 12792 7288 12804
rect 7340 12792 7346 12844
rect 7469 12835 7527 12841
rect 7469 12801 7481 12835
rect 7515 12832 7527 12835
rect 7742 12832 7748 12844
rect 7515 12804 7748 12832
rect 7515 12801 7527 12804
rect 7469 12795 7527 12801
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 8202 12792 8208 12844
rect 8260 12832 8266 12844
rect 8941 12835 8999 12841
rect 8941 12832 8953 12835
rect 8260 12804 8953 12832
rect 8260 12792 8266 12804
rect 8941 12801 8953 12804
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 9306 12792 9312 12844
rect 9364 12832 9370 12844
rect 10134 12832 10140 12844
rect 9364 12804 10140 12832
rect 9364 12792 9370 12804
rect 10134 12792 10140 12804
rect 10192 12792 10198 12844
rect 11532 12832 11560 12931
rect 11882 12928 11888 12980
rect 11940 12968 11946 12980
rect 11940 12940 20208 12968
rect 11940 12928 11946 12940
rect 13630 12860 13636 12912
rect 13688 12900 13694 12912
rect 13817 12903 13875 12909
rect 13817 12900 13829 12903
rect 13688 12872 13829 12900
rect 13688 12860 13694 12872
rect 13817 12869 13829 12872
rect 13863 12869 13875 12903
rect 16022 12900 16028 12912
rect 15983 12872 16028 12900
rect 13817 12863 13875 12869
rect 16022 12860 16028 12872
rect 16080 12860 16086 12912
rect 17034 12900 17040 12912
rect 16995 12872 17040 12900
rect 17034 12860 17040 12872
rect 17092 12860 17098 12912
rect 17770 12860 17776 12912
rect 17828 12900 17834 12912
rect 18049 12903 18107 12909
rect 18049 12900 18061 12903
rect 17828 12872 18061 12900
rect 17828 12860 17834 12872
rect 18049 12869 18061 12872
rect 18095 12869 18107 12903
rect 18049 12863 18107 12869
rect 18598 12832 18604 12844
rect 11532 12804 12572 12832
rect 18559 12804 18604 12832
rect 1679 12767 1737 12773
rect 1679 12733 1691 12767
rect 1725 12733 1737 12767
rect 3142 12764 3148 12776
rect 3103 12736 3148 12764
rect 1679 12727 1737 12733
rect 1688 12696 1716 12727
rect 3142 12724 3148 12736
rect 3200 12724 3206 12776
rect 6641 12767 6699 12773
rect 6641 12733 6653 12767
rect 6687 12764 6699 12767
rect 8757 12767 8815 12773
rect 6687 12736 8708 12764
rect 6687 12733 6699 12736
rect 6641 12727 6699 12733
rect 5350 12696 5356 12708
rect 1688 12668 5356 12696
rect 5350 12656 5356 12668
rect 5408 12656 5414 12708
rect 7193 12699 7251 12705
rect 7193 12665 7205 12699
rect 7239 12696 7251 12699
rect 8680 12696 8708 12736
rect 8757 12733 8769 12767
rect 8803 12764 8815 12767
rect 9953 12767 10011 12773
rect 9953 12764 9965 12767
rect 8803 12736 9965 12764
rect 8803 12733 8815 12736
rect 8757 12727 8815 12733
rect 9953 12733 9965 12736
rect 9999 12733 10011 12767
rect 9953 12727 10011 12733
rect 10042 12724 10048 12776
rect 10100 12764 10106 12776
rect 10393 12767 10451 12773
rect 10393 12764 10405 12767
rect 10100 12736 10405 12764
rect 10100 12724 10106 12736
rect 10393 12733 10405 12736
rect 10439 12733 10451 12767
rect 12434 12764 12440 12776
rect 12347 12736 12440 12764
rect 10393 12727 10451 12733
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 12544 12764 12572 12804
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 20180 12841 20208 12940
rect 20165 12835 20223 12841
rect 20165 12801 20177 12835
rect 20211 12801 20223 12835
rect 20165 12795 20223 12801
rect 12693 12767 12751 12773
rect 12693 12764 12705 12767
rect 12544 12736 12705 12764
rect 12693 12733 12705 12736
rect 12739 12733 12751 12767
rect 12693 12727 12751 12733
rect 14645 12767 14703 12773
rect 14645 12733 14657 12767
rect 14691 12733 14703 12767
rect 14645 12727 14703 12733
rect 16853 12767 16911 12773
rect 16853 12733 16865 12767
rect 16899 12764 16911 12767
rect 17954 12764 17960 12776
rect 16899 12736 17960 12764
rect 16899 12733 16911 12736
rect 16853 12727 16911 12733
rect 7239 12668 8432 12696
rect 8680 12668 9536 12696
rect 7239 12665 7251 12668
rect 7193 12659 7251 12665
rect 1857 12631 1915 12637
rect 1857 12597 1869 12631
rect 1903 12628 1915 12631
rect 2958 12628 2964 12640
rect 1903 12600 2964 12628
rect 1903 12597 1915 12600
rect 1857 12591 1915 12597
rect 2958 12588 2964 12600
rect 3016 12588 3022 12640
rect 3142 12588 3148 12640
rect 3200 12628 3206 12640
rect 3418 12628 3424 12640
rect 3200 12600 3424 12628
rect 3200 12588 3206 12600
rect 3418 12588 3424 12600
rect 3476 12588 3482 12640
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4338 12628 4344 12640
rect 4212 12600 4344 12628
rect 4212 12588 4218 12600
rect 4338 12588 4344 12600
rect 4396 12628 4402 12640
rect 4709 12631 4767 12637
rect 4709 12628 4721 12631
rect 4396 12600 4721 12628
rect 4396 12588 4402 12600
rect 4709 12597 4721 12600
rect 4755 12597 4767 12631
rect 4709 12591 4767 12597
rect 4801 12631 4859 12637
rect 4801 12597 4813 12631
rect 4847 12628 4859 12631
rect 5166 12628 5172 12640
rect 4847 12600 5172 12628
rect 4847 12597 4859 12600
rect 4801 12591 4859 12597
rect 5166 12588 5172 12600
rect 5224 12628 5230 12640
rect 8294 12628 8300 12640
rect 5224 12600 8300 12628
rect 5224 12588 5230 12600
rect 8294 12588 8300 12600
rect 8352 12588 8358 12640
rect 8404 12637 8432 12668
rect 8389 12631 8447 12637
rect 8389 12597 8401 12631
rect 8435 12597 8447 12631
rect 8846 12628 8852 12640
rect 8807 12600 8852 12628
rect 8389 12591 8447 12597
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 9508 12628 9536 12668
rect 9582 12656 9588 12708
rect 9640 12696 9646 12708
rect 12452 12696 12480 12724
rect 14660 12696 14688 12727
rect 17954 12724 17960 12736
rect 18012 12724 18018 12776
rect 18138 12724 18144 12776
rect 18196 12764 18202 12776
rect 18509 12767 18567 12773
rect 18509 12764 18521 12767
rect 18196 12736 18521 12764
rect 18196 12724 18202 12736
rect 18509 12733 18521 12736
rect 18555 12733 18567 12767
rect 18509 12727 18567 12733
rect 19610 12724 19616 12776
rect 19668 12764 19674 12776
rect 20073 12767 20131 12773
rect 20073 12764 20085 12767
rect 19668 12736 20085 12764
rect 19668 12724 19674 12736
rect 20073 12733 20085 12736
rect 20119 12733 20131 12767
rect 20073 12727 20131 12733
rect 9640 12668 11652 12696
rect 12452 12668 14688 12696
rect 9640 12656 9646 12668
rect 9766 12628 9772 12640
rect 9508 12600 9772 12628
rect 9766 12588 9772 12600
rect 9824 12588 9830 12640
rect 11624 12628 11652 12668
rect 14734 12656 14740 12708
rect 14792 12696 14798 12708
rect 14890 12699 14948 12705
rect 14890 12696 14902 12699
rect 14792 12668 14902 12696
rect 14792 12656 14798 12668
rect 14890 12665 14902 12668
rect 14936 12665 14948 12699
rect 17218 12696 17224 12708
rect 14890 12659 14948 12665
rect 16500 12668 17224 12696
rect 16500 12628 16528 12668
rect 17218 12656 17224 12668
rect 17276 12656 17282 12708
rect 17402 12656 17408 12708
rect 17460 12696 17466 12708
rect 17770 12696 17776 12708
rect 17460 12668 17776 12696
rect 17460 12656 17466 12668
rect 17770 12656 17776 12668
rect 17828 12656 17834 12708
rect 18417 12699 18475 12705
rect 18417 12665 18429 12699
rect 18463 12696 18475 12699
rect 18966 12696 18972 12708
rect 18463 12668 18972 12696
rect 18463 12665 18475 12668
rect 18417 12659 18475 12665
rect 18966 12656 18972 12668
rect 19024 12656 19030 12708
rect 11624 12600 16528 12628
rect 16574 12588 16580 12640
rect 16632 12628 16638 12640
rect 19613 12631 19671 12637
rect 19613 12628 19625 12631
rect 16632 12600 19625 12628
rect 16632 12588 16638 12600
rect 19613 12597 19625 12600
rect 19659 12597 19671 12631
rect 19613 12591 19671 12597
rect 19702 12588 19708 12640
rect 19760 12628 19766 12640
rect 19981 12631 20039 12637
rect 19981 12628 19993 12631
rect 19760 12600 19993 12628
rect 19760 12588 19766 12600
rect 19981 12597 19993 12600
rect 20027 12597 20039 12631
rect 19981 12591 20039 12597
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 1302 12384 1308 12436
rect 1360 12424 1366 12436
rect 1762 12424 1768 12436
rect 1360 12396 1768 12424
rect 1360 12384 1366 12396
rect 1762 12384 1768 12396
rect 1820 12384 1826 12436
rect 2593 12427 2651 12433
rect 2593 12393 2605 12427
rect 2639 12424 2651 12427
rect 6365 12427 6423 12433
rect 6365 12424 6377 12427
rect 2639 12396 6377 12424
rect 2639 12393 2651 12396
rect 2593 12387 2651 12393
rect 6365 12393 6377 12396
rect 6411 12393 6423 12427
rect 6365 12387 6423 12393
rect 6454 12384 6460 12436
rect 6512 12424 6518 12436
rect 8202 12424 8208 12436
rect 6512 12396 8208 12424
rect 6512 12384 6518 12396
rect 8202 12384 8208 12396
rect 8260 12384 8266 12436
rect 8294 12384 8300 12436
rect 8352 12424 8358 12436
rect 8352 12396 8397 12424
rect 8352 12384 8358 12396
rect 9674 12384 9680 12436
rect 9732 12424 9738 12436
rect 10594 12424 10600 12436
rect 9732 12396 10600 12424
rect 9732 12384 9738 12396
rect 10594 12384 10600 12396
rect 10652 12384 10658 12436
rect 10962 12384 10968 12436
rect 11020 12424 11026 12436
rect 11606 12424 11612 12436
rect 11020 12396 11612 12424
rect 11020 12384 11026 12396
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 11701 12427 11759 12433
rect 11701 12393 11713 12427
rect 11747 12424 11759 12427
rect 11790 12424 11796 12436
rect 11747 12396 11796 12424
rect 11747 12393 11759 12396
rect 11701 12387 11759 12393
rect 11790 12384 11796 12396
rect 11848 12384 11854 12436
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 12897 12427 12955 12433
rect 12897 12424 12909 12427
rect 12492 12396 12909 12424
rect 12492 12384 12498 12396
rect 12897 12393 12909 12396
rect 12943 12393 12955 12427
rect 12897 12387 12955 12393
rect 14274 12384 14280 12436
rect 14332 12424 14338 12436
rect 15289 12427 15347 12433
rect 15289 12424 15301 12427
rect 14332 12396 15301 12424
rect 14332 12384 14338 12396
rect 15289 12393 15301 12396
rect 15335 12393 15347 12427
rect 15289 12387 15347 12393
rect 15470 12384 15476 12436
rect 15528 12424 15534 12436
rect 15528 12396 18736 12424
rect 15528 12384 15534 12396
rect 2038 12316 2044 12368
rect 2096 12356 2102 12368
rect 2682 12356 2688 12368
rect 2096 12328 2688 12356
rect 2096 12316 2102 12328
rect 2682 12316 2688 12328
rect 2740 12316 2746 12368
rect 4338 12316 4344 12368
rect 4396 12356 4402 12368
rect 4798 12356 4804 12368
rect 4396 12328 4804 12356
rect 4396 12316 4402 12328
rect 4798 12316 4804 12328
rect 4856 12316 4862 12368
rect 5074 12316 5080 12368
rect 5132 12356 5138 12368
rect 5626 12356 5632 12368
rect 5132 12328 5632 12356
rect 5132 12316 5138 12328
rect 5626 12316 5632 12328
rect 5684 12316 5690 12368
rect 5902 12316 5908 12368
rect 5960 12356 5966 12368
rect 5960 12328 8515 12356
rect 5960 12316 5966 12328
rect 2130 12248 2136 12300
rect 2188 12288 2194 12300
rect 2501 12291 2559 12297
rect 2501 12288 2513 12291
rect 2188 12260 2513 12288
rect 2188 12248 2194 12260
rect 2501 12257 2513 12260
rect 2547 12257 2559 12291
rect 2501 12251 2559 12257
rect 4157 12291 4215 12297
rect 4157 12257 4169 12291
rect 4203 12257 4215 12291
rect 4157 12251 4215 12257
rect 4424 12291 4482 12297
rect 4424 12257 4436 12291
rect 4470 12288 4482 12291
rect 5258 12288 5264 12300
rect 4470 12260 5264 12288
rect 4470 12257 4482 12260
rect 4424 12251 4482 12257
rect 2682 12220 2688 12232
rect 2643 12192 2688 12220
rect 2682 12180 2688 12192
rect 2740 12180 2746 12232
rect 2774 12180 2780 12232
rect 2832 12220 2838 12232
rect 3510 12220 3516 12232
rect 2832 12192 3516 12220
rect 2832 12180 2838 12192
rect 3510 12180 3516 12192
rect 3568 12180 3574 12232
rect 4172 12164 4200 12251
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 6733 12291 6791 12297
rect 6733 12288 6745 12291
rect 5460 12260 6745 12288
rect 5460 12232 5488 12260
rect 6733 12257 6745 12260
rect 6779 12257 6791 12291
rect 7006 12288 7012 12300
rect 6733 12251 6791 12257
rect 6840 12260 7012 12288
rect 5442 12180 5448 12232
rect 5500 12180 5506 12232
rect 6546 12180 6552 12232
rect 6604 12220 6610 12232
rect 6840 12229 6868 12260
rect 7006 12248 7012 12260
rect 7064 12248 7070 12300
rect 8386 12288 8392 12300
rect 7392 12260 8392 12288
rect 7392 12232 7420 12260
rect 8386 12248 8392 12260
rect 8444 12248 8450 12300
rect 6825 12223 6883 12229
rect 6825 12220 6837 12223
rect 6604 12192 6837 12220
rect 6604 12180 6610 12192
rect 6825 12189 6837 12192
rect 6871 12189 6883 12223
rect 6825 12183 6883 12189
rect 6917 12223 6975 12229
rect 6917 12189 6929 12223
rect 6963 12189 6975 12223
rect 6917 12183 6975 12189
rect 4154 12112 4160 12164
rect 4212 12112 4218 12164
rect 6086 12112 6092 12164
rect 6144 12152 6150 12164
rect 6932 12152 6960 12183
rect 7374 12180 7380 12232
rect 7432 12180 7438 12232
rect 8487 12229 8515 12328
rect 11974 12316 11980 12368
rect 12032 12356 12038 12368
rect 12158 12356 12164 12368
rect 12032 12328 12164 12356
rect 12032 12316 12038 12328
rect 12158 12316 12164 12328
rect 12216 12316 12222 12368
rect 12526 12316 12532 12368
rect 12584 12356 12590 12368
rect 13078 12356 13084 12368
rect 12584 12328 13084 12356
rect 12584 12316 12590 12328
rect 13078 12316 13084 12328
rect 13136 12316 13142 12368
rect 13256 12359 13314 12365
rect 13256 12325 13268 12359
rect 13302 12356 13314 12359
rect 13630 12356 13636 12368
rect 13302 12328 13636 12356
rect 13302 12325 13314 12328
rect 13256 12319 13314 12325
rect 13630 12316 13636 12328
rect 13688 12316 13694 12368
rect 17304 12359 17362 12365
rect 17304 12325 17316 12359
rect 17350 12356 17362 12359
rect 18138 12356 18144 12368
rect 17350 12328 18144 12356
rect 17350 12325 17362 12328
rect 17304 12319 17362 12325
rect 18138 12316 18144 12328
rect 18196 12356 18202 12368
rect 18598 12356 18604 12368
rect 18196 12328 18604 12356
rect 18196 12316 18202 12328
rect 18598 12316 18604 12328
rect 18656 12316 18662 12368
rect 18708 12356 18736 12396
rect 19242 12384 19248 12436
rect 19300 12424 19306 12436
rect 19705 12427 19763 12433
rect 19705 12424 19717 12427
rect 19300 12396 19717 12424
rect 19300 12384 19306 12396
rect 19705 12393 19717 12396
rect 19751 12393 19763 12427
rect 19705 12387 19763 12393
rect 19613 12359 19671 12365
rect 19613 12356 19625 12359
rect 18708 12328 19625 12356
rect 19613 12325 19625 12328
rect 19659 12325 19671 12359
rect 19613 12319 19671 12325
rect 10045 12291 10103 12297
rect 10045 12257 10057 12291
rect 10091 12288 10103 12291
rect 10778 12288 10784 12300
rect 10091 12260 10784 12288
rect 10091 12257 10103 12260
rect 10045 12251 10103 12257
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 11609 12291 11667 12297
rect 11609 12257 11621 12291
rect 11655 12288 11667 12291
rect 12434 12288 12440 12300
rect 11655 12260 12440 12288
rect 11655 12257 11667 12260
rect 11609 12251 11667 12257
rect 12434 12248 12440 12260
rect 12492 12248 12498 12300
rect 12912 12260 14044 12288
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 8662 12180 8668 12232
rect 8720 12220 8726 12232
rect 9674 12220 9680 12232
rect 8720 12192 9680 12220
rect 8720 12180 8726 12192
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 10137 12223 10195 12229
rect 10137 12189 10149 12223
rect 10183 12189 10195 12223
rect 10318 12220 10324 12232
rect 10231 12192 10324 12220
rect 10137 12183 10195 12189
rect 6144 12124 6960 12152
rect 6144 12112 6150 12124
rect 7834 12112 7840 12164
rect 7892 12152 7898 12164
rect 10042 12152 10048 12164
rect 7892 12124 10048 12152
rect 7892 12112 7898 12124
rect 10042 12112 10048 12124
rect 10100 12112 10106 12164
rect 10152 12152 10180 12183
rect 10318 12180 10324 12192
rect 10376 12220 10382 12232
rect 11793 12223 11851 12229
rect 11793 12220 11805 12223
rect 10376 12192 11805 12220
rect 10376 12180 10382 12192
rect 11793 12189 11805 12192
rect 11839 12189 11851 12223
rect 11793 12183 11851 12189
rect 12912 12152 12940 12260
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12189 13047 12223
rect 14016 12220 14044 12260
rect 15102 12248 15108 12300
rect 15160 12288 15166 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 15160 12260 15669 12288
rect 15160 12248 15166 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 16758 12248 16764 12300
rect 16816 12288 16822 12300
rect 17037 12291 17095 12297
rect 17037 12288 17049 12291
rect 16816 12260 17049 12288
rect 16816 12248 16822 12260
rect 17037 12257 17049 12260
rect 17083 12257 17095 12291
rect 17037 12251 17095 12257
rect 15286 12220 15292 12232
rect 14016 12192 15292 12220
rect 12989 12183 13047 12189
rect 10152 12124 12940 12152
rect 2133 12087 2191 12093
rect 2133 12053 2145 12087
rect 2179 12084 2191 12087
rect 2958 12084 2964 12096
rect 2179 12056 2964 12084
rect 2179 12053 2191 12056
rect 2133 12047 2191 12053
rect 2958 12044 2964 12056
rect 3016 12044 3022 12096
rect 3050 12044 3056 12096
rect 3108 12084 3114 12096
rect 3418 12084 3424 12096
rect 3108 12056 3424 12084
rect 3108 12044 3114 12056
rect 3418 12044 3424 12056
rect 3476 12044 3482 12096
rect 4338 12044 4344 12096
rect 4396 12084 4402 12096
rect 5537 12087 5595 12093
rect 5537 12084 5549 12087
rect 4396 12056 5549 12084
rect 4396 12044 4402 12056
rect 5537 12053 5549 12056
rect 5583 12053 5595 12087
rect 5537 12047 5595 12053
rect 7466 12044 7472 12096
rect 7524 12084 7530 12096
rect 7929 12087 7987 12093
rect 7929 12084 7941 12087
rect 7524 12056 7941 12084
rect 7524 12044 7530 12056
rect 7929 12053 7941 12056
rect 7975 12053 7987 12087
rect 7929 12047 7987 12053
rect 9677 12087 9735 12093
rect 9677 12053 9689 12087
rect 9723 12084 9735 12087
rect 11054 12084 11060 12096
rect 9723 12056 11060 12084
rect 9723 12053 9735 12056
rect 9677 12047 9735 12053
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 11241 12087 11299 12093
rect 11241 12053 11253 12087
rect 11287 12084 11299 12087
rect 11698 12084 11704 12096
rect 11287 12056 11704 12084
rect 11287 12053 11299 12056
rect 11241 12047 11299 12053
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 12897 12087 12955 12093
rect 12897 12053 12909 12087
rect 12943 12084 12955 12087
rect 13004 12084 13032 12183
rect 15286 12180 15292 12192
rect 15344 12180 15350 12232
rect 15749 12223 15807 12229
rect 15749 12189 15761 12223
rect 15795 12189 15807 12223
rect 15749 12183 15807 12189
rect 15933 12223 15991 12229
rect 15933 12189 15945 12223
rect 15979 12220 15991 12223
rect 16022 12220 16028 12232
rect 15979 12192 16028 12220
rect 15979 12189 15991 12192
rect 15933 12183 15991 12189
rect 15764 12152 15792 12183
rect 16022 12180 16028 12192
rect 16080 12180 16086 12232
rect 19797 12223 19855 12229
rect 19797 12220 19809 12223
rect 18616 12192 19809 12220
rect 13924 12124 15792 12152
rect 12943 12056 13032 12084
rect 12943 12053 12955 12056
rect 12897 12047 12955 12053
rect 13630 12044 13636 12096
rect 13688 12084 13694 12096
rect 13924 12084 13952 12124
rect 18616 12096 18644 12192
rect 19797 12189 19809 12192
rect 19843 12189 19855 12223
rect 19797 12183 19855 12189
rect 13688 12056 13952 12084
rect 14369 12087 14427 12093
rect 13688 12044 13694 12056
rect 14369 12053 14381 12087
rect 14415 12084 14427 12087
rect 15654 12084 15660 12096
rect 14415 12056 15660 12084
rect 14415 12053 14427 12056
rect 14369 12047 14427 12053
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 18417 12087 18475 12093
rect 18417 12053 18429 12087
rect 18463 12084 18475 12087
rect 18598 12084 18604 12096
rect 18463 12056 18604 12084
rect 18463 12053 18475 12056
rect 18417 12047 18475 12053
rect 18598 12044 18604 12056
rect 18656 12044 18662 12096
rect 19242 12084 19248 12096
rect 19203 12056 19248 12084
rect 19242 12044 19248 12056
rect 19300 12044 19306 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 3050 11840 3056 11892
rect 3108 11880 3114 11892
rect 3789 11883 3847 11889
rect 3789 11880 3801 11883
rect 3108 11852 3801 11880
rect 3108 11840 3114 11852
rect 3789 11849 3801 11852
rect 3835 11880 3847 11883
rect 6086 11880 6092 11892
rect 3835 11852 6092 11880
rect 3835 11849 3847 11852
rect 3789 11843 3847 11849
rect 6086 11840 6092 11852
rect 6144 11840 6150 11892
rect 7009 11883 7067 11889
rect 7009 11849 7021 11883
rect 7055 11880 7067 11883
rect 7282 11880 7288 11892
rect 7055 11852 7288 11880
rect 7055 11849 7067 11852
rect 7009 11843 7067 11849
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 7650 11840 7656 11892
rect 7708 11880 7714 11892
rect 7926 11880 7932 11892
rect 7708 11852 7932 11880
rect 7708 11840 7714 11852
rect 7926 11840 7932 11852
rect 7984 11840 7990 11892
rect 8202 11840 8208 11892
rect 8260 11880 8266 11892
rect 8573 11883 8631 11889
rect 8573 11880 8585 11883
rect 8260 11852 8585 11880
rect 8260 11840 8266 11852
rect 8573 11849 8585 11852
rect 8619 11849 8631 11883
rect 8573 11843 8631 11849
rect 9232 11852 11744 11880
rect 8754 11772 8760 11824
rect 8812 11812 8818 11824
rect 9232 11812 9260 11852
rect 8812 11784 9260 11812
rect 8812 11772 8818 11784
rect 1397 11747 1455 11753
rect 1397 11713 1409 11747
rect 1443 11744 1455 11747
rect 1443 11716 2544 11744
rect 1443 11713 1455 11716
rect 1397 11707 1455 11713
rect 1486 11636 1492 11688
rect 1544 11676 1550 11688
rect 2409 11679 2467 11685
rect 2409 11676 2421 11679
rect 1544 11648 2421 11676
rect 1544 11636 1550 11648
rect 2409 11645 2421 11648
rect 2455 11645 2467 11679
rect 2516 11676 2544 11716
rect 3510 11704 3516 11756
rect 3568 11744 3574 11756
rect 5169 11747 5227 11753
rect 5169 11744 5181 11747
rect 3568 11716 5181 11744
rect 3568 11704 3574 11716
rect 5169 11713 5181 11716
rect 5215 11713 5227 11747
rect 5169 11707 5227 11713
rect 5258 11704 5264 11756
rect 5316 11744 5322 11756
rect 7282 11744 7288 11756
rect 5316 11716 7288 11744
rect 5316 11704 5322 11716
rect 7282 11704 7288 11716
rect 7340 11704 7346 11756
rect 7466 11744 7472 11756
rect 7427 11716 7472 11744
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 7653 11747 7711 11753
rect 7653 11713 7665 11747
rect 7699 11744 7711 11747
rect 8018 11744 8024 11756
rect 7699 11716 8024 11744
rect 7699 11713 7711 11716
rect 7653 11707 7711 11713
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 8294 11704 8300 11756
rect 8352 11704 8358 11756
rect 9232 11753 9260 11784
rect 11716 11753 11744 11852
rect 12434 11840 12440 11892
rect 12492 11880 12498 11892
rect 14001 11883 14059 11889
rect 12492 11852 12537 11880
rect 12492 11840 12498 11852
rect 14001 11849 14013 11883
rect 14047 11880 14059 11883
rect 14047 11852 14136 11880
rect 14047 11849 14059 11852
rect 14001 11843 14059 11849
rect 14108 11812 14136 11852
rect 17954 11840 17960 11892
rect 18012 11880 18018 11892
rect 19058 11880 19064 11892
rect 18012 11852 19064 11880
rect 18012 11840 18018 11852
rect 19058 11840 19064 11852
rect 19116 11840 19122 11892
rect 14274 11812 14280 11824
rect 14108 11784 14280 11812
rect 14274 11772 14280 11784
rect 14332 11772 14338 11824
rect 16942 11772 16948 11824
rect 17000 11812 17006 11824
rect 17000 11784 20024 11812
rect 17000 11772 17006 11784
rect 9217 11747 9275 11753
rect 9217 11713 9229 11747
rect 9263 11713 9275 11747
rect 9217 11707 9275 11713
rect 11701 11747 11759 11753
rect 11701 11713 11713 11747
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 12526 11704 12532 11756
rect 12584 11704 12590 11756
rect 12802 11744 12808 11756
rect 12636 11716 12808 11744
rect 4890 11676 4896 11688
rect 2516 11648 4896 11676
rect 2409 11639 2467 11645
rect 2424 11540 2452 11639
rect 4890 11636 4896 11648
rect 4948 11636 4954 11688
rect 8312 11676 8340 11704
rect 8662 11676 8668 11688
rect 8312 11648 8668 11676
rect 8662 11636 8668 11648
rect 8720 11676 8726 11688
rect 9033 11679 9091 11685
rect 9033 11676 9045 11679
rect 8720 11648 9045 11676
rect 8720 11636 8726 11648
rect 9033 11645 9045 11648
rect 9079 11645 9091 11679
rect 9033 11639 9091 11645
rect 9306 11636 9312 11688
rect 9364 11676 9370 11688
rect 9674 11676 9680 11688
rect 9364 11648 9680 11676
rect 9364 11636 9370 11648
rect 9674 11636 9680 11648
rect 9732 11676 9738 11688
rect 9944 11679 10002 11685
rect 9732 11648 9825 11676
rect 9732 11636 9738 11648
rect 9944 11645 9956 11679
rect 9990 11676 10002 11679
rect 10318 11676 10324 11688
rect 9990 11648 10324 11676
rect 9990 11645 10002 11648
rect 9944 11639 10002 11645
rect 10318 11636 10324 11648
rect 10376 11636 10382 11688
rect 11054 11636 11060 11688
rect 11112 11676 11118 11688
rect 11422 11676 11428 11688
rect 11112 11648 11428 11676
rect 11112 11636 11118 11648
rect 11422 11636 11428 11648
rect 11480 11636 11486 11688
rect 11609 11679 11667 11685
rect 11609 11645 11621 11679
rect 11655 11676 11667 11679
rect 12544 11676 12572 11704
rect 11655 11648 12572 11676
rect 11655 11645 11667 11648
rect 11609 11639 11667 11645
rect 2676 11611 2734 11617
rect 2676 11577 2688 11611
rect 2722 11608 2734 11611
rect 2866 11608 2872 11620
rect 2722 11580 2872 11608
rect 2722 11577 2734 11580
rect 2676 11571 2734 11577
rect 2866 11568 2872 11580
rect 2924 11568 2930 11620
rect 4985 11611 5043 11617
rect 4985 11577 4997 11611
rect 5031 11608 5043 11611
rect 5258 11608 5264 11620
rect 5031 11580 5264 11608
rect 5031 11577 5043 11580
rect 4985 11571 5043 11577
rect 5258 11568 5264 11580
rect 5316 11568 5322 11620
rect 7377 11611 7435 11617
rect 7377 11577 7389 11611
rect 7423 11608 7435 11611
rect 7834 11608 7840 11620
rect 7423 11580 7840 11608
rect 7423 11577 7435 11580
rect 7377 11571 7435 11577
rect 7834 11568 7840 11580
rect 7892 11568 7898 11620
rect 8294 11568 8300 11620
rect 8352 11608 8358 11620
rect 11517 11611 11575 11617
rect 8352 11580 11192 11608
rect 8352 11568 8358 11580
rect 4154 11540 4160 11552
rect 2424 11512 4160 11540
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 4617 11543 4675 11549
rect 4617 11509 4629 11543
rect 4663 11540 4675 11543
rect 4798 11540 4804 11552
rect 4663 11512 4804 11540
rect 4663 11509 4675 11512
rect 4617 11503 4675 11509
rect 4798 11500 4804 11512
rect 4856 11500 4862 11552
rect 5077 11543 5135 11549
rect 5077 11509 5089 11543
rect 5123 11540 5135 11543
rect 5166 11540 5172 11552
rect 5123 11512 5172 11540
rect 5123 11509 5135 11512
rect 5077 11503 5135 11509
rect 5166 11500 5172 11512
rect 5224 11500 5230 11552
rect 6086 11500 6092 11552
rect 6144 11540 6150 11552
rect 8941 11543 8999 11549
rect 8941 11540 8953 11543
rect 6144 11512 8953 11540
rect 6144 11500 6150 11512
rect 8941 11509 8953 11512
rect 8987 11509 8999 11543
rect 11054 11540 11060 11552
rect 11015 11512 11060 11540
rect 8941 11503 8999 11509
rect 11054 11500 11060 11512
rect 11112 11500 11118 11552
rect 11164 11549 11192 11580
rect 11517 11577 11529 11611
rect 11563 11608 11575 11611
rect 11790 11608 11796 11620
rect 11563 11580 11796 11608
rect 11563 11577 11575 11580
rect 11517 11571 11575 11577
rect 11790 11568 11796 11580
rect 11848 11568 11854 11620
rect 12526 11568 12532 11620
rect 12584 11608 12590 11620
rect 12636 11608 12664 11716
rect 12802 11704 12808 11716
rect 12860 11744 12866 11756
rect 12989 11747 13047 11753
rect 12989 11744 13001 11747
rect 12860 11716 13001 11744
rect 12860 11704 12866 11716
rect 12989 11713 13001 11716
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 13078 11704 13084 11756
rect 13136 11744 13142 11756
rect 14458 11744 14464 11756
rect 13136 11716 14464 11744
rect 13136 11704 13142 11716
rect 14458 11704 14464 11716
rect 14516 11704 14522 11756
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11744 15623 11747
rect 15838 11744 15844 11756
rect 15611 11716 15844 11744
rect 15611 11713 15623 11716
rect 15565 11707 15623 11713
rect 15838 11704 15844 11716
rect 15896 11704 15902 11756
rect 18693 11747 18751 11753
rect 15948 11716 16887 11744
rect 12897 11679 12955 11685
rect 12897 11645 12909 11679
rect 12943 11676 12955 11679
rect 13170 11676 13176 11688
rect 12943 11648 13176 11676
rect 12943 11645 12955 11648
rect 12897 11639 12955 11645
rect 13170 11636 13176 11648
rect 13228 11636 13234 11688
rect 14185 11679 14243 11685
rect 14185 11645 14197 11679
rect 14231 11676 14243 11679
rect 14274 11676 14280 11688
rect 14231 11648 14280 11676
rect 14231 11645 14243 11648
rect 14185 11639 14243 11645
rect 14274 11636 14280 11648
rect 14332 11636 14338 11688
rect 15948 11676 15976 11716
rect 14384 11648 15976 11676
rect 14384 11608 14412 11648
rect 16298 11636 16304 11688
rect 16356 11676 16362 11688
rect 16485 11679 16543 11685
rect 16485 11676 16497 11679
rect 16356 11648 16497 11676
rect 16356 11636 16362 11648
rect 16485 11645 16497 11648
rect 16531 11645 16543 11679
rect 16485 11639 16543 11645
rect 15102 11608 15108 11620
rect 12584 11580 12664 11608
rect 12820 11580 14412 11608
rect 14936 11580 15108 11608
rect 12584 11568 12590 11580
rect 12820 11552 12848 11580
rect 11149 11543 11207 11549
rect 11149 11509 11161 11543
rect 11195 11509 11207 11543
rect 12802 11540 12808 11552
rect 12763 11512 12808 11540
rect 11149 11503 11207 11509
rect 12802 11500 12808 11512
rect 12860 11500 12866 11552
rect 14936 11549 14964 11580
rect 15102 11568 15108 11580
rect 15160 11568 15166 11620
rect 15289 11611 15347 11617
rect 15289 11577 15301 11611
rect 15335 11608 15347 11611
rect 16666 11608 16672 11620
rect 15335 11580 16672 11608
rect 15335 11577 15347 11580
rect 15289 11571 15347 11577
rect 16666 11568 16672 11580
rect 16724 11568 16730 11620
rect 16761 11611 16819 11617
rect 16761 11577 16773 11611
rect 16807 11577 16819 11611
rect 16859 11608 16887 11716
rect 18693 11713 18705 11747
rect 18739 11744 18751 11747
rect 19058 11744 19064 11756
rect 18739 11716 19064 11744
rect 18739 11713 18751 11716
rect 18693 11707 18751 11713
rect 19058 11704 19064 11716
rect 19116 11704 19122 11756
rect 19242 11704 19248 11756
rect 19300 11704 19306 11756
rect 18509 11679 18567 11685
rect 18509 11645 18521 11679
rect 18555 11676 18567 11679
rect 19260 11676 19288 11704
rect 19996 11685 20024 11784
rect 20162 11744 20168 11756
rect 20123 11716 20168 11744
rect 20162 11704 20168 11716
rect 20220 11704 20226 11756
rect 18555 11648 19288 11676
rect 19981 11679 20039 11685
rect 18555 11645 18567 11648
rect 18509 11639 18567 11645
rect 19981 11645 19993 11679
rect 20027 11645 20039 11679
rect 19981 11639 20039 11645
rect 18690 11608 18696 11620
rect 16859 11580 18696 11608
rect 16761 11571 16819 11577
rect 14921 11543 14979 11549
rect 14921 11509 14933 11543
rect 14967 11509 14979 11543
rect 14921 11503 14979 11509
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 15436 11512 15481 11540
rect 15436 11500 15442 11512
rect 16022 11500 16028 11552
rect 16080 11540 16086 11552
rect 16776 11540 16804 11571
rect 18690 11568 18696 11580
rect 18748 11568 18754 11620
rect 18874 11568 18880 11620
rect 18932 11608 18938 11620
rect 20073 11611 20131 11617
rect 20073 11608 20085 11611
rect 18932 11580 20085 11608
rect 18932 11568 18938 11580
rect 20073 11577 20085 11580
rect 20119 11577 20131 11611
rect 20073 11571 20131 11577
rect 16080 11512 16804 11540
rect 16080 11500 16086 11512
rect 17218 11500 17224 11552
rect 17276 11540 17282 11552
rect 18049 11543 18107 11549
rect 18049 11540 18061 11543
rect 17276 11512 18061 11540
rect 17276 11500 17282 11512
rect 18049 11509 18061 11512
rect 18095 11509 18107 11543
rect 18049 11503 18107 11509
rect 18230 11500 18236 11552
rect 18288 11540 18294 11552
rect 18417 11543 18475 11549
rect 18417 11540 18429 11543
rect 18288 11512 18429 11540
rect 18288 11500 18294 11512
rect 18417 11509 18429 11512
rect 18463 11509 18475 11543
rect 18417 11503 18475 11509
rect 19334 11500 19340 11552
rect 19392 11540 19398 11552
rect 19613 11543 19671 11549
rect 19613 11540 19625 11543
rect 19392 11512 19625 11540
rect 19392 11500 19398 11512
rect 19613 11509 19625 11512
rect 19659 11509 19671 11543
rect 19613 11503 19671 11509
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 2409 11339 2467 11345
rect 2409 11305 2421 11339
rect 2455 11305 2467 11339
rect 2409 11299 2467 11305
rect 1486 11228 1492 11280
rect 1544 11268 1550 11280
rect 2038 11268 2044 11280
rect 1544 11240 2044 11268
rect 1544 11228 1550 11240
rect 2038 11228 2044 11240
rect 2096 11228 2102 11280
rect 2424 11268 2452 11299
rect 2590 11296 2596 11348
rect 2648 11336 2654 11348
rect 2869 11339 2927 11345
rect 2869 11336 2881 11339
rect 2648 11308 2881 11336
rect 2648 11296 2654 11308
rect 2869 11305 2881 11308
rect 2915 11336 2927 11339
rect 3970 11336 3976 11348
rect 2915 11308 3976 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 3970 11296 3976 11308
rect 4028 11296 4034 11348
rect 4614 11296 4620 11348
rect 4672 11336 4678 11348
rect 5902 11336 5908 11348
rect 4672 11308 5212 11336
rect 5863 11308 5908 11336
rect 4672 11296 4678 11308
rect 3602 11268 3608 11280
rect 2424 11240 3608 11268
rect 3602 11228 3608 11240
rect 3660 11228 3666 11280
rect 4792 11271 4850 11277
rect 4792 11237 4804 11271
rect 4838 11268 4850 11271
rect 4982 11268 4988 11280
rect 4838 11240 4988 11268
rect 4838 11237 4850 11240
rect 4792 11231 4850 11237
rect 4982 11228 4988 11240
rect 5040 11228 5046 11280
rect 2777 11203 2835 11209
rect 2777 11169 2789 11203
rect 2823 11200 2835 11203
rect 3234 11200 3240 11212
rect 2823 11172 3240 11200
rect 2823 11169 2835 11172
rect 2777 11163 2835 11169
rect 3234 11160 3240 11172
rect 3292 11160 3298 11212
rect 5184 11200 5212 11308
rect 5902 11296 5908 11308
rect 5960 11296 5966 11348
rect 7466 11296 7472 11348
rect 7524 11336 7530 11348
rect 7524 11308 11192 11336
rect 7524 11296 7530 11308
rect 6454 11228 6460 11280
rect 6512 11268 6518 11280
rect 6914 11268 6920 11280
rect 6512 11240 6920 11268
rect 6512 11228 6518 11240
rect 6914 11228 6920 11240
rect 6972 11228 6978 11280
rect 7644 11271 7702 11277
rect 7644 11237 7656 11271
rect 7690 11268 7702 11271
rect 11054 11268 11060 11280
rect 7690 11240 11060 11268
rect 7690 11237 7702 11240
rect 7644 11231 7702 11237
rect 11054 11228 11060 11240
rect 11112 11228 11118 11280
rect 7377 11203 7435 11209
rect 5184 11172 6960 11200
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11132 1455 11135
rect 2038 11132 2044 11144
rect 1443 11104 2044 11132
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 2038 11092 2044 11104
rect 2096 11092 2102 11144
rect 2314 11092 2320 11144
rect 2372 11132 2378 11144
rect 3050 11132 3056 11144
rect 2372 11104 3056 11132
rect 2372 11092 2378 11104
rect 3050 11092 3056 11104
rect 3108 11092 3114 11144
rect 4154 11092 4160 11144
rect 4212 11132 4218 11144
rect 4525 11135 4583 11141
rect 4525 11132 4537 11135
rect 4212 11104 4537 11132
rect 4212 11092 4218 11104
rect 4525 11101 4537 11104
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 4540 10996 4568 11095
rect 6270 10996 6276 11008
rect 4540 10968 6276 10996
rect 6270 10956 6276 10968
rect 6328 10996 6334 11008
rect 6822 10996 6828 11008
rect 6328 10968 6828 10996
rect 6328 10956 6334 10968
rect 6822 10956 6828 10968
rect 6880 10956 6886 11008
rect 6932 10996 6960 11172
rect 7377 11169 7389 11203
rect 7423 11200 7435 11203
rect 9674 11200 9680 11212
rect 7423 11172 9680 11200
rect 7423 11169 7435 11172
rect 7377 11163 7435 11169
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 10226 11160 10232 11212
rect 10284 11200 10290 11212
rect 10413 11203 10471 11209
rect 10413 11200 10425 11203
rect 10284 11172 10425 11200
rect 10284 11160 10290 11172
rect 10413 11169 10425 11172
rect 10459 11169 10471 11203
rect 10413 11163 10471 11169
rect 10686 11132 10692 11144
rect 8404 11104 10692 11132
rect 8404 11064 8432 11104
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 11072 11132 11100 11228
rect 11164 11200 11192 11308
rect 11698 11296 11704 11348
rect 11756 11336 11762 11348
rect 12713 11339 12771 11345
rect 12713 11336 12725 11339
rect 11756 11308 12725 11336
rect 11756 11296 11762 11308
rect 12713 11305 12725 11308
rect 12759 11305 12771 11339
rect 13630 11336 13636 11348
rect 13591 11308 13636 11336
rect 12713 11299 12771 11305
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 14090 11336 14096 11348
rect 14051 11308 14096 11336
rect 14090 11296 14096 11308
rect 14148 11296 14154 11348
rect 14458 11296 14464 11348
rect 14516 11336 14522 11348
rect 16022 11336 16028 11348
rect 14516 11308 16028 11336
rect 14516 11296 14522 11308
rect 16022 11296 16028 11308
rect 16080 11296 16086 11348
rect 18138 11336 18144 11348
rect 18099 11308 18144 11336
rect 18138 11296 18144 11308
rect 18196 11296 18202 11348
rect 18966 11336 18972 11348
rect 18927 11308 18972 11336
rect 18966 11296 18972 11308
rect 19024 11296 19030 11348
rect 19334 11336 19340 11348
rect 19295 11308 19340 11336
rect 19334 11296 19340 11308
rect 19392 11296 19398 11348
rect 11422 11228 11428 11280
rect 11480 11268 11486 11280
rect 12621 11271 12679 11277
rect 12621 11268 12633 11271
rect 11480 11240 12633 11268
rect 11480 11228 11486 11240
rect 12621 11237 12633 11240
rect 12667 11237 12679 11271
rect 13998 11268 14004 11280
rect 13959 11240 14004 11268
rect 12621 11231 12679 11237
rect 13998 11228 14004 11240
rect 14056 11228 14062 11280
rect 15194 11228 15200 11280
rect 15252 11268 15258 11280
rect 15565 11271 15623 11277
rect 15565 11268 15577 11271
rect 15252 11240 15577 11268
rect 15252 11228 15258 11240
rect 15565 11237 15577 11240
rect 15611 11237 15623 11271
rect 15565 11231 15623 11237
rect 15289 11203 15347 11209
rect 15289 11200 15301 11203
rect 11164 11172 15301 11200
rect 15289 11169 15301 11172
rect 15335 11169 15347 11203
rect 16758 11200 16764 11212
rect 16719 11172 16764 11200
rect 15289 11163 15347 11169
rect 16758 11160 16764 11172
rect 16816 11160 16822 11212
rect 17028 11203 17086 11209
rect 17028 11169 17040 11203
rect 17074 11200 17086 11203
rect 17862 11200 17868 11212
rect 17074 11172 17868 11200
rect 17074 11169 17086 11172
rect 17028 11163 17086 11169
rect 17862 11160 17868 11172
rect 17920 11200 17926 11212
rect 17920 11172 19564 11200
rect 17920 11160 17926 11172
rect 12805 11135 12863 11141
rect 12805 11132 12817 11135
rect 11072 11104 12817 11132
rect 12805 11101 12817 11104
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11132 14335 11135
rect 14734 11132 14740 11144
rect 14323 11104 14740 11132
rect 14323 11101 14335 11104
rect 14277 11095 14335 11101
rect 14734 11092 14740 11104
rect 14792 11132 14798 11144
rect 15838 11132 15844 11144
rect 14792 11104 15844 11132
rect 14792 11092 14798 11104
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 19426 11132 19432 11144
rect 19387 11104 19432 11132
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 19536 11141 19564 11172
rect 19521 11135 19579 11141
rect 19521 11101 19533 11135
rect 19567 11101 19579 11135
rect 19521 11095 19579 11101
rect 8754 11064 8760 11076
rect 8312 11036 8432 11064
rect 8715 11036 8760 11064
rect 8312 10996 8340 11036
rect 8754 11024 8760 11036
rect 8812 11024 8818 11076
rect 10778 11024 10784 11076
rect 10836 11064 10842 11076
rect 12253 11067 12311 11073
rect 12253 11064 12265 11067
rect 10836 11036 12265 11064
rect 10836 11024 10842 11036
rect 12253 11033 12265 11036
rect 12299 11033 12311 11067
rect 13906 11064 13912 11076
rect 12253 11027 12311 11033
rect 13556 11036 13912 11064
rect 6932 10968 8340 10996
rect 8386 10956 8392 11008
rect 8444 10996 8450 11008
rect 11146 10996 11152 11008
rect 8444 10968 11152 10996
rect 8444 10956 8450 10968
rect 11146 10956 11152 10968
rect 11204 10956 11210 11008
rect 11698 10996 11704 11008
rect 11659 10968 11704 10996
rect 11698 10956 11704 10968
rect 11756 10956 11762 11008
rect 11790 10956 11796 11008
rect 11848 10996 11854 11008
rect 13556 10996 13584 11036
rect 13906 11024 13912 11036
rect 13964 11024 13970 11076
rect 14826 11024 14832 11076
rect 14884 11064 14890 11076
rect 15930 11064 15936 11076
rect 14884 11036 15936 11064
rect 14884 11024 14890 11036
rect 15930 11024 15936 11036
rect 15988 11024 15994 11076
rect 11848 10968 13584 10996
rect 11848 10956 11854 10968
rect 13630 10956 13636 11008
rect 13688 10996 13694 11008
rect 18782 10996 18788 11008
rect 13688 10968 18788 10996
rect 13688 10956 13694 10968
rect 18782 10956 18788 10968
rect 18840 10956 18846 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 3050 10752 3056 10804
rect 3108 10792 3114 10804
rect 5166 10792 5172 10804
rect 3108 10764 5172 10792
rect 3108 10752 3114 10764
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 6730 10752 6736 10804
rect 6788 10792 6794 10804
rect 8386 10792 8392 10804
rect 6788 10764 8392 10792
rect 6788 10752 6794 10764
rect 8386 10752 8392 10764
rect 8444 10752 8450 10804
rect 9033 10795 9091 10801
rect 9033 10761 9045 10795
rect 9079 10792 9091 10795
rect 9766 10792 9772 10804
rect 9079 10764 9772 10792
rect 9079 10761 9091 10764
rect 9033 10755 9091 10761
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 10318 10752 10324 10804
rect 10376 10792 10382 10804
rect 10965 10795 11023 10801
rect 10965 10792 10977 10795
rect 10376 10764 10977 10792
rect 10376 10752 10382 10764
rect 10965 10761 10977 10764
rect 11011 10761 11023 10795
rect 10965 10755 11023 10761
rect 11054 10752 11060 10804
rect 11112 10792 11118 10804
rect 14090 10792 14096 10804
rect 11112 10764 14096 10792
rect 11112 10752 11118 10764
rect 14090 10752 14096 10764
rect 14148 10752 14154 10804
rect 15838 10792 15844 10804
rect 15799 10764 15844 10792
rect 15838 10752 15844 10764
rect 15896 10752 15902 10804
rect 16666 10752 16672 10804
rect 16724 10792 16730 10804
rect 18049 10795 18107 10801
rect 18049 10792 18061 10795
rect 16724 10764 18061 10792
rect 16724 10752 16730 10764
rect 18049 10761 18061 10764
rect 18095 10761 18107 10795
rect 18049 10755 18107 10761
rect 19426 10752 19432 10804
rect 19484 10792 19490 10804
rect 19613 10795 19671 10801
rect 19613 10792 19625 10795
rect 19484 10764 19625 10792
rect 19484 10752 19490 10764
rect 19613 10761 19625 10764
rect 19659 10761 19671 10795
rect 19613 10755 19671 10761
rect 3421 10727 3479 10733
rect 3421 10693 3433 10727
rect 3467 10693 3479 10727
rect 3421 10687 3479 10693
rect 3436 10656 3464 10687
rect 3970 10684 3976 10736
rect 4028 10724 4034 10736
rect 4028 10696 4936 10724
rect 4028 10684 4034 10696
rect 4801 10659 4859 10665
rect 4801 10656 4813 10659
rect 3436 10628 4813 10656
rect 2314 10597 2320 10600
rect 2041 10591 2099 10597
rect 2041 10557 2053 10591
rect 2087 10557 2099 10591
rect 2308 10588 2320 10597
rect 2275 10560 2320 10588
rect 2041 10551 2099 10557
rect 2308 10551 2320 10560
rect 2056 10520 2084 10551
rect 2314 10548 2320 10551
rect 2372 10548 2378 10600
rect 2498 10520 2504 10532
rect 2056 10492 2504 10520
rect 2498 10480 2504 10492
rect 2556 10480 2562 10532
rect 2682 10412 2688 10464
rect 2740 10452 2746 10464
rect 3436 10452 3464 10628
rect 4801 10625 4813 10628
rect 4847 10625 4859 10659
rect 4908 10656 4936 10696
rect 11146 10684 11152 10736
rect 11204 10724 11210 10736
rect 11882 10724 11888 10736
rect 11204 10696 11888 10724
rect 11204 10684 11210 10696
rect 11882 10684 11888 10696
rect 11940 10684 11946 10736
rect 12069 10727 12127 10733
rect 12069 10693 12081 10727
rect 12115 10724 12127 10727
rect 14274 10724 14280 10736
rect 12115 10696 14280 10724
rect 12115 10693 12127 10696
rect 12069 10687 12127 10693
rect 14274 10684 14280 10696
rect 14332 10684 14338 10736
rect 17494 10684 17500 10736
rect 17552 10724 17558 10736
rect 17552 10696 20300 10724
rect 17552 10684 17558 10696
rect 4908 10628 6960 10656
rect 4801 10619 4859 10625
rect 3602 10548 3608 10600
rect 3660 10588 3666 10600
rect 4617 10591 4675 10597
rect 4617 10588 4629 10591
rect 3660 10560 4629 10588
rect 3660 10548 3666 10560
rect 4617 10557 4629 10560
rect 4663 10557 4675 10591
rect 6822 10588 6828 10600
rect 6783 10560 6828 10588
rect 4617 10551 4675 10557
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 6932 10588 6960 10628
rect 9232 10628 9720 10656
rect 9232 10597 9260 10628
rect 9217 10591 9275 10597
rect 6932 10560 8340 10588
rect 4154 10480 4160 10532
rect 4212 10520 4218 10532
rect 4709 10523 4767 10529
rect 4709 10520 4721 10523
rect 4212 10492 4721 10520
rect 4212 10480 4218 10492
rect 4709 10489 4721 10492
rect 4755 10489 4767 10523
rect 4709 10483 4767 10489
rect 5534 10480 5540 10532
rect 5592 10520 5598 10532
rect 6638 10520 6644 10532
rect 5592 10492 6644 10520
rect 5592 10480 5598 10492
rect 6638 10480 6644 10492
rect 6696 10480 6702 10532
rect 7098 10529 7104 10532
rect 7092 10520 7104 10529
rect 7059 10492 7104 10520
rect 7092 10483 7104 10492
rect 7098 10480 7104 10483
rect 7156 10480 7162 10532
rect 2740 10424 3464 10452
rect 2740 10412 2746 10424
rect 3602 10412 3608 10464
rect 3660 10452 3666 10464
rect 4249 10455 4307 10461
rect 4249 10452 4261 10455
rect 3660 10424 4261 10452
rect 3660 10412 3666 10424
rect 4249 10421 4261 10424
rect 4295 10421 4307 10455
rect 4249 10415 4307 10421
rect 6270 10412 6276 10464
rect 6328 10452 6334 10464
rect 8205 10455 8263 10461
rect 8205 10452 8217 10455
rect 6328 10424 8217 10452
rect 6328 10412 6334 10424
rect 8205 10421 8217 10424
rect 8251 10421 8263 10455
rect 8312 10452 8340 10560
rect 9217 10557 9229 10591
rect 9263 10557 9275 10591
rect 9217 10551 9275 10557
rect 9585 10591 9643 10597
rect 9585 10557 9597 10591
rect 9631 10557 9643 10591
rect 9692 10588 9720 10628
rect 11422 10616 11428 10668
rect 11480 10656 11486 10668
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 11480 10628 13001 10656
rect 11480 10616 11486 10628
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 15562 10616 15568 10668
rect 15620 10656 15626 10668
rect 15838 10656 15844 10668
rect 15620 10628 15844 10656
rect 15620 10616 15626 10628
rect 15838 10616 15844 10628
rect 15896 10616 15902 10668
rect 16022 10616 16028 10668
rect 16080 10656 16086 10668
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 16080 10628 18613 10656
rect 16080 10616 16086 10628
rect 18601 10625 18613 10628
rect 18647 10625 18659 10659
rect 20162 10656 20168 10668
rect 20123 10628 20168 10656
rect 18601 10619 18659 10625
rect 20162 10616 20168 10628
rect 20220 10616 20226 10668
rect 11698 10588 11704 10600
rect 9692 10560 11704 10588
rect 9585 10551 9643 10557
rect 9600 10520 9628 10551
rect 11698 10548 11704 10560
rect 11756 10588 11762 10600
rect 12253 10591 12311 10597
rect 12253 10588 12265 10591
rect 11756 10560 12265 10588
rect 11756 10548 11762 10560
rect 12253 10557 12265 10560
rect 12299 10557 12311 10591
rect 14458 10588 14464 10600
rect 14419 10560 14464 10588
rect 12253 10551 12311 10557
rect 14458 10548 14464 10560
rect 14516 10548 14522 10600
rect 16669 10591 16727 10597
rect 16669 10588 16681 10591
rect 14568 10560 16681 10588
rect 9674 10520 9680 10532
rect 9600 10492 9680 10520
rect 9674 10480 9680 10492
rect 9732 10480 9738 10532
rect 9852 10523 9910 10529
rect 9852 10489 9864 10523
rect 9898 10520 9910 10523
rect 11146 10520 11152 10532
rect 9898 10492 11152 10520
rect 9898 10489 9910 10492
rect 9852 10483 9910 10489
rect 11146 10480 11152 10492
rect 11204 10480 11210 10532
rect 11330 10480 11336 10532
rect 11388 10520 11394 10532
rect 12897 10523 12955 10529
rect 12897 10520 12909 10523
rect 11388 10492 12909 10520
rect 11388 10480 11394 10492
rect 12897 10489 12909 10492
rect 12943 10489 12955 10523
rect 12897 10483 12955 10489
rect 13078 10480 13084 10532
rect 13136 10520 13142 10532
rect 14568 10520 14596 10560
rect 16669 10557 16681 10560
rect 16715 10557 16727 10591
rect 16669 10551 16727 10557
rect 16758 10548 16764 10600
rect 16816 10588 16822 10600
rect 19429 10591 19487 10597
rect 19429 10588 19441 10591
rect 16816 10560 19441 10588
rect 16816 10548 16822 10560
rect 19429 10557 19441 10560
rect 19475 10588 19487 10591
rect 19981 10591 20039 10597
rect 19981 10588 19993 10591
rect 19475 10560 19993 10588
rect 19475 10557 19487 10560
rect 19429 10551 19487 10557
rect 19981 10557 19993 10560
rect 20027 10557 20039 10591
rect 19981 10551 20039 10557
rect 20073 10591 20131 10597
rect 20073 10557 20085 10591
rect 20119 10588 20131 10591
rect 20272 10588 20300 10696
rect 20441 10591 20499 10597
rect 20441 10588 20453 10591
rect 20119 10560 20453 10588
rect 20119 10557 20131 10560
rect 20073 10551 20131 10557
rect 20441 10557 20453 10560
rect 20487 10557 20499 10591
rect 20441 10551 20499 10557
rect 13136 10492 14596 10520
rect 14728 10523 14786 10529
rect 13136 10480 13142 10492
rect 14728 10489 14740 10523
rect 14774 10520 14786 10523
rect 15654 10520 15660 10532
rect 14774 10492 15660 10520
rect 14774 10489 14786 10492
rect 14728 10483 14786 10489
rect 15654 10480 15660 10492
rect 15712 10520 15718 10532
rect 16022 10520 16028 10532
rect 15712 10492 16028 10520
rect 15712 10480 15718 10492
rect 16022 10480 16028 10492
rect 16080 10480 16086 10532
rect 16850 10480 16856 10532
rect 16908 10520 16914 10532
rect 16945 10523 17003 10529
rect 16945 10520 16957 10523
rect 16908 10492 16957 10520
rect 16908 10480 16914 10492
rect 16945 10489 16957 10492
rect 16991 10489 17003 10523
rect 16945 10483 17003 10489
rect 17954 10480 17960 10532
rect 18012 10520 18018 10532
rect 18417 10523 18475 10529
rect 18417 10520 18429 10523
rect 18012 10492 18429 10520
rect 18012 10480 18018 10492
rect 18417 10489 18429 10492
rect 18463 10489 18475 10523
rect 18417 10483 18475 10489
rect 11054 10452 11060 10464
rect 8312 10424 11060 10452
rect 8205 10415 8263 10421
rect 11054 10412 11060 10424
rect 11112 10412 11118 10464
rect 11514 10412 11520 10464
rect 11572 10452 11578 10464
rect 12437 10455 12495 10461
rect 12437 10452 12449 10455
rect 11572 10424 12449 10452
rect 11572 10412 11578 10424
rect 12437 10421 12449 10424
rect 12483 10421 12495 10455
rect 12802 10452 12808 10464
rect 12763 10424 12808 10452
rect 12437 10415 12495 10421
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 14090 10412 14096 10464
rect 14148 10452 14154 10464
rect 15930 10452 15936 10464
rect 14148 10424 15936 10452
rect 14148 10412 14154 10424
rect 15930 10412 15936 10424
rect 15988 10412 15994 10464
rect 17678 10412 17684 10464
rect 17736 10452 17742 10464
rect 18509 10455 18567 10461
rect 18509 10452 18521 10455
rect 17736 10424 18521 10452
rect 17736 10412 17742 10424
rect 18509 10421 18521 10424
rect 18555 10452 18567 10455
rect 18877 10455 18935 10461
rect 18877 10452 18889 10455
rect 18555 10424 18889 10452
rect 18555 10421 18567 10424
rect 18509 10415 18567 10421
rect 18877 10421 18889 10424
rect 18923 10452 18935 10455
rect 19978 10452 19984 10464
rect 18923 10424 19984 10452
rect 18923 10421 18935 10424
rect 18877 10415 18935 10421
rect 19978 10412 19984 10424
rect 20036 10412 20042 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 1854 10208 1860 10260
rect 1912 10248 1918 10260
rect 7466 10248 7472 10260
rect 1912 10220 7472 10248
rect 1912 10208 1918 10220
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 7929 10251 7987 10257
rect 7929 10217 7941 10251
rect 7975 10248 7987 10251
rect 8202 10248 8208 10260
rect 7975 10220 8208 10248
rect 7975 10217 7987 10220
rect 7929 10211 7987 10217
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 11330 10248 11336 10260
rect 8444 10220 11336 10248
rect 8444 10208 8450 10220
rect 11330 10208 11336 10220
rect 11388 10208 11394 10260
rect 11882 10208 11888 10260
rect 11940 10248 11946 10260
rect 15289 10251 15347 10257
rect 11940 10220 13492 10248
rect 11940 10208 11946 10220
rect 1756 10183 1814 10189
rect 1756 10149 1768 10183
rect 1802 10180 1814 10183
rect 2682 10180 2688 10192
rect 1802 10152 2688 10180
rect 1802 10149 1814 10152
rect 1756 10143 1814 10149
rect 2682 10140 2688 10152
rect 2740 10140 2746 10192
rect 4246 10140 4252 10192
rect 4304 10180 4310 10192
rect 4341 10183 4399 10189
rect 4341 10180 4353 10183
rect 4304 10152 4353 10180
rect 4304 10140 4310 10152
rect 4341 10149 4353 10152
rect 4387 10149 4399 10183
rect 4341 10143 4399 10149
rect 8021 10183 8079 10189
rect 8021 10149 8033 10183
rect 8067 10180 8079 10183
rect 8294 10180 8300 10192
rect 8067 10152 8300 10180
rect 8067 10149 8079 10152
rect 8021 10143 8079 10149
rect 8294 10140 8300 10152
rect 8352 10140 8358 10192
rect 10496 10183 10554 10189
rect 10496 10149 10508 10183
rect 10542 10180 10554 10183
rect 13170 10180 13176 10192
rect 10542 10152 13176 10180
rect 10542 10149 10554 10152
rect 10496 10143 10554 10149
rect 13170 10140 13176 10152
rect 13228 10140 13234 10192
rect 1489 10115 1547 10121
rect 1489 10081 1501 10115
rect 1535 10112 1547 10115
rect 4062 10112 4068 10124
rect 1535 10084 2544 10112
rect 4023 10084 4068 10112
rect 1535 10081 1547 10084
rect 1489 10075 1547 10081
rect 2516 10056 2544 10084
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 5620 10115 5678 10121
rect 5620 10081 5632 10115
rect 5666 10112 5678 10115
rect 5902 10112 5908 10124
rect 5666 10084 5908 10112
rect 5666 10081 5678 10084
rect 5620 10075 5678 10081
rect 5902 10072 5908 10084
rect 5960 10112 5966 10124
rect 6086 10112 6092 10124
rect 5960 10084 6092 10112
rect 5960 10072 5966 10084
rect 6086 10072 6092 10084
rect 6144 10072 6150 10124
rect 7558 10072 7564 10124
rect 7616 10112 7622 10124
rect 7834 10112 7840 10124
rect 7616 10084 7840 10112
rect 7616 10072 7622 10084
rect 7834 10072 7840 10084
rect 7892 10072 7898 10124
rect 7926 10072 7932 10124
rect 7984 10112 7990 10124
rect 12342 10112 12348 10124
rect 7984 10084 12348 10112
rect 7984 10072 7990 10084
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 12526 10072 12532 10124
rect 12584 10112 12590 10124
rect 12693 10115 12751 10121
rect 12693 10112 12705 10115
rect 12584 10084 12705 10112
rect 12584 10072 12590 10084
rect 12693 10081 12705 10084
rect 12739 10081 12751 10115
rect 12693 10075 12751 10081
rect 2498 10004 2504 10056
rect 2556 10044 2562 10056
rect 5353 10047 5411 10053
rect 5353 10044 5365 10047
rect 2556 10016 5365 10044
rect 2556 10004 2562 10016
rect 5353 10013 5365 10016
rect 5399 10013 5411 10047
rect 5353 10007 5411 10013
rect 6822 10004 6828 10056
rect 6880 10044 6886 10056
rect 8018 10044 8024 10056
rect 6880 10016 8024 10044
rect 6880 10004 6886 10016
rect 8018 10004 8024 10016
rect 8076 10004 8082 10056
rect 8113 10047 8171 10053
rect 8113 10013 8125 10047
rect 8159 10013 8171 10047
rect 8113 10007 8171 10013
rect 6733 9979 6791 9985
rect 6733 9945 6745 9979
rect 6779 9976 6791 9979
rect 7098 9976 7104 9988
rect 6779 9948 7104 9976
rect 6779 9945 6791 9948
rect 6733 9939 6791 9945
rect 7098 9936 7104 9948
rect 7156 9976 7162 9988
rect 8128 9976 8156 10007
rect 9674 10004 9680 10056
rect 9732 10044 9738 10056
rect 10229 10047 10287 10053
rect 10229 10044 10241 10047
rect 9732 10016 10241 10044
rect 9732 10004 9738 10016
rect 10229 10013 10241 10016
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 11974 10004 11980 10056
rect 12032 10044 12038 10056
rect 12437 10047 12495 10053
rect 12437 10044 12449 10047
rect 12032 10016 12449 10044
rect 12032 10004 12038 10016
rect 12437 10013 12449 10016
rect 12483 10013 12495 10047
rect 12437 10007 12495 10013
rect 7156 9948 8432 9976
rect 7156 9936 7162 9948
rect 2866 9908 2872 9920
rect 2827 9880 2872 9908
rect 2866 9868 2872 9880
rect 2924 9868 2930 9920
rect 3602 9868 3608 9920
rect 3660 9908 3666 9920
rect 4338 9908 4344 9920
rect 3660 9880 4344 9908
rect 3660 9868 3666 9880
rect 4338 9868 4344 9880
rect 4396 9868 4402 9920
rect 6822 9868 6828 9920
rect 6880 9908 6886 9920
rect 7561 9911 7619 9917
rect 7561 9908 7573 9911
rect 6880 9880 7573 9908
rect 6880 9868 6886 9880
rect 7561 9877 7573 9880
rect 7607 9877 7619 9911
rect 7561 9871 7619 9877
rect 7650 9868 7656 9920
rect 7708 9908 7714 9920
rect 7834 9908 7840 9920
rect 7708 9880 7840 9908
rect 7708 9868 7714 9880
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 8404 9908 8432 9948
rect 8754 9936 8760 9988
rect 8812 9976 8818 9988
rect 9398 9976 9404 9988
rect 8812 9948 9404 9976
rect 8812 9936 8818 9948
rect 9398 9936 9404 9948
rect 9456 9936 9462 9988
rect 11422 9936 11428 9988
rect 11480 9936 11486 9988
rect 11514 9936 11520 9988
rect 11572 9976 11578 9988
rect 11609 9979 11667 9985
rect 11609 9976 11621 9979
rect 11572 9948 11621 9976
rect 11572 9936 11578 9948
rect 11609 9945 11621 9948
rect 11655 9945 11667 9979
rect 13464 9976 13492 10220
rect 15289 10217 15301 10251
rect 15335 10248 15347 10251
rect 15378 10248 15384 10260
rect 15335 10220 15384 10248
rect 15335 10217 15347 10220
rect 15289 10211 15347 10217
rect 15378 10208 15384 10220
rect 15436 10208 15442 10260
rect 15562 10208 15568 10260
rect 15620 10248 15626 10260
rect 15749 10251 15807 10257
rect 15749 10248 15761 10251
rect 15620 10220 15761 10248
rect 15620 10208 15626 10220
rect 15749 10217 15761 10220
rect 15795 10217 15807 10251
rect 18417 10251 18475 10257
rect 18417 10248 18429 10251
rect 15749 10211 15807 10217
rect 15856 10220 18429 10248
rect 15654 10140 15660 10192
rect 15712 10180 15718 10192
rect 15712 10152 15757 10180
rect 15712 10140 15718 10152
rect 15856 10112 15884 10220
rect 18417 10217 18429 10220
rect 18463 10217 18475 10251
rect 18782 10248 18788 10260
rect 18743 10220 18788 10248
rect 18417 10211 18475 10217
rect 18782 10208 18788 10220
rect 18840 10208 18846 10260
rect 15930 10140 15936 10192
rect 15988 10180 15994 10192
rect 18877 10183 18935 10189
rect 18877 10180 18889 10183
rect 15988 10152 18889 10180
rect 15988 10140 15994 10152
rect 18877 10149 18889 10152
rect 18923 10149 18935 10183
rect 18877 10143 18935 10149
rect 15764 10084 15884 10112
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 15764 10044 15792 10084
rect 16114 10072 16120 10124
rect 16172 10112 16178 10124
rect 17221 10115 17279 10121
rect 17221 10112 17233 10115
rect 16172 10084 17233 10112
rect 16172 10072 16178 10084
rect 17221 10081 17233 10084
rect 17267 10081 17279 10115
rect 17221 10075 17279 10081
rect 13872 10016 15792 10044
rect 15933 10047 15991 10053
rect 13872 10004 13878 10016
rect 15933 10013 15945 10047
rect 15979 10044 15991 10047
rect 16022 10044 16028 10056
rect 15979 10016 16028 10044
rect 15979 10013 15991 10016
rect 15933 10007 15991 10013
rect 16022 10004 16028 10016
rect 16080 10004 16086 10056
rect 17313 10047 17371 10053
rect 17313 10013 17325 10047
rect 17359 10013 17371 10047
rect 17313 10007 17371 10013
rect 17328 9976 17356 10007
rect 17402 10004 17408 10056
rect 17460 10044 17466 10056
rect 17460 10016 17505 10044
rect 17460 10004 17466 10016
rect 18598 10004 18604 10056
rect 18656 10044 18662 10056
rect 18782 10044 18788 10056
rect 18656 10016 18788 10044
rect 18656 10004 18662 10016
rect 18782 10004 18788 10016
rect 18840 10044 18846 10056
rect 18969 10047 19027 10053
rect 18969 10044 18981 10047
rect 18840 10016 18981 10044
rect 18840 10004 18846 10016
rect 18969 10013 18981 10016
rect 19015 10013 19027 10047
rect 18969 10007 19027 10013
rect 13464 9948 17356 9976
rect 11609 9939 11667 9945
rect 11440 9908 11468 9936
rect 8404 9880 11468 9908
rect 13170 9868 13176 9920
rect 13228 9908 13234 9920
rect 13817 9911 13875 9917
rect 13817 9908 13829 9911
rect 13228 9880 13829 9908
rect 13228 9868 13234 9880
rect 13817 9877 13829 9880
rect 13863 9877 13875 9911
rect 13817 9871 13875 9877
rect 13906 9868 13912 9920
rect 13964 9908 13970 9920
rect 14182 9908 14188 9920
rect 13964 9880 14188 9908
rect 13964 9868 13970 9880
rect 14182 9868 14188 9880
rect 14240 9868 14246 9920
rect 15286 9868 15292 9920
rect 15344 9908 15350 9920
rect 16853 9911 16911 9917
rect 16853 9908 16865 9911
rect 15344 9880 16865 9908
rect 15344 9868 15350 9880
rect 16853 9877 16865 9880
rect 16899 9877 16911 9911
rect 16853 9871 16911 9877
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 1946 9704 1952 9716
rect 1907 9676 1952 9704
rect 1946 9664 1952 9676
rect 2004 9664 2010 9716
rect 5902 9664 5908 9716
rect 5960 9704 5966 9716
rect 8386 9704 8392 9716
rect 5960 9676 8392 9704
rect 5960 9664 5966 9676
rect 8386 9664 8392 9676
rect 8444 9664 8450 9716
rect 8478 9664 8484 9716
rect 8536 9704 8542 9716
rect 9306 9704 9312 9716
rect 8536 9676 9312 9704
rect 8536 9664 8542 9676
rect 9306 9664 9312 9676
rect 9364 9664 9370 9716
rect 9950 9664 9956 9716
rect 10008 9664 10014 9716
rect 10226 9664 10232 9716
rect 10284 9704 10290 9716
rect 12342 9704 12348 9716
rect 10284 9676 12348 9704
rect 10284 9664 10290 9676
rect 12342 9664 12348 9676
rect 12400 9664 12406 9716
rect 13078 9704 13084 9716
rect 12452 9676 13084 9704
rect 2590 9636 2596 9648
rect 1412 9608 2596 9636
rect 1412 9509 1440 9608
rect 2590 9596 2596 9608
rect 2648 9596 2654 9648
rect 3234 9596 3240 9648
rect 3292 9636 3298 9648
rect 7006 9636 7012 9648
rect 3292 9608 6776 9636
rect 6967 9608 7012 9636
rect 3292 9596 3298 9608
rect 2332 9540 2544 9568
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9469 1455 9503
rect 1397 9463 1455 9469
rect 1765 9503 1823 9509
rect 1765 9469 1777 9503
rect 1811 9469 1823 9503
rect 1765 9463 1823 9469
rect 1210 9392 1216 9444
rect 1268 9432 1274 9444
rect 1486 9432 1492 9444
rect 1268 9404 1492 9432
rect 1268 9392 1274 9404
rect 1486 9392 1492 9404
rect 1544 9392 1550 9444
rect 1780 9432 1808 9463
rect 2038 9460 2044 9512
rect 2096 9500 2102 9512
rect 2332 9500 2360 9540
rect 2516 9509 2544 9540
rect 2682 9528 2688 9580
rect 2740 9568 2746 9580
rect 2777 9571 2835 9577
rect 2777 9568 2789 9571
rect 2740 9540 2789 9568
rect 2740 9528 2746 9540
rect 2777 9537 2789 9540
rect 2823 9568 2835 9571
rect 4249 9571 4307 9577
rect 4249 9568 4261 9571
rect 2823 9540 4261 9568
rect 2823 9537 2835 9540
rect 2777 9531 2835 9537
rect 4249 9537 4261 9540
rect 4295 9537 4307 9571
rect 5445 9571 5503 9577
rect 5445 9568 5457 9571
rect 4249 9531 4307 9537
rect 4356 9540 5457 9568
rect 2096 9472 2360 9500
rect 2501 9503 2559 9509
rect 2096 9460 2102 9472
rect 2501 9469 2513 9503
rect 2547 9469 2559 9503
rect 2501 9463 2559 9469
rect 3878 9460 3884 9512
rect 3936 9500 3942 9512
rect 4356 9500 4384 9540
rect 5445 9537 5457 9540
rect 5491 9537 5503 9571
rect 5445 9531 5503 9537
rect 3936 9472 4384 9500
rect 5292 9503 5350 9509
rect 3936 9460 3942 9472
rect 5292 9469 5304 9503
rect 5338 9500 5350 9503
rect 6748 9500 6776 9608
rect 7006 9596 7012 9608
rect 7064 9596 7070 9648
rect 7098 9596 7104 9648
rect 7156 9636 7162 9648
rect 9968 9636 9996 9664
rect 7156 9608 9996 9636
rect 7156 9596 7162 9608
rect 8573 9571 8631 9577
rect 7668 9540 8524 9568
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 5338 9472 6123 9500
rect 6748 9472 6837 9500
rect 5338 9469 5350 9472
rect 5292 9463 5350 9469
rect 2314 9432 2320 9444
rect 1780 9404 2320 9432
rect 2314 9392 2320 9404
rect 2372 9392 2378 9444
rect 4157 9435 4215 9441
rect 4157 9401 4169 9435
rect 4203 9432 4215 9435
rect 5534 9432 5540 9444
rect 4203 9404 5540 9432
rect 4203 9401 4215 9404
rect 4157 9395 4215 9401
rect 5534 9392 5540 9404
rect 5592 9392 5598 9444
rect 6095 9432 6123 9472
rect 6825 9469 6837 9472
rect 6871 9469 6883 9503
rect 6825 9463 6883 9469
rect 7006 9460 7012 9512
rect 7064 9500 7070 9512
rect 7558 9500 7564 9512
rect 7064 9472 7564 9500
rect 7064 9460 7070 9472
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 7668 9432 7696 9540
rect 7742 9460 7748 9512
rect 7800 9460 7806 9512
rect 8018 9460 8024 9512
rect 8076 9500 8082 9512
rect 8297 9503 8355 9509
rect 8297 9500 8309 9503
rect 8076 9472 8309 9500
rect 8076 9460 8082 9472
rect 8297 9469 8309 9472
rect 8343 9469 8355 9503
rect 8297 9463 8355 9469
rect 6095 9404 7696 9432
rect 7760 9432 7788 9460
rect 8386 9432 8392 9444
rect 7760 9404 8392 9432
rect 8386 9392 8392 9404
rect 8444 9392 8450 9444
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9364 1639 9367
rect 1854 9364 1860 9376
rect 1627 9336 1860 9364
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 1854 9324 1860 9336
rect 1912 9324 1918 9376
rect 2130 9324 2136 9376
rect 2188 9364 2194 9376
rect 2590 9364 2596 9376
rect 2188 9336 2233 9364
rect 2551 9336 2596 9364
rect 2188 9324 2194 9336
rect 2590 9324 2596 9336
rect 2648 9324 2654 9376
rect 3602 9324 3608 9376
rect 3660 9364 3666 9376
rect 3697 9367 3755 9373
rect 3697 9364 3709 9367
rect 3660 9336 3709 9364
rect 3660 9324 3666 9336
rect 3697 9333 3709 9336
rect 3743 9333 3755 9367
rect 3697 9327 3755 9333
rect 3878 9324 3884 9376
rect 3936 9364 3942 9376
rect 4065 9367 4123 9373
rect 4065 9364 4077 9367
rect 3936 9336 4077 9364
rect 3936 9324 3942 9336
rect 4065 9333 4077 9336
rect 4111 9333 4123 9367
rect 4065 9327 4123 9333
rect 4614 9324 4620 9376
rect 4672 9364 4678 9376
rect 6454 9364 6460 9376
rect 4672 9336 6460 9364
rect 4672 9324 4678 9336
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 7742 9324 7748 9376
rect 7800 9364 7806 9376
rect 7929 9367 7987 9373
rect 7929 9364 7941 9367
rect 7800 9336 7941 9364
rect 7800 9324 7806 9336
rect 7929 9333 7941 9336
rect 7975 9333 7987 9367
rect 8496 9364 8524 9540
rect 8573 9537 8585 9571
rect 8619 9568 8631 9571
rect 8938 9568 8944 9580
rect 8619 9540 8944 9568
rect 8619 9537 8631 9540
rect 8573 9531 8631 9537
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 9490 9528 9496 9580
rect 9548 9568 9554 9580
rect 9548 9540 9904 9568
rect 9548 9528 9554 9540
rect 9677 9503 9735 9509
rect 8680 9472 8892 9500
rect 8570 9392 8576 9444
rect 8628 9432 8634 9444
rect 8680 9432 8708 9472
rect 8628 9404 8708 9432
rect 8864 9432 8892 9472
rect 9677 9469 9689 9503
rect 9723 9500 9735 9503
rect 9766 9500 9772 9512
rect 9723 9472 9772 9500
rect 9723 9469 9735 9472
rect 9677 9463 9735 9469
rect 9766 9460 9772 9472
rect 9824 9460 9830 9512
rect 9876 9500 9904 9540
rect 9950 9528 9956 9580
rect 10008 9568 10014 9580
rect 10321 9571 10379 9577
rect 10321 9568 10333 9571
rect 10008 9540 10333 9568
rect 10008 9528 10014 9540
rect 10321 9537 10333 9540
rect 10367 9537 10379 9571
rect 10502 9568 10508 9580
rect 10463 9540 10508 9568
rect 10321 9531 10379 9537
rect 10502 9528 10508 9540
rect 10560 9528 10566 9580
rect 12452 9568 12480 9676
rect 13078 9664 13084 9676
rect 13136 9704 13142 9716
rect 13630 9704 13636 9716
rect 13136 9676 13636 9704
rect 13136 9664 13142 9676
rect 13630 9664 13636 9676
rect 13688 9664 13694 9716
rect 13906 9704 13912 9716
rect 13832 9676 13912 9704
rect 12529 9639 12587 9645
rect 12529 9605 12541 9639
rect 12575 9636 12587 9639
rect 12894 9636 12900 9648
rect 12575 9608 12900 9636
rect 12575 9605 12587 9608
rect 12529 9599 12587 9605
rect 12894 9596 12900 9608
rect 12952 9596 12958 9648
rect 13170 9568 13176 9580
rect 10612 9540 12480 9568
rect 13131 9540 13176 9568
rect 10612 9500 10640 9540
rect 13170 9528 13176 9540
rect 13228 9528 13234 9580
rect 13832 9500 13860 9676
rect 13906 9664 13912 9676
rect 13964 9664 13970 9716
rect 13998 9664 14004 9716
rect 14056 9704 14062 9716
rect 14182 9704 14188 9716
rect 14056 9676 14188 9704
rect 14056 9664 14062 9676
rect 14182 9664 14188 9676
rect 14240 9664 14246 9716
rect 16114 9704 16120 9716
rect 14752 9676 15700 9704
rect 16075 9676 16120 9704
rect 14752 9636 14780 9676
rect 9876 9472 10640 9500
rect 11716 9472 13860 9500
rect 13924 9608 14780 9636
rect 15672 9636 15700 9676
rect 16114 9664 16120 9676
rect 16172 9664 16178 9716
rect 17494 9664 17500 9716
rect 17552 9704 17558 9716
rect 17862 9704 17868 9716
rect 17552 9676 17868 9704
rect 17552 9664 17558 9676
rect 17862 9664 17868 9676
rect 17920 9664 17926 9716
rect 17218 9636 17224 9648
rect 15672 9608 17224 9636
rect 8864 9404 10364 9432
rect 8628 9392 8634 9404
rect 9122 9364 9128 9376
rect 8496 9336 9128 9364
rect 7929 9327 7987 9333
rect 9122 9324 9128 9336
rect 9180 9324 9186 9376
rect 9490 9364 9496 9376
rect 9451 9336 9496 9364
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 9858 9364 9864 9376
rect 9819 9336 9864 9364
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 10226 9364 10232 9376
rect 10187 9336 10232 9364
rect 10226 9324 10232 9336
rect 10284 9324 10290 9376
rect 10336 9364 10364 9404
rect 11716 9364 11744 9472
rect 12897 9435 12955 9441
rect 12897 9432 12909 9435
rect 12544 9404 12909 9432
rect 10336 9336 11744 9364
rect 12342 9324 12348 9376
rect 12400 9364 12406 9376
rect 12544 9364 12572 9404
rect 12897 9401 12909 9404
rect 12943 9401 12955 9435
rect 12897 9395 12955 9401
rect 12400 9336 12572 9364
rect 12989 9367 13047 9373
rect 12400 9324 12406 9336
rect 12989 9333 13001 9367
rect 13035 9364 13047 9367
rect 13924 9364 13952 9608
rect 17218 9596 17224 9608
rect 17276 9596 17282 9648
rect 14458 9528 14464 9580
rect 14516 9568 14522 9580
rect 14737 9571 14795 9577
rect 14737 9568 14749 9571
rect 14516 9540 14749 9568
rect 14516 9528 14522 9540
rect 14737 9537 14749 9540
rect 14783 9537 14795 9571
rect 14737 9531 14795 9537
rect 16945 9571 17003 9577
rect 16945 9537 16957 9571
rect 16991 9568 17003 9571
rect 17954 9568 17960 9580
rect 16991 9540 17960 9568
rect 16991 9537 17003 9540
rect 16945 9531 17003 9537
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 14274 9500 14280 9512
rect 14235 9472 14280 9500
rect 14274 9460 14280 9472
rect 14332 9460 14338 9512
rect 15562 9460 15568 9512
rect 15620 9500 15626 9512
rect 16206 9500 16212 9512
rect 15620 9472 16212 9500
rect 15620 9460 15626 9472
rect 16206 9460 16212 9472
rect 16264 9460 16270 9512
rect 16666 9460 16672 9512
rect 16724 9500 16730 9512
rect 16724 9472 17172 9500
rect 16724 9460 16730 9472
rect 15004 9435 15062 9441
rect 15004 9401 15016 9435
rect 15050 9432 15062 9435
rect 15470 9432 15476 9444
rect 15050 9404 15476 9432
rect 15050 9401 15062 9404
rect 15004 9395 15062 9401
rect 15470 9392 15476 9404
rect 15528 9392 15534 9444
rect 15746 9392 15752 9444
rect 15804 9432 15810 9444
rect 17034 9432 17040 9444
rect 15804 9404 17040 9432
rect 15804 9392 15810 9404
rect 17034 9392 17040 9404
rect 17092 9392 17098 9444
rect 17144 9432 17172 9472
rect 17862 9460 17868 9512
rect 17920 9500 17926 9512
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 17920 9472 18061 9500
rect 17920 9460 17926 9472
rect 18049 9469 18061 9472
rect 18095 9469 18107 9503
rect 18049 9463 18107 9469
rect 18598 9460 18604 9512
rect 18656 9500 18662 9512
rect 20257 9503 20315 9509
rect 20257 9500 20269 9503
rect 18656 9472 20269 9500
rect 18656 9460 18662 9472
rect 20257 9469 20269 9472
rect 20303 9469 20315 9503
rect 20257 9463 20315 9469
rect 18294 9435 18352 9441
rect 18294 9432 18306 9435
rect 17144 9404 18306 9432
rect 18294 9401 18306 9404
rect 18340 9432 18352 9435
rect 18782 9432 18788 9444
rect 18340 9404 18788 9432
rect 18340 9401 18352 9404
rect 18294 9395 18352 9401
rect 18782 9392 18788 9404
rect 18840 9392 18846 9444
rect 13035 9336 13952 9364
rect 13035 9333 13047 9336
rect 12989 9327 13047 9333
rect 13998 9324 14004 9376
rect 14056 9364 14062 9376
rect 14093 9367 14151 9373
rect 14093 9364 14105 9367
rect 14056 9336 14105 9364
rect 14056 9324 14062 9336
rect 14093 9333 14105 9336
rect 14139 9333 14151 9367
rect 14093 9327 14151 9333
rect 14274 9324 14280 9376
rect 14332 9364 14338 9376
rect 19242 9364 19248 9376
rect 14332 9336 19248 9364
rect 14332 9324 14338 9336
rect 19242 9324 19248 9336
rect 19300 9324 19306 9376
rect 19426 9364 19432 9376
rect 19387 9336 19432 9364
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 1397 9163 1455 9169
rect 1397 9129 1409 9163
rect 1443 9160 1455 9163
rect 1578 9160 1584 9172
rect 1443 9132 1584 9160
rect 1443 9129 1455 9132
rect 1397 9123 1455 9129
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 3237 9163 3295 9169
rect 3237 9129 3249 9163
rect 3283 9160 3295 9163
rect 3326 9160 3332 9172
rect 3283 9132 3332 9160
rect 3283 9129 3295 9132
rect 3237 9123 3295 9129
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 3602 9120 3608 9172
rect 3660 9160 3666 9172
rect 4154 9160 4160 9172
rect 3660 9132 4160 9160
rect 3660 9120 3666 9132
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 4433 9163 4491 9169
rect 4433 9129 4445 9163
rect 4479 9160 4491 9163
rect 4706 9160 4712 9172
rect 4479 9132 4712 9160
rect 4479 9129 4491 9132
rect 4433 9123 4491 9129
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9129 5503 9163
rect 5445 9123 5503 9129
rect 5813 9163 5871 9169
rect 5813 9129 5825 9163
rect 5859 9160 5871 9163
rect 6178 9160 6184 9172
rect 5859 9132 6184 9160
rect 5859 9129 5871 9132
rect 5813 9123 5871 9129
rect 1302 9052 1308 9104
rect 1360 9092 1366 9104
rect 2590 9092 2596 9104
rect 1360 9064 2596 9092
rect 1360 9052 1366 9064
rect 2590 9052 2596 9064
rect 2648 9052 2654 9104
rect 2869 9095 2927 9101
rect 2869 9061 2881 9095
rect 2915 9092 2927 9095
rect 4614 9092 4620 9104
rect 2915 9064 4620 9092
rect 2915 9061 2927 9064
rect 2869 9055 2927 9061
rect 4614 9052 4620 9064
rect 4672 9052 4678 9104
rect 5460 9092 5488 9123
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 7650 9120 7656 9172
rect 7708 9160 7714 9172
rect 9766 9160 9772 9172
rect 7708 9132 9772 9160
rect 7708 9120 7714 9132
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 9861 9163 9919 9169
rect 9861 9129 9873 9163
rect 9907 9160 9919 9163
rect 10226 9160 10232 9172
rect 9907 9132 10232 9160
rect 9907 9129 9919 9132
rect 9861 9123 9919 9129
rect 10226 9120 10232 9132
rect 10284 9120 10290 9172
rect 12342 9160 12348 9172
rect 10336 9132 11468 9160
rect 12303 9132 12348 9160
rect 5902 9092 5908 9104
rect 5460 9064 5908 9092
rect 5902 9052 5908 9064
rect 5960 9052 5966 9104
rect 6012 9064 6224 9092
rect 1762 9024 1768 9036
rect 1723 8996 1768 9024
rect 1762 8984 1768 8996
rect 1820 8984 1826 9036
rect 1854 8984 1860 9036
rect 1912 9024 1918 9036
rect 1912 8996 1957 9024
rect 1912 8984 1918 8996
rect 2774 8984 2780 9036
rect 2832 9024 2838 9036
rect 3602 9024 3608 9036
rect 2832 8996 2877 9024
rect 2976 8996 3608 9024
rect 2832 8984 2838 8996
rect 2041 8959 2099 8965
rect 2041 8925 2053 8959
rect 2087 8956 2099 8959
rect 2130 8956 2136 8968
rect 2087 8928 2136 8956
rect 2087 8925 2099 8928
rect 2041 8919 2099 8925
rect 2130 8916 2136 8928
rect 2188 8916 2194 8968
rect 2682 8916 2688 8968
rect 2740 8956 2746 8968
rect 2976 8956 3004 8996
rect 3602 8984 3608 8996
rect 3660 8984 3666 9036
rect 4430 8984 4436 9036
rect 4488 9024 4494 9036
rect 4893 9027 4951 9033
rect 4893 9024 4905 9027
rect 4488 8996 4905 9024
rect 4488 8984 4494 8996
rect 4893 8993 4905 8996
rect 4939 8993 4951 9027
rect 5166 9024 5172 9036
rect 4893 8987 4951 8993
rect 5000 8996 5172 9024
rect 2740 8928 3004 8956
rect 3053 8959 3111 8965
rect 2740 8916 2746 8928
rect 3053 8925 3065 8959
rect 3099 8956 3111 8959
rect 4522 8956 4528 8968
rect 3099 8928 4384 8956
rect 4483 8928 4528 8956
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 1854 8848 1860 8900
rect 1912 8888 1918 8900
rect 3970 8888 3976 8900
rect 1912 8860 3976 8888
rect 1912 8848 1918 8860
rect 3970 8848 3976 8860
rect 4028 8848 4034 8900
rect 4065 8891 4123 8897
rect 4065 8857 4077 8891
rect 4111 8888 4123 8891
rect 4154 8888 4160 8900
rect 4111 8860 4160 8888
rect 4111 8857 4123 8860
rect 4065 8851 4123 8857
rect 4154 8848 4160 8860
rect 4212 8848 4218 8900
rect 4356 8888 4384 8928
rect 4522 8916 4528 8928
rect 4580 8916 4586 8968
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8956 4767 8959
rect 5000 8956 5028 8996
rect 5166 8984 5172 8996
rect 5224 8984 5230 9036
rect 6012 9024 6040 9064
rect 5460 8996 6040 9024
rect 4755 8928 5028 8956
rect 5077 8959 5135 8965
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5350 8956 5356 8968
rect 5123 8928 5356 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5350 8916 5356 8928
rect 5408 8916 5414 8968
rect 4982 8888 4988 8900
rect 4356 8860 4988 8888
rect 4982 8848 4988 8860
rect 5040 8848 5046 8900
rect 5166 8848 5172 8900
rect 5224 8888 5230 8900
rect 5460 8888 5488 8996
rect 6086 8984 6092 9036
rect 6144 8984 6150 9036
rect 6196 9024 6224 9064
rect 6270 9052 6276 9104
rect 6328 9092 6334 9104
rect 6546 9092 6552 9104
rect 6328 9064 6552 9092
rect 6328 9052 6334 9064
rect 6546 9052 6552 9064
rect 6604 9052 6610 9104
rect 6730 9052 6736 9104
rect 6788 9092 6794 9104
rect 7469 9095 7527 9101
rect 7469 9092 7481 9095
rect 6788 9064 7481 9092
rect 6788 9052 6794 9064
rect 7469 9061 7481 9064
rect 7515 9061 7527 9095
rect 7469 9055 7527 9061
rect 7558 9052 7564 9104
rect 7616 9092 7622 9104
rect 7926 9092 7932 9104
rect 7616 9064 7932 9092
rect 7616 9052 7622 9064
rect 7926 9052 7932 9064
rect 7984 9052 7990 9104
rect 8570 9092 8576 9104
rect 8531 9064 8576 9092
rect 8570 9052 8576 9064
rect 8628 9052 8634 9104
rect 9122 9052 9128 9104
rect 9180 9092 9186 9104
rect 10336 9092 10364 9132
rect 9180 9064 10364 9092
rect 9180 9052 9186 9064
rect 10594 9052 10600 9104
rect 10652 9052 10658 9104
rect 7377 9027 7435 9033
rect 6196 8996 7225 9024
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 5997 8959 6055 8965
rect 5997 8925 6009 8959
rect 6043 8956 6055 8959
rect 6104 8956 6132 8984
rect 7197 8956 7225 8996
rect 7377 8993 7389 9027
rect 7423 9024 7435 9027
rect 8938 9024 8944 9036
rect 7423 8996 8944 9024
rect 7423 8993 7435 8996
rect 7377 8987 7435 8993
rect 8938 8984 8944 8996
rect 8996 8984 9002 9036
rect 10226 9024 10232 9036
rect 10187 8996 10232 9024
rect 10226 8984 10232 8996
rect 10284 8984 10290 9036
rect 10321 9027 10379 9033
rect 10321 8993 10333 9027
rect 10367 9024 10379 9027
rect 10612 9024 10640 9052
rect 11146 9024 11152 9036
rect 10367 8996 11152 9024
rect 10367 8993 10379 8996
rect 10321 8987 10379 8993
rect 11146 8984 11152 8996
rect 11204 8984 11210 9036
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 6043 8928 6132 8956
rect 6196 8928 7135 8956
rect 7197 8928 7573 8956
rect 6043 8925 6055 8928
rect 5997 8919 6055 8925
rect 5224 8860 5488 8888
rect 5224 8848 5230 8860
rect 2409 8823 2467 8829
rect 2409 8789 2421 8823
rect 2455 8820 2467 8823
rect 2682 8820 2688 8832
rect 2455 8792 2688 8820
rect 2455 8789 2467 8792
rect 2409 8783 2467 8789
rect 2682 8780 2688 8792
rect 2740 8780 2746 8832
rect 3988 8820 4016 8848
rect 5920 8820 5948 8919
rect 6196 8888 6224 8928
rect 6012 8860 6224 8888
rect 6012 8832 6040 8860
rect 6454 8848 6460 8900
rect 6512 8888 6518 8900
rect 7009 8891 7067 8897
rect 7009 8888 7021 8891
rect 6512 8860 7021 8888
rect 6512 8848 6518 8860
rect 7009 8857 7021 8860
rect 7055 8857 7067 8891
rect 7107 8888 7135 8928
rect 7561 8925 7573 8928
rect 7607 8925 7619 8959
rect 7561 8919 7619 8925
rect 7834 8916 7840 8968
rect 7892 8956 7898 8968
rect 8386 8956 8392 8968
rect 7892 8928 8392 8956
rect 7892 8916 7898 8928
rect 8386 8916 8392 8928
rect 8444 8916 8450 8968
rect 8570 8916 8576 8968
rect 8628 8956 8634 8968
rect 9950 8956 9956 8968
rect 8628 8928 9956 8956
rect 8628 8916 8634 8928
rect 9950 8916 9956 8928
rect 10008 8916 10014 8968
rect 10505 8959 10563 8965
rect 10505 8925 10517 8959
rect 10551 8956 10563 8959
rect 10594 8956 10600 8968
rect 10551 8928 10600 8956
rect 10551 8925 10563 8928
rect 10505 8919 10563 8925
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 11440 8956 11468 9132
rect 12342 9120 12348 9132
rect 12400 9120 12406 9172
rect 12805 9163 12863 9169
rect 12805 9129 12817 9163
rect 12851 9160 12863 9163
rect 13814 9160 13820 9172
rect 12851 9132 13820 9160
rect 12851 9129 12863 9132
rect 12805 9123 12863 9129
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 13909 9163 13967 9169
rect 13909 9129 13921 9163
rect 13955 9160 13967 9163
rect 14090 9160 14096 9172
rect 13955 9132 14096 9160
rect 13955 9129 13967 9132
rect 13909 9123 13967 9129
rect 14090 9120 14096 9132
rect 14148 9120 14154 9172
rect 14185 9163 14243 9169
rect 14185 9129 14197 9163
rect 14231 9160 14243 9163
rect 14231 9132 14320 9160
rect 14231 9129 14243 9132
rect 14185 9123 14243 9129
rect 13998 9092 14004 9104
rect 11900 9064 14004 9092
rect 11900 9033 11928 9064
rect 13998 9052 14004 9064
rect 14056 9092 14062 9104
rect 14056 9064 14136 9092
rect 14056 9052 14062 9064
rect 14108 9033 14136 9064
rect 11885 9027 11943 9033
rect 11885 8993 11897 9027
rect 11931 8993 11943 9027
rect 11885 8987 11943 8993
rect 12713 9027 12771 9033
rect 12713 8993 12725 9027
rect 12759 8993 12771 9027
rect 12713 8987 12771 8993
rect 14085 9027 14143 9033
rect 14085 8993 14097 9027
rect 14131 8993 14143 9027
rect 14292 9024 14320 9132
rect 14458 9120 14464 9172
rect 14516 9160 14522 9172
rect 16206 9160 16212 9172
rect 14516 9132 16212 9160
rect 14516 9120 14522 9132
rect 16206 9120 16212 9132
rect 16264 9160 16270 9172
rect 17862 9160 17868 9172
rect 16264 9132 17868 9160
rect 16264 9120 16270 9132
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 18874 9160 18880 9172
rect 18835 9132 18880 9160
rect 18874 9120 18880 9132
rect 18932 9120 18938 9172
rect 14734 9052 14740 9104
rect 14792 9092 14798 9104
rect 19058 9092 19064 9104
rect 14792 9064 19064 9092
rect 14792 9052 14798 9064
rect 19058 9052 19064 9064
rect 19116 9092 19122 9104
rect 19426 9092 19432 9104
rect 19116 9064 19432 9092
rect 19116 9052 19122 9064
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 14292 8996 15516 9024
rect 14085 8987 14143 8993
rect 12728 8956 12756 8987
rect 11440 8928 12756 8956
rect 12897 8959 12955 8965
rect 12897 8925 12909 8959
rect 12943 8956 12955 8959
rect 13814 8956 13820 8968
rect 12943 8928 13820 8956
rect 12943 8925 12955 8928
rect 12897 8919 12955 8925
rect 7107 8860 12480 8888
rect 7009 8851 7067 8857
rect 3988 8792 5948 8820
rect 5994 8780 6000 8832
rect 6052 8780 6058 8832
rect 6086 8780 6092 8832
rect 6144 8820 6150 8832
rect 8294 8820 8300 8832
rect 6144 8792 8300 8820
rect 6144 8780 6150 8792
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 8386 8780 8392 8832
rect 8444 8820 8450 8832
rect 9122 8820 9128 8832
rect 8444 8792 9128 8820
rect 8444 8780 8450 8792
rect 9122 8780 9128 8792
rect 9180 8780 9186 8832
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 11701 8823 11759 8829
rect 11701 8820 11713 8823
rect 9732 8792 11713 8820
rect 9732 8780 9738 8792
rect 11701 8789 11713 8792
rect 11747 8820 11759 8823
rect 11974 8820 11980 8832
rect 11747 8792 11980 8820
rect 11747 8789 11759 8792
rect 11701 8783 11759 8789
rect 11974 8780 11980 8792
rect 12032 8820 12038 8832
rect 12342 8820 12348 8832
rect 12032 8792 12348 8820
rect 12032 8780 12038 8792
rect 12342 8780 12348 8792
rect 12400 8780 12406 8832
rect 12452 8820 12480 8860
rect 12526 8848 12532 8900
rect 12584 8888 12590 8900
rect 12912 8888 12940 8919
rect 13814 8916 13820 8928
rect 13872 8916 13878 8968
rect 15378 8956 15384 8968
rect 15304 8928 15384 8956
rect 15304 8897 15332 8928
rect 15378 8916 15384 8928
rect 15436 8916 15442 8968
rect 12584 8860 12940 8888
rect 15289 8891 15347 8897
rect 12584 8848 12590 8860
rect 15289 8857 15301 8891
rect 15335 8857 15347 8891
rect 15488 8888 15516 8996
rect 15562 8984 15568 9036
rect 15620 9024 15626 9036
rect 15657 9027 15715 9033
rect 15657 9024 15669 9027
rect 15620 8996 15669 9024
rect 15620 8984 15626 8996
rect 15657 8993 15669 8996
rect 15703 8993 15715 9027
rect 16390 9024 16396 9036
rect 15657 8987 15715 8993
rect 15856 8996 16396 9024
rect 15856 8968 15884 8996
rect 16390 8984 16396 8996
rect 16448 8984 16454 9036
rect 17405 9027 17463 9033
rect 17405 8993 17417 9027
rect 17451 9024 17463 9027
rect 18785 9027 18843 9033
rect 18785 9024 18797 9027
rect 17451 8996 18797 9024
rect 17451 8993 17463 8996
rect 17405 8987 17463 8993
rect 18785 8993 18797 8996
rect 18831 8993 18843 9027
rect 18785 8987 18843 8993
rect 15749 8959 15807 8965
rect 15749 8925 15761 8959
rect 15795 8956 15807 8959
rect 15838 8956 15844 8968
rect 15795 8928 15844 8956
rect 15795 8925 15807 8928
rect 15749 8919 15807 8925
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 15933 8959 15991 8965
rect 15933 8925 15945 8959
rect 15979 8956 15991 8959
rect 16022 8956 16028 8968
rect 15979 8928 16028 8956
rect 15979 8925 15991 8928
rect 15933 8919 15991 8925
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 18966 8956 18972 8968
rect 18927 8928 18972 8956
rect 18966 8916 18972 8928
rect 19024 8916 19030 8968
rect 16482 8888 16488 8900
rect 15488 8860 16488 8888
rect 15289 8851 15347 8857
rect 16482 8848 16488 8860
rect 16540 8848 16546 8900
rect 15746 8820 15752 8832
rect 12452 8792 15752 8820
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 16758 8780 16764 8832
rect 16816 8820 16822 8832
rect 18417 8823 18475 8829
rect 18417 8820 18429 8823
rect 16816 8792 18429 8820
rect 16816 8780 16822 8792
rect 18417 8789 18429 8792
rect 18463 8789 18475 8823
rect 18417 8783 18475 8789
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 1118 8576 1124 8628
rect 1176 8616 1182 8628
rect 1176 8588 4936 8616
rect 1176 8576 1182 8588
rect 2869 8551 2927 8557
rect 2869 8517 2881 8551
rect 2915 8548 2927 8551
rect 3602 8548 3608 8560
rect 2915 8520 3608 8548
rect 2915 8517 2927 8520
rect 2869 8511 2927 8517
rect 3602 8508 3608 8520
rect 3660 8508 3666 8560
rect 2590 8440 2596 8492
rect 2648 8480 2654 8492
rect 3145 8483 3203 8489
rect 3145 8480 3157 8483
rect 2648 8452 3157 8480
rect 2648 8440 2654 8452
rect 3145 8449 3157 8452
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 1489 8415 1547 8421
rect 1489 8381 1501 8415
rect 1535 8381 1547 8415
rect 1489 8375 1547 8381
rect 1756 8415 1814 8421
rect 1756 8381 1768 8415
rect 1802 8412 1814 8415
rect 2866 8412 2872 8424
rect 1802 8384 2872 8412
rect 1802 8381 1814 8384
rect 1756 8375 1814 8381
rect 1504 8276 1532 8375
rect 2866 8372 2872 8384
rect 2924 8372 2930 8424
rect 2961 8415 3019 8421
rect 2961 8381 2973 8415
rect 3007 8381 3019 8415
rect 2961 8375 3019 8381
rect 2976 8344 3004 8375
rect 3326 8372 3332 8424
rect 3384 8412 3390 8424
rect 3697 8415 3755 8421
rect 3697 8412 3709 8415
rect 3384 8384 3709 8412
rect 3384 8372 3390 8384
rect 3697 8381 3709 8384
rect 3743 8381 3755 8415
rect 4908 8412 4936 8588
rect 4982 8576 4988 8628
rect 5040 8616 5046 8628
rect 5077 8619 5135 8625
rect 5077 8616 5089 8619
rect 5040 8588 5089 8616
rect 5040 8576 5046 8588
rect 5077 8585 5089 8588
rect 5123 8585 5135 8619
rect 5626 8616 5632 8628
rect 5077 8579 5135 8585
rect 5184 8588 5632 8616
rect 4982 8440 4988 8492
rect 5040 8480 5046 8492
rect 5184 8480 5212 8588
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 5721 8619 5779 8625
rect 5721 8585 5733 8619
rect 5767 8616 5779 8619
rect 5994 8616 6000 8628
rect 5767 8588 6000 8616
rect 5767 8585 5779 8588
rect 5721 8579 5779 8585
rect 5994 8576 6000 8588
rect 6052 8576 6058 8628
rect 6546 8576 6552 8628
rect 6604 8616 6610 8628
rect 6604 8588 8432 8616
rect 6604 8576 6610 8588
rect 5258 8508 5264 8560
rect 5316 8548 5322 8560
rect 5445 8551 5503 8557
rect 5445 8548 5457 8551
rect 5316 8520 5457 8548
rect 5316 8508 5322 8520
rect 5445 8517 5457 8520
rect 5491 8517 5503 8551
rect 6270 8548 6276 8560
rect 5445 8511 5503 8517
rect 5552 8520 6276 8548
rect 5040 8452 5212 8480
rect 5040 8440 5046 8452
rect 5552 8412 5580 8520
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 7466 8508 7472 8560
rect 7524 8548 7530 8560
rect 7561 8551 7619 8557
rect 7561 8548 7573 8551
rect 7524 8520 7573 8548
rect 7524 8508 7530 8520
rect 7561 8517 7573 8520
rect 7607 8517 7619 8551
rect 7561 8511 7619 8517
rect 7659 8520 8340 8548
rect 6362 8480 6368 8492
rect 5920 8452 6368 8480
rect 5920 8424 5948 8452
rect 6362 8440 6368 8452
rect 6420 8440 6426 8492
rect 6546 8440 6552 8492
rect 6604 8480 6610 8492
rect 7659 8480 7687 8520
rect 6604 8452 7687 8480
rect 6604 8440 6610 8452
rect 7742 8440 7748 8492
rect 7800 8480 7806 8492
rect 8021 8483 8079 8489
rect 8021 8480 8033 8483
rect 7800 8452 8033 8480
rect 7800 8440 7806 8452
rect 8021 8449 8033 8452
rect 8067 8449 8079 8483
rect 8202 8480 8208 8492
rect 8163 8452 8208 8480
rect 8021 8443 8079 8449
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 4908 8384 5580 8412
rect 5629 8415 5687 8421
rect 3697 8375 3755 8381
rect 5629 8381 5641 8415
rect 5675 8381 5687 8415
rect 5629 8375 5687 8381
rect 3964 8347 4022 8353
rect 2976 8316 3924 8344
rect 2498 8276 2504 8288
rect 1504 8248 2504 8276
rect 2498 8236 2504 8248
rect 2556 8276 2562 8288
rect 3326 8276 3332 8288
rect 2556 8248 3332 8276
rect 2556 8236 2562 8248
rect 3326 8236 3332 8248
rect 3384 8236 3390 8288
rect 3896 8276 3924 8316
rect 3964 8313 3976 8347
rect 4010 8344 4022 8347
rect 4430 8344 4436 8356
rect 4010 8316 4436 8344
rect 4010 8313 4022 8316
rect 3964 8307 4022 8313
rect 4430 8304 4436 8316
rect 4488 8344 4494 8356
rect 5166 8344 5172 8356
rect 4488 8316 5172 8344
rect 4488 8304 4494 8316
rect 5166 8304 5172 8316
rect 5224 8304 5230 8356
rect 5644 8344 5672 8375
rect 5902 8372 5908 8424
rect 5960 8372 5966 8424
rect 6089 8415 6147 8421
rect 6089 8381 6101 8415
rect 6135 8412 6147 8415
rect 7098 8412 7104 8424
rect 6135 8384 7104 8412
rect 6135 8381 6147 8384
rect 6089 8375 6147 8381
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 7926 8412 7932 8424
rect 7887 8384 7932 8412
rect 7926 8372 7932 8384
rect 7984 8372 7990 8424
rect 8312 8412 8340 8520
rect 8404 8480 8432 8588
rect 9122 8576 9128 8628
rect 9180 8616 9186 8628
rect 9766 8616 9772 8628
rect 9180 8588 9772 8616
rect 9180 8576 9186 8588
rect 9766 8576 9772 8588
rect 9824 8576 9830 8628
rect 9950 8576 9956 8628
rect 10008 8616 10014 8628
rect 10594 8616 10600 8628
rect 10008 8588 10600 8616
rect 10008 8576 10014 8588
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 14001 8619 14059 8625
rect 14001 8585 14013 8619
rect 14047 8616 14059 8619
rect 14274 8616 14280 8628
rect 14047 8588 14280 8616
rect 14047 8585 14059 8588
rect 14001 8579 14059 8585
rect 14274 8576 14280 8588
rect 14332 8576 14338 8628
rect 15470 8616 15476 8628
rect 15431 8588 15476 8616
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 19429 8619 19487 8625
rect 19429 8616 19441 8619
rect 18064 8588 19441 8616
rect 12526 8548 12532 8560
rect 9232 8520 12532 8548
rect 9232 8489 9260 8520
rect 12526 8508 12532 8520
rect 12584 8508 12590 8560
rect 12618 8508 12624 8560
rect 12676 8548 12682 8560
rect 16393 8551 16451 8557
rect 12676 8520 14136 8548
rect 12676 8508 12682 8520
rect 9125 8483 9183 8489
rect 9125 8480 9137 8483
rect 8404 8452 9137 8480
rect 9125 8449 9137 8452
rect 9171 8449 9183 8483
rect 9125 8443 9183 8449
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8449 9275 8483
rect 10226 8480 10232 8492
rect 10187 8452 10232 8480
rect 9217 8443 9275 8449
rect 10226 8440 10232 8452
rect 10284 8440 10290 8492
rect 14108 8489 14136 8520
rect 16393 8517 16405 8551
rect 16439 8548 16451 8551
rect 17954 8548 17960 8560
rect 16439 8520 17960 8548
rect 16439 8517 16451 8520
rect 16393 8511 16451 8517
rect 17954 8508 17960 8520
rect 18012 8508 18018 8560
rect 14001 8483 14059 8489
rect 14001 8480 14013 8483
rect 10336 8452 14013 8480
rect 8312 8384 9628 8412
rect 9490 8344 9496 8356
rect 5644 8316 9496 8344
rect 9490 8304 9496 8316
rect 9548 8304 9554 8356
rect 9600 8344 9628 8384
rect 9766 8372 9772 8424
rect 9824 8412 9830 8424
rect 10336 8412 10364 8452
rect 14001 8449 14013 8452
rect 14047 8449 14059 8483
rect 14001 8443 14059 8449
rect 14093 8483 14151 8489
rect 14093 8449 14105 8483
rect 14139 8449 14151 8483
rect 16942 8480 16948 8492
rect 16903 8452 16948 8480
rect 14093 8443 14151 8449
rect 16942 8440 16948 8452
rect 17000 8480 17006 8492
rect 17862 8480 17868 8492
rect 17000 8452 17868 8480
rect 17000 8440 17006 8452
rect 17862 8440 17868 8452
rect 17920 8480 17926 8492
rect 18064 8480 18092 8588
rect 19429 8585 19441 8588
rect 19475 8585 19487 8619
rect 19429 8579 19487 8585
rect 17920 8452 18092 8480
rect 17920 8440 17926 8452
rect 9824 8384 10364 8412
rect 9824 8372 9830 8384
rect 10594 8372 10600 8424
rect 10652 8412 10658 8424
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 10652 8384 12909 8412
rect 10652 8372 10658 8384
rect 12897 8381 12909 8384
rect 12943 8381 12955 8415
rect 16758 8412 16764 8424
rect 12897 8375 12955 8381
rect 14200 8384 14504 8412
rect 16719 8384 16764 8412
rect 11333 8347 11391 8353
rect 11333 8344 11345 8347
rect 9600 8316 11345 8344
rect 11333 8313 11345 8316
rect 11379 8313 11391 8347
rect 11333 8307 11391 8313
rect 11422 8304 11428 8356
rect 11480 8344 11486 8356
rect 14200 8344 14228 8384
rect 11480 8316 14228 8344
rect 11480 8304 11486 8316
rect 14274 8304 14280 8356
rect 14332 8353 14338 8356
rect 14332 8347 14396 8353
rect 14332 8313 14350 8347
rect 14384 8313 14396 8347
rect 14476 8344 14504 8384
rect 16758 8372 16764 8384
rect 16816 8372 16822 8424
rect 18046 8412 18052 8424
rect 18007 8384 18052 8412
rect 18046 8372 18052 8384
rect 18104 8372 18110 8424
rect 16853 8347 16911 8353
rect 16853 8344 16865 8347
rect 14476 8316 16865 8344
rect 14332 8307 14396 8313
rect 16853 8313 16865 8316
rect 16899 8313 16911 8347
rect 16853 8307 16911 8313
rect 14332 8304 14338 8307
rect 17218 8304 17224 8356
rect 17276 8344 17282 8356
rect 18294 8347 18352 8353
rect 18294 8344 18306 8347
rect 17276 8316 18306 8344
rect 17276 8304 17282 8316
rect 18294 8313 18306 8316
rect 18340 8344 18352 8347
rect 18966 8344 18972 8356
rect 18340 8316 18972 8344
rect 18340 8313 18352 8316
rect 18294 8307 18352 8313
rect 18966 8304 18972 8316
rect 19024 8304 19030 8356
rect 20254 8344 20260 8356
rect 20215 8316 20260 8344
rect 20254 8304 20260 8316
rect 20312 8304 20318 8356
rect 4706 8276 4712 8288
rect 3896 8248 4712 8276
rect 4706 8236 4712 8248
rect 4764 8236 4770 8288
rect 5074 8236 5080 8288
rect 5132 8276 5138 8288
rect 6086 8276 6092 8288
rect 5132 8248 6092 8276
rect 5132 8236 5138 8248
rect 6086 8236 6092 8248
rect 6144 8236 6150 8288
rect 6181 8279 6239 8285
rect 6181 8245 6193 8279
rect 6227 8276 6239 8279
rect 6822 8276 6828 8288
rect 6227 8248 6828 8276
rect 6227 8245 6239 8248
rect 6181 8239 6239 8245
rect 6822 8236 6828 8248
rect 6880 8236 6886 8288
rect 7098 8236 7104 8288
rect 7156 8276 7162 8288
rect 8570 8276 8576 8288
rect 7156 8248 8576 8276
rect 7156 8236 7162 8248
rect 8570 8236 8576 8248
rect 8628 8236 8634 8288
rect 9125 8279 9183 8285
rect 9125 8245 9137 8279
rect 9171 8276 9183 8279
rect 15654 8276 15660 8288
rect 9171 8248 15660 8276
rect 9171 8245 9183 8248
rect 9125 8239 9183 8245
rect 15654 8236 15660 8248
rect 15712 8236 15718 8288
rect 16758 8236 16764 8288
rect 16816 8276 16822 8288
rect 18598 8276 18604 8288
rect 16816 8248 18604 8276
rect 16816 8236 16822 8248
rect 18598 8236 18604 8248
rect 18656 8236 18662 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 1946 8032 1952 8084
rect 2004 8072 2010 8084
rect 2409 8075 2467 8081
rect 2409 8072 2421 8075
rect 2004 8044 2421 8072
rect 2004 8032 2010 8044
rect 2409 8041 2421 8044
rect 2455 8041 2467 8075
rect 2409 8035 2467 8041
rect 2869 8075 2927 8081
rect 2869 8041 2881 8075
rect 2915 8072 2927 8075
rect 4338 8072 4344 8084
rect 2915 8044 4344 8072
rect 2915 8041 2927 8044
rect 2869 8035 2927 8041
rect 4338 8032 4344 8044
rect 4396 8032 4402 8084
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 4798 8072 4804 8084
rect 4571 8044 4804 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 4798 8032 4804 8044
rect 4856 8032 4862 8084
rect 4893 8075 4951 8081
rect 4893 8041 4905 8075
rect 4939 8072 4951 8075
rect 5258 8072 5264 8084
rect 4939 8044 5264 8072
rect 4939 8041 4951 8044
rect 4893 8035 4951 8041
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 6638 8072 6644 8084
rect 6599 8044 6644 8072
rect 6638 8032 6644 8044
rect 6696 8032 6702 8084
rect 6730 8032 6736 8084
rect 6788 8072 6794 8084
rect 7193 8075 7251 8081
rect 7193 8072 7205 8075
rect 6788 8044 7205 8072
rect 6788 8032 6794 8044
rect 7193 8041 7205 8044
rect 7239 8041 7251 8075
rect 7193 8035 7251 8041
rect 10502 8032 10508 8084
rect 10560 8072 10566 8084
rect 11057 8075 11115 8081
rect 11057 8072 11069 8075
rect 10560 8044 11069 8072
rect 10560 8032 10566 8044
rect 11057 8041 11069 8044
rect 11103 8041 11115 8075
rect 11057 8035 11115 8041
rect 11977 8075 12035 8081
rect 11977 8041 11989 8075
rect 12023 8072 12035 8075
rect 12158 8072 12164 8084
rect 12023 8044 12164 8072
rect 12023 8041 12035 8044
rect 11977 8035 12035 8041
rect 12158 8032 12164 8044
rect 12216 8072 12222 8084
rect 12342 8072 12348 8084
rect 12216 8044 12348 8072
rect 12216 8032 12222 8044
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 12529 8075 12587 8081
rect 12529 8041 12541 8075
rect 12575 8072 12587 8075
rect 13078 8072 13084 8084
rect 12575 8044 13084 8072
rect 12575 8041 12587 8044
rect 12529 8035 12587 8041
rect 13078 8032 13084 8044
rect 13136 8032 13142 8084
rect 13630 8072 13636 8084
rect 13591 8044 13636 8072
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 13814 8032 13820 8084
rect 13872 8072 13878 8084
rect 14734 8072 14740 8084
rect 13872 8044 14740 8072
rect 13872 8032 13878 8044
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 15378 8032 15384 8084
rect 15436 8072 15442 8084
rect 15749 8075 15807 8081
rect 15749 8072 15761 8075
rect 15436 8044 15761 8072
rect 15436 8032 15442 8044
rect 15749 8041 15761 8044
rect 15795 8041 15807 8075
rect 18046 8072 18052 8084
rect 15749 8035 15807 8041
rect 17512 8044 18052 8072
rect 2777 8007 2835 8013
rect 2777 7973 2789 8007
rect 2823 8004 2835 8007
rect 2958 8004 2964 8016
rect 2823 7976 2964 8004
rect 2823 7973 2835 7976
rect 2777 7967 2835 7973
rect 2958 7964 2964 7976
rect 3016 7964 3022 8016
rect 14001 8007 14059 8013
rect 3068 7976 13952 8004
rect 1765 7939 1823 7945
rect 1765 7905 1777 7939
rect 1811 7936 1823 7939
rect 2314 7936 2320 7948
rect 1811 7908 2320 7936
rect 1811 7905 1823 7908
rect 1765 7899 1823 7905
rect 2314 7896 2320 7908
rect 2372 7896 2378 7948
rect 3068 7936 3096 7976
rect 4433 7939 4491 7945
rect 2792 7908 3096 7936
rect 3140 7908 4384 7936
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7837 1915 7871
rect 1857 7831 1915 7837
rect 2041 7871 2099 7877
rect 2041 7837 2053 7871
rect 2087 7868 2099 7871
rect 2792 7868 2820 7908
rect 2087 7840 2820 7868
rect 2087 7837 2099 7840
rect 2041 7831 2099 7837
rect 1872 7800 1900 7831
rect 2866 7828 2872 7880
rect 2924 7868 2930 7880
rect 2961 7871 3019 7877
rect 2961 7868 2973 7871
rect 2924 7840 2973 7868
rect 2924 7828 2930 7840
rect 2961 7837 2973 7840
rect 3007 7837 3019 7871
rect 2961 7831 3019 7837
rect 2317 7803 2375 7809
rect 2317 7800 2329 7803
rect 1872 7772 2329 7800
rect 2317 7769 2329 7772
rect 2363 7800 2375 7803
rect 2498 7800 2504 7812
rect 2363 7772 2504 7800
rect 2363 7769 2375 7772
rect 2317 7763 2375 7769
rect 2498 7760 2504 7772
rect 2556 7760 2562 7812
rect 1394 7732 1400 7744
rect 1355 7704 1400 7732
rect 1394 7692 1400 7704
rect 1452 7692 1458 7744
rect 1578 7692 1584 7744
rect 1636 7732 1642 7744
rect 2590 7732 2596 7744
rect 1636 7704 2596 7732
rect 1636 7692 1642 7704
rect 2590 7692 2596 7704
rect 2648 7692 2654 7744
rect 2958 7692 2964 7744
rect 3016 7732 3022 7744
rect 3140 7732 3168 7908
rect 4356 7868 4384 7908
rect 4433 7905 4445 7939
rect 4479 7936 4491 7939
rect 4614 7936 4620 7948
rect 4479 7908 4620 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 4614 7896 4620 7908
rect 4672 7896 4678 7948
rect 4890 7896 4896 7948
rect 4948 7936 4954 7948
rect 5074 7936 5080 7948
rect 4948 7908 5080 7936
rect 4948 7896 4954 7908
rect 5074 7896 5080 7908
rect 5132 7936 5138 7948
rect 5241 7939 5299 7945
rect 5241 7936 5253 7939
rect 5132 7908 5253 7936
rect 5132 7896 5138 7908
rect 5241 7905 5253 7908
rect 5287 7905 5299 7939
rect 5241 7899 5299 7905
rect 5810 7896 5816 7948
rect 5868 7936 5874 7948
rect 6457 7939 6515 7945
rect 5868 7908 6040 7936
rect 5868 7896 5874 7908
rect 4709 7871 4767 7877
rect 4709 7868 4721 7871
rect 4356 7840 4721 7868
rect 4709 7837 4721 7840
rect 4755 7837 4767 7871
rect 4709 7831 4767 7837
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7837 5043 7871
rect 6012 7868 6040 7908
rect 6457 7905 6469 7939
rect 6503 7905 6515 7939
rect 6457 7899 6515 7905
rect 6472 7868 6500 7899
rect 6822 7896 6828 7948
rect 6880 7936 6886 7948
rect 7098 7936 7104 7948
rect 6880 7908 7104 7936
rect 6880 7896 6886 7908
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 7558 7936 7564 7948
rect 7519 7908 7564 7936
rect 7558 7896 7564 7908
rect 7616 7896 7622 7948
rect 7653 7939 7711 7945
rect 7653 7905 7665 7939
rect 7699 7936 7711 7939
rect 8941 7939 8999 7945
rect 7699 7908 7880 7936
rect 7699 7905 7711 7908
rect 7653 7899 7711 7905
rect 7745 7871 7803 7877
rect 7745 7868 7757 7871
rect 6012 7840 6500 7868
rect 6564 7840 7757 7868
rect 4985 7831 5043 7837
rect 3326 7760 3332 7812
rect 3384 7800 3390 7812
rect 4893 7803 4951 7809
rect 4893 7800 4905 7803
rect 3384 7772 4905 7800
rect 3384 7760 3390 7772
rect 4893 7769 4905 7772
rect 4939 7800 4951 7803
rect 5000 7800 5028 7831
rect 4939 7772 5028 7800
rect 4939 7769 4951 7772
rect 4893 7763 4951 7769
rect 3016 7704 3168 7732
rect 4065 7735 4123 7741
rect 3016 7692 3022 7704
rect 4065 7701 4077 7735
rect 4111 7732 4123 7735
rect 6086 7732 6092 7744
rect 4111 7704 6092 7732
rect 4111 7701 4123 7704
rect 4065 7695 4123 7701
rect 6086 7692 6092 7704
rect 6144 7692 6150 7744
rect 6365 7735 6423 7741
rect 6365 7701 6377 7735
rect 6411 7732 6423 7735
rect 6454 7732 6460 7744
rect 6411 7704 6460 7732
rect 6411 7701 6423 7704
rect 6365 7695 6423 7701
rect 6454 7692 6460 7704
rect 6512 7732 6518 7744
rect 6564 7732 6592 7840
rect 7745 7837 7757 7840
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 7852 7800 7880 7908
rect 8941 7905 8953 7939
rect 8987 7936 8999 7939
rect 9490 7936 9496 7948
rect 8987 7908 9496 7936
rect 8987 7905 8999 7908
rect 8941 7899 8999 7905
rect 9490 7896 9496 7908
rect 9548 7896 9554 7948
rect 9674 7936 9680 7948
rect 9635 7908 9680 7936
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 9950 7945 9956 7948
rect 9944 7936 9956 7945
rect 9911 7908 9956 7936
rect 9944 7899 9956 7908
rect 9950 7896 9956 7899
rect 10008 7896 10014 7948
rect 11974 7896 11980 7948
rect 12032 7936 12038 7948
rect 12437 7939 12495 7945
rect 12437 7936 12449 7939
rect 12032 7908 12449 7936
rect 12032 7896 12038 7908
rect 12437 7905 12449 7908
rect 12483 7905 12495 7939
rect 13814 7936 13820 7948
rect 12437 7899 12495 7905
rect 12636 7908 13820 7936
rect 7926 7828 7932 7880
rect 7984 7868 7990 7880
rect 12526 7868 12532 7880
rect 7984 7840 8800 7868
rect 7984 7828 7990 7840
rect 8110 7800 8116 7812
rect 7852 7772 8116 7800
rect 8110 7760 8116 7772
rect 8168 7760 8174 7812
rect 8772 7809 8800 7840
rect 10980 7840 12532 7868
rect 10980 7812 11008 7840
rect 12526 7828 12532 7840
rect 12584 7828 12590 7880
rect 8757 7803 8815 7809
rect 8757 7769 8769 7803
rect 8803 7769 8815 7803
rect 8757 7763 8815 7769
rect 10962 7760 10968 7812
rect 11020 7760 11026 7812
rect 11977 7803 12035 7809
rect 11977 7800 11989 7803
rect 11072 7772 11989 7800
rect 6512 7704 6592 7732
rect 6512 7692 6518 7704
rect 6730 7692 6736 7744
rect 6788 7732 6794 7744
rect 8846 7732 8852 7744
rect 6788 7704 8852 7732
rect 6788 7692 6794 7704
rect 8846 7692 8852 7704
rect 8904 7692 8910 7744
rect 9858 7692 9864 7744
rect 9916 7732 9922 7744
rect 11072 7732 11100 7772
rect 11977 7769 11989 7772
rect 12023 7769 12035 7803
rect 11977 7763 12035 7769
rect 12069 7803 12127 7809
rect 12069 7769 12081 7803
rect 12115 7800 12127 7803
rect 12636 7800 12664 7908
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 13924 7936 13952 7976
rect 14001 7973 14013 8007
rect 14047 8004 14059 8007
rect 14090 8004 14096 8016
rect 14047 7976 14096 8004
rect 14047 7973 14059 7976
rect 14001 7967 14059 7973
rect 14090 7964 14096 7976
rect 14148 7964 14154 8016
rect 16942 8004 16948 8016
rect 15580 7976 16948 8004
rect 15580 7936 15608 7976
rect 16942 7964 16948 7976
rect 17000 7964 17006 8016
rect 13924 7908 15608 7936
rect 15654 7896 15660 7948
rect 15712 7936 15718 7948
rect 17512 7945 17540 8044
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 18690 8004 18696 8016
rect 17604 7976 18696 8004
rect 17497 7939 17555 7945
rect 15712 7908 15757 7936
rect 15712 7896 15718 7908
rect 17497 7905 17509 7939
rect 17543 7905 17555 7939
rect 17497 7899 17555 7905
rect 12713 7871 12771 7877
rect 12713 7837 12725 7871
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 12115 7772 12664 7800
rect 12728 7800 12756 7831
rect 12986 7828 12992 7880
rect 13044 7868 13050 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 13044 7840 14105 7868
rect 13044 7828 13050 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7868 14335 7871
rect 14366 7868 14372 7880
rect 14323 7840 14372 7868
rect 14323 7837 14335 7840
rect 14277 7831 14335 7837
rect 14366 7828 14372 7840
rect 14424 7828 14430 7880
rect 15470 7828 15476 7880
rect 15528 7868 15534 7880
rect 15841 7871 15899 7877
rect 15841 7868 15853 7871
rect 15528 7840 15853 7868
rect 15528 7828 15534 7840
rect 15841 7837 15853 7840
rect 15887 7837 15899 7871
rect 17604 7868 17632 7976
rect 18690 7964 18696 7976
rect 18748 7964 18754 8016
rect 17764 7939 17822 7945
rect 17764 7905 17776 7939
rect 17810 7936 17822 7939
rect 18046 7936 18052 7948
rect 17810 7908 18052 7936
rect 17810 7905 17822 7908
rect 17764 7899 17822 7905
rect 18046 7896 18052 7908
rect 18104 7896 18110 7948
rect 18598 7896 18604 7948
rect 18656 7936 18662 7948
rect 19705 7939 19763 7945
rect 19705 7936 19717 7939
rect 18656 7908 19717 7936
rect 18656 7896 18662 7908
rect 19705 7905 19717 7908
rect 19751 7905 19763 7939
rect 19705 7899 19763 7905
rect 15841 7831 15899 7837
rect 15948 7840 17632 7868
rect 13078 7800 13084 7812
rect 12728 7772 13084 7800
rect 12115 7769 12127 7772
rect 12069 7763 12127 7769
rect 13078 7760 13084 7772
rect 13136 7760 13142 7812
rect 15948 7800 15976 7840
rect 14292 7772 15976 7800
rect 9916 7704 11100 7732
rect 9916 7692 9922 7704
rect 12526 7692 12532 7744
rect 12584 7732 12590 7744
rect 14292 7732 14320 7772
rect 12584 7704 14320 7732
rect 15289 7735 15347 7741
rect 12584 7692 12590 7704
rect 15289 7701 15301 7735
rect 15335 7732 15347 7735
rect 15378 7732 15384 7744
rect 15335 7704 15384 7732
rect 15335 7701 15347 7704
rect 15289 7695 15347 7701
rect 15378 7692 15384 7704
rect 15436 7692 15442 7744
rect 16022 7692 16028 7744
rect 16080 7732 16086 7744
rect 17034 7732 17040 7744
rect 16080 7704 17040 7732
rect 16080 7692 16086 7704
rect 17034 7692 17040 7704
rect 17092 7732 17098 7744
rect 18877 7735 18935 7741
rect 18877 7732 18889 7735
rect 17092 7704 18889 7732
rect 17092 7692 17098 7704
rect 18877 7701 18889 7704
rect 18923 7701 18935 7735
rect 18877 7695 18935 7701
rect 18966 7692 18972 7744
rect 19024 7732 19030 7744
rect 19889 7735 19947 7741
rect 19889 7732 19901 7735
rect 19024 7704 19901 7732
rect 19024 7692 19030 7704
rect 19889 7701 19901 7704
rect 19935 7701 19947 7735
rect 19889 7695 19947 7701
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 1762 7488 1768 7540
rect 1820 7528 1826 7540
rect 2130 7528 2136 7540
rect 1820 7500 2136 7528
rect 1820 7488 1826 7500
rect 2130 7488 2136 7500
rect 2188 7488 2194 7540
rect 2225 7531 2283 7537
rect 2225 7497 2237 7531
rect 2271 7528 2283 7531
rect 2406 7528 2412 7540
rect 2271 7500 2412 7528
rect 2271 7497 2283 7500
rect 2225 7491 2283 7497
rect 2406 7488 2412 7500
rect 2464 7488 2470 7540
rect 2774 7488 2780 7540
rect 2832 7528 2838 7540
rect 4065 7531 4123 7537
rect 4065 7528 4077 7531
rect 2832 7500 4077 7528
rect 2832 7488 2838 7500
rect 4065 7497 4077 7500
rect 4111 7497 4123 7531
rect 4065 7491 4123 7497
rect 5626 7488 5632 7540
rect 5684 7528 5690 7540
rect 5721 7531 5779 7537
rect 5721 7528 5733 7531
rect 5684 7500 5733 7528
rect 5684 7488 5690 7500
rect 5721 7497 5733 7500
rect 5767 7497 5779 7531
rect 13078 7528 13084 7540
rect 5721 7491 5779 7497
rect 5828 7500 13084 7528
rect 5828 7460 5856 7500
rect 13078 7488 13084 7500
rect 13136 7488 13142 7540
rect 13170 7488 13176 7540
rect 13228 7528 13234 7540
rect 13446 7528 13452 7540
rect 13228 7500 13452 7528
rect 13228 7488 13234 7500
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 15746 7488 15752 7540
rect 15804 7528 15810 7540
rect 19429 7531 19487 7537
rect 19429 7528 19441 7531
rect 15804 7500 19441 7528
rect 15804 7488 15810 7500
rect 19429 7497 19441 7500
rect 19475 7528 19487 7531
rect 19475 7500 20116 7528
rect 19475 7497 19487 7500
rect 19429 7491 19487 7497
rect 2056 7432 5856 7460
rect 2056 7401 2084 7432
rect 6454 7420 6460 7472
rect 6512 7460 6518 7472
rect 6638 7460 6644 7472
rect 6512 7432 6644 7460
rect 6512 7420 6518 7432
rect 6638 7420 6644 7432
rect 6696 7420 6702 7472
rect 7834 7420 7840 7472
rect 7892 7460 7898 7472
rect 8205 7463 8263 7469
rect 8205 7460 8217 7463
rect 7892 7432 8217 7460
rect 7892 7420 7898 7432
rect 8205 7429 8217 7432
rect 8251 7429 8263 7463
rect 8205 7423 8263 7429
rect 8294 7420 8300 7472
rect 8352 7460 8358 7472
rect 9490 7460 9496 7472
rect 8352 7432 9496 7460
rect 8352 7420 8358 7432
rect 9490 7420 9496 7432
rect 9548 7420 9554 7472
rect 11517 7463 11575 7469
rect 11517 7429 11529 7463
rect 11563 7460 11575 7463
rect 12158 7460 12164 7472
rect 11563 7432 12164 7460
rect 11563 7429 11575 7432
rect 11517 7423 11575 7429
rect 12158 7420 12164 7432
rect 12216 7420 12222 7472
rect 15013 7463 15071 7469
rect 15013 7429 15025 7463
rect 15059 7460 15071 7463
rect 15059 7432 16620 7460
rect 15059 7429 15071 7432
rect 15013 7423 15071 7429
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7361 2099 7395
rect 2041 7355 2099 7361
rect 2590 7352 2596 7404
rect 2648 7392 2654 7404
rect 2685 7395 2743 7401
rect 2685 7392 2697 7395
rect 2648 7364 2697 7392
rect 2648 7352 2654 7364
rect 2685 7361 2697 7364
rect 2731 7361 2743 7395
rect 2685 7355 2743 7361
rect 2869 7395 2927 7401
rect 2869 7361 2881 7395
rect 2915 7392 2927 7395
rect 4246 7392 4252 7404
rect 2915 7364 4252 7392
rect 2915 7361 2927 7364
rect 2869 7355 2927 7361
rect 4246 7352 4252 7364
rect 4304 7352 4310 7404
rect 4338 7352 4344 7404
rect 4396 7392 4402 7404
rect 4617 7395 4675 7401
rect 4617 7392 4629 7395
rect 4396 7364 4629 7392
rect 4396 7352 4402 7364
rect 4617 7361 4629 7364
rect 4663 7361 4675 7395
rect 5258 7392 5264 7404
rect 4617 7355 4675 7361
rect 5256 7352 5264 7392
rect 5316 7352 5322 7404
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7392 5503 7395
rect 5491 7364 5948 7392
rect 5491 7361 5503 7364
rect 5445 7355 5503 7361
rect 1762 7324 1768 7336
rect 1723 7296 1768 7324
rect 1762 7284 1768 7296
rect 1820 7284 1826 7336
rect 3789 7327 3847 7333
rect 3789 7324 3801 7327
rect 2332 7296 3801 7324
rect 1026 7216 1032 7268
rect 1084 7256 1090 7268
rect 2332 7256 2360 7296
rect 3789 7293 3801 7296
rect 3835 7293 3847 7327
rect 3789 7287 3847 7293
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7324 4031 7327
rect 4433 7327 4491 7333
rect 4433 7324 4445 7327
rect 4019 7296 4445 7324
rect 4019 7293 4031 7296
rect 3973 7287 4031 7293
rect 4433 7293 4445 7296
rect 4479 7324 4491 7327
rect 5256 7324 5284 7352
rect 4479 7296 5284 7324
rect 5920 7324 5948 7364
rect 5994 7352 6000 7404
rect 6052 7392 6058 7404
rect 6181 7395 6239 7401
rect 6181 7392 6193 7395
rect 6052 7364 6193 7392
rect 6052 7352 6058 7364
rect 6181 7361 6193 7364
rect 6227 7361 6239 7395
rect 6181 7355 6239 7361
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7392 6423 7395
rect 6730 7392 6736 7404
rect 6411 7364 6736 7392
rect 6411 7361 6423 7364
rect 6365 7355 6423 7361
rect 6730 7352 6736 7364
rect 6788 7352 6794 7404
rect 8018 7352 8024 7404
rect 8076 7392 8082 7404
rect 9033 7395 9091 7401
rect 8076 7364 8984 7392
rect 8076 7352 8082 7364
rect 6638 7324 6644 7336
rect 5920 7296 6644 7324
rect 4479 7293 4491 7296
rect 4433 7287 4491 7293
rect 6638 7284 6644 7296
rect 6696 7284 6702 7336
rect 6825 7327 6883 7333
rect 6825 7293 6837 7327
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 7092 7327 7150 7333
rect 7092 7293 7104 7327
rect 7138 7324 7150 7327
rect 8202 7324 8208 7336
rect 7138 7296 8208 7324
rect 7138 7293 7150 7296
rect 7092 7287 7150 7293
rect 1084 7228 2360 7256
rect 1084 7216 1090 7228
rect 2406 7216 2412 7268
rect 2464 7256 2470 7268
rect 3234 7256 3240 7268
rect 2464 7228 3240 7256
rect 2464 7216 2470 7228
rect 3234 7216 3240 7228
rect 3292 7256 3298 7268
rect 4525 7259 4583 7265
rect 4525 7256 4537 7259
rect 3292 7228 4537 7256
rect 3292 7216 3298 7228
rect 4525 7225 4537 7228
rect 4571 7225 4583 7259
rect 5074 7256 5080 7268
rect 4525 7219 4583 7225
rect 4623 7228 5080 7256
rect 1302 7148 1308 7200
rect 1360 7188 1366 7200
rect 1397 7191 1455 7197
rect 1397 7188 1409 7191
rect 1360 7160 1409 7188
rect 1360 7148 1366 7160
rect 1397 7157 1409 7160
rect 1443 7157 1455 7191
rect 1854 7188 1860 7200
rect 1815 7160 1860 7188
rect 1397 7151 1455 7157
rect 1854 7148 1860 7160
rect 1912 7148 1918 7200
rect 2038 7148 2044 7200
rect 2096 7188 2102 7200
rect 2593 7191 2651 7197
rect 2593 7188 2605 7191
rect 2096 7160 2605 7188
rect 2096 7148 2102 7160
rect 2593 7157 2605 7160
rect 2639 7157 2651 7191
rect 2593 7151 2651 7157
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 3602 7188 3608 7200
rect 2832 7160 3608 7188
rect 2832 7148 2838 7160
rect 3602 7148 3608 7160
rect 3660 7148 3666 7200
rect 3789 7191 3847 7197
rect 3789 7157 3801 7191
rect 3835 7188 3847 7191
rect 4623 7188 4651 7228
rect 5074 7216 5080 7228
rect 5132 7256 5138 7268
rect 5261 7259 5319 7265
rect 5261 7256 5273 7259
rect 5132 7228 5273 7256
rect 5132 7216 5138 7228
rect 5261 7225 5273 7228
rect 5307 7225 5319 7259
rect 5261 7219 5319 7225
rect 5353 7259 5411 7265
rect 5353 7225 5365 7259
rect 5399 7256 5411 7259
rect 5718 7256 5724 7268
rect 5399 7228 5724 7256
rect 5399 7225 5411 7228
rect 5353 7219 5411 7225
rect 5718 7216 5724 7228
rect 5776 7216 5782 7268
rect 6086 7256 6092 7268
rect 6047 7228 6092 7256
rect 6086 7216 6092 7228
rect 6144 7216 6150 7268
rect 6840 7256 6868 7287
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 7558 7256 7564 7268
rect 6840 7228 7564 7256
rect 7558 7216 7564 7228
rect 7616 7256 7622 7268
rect 7926 7256 7932 7268
rect 7616 7228 7932 7256
rect 7616 7216 7622 7228
rect 7926 7216 7932 7228
rect 7984 7216 7990 7268
rect 8110 7216 8116 7268
rect 8168 7256 8174 7268
rect 8294 7256 8300 7268
rect 8168 7228 8300 7256
rect 8168 7216 8174 7228
rect 8294 7216 8300 7228
rect 8352 7216 8358 7268
rect 8846 7216 8852 7268
rect 8904 7256 8910 7268
rect 8956 7256 8984 7364
rect 9033 7361 9045 7395
rect 9079 7392 9091 7395
rect 10045 7395 10103 7401
rect 10045 7392 10057 7395
rect 9079 7364 10057 7392
rect 9079 7361 9091 7364
rect 9033 7355 9091 7361
rect 10045 7361 10057 7364
rect 10091 7361 10103 7395
rect 10045 7355 10103 7361
rect 11422 7352 11428 7404
rect 11480 7392 11486 7404
rect 15657 7395 15715 7401
rect 11480 7364 12572 7392
rect 11480 7352 11486 7364
rect 9674 7284 9680 7336
rect 9732 7324 9738 7336
rect 10410 7333 10416 7336
rect 10137 7327 10195 7333
rect 10137 7324 10149 7327
rect 9732 7296 10149 7324
rect 9732 7284 9738 7296
rect 10137 7293 10149 7296
rect 10183 7293 10195 7327
rect 10404 7324 10416 7333
rect 10371 7296 10416 7324
rect 10137 7287 10195 7293
rect 10404 7287 10416 7296
rect 10468 7324 10474 7336
rect 11330 7324 11336 7336
rect 10468 7296 11336 7324
rect 10410 7284 10416 7287
rect 10468 7284 10474 7296
rect 11330 7284 11336 7296
rect 11388 7284 11394 7336
rect 12434 7324 12440 7336
rect 12395 7296 12440 7324
rect 12434 7284 12440 7296
rect 12492 7284 12498 7336
rect 12544 7324 12572 7364
rect 15657 7361 15669 7395
rect 15703 7392 15715 7395
rect 16114 7392 16120 7404
rect 15703 7364 16120 7392
rect 15703 7361 15715 7364
rect 15657 7355 15715 7361
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 13722 7324 13728 7336
rect 12544 7296 13728 7324
rect 13722 7284 13728 7296
rect 13780 7284 13786 7336
rect 15378 7324 15384 7336
rect 15339 7296 15384 7324
rect 15378 7284 15384 7296
rect 15436 7284 15442 7336
rect 16592 7333 16620 7432
rect 18690 7420 18696 7472
rect 18748 7460 18754 7472
rect 19613 7463 19671 7469
rect 19613 7460 19625 7463
rect 18748 7432 19625 7460
rect 18748 7420 18754 7432
rect 19613 7429 19625 7432
rect 19659 7429 19671 7463
rect 19613 7423 19671 7429
rect 18598 7392 18604 7404
rect 18559 7364 18604 7392
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 20088 7401 20116 7500
rect 20073 7395 20131 7401
rect 20073 7361 20085 7395
rect 20119 7361 20131 7395
rect 20073 7355 20131 7361
rect 20165 7395 20223 7401
rect 20165 7361 20177 7395
rect 20211 7361 20223 7395
rect 20165 7355 20223 7361
rect 16577 7327 16635 7333
rect 16577 7293 16589 7327
rect 16623 7293 16635 7327
rect 16577 7287 16635 7293
rect 18138 7284 18144 7336
rect 18196 7324 18202 7336
rect 18325 7327 18383 7333
rect 18325 7324 18337 7327
rect 18196 7296 18337 7324
rect 18196 7284 18202 7296
rect 18325 7293 18337 7296
rect 18371 7293 18383 7327
rect 19978 7324 19984 7336
rect 19939 7296 19984 7324
rect 18325 7287 18383 7293
rect 19978 7284 19984 7296
rect 20036 7284 20042 7336
rect 20180 7324 20208 7355
rect 20088 7296 20208 7324
rect 11974 7256 11980 7268
rect 8904 7228 11980 7256
rect 8904 7216 8910 7228
rect 11974 7216 11980 7228
rect 12032 7216 12038 7268
rect 12158 7216 12164 7268
rect 12216 7256 12222 7268
rect 12682 7259 12740 7265
rect 12682 7256 12694 7259
rect 12216 7228 12694 7256
rect 12216 7216 12222 7228
rect 12682 7225 12694 7228
rect 12728 7225 12740 7259
rect 12682 7219 12740 7225
rect 12894 7216 12900 7268
rect 12952 7256 12958 7268
rect 12952 7228 15608 7256
rect 12952 7216 12958 7228
rect 3835 7160 4651 7188
rect 4893 7191 4951 7197
rect 3835 7157 3847 7160
rect 3789 7151 3847 7157
rect 4893 7157 4905 7191
rect 4939 7188 4951 7191
rect 9030 7188 9036 7200
rect 4939 7160 9036 7188
rect 4939 7157 4951 7160
rect 4893 7151 4951 7157
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 9674 7148 9680 7200
rect 9732 7188 9738 7200
rect 9858 7188 9864 7200
rect 9732 7160 9864 7188
rect 9732 7148 9738 7160
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 10045 7191 10103 7197
rect 10045 7157 10057 7191
rect 10091 7188 10103 7191
rect 12802 7188 12808 7200
rect 10091 7160 12808 7188
rect 10091 7157 10103 7160
rect 10045 7151 10103 7157
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 13078 7148 13084 7200
rect 13136 7188 13142 7200
rect 13817 7191 13875 7197
rect 13817 7188 13829 7191
rect 13136 7160 13829 7188
rect 13136 7148 13142 7160
rect 13817 7157 13829 7160
rect 13863 7157 13875 7191
rect 15470 7188 15476 7200
rect 15431 7160 15476 7188
rect 13817 7151 13875 7157
rect 15470 7148 15476 7160
rect 15528 7148 15534 7200
rect 15580 7188 15608 7228
rect 16666 7216 16672 7268
rect 16724 7256 16730 7268
rect 16853 7259 16911 7265
rect 16853 7256 16865 7259
rect 16724 7228 16865 7256
rect 16724 7216 16730 7228
rect 16853 7225 16865 7228
rect 16899 7225 16911 7259
rect 16853 7219 16911 7225
rect 17586 7216 17592 7268
rect 17644 7256 17650 7268
rect 20088 7256 20116 7296
rect 17644 7228 20116 7256
rect 17644 7216 17650 7228
rect 17126 7188 17132 7200
rect 15580 7160 17132 7188
rect 17126 7148 17132 7160
rect 17184 7148 17190 7200
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 1302 6944 1308 6996
rect 1360 6984 1366 6996
rect 3329 6987 3387 6993
rect 3329 6984 3341 6987
rect 1360 6956 3341 6984
rect 1360 6944 1366 6956
rect 3329 6953 3341 6956
rect 3375 6953 3387 6987
rect 3602 6984 3608 6996
rect 3329 6947 3387 6953
rect 3436 6956 3608 6984
rect 3237 6919 3295 6925
rect 3237 6885 3249 6919
rect 3283 6916 3295 6919
rect 3436 6916 3464 6956
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 4433 6987 4491 6993
rect 4433 6953 4445 6987
rect 4479 6984 4491 6987
rect 4982 6984 4988 6996
rect 4479 6956 4988 6984
rect 4479 6953 4491 6956
rect 4433 6947 4491 6953
rect 4982 6944 4988 6956
rect 5040 6944 5046 6996
rect 5258 6984 5264 6996
rect 5219 6956 5264 6984
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 5353 6987 5411 6993
rect 5353 6953 5365 6987
rect 5399 6984 5411 6987
rect 5626 6984 5632 6996
rect 5399 6956 5632 6984
rect 5399 6953 5411 6956
rect 5353 6947 5411 6953
rect 5626 6944 5632 6956
rect 5684 6944 5690 6996
rect 5721 6987 5779 6993
rect 5721 6953 5733 6987
rect 5767 6953 5779 6987
rect 5721 6947 5779 6953
rect 6089 6987 6147 6993
rect 6089 6953 6101 6987
rect 6135 6984 6147 6987
rect 6270 6984 6276 6996
rect 6135 6956 6276 6984
rect 6135 6953 6147 6956
rect 6089 6947 6147 6953
rect 3283 6888 3464 6916
rect 3283 6885 3295 6888
rect 3237 6879 3295 6885
rect 4798 6876 4804 6928
rect 4856 6916 4862 6928
rect 5736 6916 5764 6947
rect 6270 6944 6276 6956
rect 6328 6944 6334 6996
rect 6362 6944 6368 6996
rect 6420 6984 6426 6996
rect 11422 6984 11428 6996
rect 6420 6956 11428 6984
rect 6420 6944 6426 6956
rect 11422 6944 11428 6956
rect 11480 6944 11486 6996
rect 11514 6944 11520 6996
rect 11572 6984 11578 6996
rect 12069 6987 12127 6993
rect 12069 6984 12081 6987
rect 11572 6956 12081 6984
rect 11572 6944 11578 6956
rect 12069 6953 12081 6956
rect 12115 6953 12127 6987
rect 12069 6947 12127 6953
rect 4856 6888 5764 6916
rect 5828 6888 6316 6916
rect 4856 6876 4862 6888
rect 1664 6851 1722 6857
rect 1664 6817 1676 6851
rect 1710 6848 1722 6851
rect 2958 6848 2964 6860
rect 1710 6820 2964 6848
rect 1710 6817 1722 6820
rect 1664 6811 1722 6817
rect 2958 6808 2964 6820
rect 3016 6848 3022 6860
rect 3326 6848 3332 6860
rect 3016 6820 3332 6848
rect 3016 6808 3022 6820
rect 3326 6808 3332 6820
rect 3384 6808 3390 6860
rect 5828 6848 5856 6888
rect 3436 6820 5856 6848
rect 6181 6851 6239 6857
rect 1302 6740 1308 6792
rect 1360 6780 1366 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 1360 6752 1409 6780
rect 1360 6740 1366 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 3436 6780 3464 6820
rect 6181 6817 6193 6851
rect 6227 6817 6239 6851
rect 6181 6811 6239 6817
rect 2832 6752 3464 6780
rect 3513 6783 3571 6789
rect 2832 6740 2838 6752
rect 3513 6749 3525 6783
rect 3559 6780 3571 6783
rect 3694 6780 3700 6792
rect 3559 6752 3700 6780
rect 3559 6749 3571 6752
rect 3513 6743 3571 6749
rect 3694 6740 3700 6752
rect 3752 6740 3758 6792
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6780 4767 6783
rect 4982 6780 4988 6792
rect 4755 6752 4988 6780
rect 4755 6749 4767 6752
rect 4709 6743 4767 6749
rect 4540 6712 4568 6743
rect 2608 6684 4568 6712
rect 1210 6604 1216 6656
rect 1268 6644 1274 6656
rect 2608 6644 2636 6684
rect 2774 6644 2780 6656
rect 1268 6616 2636 6644
rect 2735 6616 2780 6644
rect 1268 6604 1274 6616
rect 2774 6604 2780 6616
rect 2832 6604 2838 6656
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 3234 6644 3240 6656
rect 2915 6616 3240 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 4062 6644 4068 6656
rect 4023 6616 4068 6644
rect 4062 6604 4068 6616
rect 4120 6604 4126 6656
rect 4154 6604 4160 6656
rect 4212 6644 4218 6656
rect 4724 6644 4752 6743
rect 4982 6740 4988 6752
rect 5040 6740 5046 6792
rect 5350 6740 5356 6792
rect 5408 6780 5414 6792
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 5408 6752 5457 6780
rect 5408 6740 5414 6752
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 6196 6780 6224 6811
rect 6288 6789 6316 6888
rect 6638 6876 6644 6928
rect 6696 6916 6702 6928
rect 7190 6916 7196 6928
rect 6696 6888 7196 6916
rect 6696 6876 6702 6888
rect 7190 6876 7196 6888
rect 7248 6876 7254 6928
rect 7466 6876 7472 6928
rect 7524 6916 7530 6928
rect 7653 6919 7711 6925
rect 7653 6916 7665 6919
rect 7524 6888 7665 6916
rect 7524 6876 7530 6888
rect 7653 6885 7665 6888
rect 7699 6885 7711 6919
rect 7653 6879 7711 6885
rect 7745 6919 7803 6925
rect 7745 6885 7757 6919
rect 7791 6916 7803 6919
rect 7926 6916 7932 6928
rect 7791 6888 7932 6916
rect 7791 6885 7803 6888
rect 7745 6879 7803 6885
rect 7926 6876 7932 6888
rect 7984 6876 7990 6928
rect 11698 6916 11704 6928
rect 8036 6888 11704 6916
rect 8036 6848 8064 6888
rect 11698 6876 11704 6888
rect 11756 6876 11762 6928
rect 11977 6919 12035 6925
rect 11977 6916 11989 6919
rect 11900 6888 11989 6916
rect 10410 6848 10416 6860
rect 6380 6820 8064 6848
rect 10371 6820 10416 6848
rect 6380 6792 6408 6820
rect 10410 6808 10416 6820
rect 10468 6808 10474 6860
rect 10962 6808 10968 6860
rect 11020 6848 11026 6860
rect 11900 6848 11928 6888
rect 11977 6885 11989 6888
rect 12023 6885 12035 6919
rect 11977 6879 12035 6885
rect 16114 6876 16120 6928
rect 16172 6916 16178 6928
rect 16454 6919 16512 6925
rect 16454 6916 16466 6919
rect 16172 6888 16466 6916
rect 16172 6876 16178 6888
rect 16454 6885 16466 6888
rect 16500 6885 16512 6919
rect 16454 6879 16512 6885
rect 11020 6820 11928 6848
rect 12176 6820 12480 6848
rect 11020 6808 11026 6820
rect 5445 6743 5503 6749
rect 5552 6752 6224 6780
rect 6273 6783 6331 6789
rect 4893 6715 4951 6721
rect 4893 6681 4905 6715
rect 4939 6712 4951 6715
rect 5552 6712 5580 6752
rect 6273 6749 6285 6783
rect 6319 6749 6331 6783
rect 6273 6743 6331 6749
rect 6362 6740 6368 6792
rect 6420 6740 6426 6792
rect 6546 6780 6552 6792
rect 6507 6752 6552 6780
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 7742 6740 7748 6792
rect 7800 6780 7806 6792
rect 7837 6783 7895 6789
rect 7837 6780 7849 6783
rect 7800 6752 7849 6780
rect 7800 6740 7806 6752
rect 7837 6749 7849 6752
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 9122 6740 9128 6792
rect 9180 6780 9186 6792
rect 9858 6780 9864 6792
rect 9180 6752 9864 6780
rect 9180 6740 9186 6752
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 10502 6780 10508 6792
rect 10463 6752 10508 6780
rect 10502 6740 10508 6752
rect 10560 6740 10566 6792
rect 10689 6783 10747 6789
rect 10689 6749 10701 6783
rect 10735 6780 10747 6783
rect 11330 6780 11336 6792
rect 10735 6752 11336 6780
rect 10735 6749 10747 6752
rect 10689 6743 10747 6749
rect 11330 6740 11336 6752
rect 11388 6740 11394 6792
rect 11698 6740 11704 6792
rect 11756 6780 11762 6792
rect 12176 6780 12204 6820
rect 11756 6752 12204 6780
rect 12253 6783 12311 6789
rect 11756 6740 11762 6752
rect 12253 6749 12265 6783
rect 12299 6749 12311 6783
rect 12452 6780 12480 6820
rect 12526 6808 12532 6860
rect 12584 6848 12590 6860
rect 14001 6851 14059 6857
rect 14001 6848 14013 6851
rect 12584 6820 14013 6848
rect 12584 6808 12590 6820
rect 14001 6817 14013 6820
rect 14047 6817 14059 6851
rect 14001 6811 14059 6817
rect 14093 6851 14151 6857
rect 14093 6817 14105 6851
rect 14139 6848 14151 6851
rect 14734 6848 14740 6860
rect 14139 6820 14740 6848
rect 14139 6817 14151 6820
rect 14093 6811 14151 6817
rect 14734 6808 14740 6820
rect 14792 6808 14798 6860
rect 15838 6808 15844 6860
rect 15896 6848 15902 6860
rect 16206 6848 16212 6860
rect 15896 6820 16212 6848
rect 15896 6808 15902 6820
rect 16206 6808 16212 6820
rect 16264 6848 16270 6860
rect 16264 6820 17264 6848
rect 16264 6808 16270 6820
rect 14185 6783 14243 6789
rect 14185 6780 14197 6783
rect 12452 6752 14197 6780
rect 12253 6743 12311 6749
rect 14185 6749 14197 6752
rect 14231 6780 14243 6783
rect 14274 6780 14280 6792
rect 14231 6752 14280 6780
rect 14231 6749 14243 6752
rect 14185 6743 14243 6749
rect 4939 6684 5580 6712
rect 4939 6681 4951 6684
rect 4893 6675 4951 6681
rect 6178 6672 6184 6724
rect 6236 6712 6242 6724
rect 10045 6715 10103 6721
rect 6236 6684 9895 6712
rect 6236 6672 6242 6684
rect 9867 6656 9895 6684
rect 10045 6681 10057 6715
rect 10091 6712 10103 6715
rect 11514 6712 11520 6724
rect 10091 6684 11520 6712
rect 10091 6681 10103 6684
rect 10045 6675 10103 6681
rect 11514 6672 11520 6684
rect 11572 6672 11578 6724
rect 12158 6672 12164 6724
rect 12216 6712 12222 6724
rect 12268 6712 12296 6743
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 17236 6780 17264 6820
rect 17862 6808 17868 6860
rect 17920 6848 17926 6860
rect 18673 6851 18731 6857
rect 18673 6848 18685 6851
rect 17920 6820 18685 6848
rect 17920 6808 17926 6820
rect 18673 6817 18685 6820
rect 18719 6817 18731 6851
rect 18673 6811 18731 6817
rect 18417 6783 18475 6789
rect 18417 6780 18429 6783
rect 17236 6752 18429 6780
rect 17880 6724 17908 6752
rect 18417 6749 18429 6752
rect 18463 6749 18475 6783
rect 18417 6743 18475 6749
rect 12216 6684 12296 6712
rect 12216 6672 12222 6684
rect 17862 6672 17868 6724
rect 17920 6672 17926 6724
rect 4212 6616 4752 6644
rect 4212 6604 4218 6616
rect 4798 6604 4804 6656
rect 4856 6644 4862 6656
rect 5350 6644 5356 6656
rect 4856 6616 5356 6644
rect 4856 6604 4862 6616
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 5810 6604 5816 6656
rect 5868 6644 5874 6656
rect 7006 6644 7012 6656
rect 5868 6616 7012 6644
rect 5868 6604 5874 6616
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 7285 6647 7343 6653
rect 7285 6613 7297 6647
rect 7331 6644 7343 6647
rect 7650 6644 7656 6656
rect 7331 6616 7656 6644
rect 7331 6613 7343 6616
rect 7285 6607 7343 6613
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 9849 6604 9855 6656
rect 9907 6604 9913 6656
rect 11054 6604 11060 6656
rect 11112 6644 11118 6656
rect 11609 6647 11667 6653
rect 11609 6644 11621 6647
rect 11112 6616 11621 6644
rect 11112 6604 11118 6616
rect 11609 6613 11621 6616
rect 11655 6613 11667 6647
rect 11609 6607 11667 6613
rect 13633 6647 13691 6653
rect 13633 6613 13645 6647
rect 13679 6644 13691 6647
rect 15010 6644 15016 6656
rect 13679 6616 15016 6644
rect 13679 6613 13691 6616
rect 13633 6607 13691 6613
rect 15010 6604 15016 6616
rect 15068 6604 15074 6656
rect 17586 6644 17592 6656
rect 17547 6616 17592 6644
rect 17586 6604 17592 6616
rect 17644 6604 17650 6656
rect 18046 6604 18052 6656
rect 18104 6644 18110 6656
rect 19797 6647 19855 6653
rect 19797 6644 19809 6647
rect 18104 6616 19809 6644
rect 18104 6604 18110 6616
rect 19797 6613 19809 6616
rect 19843 6613 19855 6647
rect 19797 6607 19855 6613
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 1302 6400 1308 6452
rect 1360 6440 1366 6452
rect 1949 6443 2007 6449
rect 1949 6440 1961 6443
rect 1360 6412 1961 6440
rect 1360 6400 1366 6412
rect 1949 6409 1961 6412
rect 1995 6440 2007 6443
rect 1995 6412 3004 6440
rect 1995 6409 2007 6412
rect 1949 6403 2007 6409
rect 2976 6372 3004 6412
rect 3326 6400 3332 6452
rect 3384 6440 3390 6452
rect 3421 6443 3479 6449
rect 3421 6440 3433 6443
rect 3384 6412 3433 6440
rect 3384 6400 3390 6412
rect 3421 6409 3433 6412
rect 3467 6440 3479 6443
rect 4798 6440 4804 6452
rect 3467 6412 4804 6440
rect 3467 6409 3479 6412
rect 3421 6403 3479 6409
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 5166 6400 5172 6452
rect 5224 6440 5230 6452
rect 5905 6443 5963 6449
rect 5905 6440 5917 6443
rect 5224 6412 5917 6440
rect 5224 6400 5230 6412
rect 5905 6409 5917 6412
rect 5951 6409 5963 6443
rect 5905 6403 5963 6409
rect 6181 6443 6239 6449
rect 6181 6409 6193 6443
rect 6227 6440 6239 6443
rect 6270 6440 6276 6452
rect 6227 6412 6276 6440
rect 6227 6409 6239 6412
rect 6181 6403 6239 6409
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 6454 6400 6460 6452
rect 6512 6440 6518 6452
rect 6549 6443 6607 6449
rect 6549 6440 6561 6443
rect 6512 6412 6561 6440
rect 6512 6400 6518 6412
rect 6549 6409 6561 6412
rect 6595 6409 6607 6443
rect 7558 6440 7564 6452
rect 6549 6403 6607 6409
rect 6932 6412 7564 6440
rect 2976 6344 4568 6372
rect 4540 6316 4568 6344
rect 5534 6332 5540 6384
rect 5592 6372 5598 6384
rect 5592 6344 6408 6372
rect 5592 6332 5598 6344
rect 1412 6276 2176 6304
rect 1412 6245 1440 6276
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6205 1455 6239
rect 1946 6236 1952 6248
rect 1859 6208 1952 6236
rect 1397 6199 1455 6205
rect 1946 6196 1952 6208
rect 2004 6236 2010 6248
rect 2041 6239 2099 6245
rect 2041 6236 2053 6239
rect 2004 6208 2053 6236
rect 2004 6196 2010 6208
rect 2041 6205 2053 6208
rect 2087 6205 2099 6239
rect 2148 6236 2176 6276
rect 3694 6264 3700 6316
rect 3752 6304 3758 6316
rect 4157 6307 4215 6313
rect 4157 6304 4169 6307
rect 3752 6276 4169 6304
rect 3752 6264 3758 6276
rect 4157 6273 4169 6276
rect 4203 6304 4215 6307
rect 4203 6276 4476 6304
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 4338 6236 4344 6248
rect 2148 6208 4344 6236
rect 2041 6199 2099 6205
rect 4338 6196 4344 6208
rect 4396 6196 4402 6248
rect 4448 6236 4476 6276
rect 4522 6264 4528 6316
rect 4580 6304 4586 6316
rect 6270 6304 6276 6316
rect 4580 6276 4625 6304
rect 5644 6276 6276 6304
rect 4580 6264 4586 6276
rect 5644 6236 5672 6276
rect 6270 6264 6276 6276
rect 6328 6264 6334 6316
rect 6380 6245 6408 6344
rect 6932 6313 6960 6412
rect 7558 6400 7564 6412
rect 7616 6400 7622 6452
rect 8202 6400 8208 6452
rect 8260 6440 8266 6452
rect 8297 6443 8355 6449
rect 8297 6440 8309 6443
rect 8260 6412 8309 6440
rect 8260 6400 8266 6412
rect 8297 6409 8309 6412
rect 8343 6409 8355 6443
rect 8297 6403 8355 6409
rect 8386 6400 8392 6452
rect 8444 6440 8450 6452
rect 9401 6443 9459 6449
rect 8444 6412 8489 6440
rect 8444 6400 8450 6412
rect 9401 6409 9413 6443
rect 9447 6440 9459 6443
rect 10137 6443 10195 6449
rect 9447 6412 10088 6440
rect 9447 6409 9459 6412
rect 9401 6403 9459 6409
rect 9766 6372 9772 6384
rect 8956 6344 9772 6372
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6273 6975 6307
rect 8846 6304 8852 6316
rect 8807 6276 8852 6304
rect 6917 6267 6975 6273
rect 8846 6264 8852 6276
rect 8904 6264 8910 6316
rect 4448 6208 5672 6236
rect 5997 6239 6055 6245
rect 5997 6205 6009 6239
rect 6043 6236 6055 6239
rect 6365 6239 6423 6245
rect 6043 6208 6316 6236
rect 6043 6205 6055 6208
rect 5997 6199 6055 6205
rect 1673 6171 1731 6177
rect 1673 6137 1685 6171
rect 1719 6168 1731 6171
rect 2130 6168 2136 6180
rect 1719 6140 2136 6168
rect 1719 6137 1731 6140
rect 1673 6131 1731 6137
rect 2130 6128 2136 6140
rect 2188 6128 2194 6180
rect 2308 6171 2366 6177
rect 2308 6137 2320 6171
rect 2354 6168 2366 6171
rect 2682 6168 2688 6180
rect 2354 6140 2688 6168
rect 2354 6137 2366 6140
rect 2308 6131 2366 6137
rect 2682 6128 2688 6140
rect 2740 6128 2746 6180
rect 3973 6171 4031 6177
rect 3973 6137 3985 6171
rect 4019 6168 4031 6171
rect 4614 6168 4620 6180
rect 4019 6140 4620 6168
rect 4019 6137 4031 6140
rect 3973 6131 4031 6137
rect 4614 6128 4620 6140
rect 4672 6128 4678 6180
rect 4792 6171 4850 6177
rect 4792 6137 4804 6171
rect 4838 6168 4850 6171
rect 5350 6168 5356 6180
rect 4838 6140 5356 6168
rect 4838 6137 4850 6140
rect 4792 6131 4850 6137
rect 5350 6128 5356 6140
rect 5408 6128 5414 6180
rect 6288 6168 6316 6208
rect 6365 6205 6377 6239
rect 6411 6236 6423 6239
rect 6638 6236 6644 6248
rect 6411 6208 6644 6236
rect 6411 6205 6423 6208
rect 6365 6199 6423 6205
rect 6638 6196 6644 6208
rect 6696 6196 6702 6248
rect 8757 6239 8815 6245
rect 7107 6208 8524 6236
rect 7107 6168 7135 6208
rect 6288 6140 7135 6168
rect 7184 6171 7242 6177
rect 7184 6137 7196 6171
rect 7230 6168 7242 6171
rect 8386 6168 8392 6180
rect 7230 6140 8392 6168
rect 7230 6137 7242 6140
rect 7184 6131 7242 6137
rect 8386 6128 8392 6140
rect 8444 6128 8450 6180
rect 8496 6168 8524 6208
rect 8757 6205 8769 6239
rect 8803 6236 8815 6239
rect 8956 6236 8984 6344
rect 9766 6332 9772 6344
rect 9824 6332 9830 6384
rect 10060 6372 10088 6412
rect 10137 6409 10149 6443
rect 10183 6440 10195 6443
rect 10183 6412 11652 6440
rect 10183 6409 10195 6412
rect 10137 6403 10195 6409
rect 11624 6384 11652 6412
rect 12342 6400 12348 6452
rect 12400 6440 12406 6452
rect 14645 6443 14703 6449
rect 12400 6412 13400 6440
rect 12400 6400 12406 6412
rect 10229 6375 10287 6381
rect 10060 6344 10180 6372
rect 9033 6307 9091 6313
rect 9033 6273 9045 6307
rect 9079 6304 9091 6307
rect 9122 6304 9128 6316
rect 9079 6276 9128 6304
rect 9079 6273 9091 6276
rect 9033 6267 9091 6273
rect 9122 6264 9128 6276
rect 9180 6264 9186 6316
rect 9674 6304 9680 6316
rect 9232 6276 9680 6304
rect 9232 6245 9260 6276
rect 9674 6264 9680 6276
rect 9732 6264 9738 6316
rect 10152 6304 10180 6344
rect 10229 6341 10241 6375
rect 10275 6372 10287 6375
rect 10410 6372 10416 6384
rect 10275 6344 10416 6372
rect 10275 6341 10287 6344
rect 10229 6335 10287 6341
rect 10410 6332 10416 6344
rect 10468 6332 10474 6384
rect 10796 6344 11560 6372
rect 10796 6304 10824 6344
rect 10152 6276 10824 6304
rect 10873 6307 10931 6313
rect 10873 6273 10885 6307
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 8803 6208 8984 6236
rect 9217 6239 9275 6245
rect 8803 6205 8815 6208
rect 8757 6199 8815 6205
rect 9217 6205 9229 6239
rect 9263 6205 9275 6239
rect 9217 6199 9275 6205
rect 9766 6196 9772 6248
rect 9824 6236 9830 6248
rect 9824 6208 10272 6236
rect 9824 6196 9830 6208
rect 9674 6168 9680 6180
rect 8496 6140 9680 6168
rect 9674 6128 9680 6140
rect 9732 6128 9738 6180
rect 3513 6103 3571 6109
rect 3513 6069 3525 6103
rect 3559 6100 3571 6103
rect 3786 6100 3792 6112
rect 3559 6072 3792 6100
rect 3559 6069 3571 6072
rect 3513 6063 3571 6069
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 3881 6103 3939 6109
rect 3881 6069 3893 6103
rect 3927 6100 3939 6103
rect 6178 6100 6184 6112
rect 3927 6072 6184 6100
rect 3927 6069 3939 6072
rect 3881 6063 3939 6069
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 6270 6060 6276 6112
rect 6328 6100 6334 6112
rect 10137 6103 10195 6109
rect 10137 6100 10149 6103
rect 6328 6072 10149 6100
rect 6328 6060 6334 6072
rect 10137 6069 10149 6072
rect 10183 6069 10195 6103
rect 10244 6100 10272 6208
rect 10594 6196 10600 6248
rect 10652 6196 10658 6248
rect 10689 6239 10747 6245
rect 10689 6205 10701 6239
rect 10735 6236 10747 6239
rect 10888 6236 10916 6267
rect 11146 6264 11152 6316
rect 11204 6304 11210 6316
rect 11422 6304 11428 6316
rect 11204 6276 11428 6304
rect 11204 6264 11210 6276
rect 11422 6264 11428 6276
rect 11480 6264 11486 6316
rect 11532 6304 11560 6344
rect 11606 6332 11612 6384
rect 11664 6332 11670 6384
rect 13372 6372 13400 6412
rect 14645 6409 14657 6443
rect 14691 6440 14703 6443
rect 15470 6440 15476 6452
rect 14691 6412 15476 6440
rect 14691 6409 14703 6412
rect 14645 6403 14703 6409
rect 15470 6400 15476 6412
rect 15528 6400 15534 6452
rect 16114 6400 16120 6452
rect 16172 6440 16178 6452
rect 17494 6440 17500 6452
rect 16172 6412 17500 6440
rect 16172 6400 16178 6412
rect 17494 6400 17500 6412
rect 17552 6400 17558 6452
rect 19610 6440 19616 6452
rect 19571 6412 19616 6440
rect 19610 6400 19616 6412
rect 19668 6400 19674 6452
rect 13372 6344 16620 6372
rect 12158 6304 12164 6316
rect 11532 6276 12164 6304
rect 12158 6264 12164 6276
rect 12216 6264 12222 6316
rect 12434 6304 12440 6316
rect 12395 6276 12440 6304
rect 12434 6264 12440 6276
rect 12492 6264 12498 6316
rect 15289 6307 15347 6313
rect 15289 6273 15301 6307
rect 15335 6304 15347 6307
rect 15562 6304 15568 6316
rect 15335 6276 15568 6304
rect 15335 6273 15347 6276
rect 15289 6267 15347 6273
rect 15562 6264 15568 6276
rect 15620 6264 15626 6316
rect 11330 6236 11336 6248
rect 10735 6208 10824 6236
rect 10888 6208 11336 6236
rect 10735 6205 10747 6208
rect 10689 6199 10747 6205
rect 10612 6168 10640 6196
rect 10796 6168 10824 6208
rect 11330 6196 11336 6208
rect 11388 6196 11394 6248
rect 12704 6239 12762 6245
rect 12704 6205 12716 6239
rect 12750 6236 12762 6239
rect 13078 6236 13084 6248
rect 12750 6208 13084 6236
rect 12750 6205 12762 6208
rect 12704 6199 12762 6205
rect 12526 6168 12532 6180
rect 10612 6140 10732 6168
rect 10796 6140 12532 6168
rect 10597 6103 10655 6109
rect 10597 6100 10609 6103
rect 10244 6072 10609 6100
rect 10137 6063 10195 6069
rect 10597 6069 10609 6072
rect 10643 6069 10655 6103
rect 10704 6100 10732 6140
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 12618 6128 12624 6180
rect 12676 6168 12682 6180
rect 12719 6168 12747 6199
rect 13078 6196 13084 6208
rect 13136 6196 13142 6248
rect 13446 6196 13452 6248
rect 13504 6236 13510 6248
rect 13906 6236 13912 6248
rect 13504 6208 13912 6236
rect 13504 6196 13510 6208
rect 13906 6196 13912 6208
rect 13964 6196 13970 6248
rect 15010 6236 15016 6248
rect 14971 6208 15016 6236
rect 15010 6196 15016 6208
rect 15068 6196 15074 6248
rect 16592 6245 16620 6344
rect 16853 6307 16911 6313
rect 16853 6273 16865 6307
rect 16899 6304 16911 6307
rect 17034 6304 17040 6316
rect 16899 6276 17040 6304
rect 16899 6273 16911 6276
rect 16853 6267 16911 6273
rect 17034 6264 17040 6276
rect 17092 6264 17098 6316
rect 18046 6264 18052 6316
rect 18104 6304 18110 6316
rect 18601 6307 18659 6313
rect 18601 6304 18613 6307
rect 18104 6276 18613 6304
rect 18104 6264 18110 6276
rect 18601 6273 18613 6276
rect 18647 6273 18659 6307
rect 18601 6267 18659 6273
rect 20165 6307 20223 6313
rect 20165 6273 20177 6307
rect 20211 6273 20223 6307
rect 20165 6267 20223 6273
rect 16577 6239 16635 6245
rect 16577 6205 16589 6239
rect 16623 6205 16635 6239
rect 16577 6199 16635 6205
rect 16669 6239 16727 6245
rect 16669 6205 16681 6239
rect 16715 6236 16727 6239
rect 16942 6236 16948 6248
rect 16715 6208 16948 6236
rect 16715 6205 16727 6208
rect 16669 6199 16727 6205
rect 16942 6196 16948 6208
rect 17000 6236 17006 6248
rect 17770 6236 17776 6248
rect 17000 6208 17776 6236
rect 17000 6196 17006 6208
rect 17770 6196 17776 6208
rect 17828 6196 17834 6248
rect 17954 6196 17960 6248
rect 18012 6236 18018 6248
rect 18417 6239 18475 6245
rect 18417 6236 18429 6239
rect 18012 6208 18429 6236
rect 18012 6196 18018 6208
rect 18417 6205 18429 6208
rect 18463 6205 18475 6239
rect 18417 6199 18475 6205
rect 18506 6196 18512 6248
rect 18564 6236 18570 6248
rect 18564 6208 18609 6236
rect 18564 6196 18570 6208
rect 19886 6196 19892 6248
rect 19944 6236 19950 6248
rect 19981 6239 20039 6245
rect 19981 6236 19993 6239
rect 19944 6208 19993 6236
rect 19944 6196 19950 6208
rect 19981 6205 19993 6208
rect 20027 6205 20039 6239
rect 19981 6199 20039 6205
rect 12676 6140 12747 6168
rect 12676 6128 12682 6140
rect 12894 6128 12900 6180
rect 12952 6168 12958 6180
rect 20180 6168 20208 6267
rect 12952 6140 20208 6168
rect 12952 6128 12958 6140
rect 13722 6100 13728 6112
rect 10704 6072 13728 6100
rect 10597 6063 10655 6069
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 13817 6103 13875 6109
rect 13817 6069 13829 6103
rect 13863 6100 13875 6103
rect 13906 6100 13912 6112
rect 13863 6072 13912 6100
rect 13863 6069 13875 6072
rect 13817 6063 13875 6069
rect 13906 6060 13912 6072
rect 13964 6060 13970 6112
rect 15105 6103 15163 6109
rect 15105 6069 15117 6103
rect 15151 6100 15163 6103
rect 16209 6103 16267 6109
rect 16209 6100 16221 6103
rect 15151 6072 16221 6100
rect 15151 6069 15163 6072
rect 15105 6063 15163 6069
rect 16209 6069 16221 6072
rect 16255 6069 16267 6103
rect 18046 6100 18052 6112
rect 18007 6072 18052 6100
rect 16209 6063 16267 6069
rect 18046 6060 18052 6072
rect 18104 6060 18110 6112
rect 20070 6100 20076 6112
rect 20031 6072 20076 6100
rect 20070 6060 20076 6072
rect 20128 6060 20134 6112
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 2869 5899 2927 5905
rect 2869 5865 2881 5899
rect 2915 5896 2927 5899
rect 2958 5896 2964 5908
rect 2915 5868 2964 5896
rect 2915 5865 2927 5868
rect 2869 5859 2927 5865
rect 2958 5856 2964 5868
rect 3016 5856 3022 5908
rect 5350 5896 5356 5908
rect 3528 5868 5356 5896
rect 1670 5837 1676 5840
rect 1664 5828 1676 5837
rect 1631 5800 1676 5828
rect 1664 5791 1676 5800
rect 1670 5788 1676 5791
rect 1728 5788 1734 5840
rect 3234 5760 3240 5772
rect 3195 5732 3240 5760
rect 3234 5720 3240 5732
rect 3292 5720 3298 5772
rect 3326 5692 3332 5704
rect 3287 5664 3332 5692
rect 3326 5652 3332 5664
rect 3384 5652 3390 5704
rect 3528 5701 3556 5868
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 5721 5899 5779 5905
rect 5721 5896 5733 5899
rect 5592 5868 5733 5896
rect 5592 5856 5598 5868
rect 5721 5865 5733 5868
rect 5767 5865 5779 5899
rect 5721 5859 5779 5865
rect 6181 5899 6239 5905
rect 6181 5865 6193 5899
rect 6227 5896 6239 5899
rect 6822 5896 6828 5908
rect 6227 5868 6828 5896
rect 6227 5865 6239 5868
rect 6181 5859 6239 5865
rect 3786 5788 3792 5840
rect 3844 5828 3850 5840
rect 5074 5828 5080 5840
rect 3844 5800 5080 5828
rect 3844 5788 3850 5800
rect 5074 5788 5080 5800
rect 5132 5788 5138 5840
rect 5166 5788 5172 5840
rect 5224 5828 5230 5840
rect 6196 5828 6224 5859
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 7009 5899 7067 5905
rect 7009 5865 7021 5899
rect 7055 5896 7067 5899
rect 7098 5896 7104 5908
rect 7055 5868 7104 5896
rect 7055 5865 7067 5868
rect 7009 5859 7067 5865
rect 7098 5856 7104 5868
rect 7156 5856 7162 5908
rect 7469 5899 7527 5905
rect 7469 5865 7481 5899
rect 7515 5896 7527 5899
rect 7650 5896 7656 5908
rect 7515 5868 7656 5896
rect 7515 5865 7527 5868
rect 7469 5859 7527 5865
rect 7650 5856 7656 5868
rect 7708 5856 7714 5908
rect 7742 5856 7748 5908
rect 7800 5896 7806 5908
rect 8754 5896 8760 5908
rect 7800 5868 8760 5896
rect 7800 5856 7806 5868
rect 8754 5856 8760 5868
rect 8812 5856 8818 5908
rect 8941 5899 8999 5905
rect 8941 5865 8953 5899
rect 8987 5896 8999 5899
rect 9214 5896 9220 5908
rect 8987 5868 9220 5896
rect 8987 5865 8999 5868
rect 8941 5859 8999 5865
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 9674 5856 9680 5908
rect 9732 5896 9738 5908
rect 11146 5896 11152 5908
rect 9732 5868 11152 5896
rect 9732 5856 9738 5868
rect 11146 5856 11152 5868
rect 11204 5856 11210 5908
rect 12894 5896 12900 5908
rect 11256 5868 12900 5896
rect 7374 5828 7380 5840
rect 5224 5800 6224 5828
rect 6748 5800 7380 5828
rect 5224 5788 5230 5800
rect 4249 5763 4307 5769
rect 4249 5729 4261 5763
rect 4295 5760 4307 5763
rect 4338 5760 4344 5772
rect 4295 5732 4344 5760
rect 4295 5729 4307 5732
rect 4249 5723 4307 5729
rect 4338 5720 4344 5732
rect 4396 5720 4402 5772
rect 4516 5763 4574 5769
rect 4516 5729 4528 5763
rect 4562 5760 4574 5763
rect 4562 5732 5488 5760
rect 4562 5729 4574 5732
rect 4516 5723 4574 5729
rect 3513 5695 3571 5701
rect 3513 5661 3525 5695
rect 3559 5661 3571 5695
rect 5460 5692 5488 5732
rect 5534 5720 5540 5772
rect 5592 5760 5598 5772
rect 6089 5763 6147 5769
rect 6089 5760 6101 5763
rect 5592 5732 6101 5760
rect 5592 5720 5598 5732
rect 6089 5729 6101 5732
rect 6135 5729 6147 5763
rect 6748 5760 6776 5800
rect 7374 5788 7380 5800
rect 7432 5788 7438 5840
rect 9490 5828 9496 5840
rect 7760 5800 9496 5828
rect 6089 5723 6147 5729
rect 6196 5732 6776 5760
rect 5626 5692 5632 5704
rect 5460 5664 5632 5692
rect 3513 5655 3571 5661
rect 5626 5652 5632 5664
rect 5684 5652 5690 5704
rect 5810 5652 5816 5704
rect 5868 5692 5874 5704
rect 6196 5692 6224 5732
rect 6822 5720 6828 5772
rect 6880 5760 6886 5772
rect 6917 5763 6975 5769
rect 6917 5760 6929 5763
rect 6880 5732 6929 5760
rect 6880 5720 6886 5732
rect 6917 5729 6929 5732
rect 6963 5729 6975 5763
rect 7760 5760 7788 5800
rect 9490 5788 9496 5800
rect 9548 5788 9554 5840
rect 11256 5828 11284 5868
rect 12894 5856 12900 5868
rect 12952 5856 12958 5908
rect 13814 5856 13820 5908
rect 13872 5896 13878 5908
rect 13909 5899 13967 5905
rect 13909 5896 13921 5899
rect 13872 5868 13921 5896
rect 13872 5856 13878 5868
rect 13909 5865 13921 5868
rect 13955 5865 13967 5899
rect 13909 5859 13967 5865
rect 9600 5800 11284 5828
rect 6917 5723 6975 5729
rect 7024 5732 7788 5760
rect 7837 5763 7895 5769
rect 5868 5664 6224 5692
rect 6365 5695 6423 5701
rect 5868 5652 5874 5664
rect 6365 5661 6377 5695
rect 6411 5692 6423 5695
rect 7024 5692 7052 5732
rect 7837 5729 7849 5763
rect 7883 5760 7895 5763
rect 9600 5760 9628 5800
rect 11974 5788 11980 5840
rect 12032 5828 12038 5840
rect 12253 5831 12311 5837
rect 12253 5828 12265 5831
rect 12032 5800 12265 5828
rect 12032 5788 12038 5800
rect 12253 5797 12265 5800
rect 12299 5828 12311 5831
rect 12802 5828 12808 5840
rect 12299 5800 12808 5828
rect 12299 5797 12311 5800
rect 12253 5791 12311 5797
rect 12802 5788 12808 5800
rect 12860 5788 12866 5840
rect 20254 5828 20260 5840
rect 13832 5800 20260 5828
rect 7883 5732 8064 5760
rect 7883 5729 7895 5732
rect 7837 5723 7895 5729
rect 8036 5704 8064 5732
rect 8312 5732 9628 5760
rect 9944 5763 10002 5769
rect 7190 5692 7196 5704
rect 6411 5664 6500 5692
rect 6411 5661 6423 5664
rect 6365 5655 6423 5661
rect 2777 5627 2835 5633
rect 2777 5593 2789 5627
rect 2823 5624 2835 5627
rect 4154 5624 4160 5636
rect 2823 5596 4160 5624
rect 2823 5593 2835 5596
rect 2777 5587 2835 5593
rect 4154 5584 4160 5596
rect 4212 5584 4218 5636
rect 6472 5624 6500 5664
rect 6564 5664 7052 5692
rect 7103 5664 7196 5692
rect 6564 5633 6592 5664
rect 7190 5652 7196 5664
rect 7248 5692 7254 5704
rect 7374 5692 7380 5704
rect 7248 5664 7380 5692
rect 7248 5652 7254 5664
rect 7374 5652 7380 5664
rect 7432 5652 7438 5704
rect 7742 5652 7748 5704
rect 7800 5692 7806 5704
rect 7929 5695 7987 5701
rect 7929 5692 7941 5695
rect 7800 5664 7941 5692
rect 7800 5652 7806 5664
rect 7929 5661 7941 5664
rect 7975 5661 7987 5695
rect 7929 5655 7987 5661
rect 8018 5652 8024 5704
rect 8076 5652 8082 5704
rect 8113 5695 8171 5701
rect 8113 5661 8125 5695
rect 8159 5692 8171 5695
rect 8202 5692 8208 5704
rect 8159 5664 8208 5692
rect 8159 5661 8171 5664
rect 8113 5655 8171 5661
rect 8202 5652 8208 5664
rect 8260 5652 8266 5704
rect 5184 5596 6500 5624
rect 2682 5516 2688 5568
rect 2740 5556 2746 5568
rect 5184 5556 5212 5596
rect 2740 5528 5212 5556
rect 2740 5516 2746 5528
rect 5258 5516 5264 5568
rect 5316 5556 5322 5568
rect 5629 5559 5687 5565
rect 5629 5556 5641 5559
rect 5316 5528 5641 5556
rect 5316 5516 5322 5528
rect 5629 5525 5641 5528
rect 5675 5525 5687 5559
rect 6472 5556 6500 5596
rect 6549 5627 6607 5633
rect 6549 5593 6561 5627
rect 6595 5593 6607 5627
rect 8312 5624 8340 5732
rect 9944 5729 9956 5763
rect 9990 5760 10002 5763
rect 11698 5760 11704 5772
rect 9990 5732 11704 5760
rect 9990 5729 10002 5732
rect 9944 5723 10002 5729
rect 11698 5720 11704 5732
rect 11756 5760 11762 5772
rect 13832 5769 13860 5800
rect 20254 5788 20260 5800
rect 20312 5788 20318 5840
rect 13817 5763 13875 5769
rect 11756 5732 12480 5760
rect 11756 5720 11762 5732
rect 8754 5652 8760 5704
rect 8812 5692 8818 5704
rect 9033 5695 9091 5701
rect 9033 5692 9045 5695
rect 8812 5664 9045 5692
rect 8812 5652 8818 5664
rect 9033 5661 9045 5664
rect 9079 5661 9091 5695
rect 9033 5655 9091 5661
rect 9122 5652 9128 5704
rect 9180 5692 9186 5704
rect 9217 5695 9275 5701
rect 9217 5692 9229 5695
rect 9180 5664 9229 5692
rect 9180 5652 9186 5664
rect 9217 5661 9229 5664
rect 9263 5692 9275 5695
rect 9401 5695 9459 5701
rect 9401 5692 9413 5695
rect 9263 5664 9413 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 9401 5661 9413 5664
rect 9447 5661 9459 5695
rect 9401 5655 9459 5661
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5661 9735 5695
rect 11330 5692 11336 5704
rect 9677 5655 9735 5661
rect 11072 5664 11336 5692
rect 6549 5587 6607 5593
rect 7197 5596 8340 5624
rect 8573 5627 8631 5633
rect 7197 5556 7225 5596
rect 8573 5593 8585 5627
rect 8619 5624 8631 5627
rect 8662 5624 8668 5636
rect 8619 5596 8668 5624
rect 8619 5593 8631 5596
rect 8573 5587 8631 5593
rect 8662 5584 8668 5596
rect 8720 5584 8726 5636
rect 9692 5624 9720 5655
rect 9324 5596 9720 5624
rect 6472 5528 7225 5556
rect 5629 5519 5687 5525
rect 7558 5516 7564 5568
rect 7616 5556 7622 5568
rect 9324 5556 9352 5596
rect 10962 5584 10968 5636
rect 11020 5624 11026 5636
rect 11072 5633 11100 5664
rect 11330 5652 11336 5664
rect 11388 5652 11394 5704
rect 11606 5652 11612 5704
rect 11664 5692 11670 5704
rect 11974 5692 11980 5704
rect 11664 5664 11980 5692
rect 11664 5652 11670 5664
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 12342 5692 12348 5704
rect 12303 5664 12348 5692
rect 12342 5652 12348 5664
rect 12400 5652 12406 5704
rect 12452 5701 12480 5732
rect 13817 5729 13829 5763
rect 13863 5729 13875 5763
rect 15838 5760 15844 5772
rect 15799 5732 15844 5760
rect 13817 5723 13875 5729
rect 15838 5720 15844 5732
rect 15896 5720 15902 5772
rect 16108 5763 16166 5769
rect 16108 5729 16120 5763
rect 16154 5760 16166 5763
rect 16390 5760 16396 5772
rect 16154 5732 16396 5760
rect 16154 5729 16166 5732
rect 16108 5723 16166 5729
rect 16390 5720 16396 5732
rect 16448 5720 16454 5772
rect 17862 5760 17868 5772
rect 17420 5732 17868 5760
rect 17420 5704 17448 5732
rect 17862 5720 17868 5732
rect 17920 5760 17926 5772
rect 18598 5769 18604 5772
rect 18325 5763 18383 5769
rect 18325 5760 18337 5763
rect 17920 5732 18337 5760
rect 17920 5720 17926 5732
rect 18325 5729 18337 5732
rect 18371 5729 18383 5763
rect 18592 5760 18604 5769
rect 18559 5732 18604 5760
rect 18325 5723 18383 5729
rect 18592 5723 18604 5732
rect 18598 5720 18604 5723
rect 18656 5720 18662 5772
rect 12437 5695 12495 5701
rect 12437 5661 12449 5695
rect 12483 5661 12495 5695
rect 12437 5655 12495 5661
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 14001 5695 14059 5701
rect 14001 5692 14013 5695
rect 13964 5664 14013 5692
rect 13964 5652 13970 5664
rect 14001 5661 14013 5664
rect 14047 5661 14059 5695
rect 14001 5655 14059 5661
rect 17402 5652 17408 5704
rect 17460 5652 17466 5704
rect 11057 5627 11115 5633
rect 11057 5624 11069 5627
rect 11020 5596 11069 5624
rect 11020 5584 11026 5596
rect 11057 5593 11069 5596
rect 11103 5593 11115 5627
rect 14458 5624 14464 5636
rect 11057 5587 11115 5593
rect 11164 5596 14464 5624
rect 7616 5528 9352 5556
rect 9401 5559 9459 5565
rect 7616 5516 7622 5528
rect 9401 5525 9413 5559
rect 9447 5556 9459 5559
rect 11164 5556 11192 5596
rect 14458 5584 14464 5596
rect 14516 5584 14522 5636
rect 19426 5584 19432 5636
rect 19484 5624 19490 5636
rect 19705 5627 19763 5633
rect 19705 5624 19717 5627
rect 19484 5596 19717 5624
rect 19484 5584 19490 5596
rect 19705 5593 19717 5596
rect 19751 5593 19763 5627
rect 19705 5587 19763 5593
rect 11882 5556 11888 5568
rect 9447 5528 11192 5556
rect 11843 5528 11888 5556
rect 9447 5525 9459 5528
rect 9401 5519 9459 5525
rect 11882 5516 11888 5528
rect 11940 5516 11946 5568
rect 12158 5516 12164 5568
rect 12216 5556 12222 5568
rect 13449 5559 13507 5565
rect 13449 5556 13461 5559
rect 12216 5528 13461 5556
rect 12216 5516 12222 5528
rect 13449 5525 13461 5528
rect 13495 5525 13507 5559
rect 13449 5519 13507 5525
rect 13538 5516 13544 5568
rect 13596 5556 13602 5568
rect 16574 5556 16580 5568
rect 13596 5528 16580 5556
rect 13596 5516 13602 5528
rect 16574 5516 16580 5528
rect 16632 5516 16638 5568
rect 17218 5556 17224 5568
rect 17131 5528 17224 5556
rect 17218 5516 17224 5528
rect 17276 5556 17282 5568
rect 17770 5556 17776 5568
rect 17276 5528 17776 5556
rect 17276 5516 17282 5528
rect 17770 5516 17776 5528
rect 17828 5516 17834 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 2406 5312 2412 5364
rect 2464 5352 2470 5364
rect 7745 5355 7803 5361
rect 2464 5324 6488 5352
rect 2464 5312 2470 5324
rect 4062 5244 4068 5296
rect 4120 5244 4126 5296
rect 4154 5244 4160 5296
rect 4212 5284 4218 5296
rect 4249 5287 4307 5293
rect 4249 5284 4261 5287
rect 4212 5256 4261 5284
rect 4212 5244 4218 5256
rect 4249 5253 4261 5256
rect 4295 5253 4307 5287
rect 4249 5247 4307 5253
rect 2774 5176 2780 5228
rect 2832 5216 2838 5228
rect 4080 5216 4108 5244
rect 6362 5216 6368 5228
rect 2832 5188 3004 5216
rect 4080 5188 4476 5216
rect 6323 5188 6368 5216
rect 2832 5176 2838 5188
rect 2866 5148 2872 5160
rect 2779 5120 2872 5148
rect 2866 5108 2872 5120
rect 2924 5108 2930 5160
rect 2976 5148 3004 5188
rect 3125 5151 3183 5157
rect 3125 5148 3137 5151
rect 2976 5120 3137 5148
rect 3125 5117 3137 5120
rect 3171 5117 3183 5151
rect 3125 5111 3183 5117
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 4341 5151 4399 5157
rect 4341 5148 4353 5151
rect 4120 5120 4353 5148
rect 4120 5108 4126 5120
rect 4341 5117 4353 5120
rect 4387 5117 4399 5151
rect 4341 5111 4399 5117
rect 1670 5089 1676 5092
rect 1664 5080 1676 5089
rect 1631 5052 1676 5080
rect 1664 5043 1676 5052
rect 1670 5040 1676 5043
rect 1728 5040 1734 5092
rect 2884 5080 2912 5108
rect 4080 5080 4108 5108
rect 2884 5052 4108 5080
rect 4448 5080 4476 5188
rect 6362 5176 6368 5188
rect 6420 5176 6426 5228
rect 4608 5151 4666 5157
rect 4608 5117 4620 5151
rect 4654 5148 4666 5151
rect 5350 5148 5356 5160
rect 4654 5120 5356 5148
rect 4654 5117 4666 5120
rect 4608 5111 4666 5117
rect 5350 5108 5356 5120
rect 5408 5108 5414 5160
rect 6181 5151 6239 5157
rect 6181 5117 6193 5151
rect 6227 5148 6239 5151
rect 6270 5148 6276 5160
rect 6227 5120 6276 5148
rect 6227 5117 6239 5120
rect 6181 5111 6239 5117
rect 6270 5108 6276 5120
rect 6328 5108 6334 5160
rect 6460 5148 6488 5324
rect 7745 5321 7757 5355
rect 7791 5352 7803 5355
rect 7834 5352 7840 5364
rect 7791 5324 7840 5352
rect 7791 5321 7803 5324
rect 7745 5315 7803 5321
rect 7834 5312 7840 5324
rect 7892 5312 7898 5364
rect 11882 5352 11888 5364
rect 7944 5324 9352 5352
rect 7944 5284 7972 5324
rect 8294 5284 8300 5296
rect 6840 5256 7972 5284
rect 8220 5256 8300 5284
rect 6730 5176 6736 5228
rect 6788 5216 6794 5228
rect 6840 5216 6868 5256
rect 6788 5188 6868 5216
rect 6788 5176 6794 5188
rect 6914 5176 6920 5228
rect 6972 5216 6978 5228
rect 7285 5219 7343 5225
rect 7285 5216 7297 5219
rect 6972 5188 7297 5216
rect 6972 5176 6978 5188
rect 7285 5185 7297 5188
rect 7331 5185 7343 5219
rect 7285 5179 7343 5185
rect 7374 5176 7380 5228
rect 7432 5216 7438 5228
rect 7469 5219 7527 5225
rect 7469 5216 7481 5219
rect 7432 5188 7481 5216
rect 7432 5176 7438 5188
rect 7469 5185 7481 5188
rect 7515 5216 7527 5219
rect 7653 5219 7711 5225
rect 7653 5216 7665 5219
rect 7515 5188 7665 5216
rect 7515 5185 7527 5188
rect 7469 5179 7527 5185
rect 7653 5185 7665 5188
rect 7699 5185 7711 5219
rect 8220 5216 8248 5256
rect 8294 5244 8300 5256
rect 8352 5244 8358 5296
rect 8662 5284 8668 5296
rect 8623 5256 8668 5284
rect 8662 5244 8668 5256
rect 8720 5244 8726 5296
rect 9030 5244 9036 5296
rect 9088 5284 9094 5296
rect 9088 5256 9168 5284
rect 9088 5244 9094 5256
rect 8386 5216 8392 5228
rect 7653 5179 7711 5185
rect 7852 5188 8248 5216
rect 8347 5188 8392 5216
rect 6460 5120 6592 5148
rect 5166 5080 5172 5092
rect 4448 5052 5172 5080
rect 5166 5040 5172 5052
rect 5224 5040 5230 5092
rect 5902 5080 5908 5092
rect 5552 5052 5908 5080
rect 2777 5015 2835 5021
rect 2777 4981 2789 5015
rect 2823 5012 2835 5015
rect 4246 5012 4252 5024
rect 2823 4984 4252 5012
rect 2823 4981 2835 4984
rect 2777 4975 2835 4981
rect 4246 4972 4252 4984
rect 4304 4972 4310 5024
rect 4430 4972 4436 5024
rect 4488 5012 4494 5024
rect 5552 5012 5580 5052
rect 5902 5040 5908 5052
rect 5960 5040 5966 5092
rect 6454 5040 6460 5092
rect 6512 5040 6518 5092
rect 6564 5080 6592 5120
rect 7098 5108 7104 5160
rect 7156 5148 7162 5160
rect 7392 5148 7420 5176
rect 7852 5148 7880 5188
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 9140 5225 9168 5256
rect 9324 5225 9352 5324
rect 11164 5324 11888 5352
rect 9674 5244 9680 5296
rect 9732 5284 9738 5296
rect 11164 5284 11192 5324
rect 11882 5312 11888 5324
rect 11940 5312 11946 5364
rect 11992 5324 14044 5352
rect 9732 5256 10272 5284
rect 9732 5244 9738 5256
rect 9125 5219 9183 5225
rect 9125 5185 9137 5219
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 9309 5219 9367 5225
rect 9309 5185 9321 5219
rect 9355 5216 9367 5219
rect 9355 5188 10088 5216
rect 9355 5185 9367 5188
rect 9309 5179 9367 5185
rect 7156 5120 7420 5148
rect 7576 5120 7880 5148
rect 7156 5108 7162 5120
rect 7193 5083 7251 5089
rect 7193 5080 7205 5083
rect 6564 5052 7205 5080
rect 7193 5049 7205 5052
rect 7239 5049 7251 5083
rect 7193 5043 7251 5049
rect 7282 5040 7288 5092
rect 7340 5080 7346 5092
rect 7576 5080 7604 5120
rect 7926 5108 7932 5160
rect 7984 5148 7990 5160
rect 8113 5151 8171 5157
rect 8113 5148 8125 5151
rect 7984 5120 8125 5148
rect 7984 5108 7990 5120
rect 8113 5117 8125 5120
rect 8159 5117 8171 5151
rect 8113 5111 8171 5117
rect 8202 5108 8208 5160
rect 8260 5148 8266 5160
rect 8662 5148 8668 5160
rect 8260 5120 8305 5148
rect 8404 5120 8668 5148
rect 8260 5108 8266 5120
rect 7340 5052 7604 5080
rect 7653 5083 7711 5089
rect 7340 5040 7346 5052
rect 7653 5049 7665 5083
rect 7699 5080 7711 5083
rect 8404 5080 8432 5120
rect 8662 5108 8668 5120
rect 8720 5108 8726 5160
rect 9033 5151 9091 5157
rect 9033 5117 9045 5151
rect 9079 5148 9091 5151
rect 9950 5148 9956 5160
rect 9079 5120 9956 5148
rect 9079 5117 9091 5120
rect 9033 5111 9091 5117
rect 9950 5108 9956 5120
rect 10008 5108 10014 5160
rect 7699 5052 8432 5080
rect 7699 5049 7711 5052
rect 7653 5043 7711 5049
rect 8478 5040 8484 5092
rect 8536 5080 8542 5092
rect 10060 5080 10088 5188
rect 10244 5157 10272 5256
rect 10336 5256 11192 5284
rect 10336 5225 10364 5256
rect 11330 5244 11336 5296
rect 11388 5284 11394 5296
rect 11992 5284 12020 5324
rect 11388 5256 12020 5284
rect 11388 5244 11394 5256
rect 10321 5219 10379 5225
rect 10321 5185 10333 5219
rect 10367 5185 10379 5219
rect 10321 5179 10379 5185
rect 10413 5219 10471 5225
rect 10413 5185 10425 5219
rect 10459 5185 10471 5219
rect 10413 5179 10471 5185
rect 10229 5151 10287 5157
rect 10229 5117 10241 5151
rect 10275 5117 10287 5151
rect 10428 5148 10456 5179
rect 10686 5176 10692 5228
rect 10744 5216 10750 5228
rect 12158 5216 12164 5228
rect 10744 5188 12164 5216
rect 10744 5176 10750 5188
rect 12158 5176 12164 5188
rect 12216 5176 12222 5228
rect 12434 5216 12440 5228
rect 12395 5188 12440 5216
rect 12434 5176 12440 5188
rect 12492 5176 12498 5228
rect 10502 5148 10508 5160
rect 10428 5120 10508 5148
rect 10229 5111 10287 5117
rect 10502 5108 10508 5120
rect 10560 5108 10566 5160
rect 10594 5108 10600 5160
rect 10652 5148 10658 5160
rect 10962 5148 10968 5160
rect 10652 5120 10968 5148
rect 10652 5108 10658 5120
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 11974 5108 11980 5160
rect 12032 5148 12038 5160
rect 12693 5151 12751 5157
rect 12693 5148 12705 5151
rect 12032 5120 12705 5148
rect 12032 5108 12038 5120
rect 12693 5117 12705 5120
rect 12739 5148 12751 5151
rect 13078 5148 13084 5160
rect 12739 5120 13084 5148
rect 12739 5117 12751 5120
rect 12693 5111 12751 5117
rect 13078 5108 13084 5120
rect 13136 5148 13142 5160
rect 13906 5148 13912 5160
rect 13136 5120 13912 5148
rect 13136 5108 13142 5120
rect 13906 5108 13912 5120
rect 13964 5108 13970 5160
rect 11882 5080 11888 5092
rect 8536 5052 8984 5080
rect 10060 5052 11888 5080
rect 8536 5040 8542 5052
rect 4488 4984 5580 5012
rect 4488 4972 4494 4984
rect 5626 4972 5632 5024
rect 5684 5012 5690 5024
rect 5721 5015 5779 5021
rect 5721 5012 5733 5015
rect 5684 4984 5733 5012
rect 5684 4972 5690 4984
rect 5721 4981 5733 4984
rect 5767 4981 5779 5015
rect 5721 4975 5779 4981
rect 5810 4972 5816 5024
rect 5868 5012 5874 5024
rect 6270 5012 6276 5024
rect 5868 4984 5913 5012
rect 6231 4984 6276 5012
rect 5868 4972 5874 4984
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 6472 5012 6500 5040
rect 6546 5012 6552 5024
rect 6472 4984 6552 5012
rect 6546 4972 6552 4984
rect 6604 4972 6610 5024
rect 6825 5015 6883 5021
rect 6825 4981 6837 5015
rect 6871 5012 6883 5015
rect 7374 5012 7380 5024
rect 6871 4984 7380 5012
rect 6871 4981 6883 4984
rect 6825 4975 6883 4981
rect 7374 4972 7380 4984
rect 7432 4972 7438 5024
rect 7558 4972 7564 5024
rect 7616 5012 7622 5024
rect 8754 5012 8760 5024
rect 7616 4984 8760 5012
rect 7616 4972 7622 4984
rect 8754 4972 8760 4984
rect 8812 4972 8818 5024
rect 8956 5012 8984 5052
rect 11882 5040 11888 5052
rect 11940 5040 11946 5092
rect 12342 5040 12348 5092
rect 12400 5040 12406 5092
rect 14016 5080 14044 5324
rect 14550 5312 14556 5364
rect 14608 5352 14614 5364
rect 14608 5324 15700 5352
rect 14608 5312 14614 5324
rect 15672 5216 15700 5324
rect 16574 5312 16580 5364
rect 16632 5352 16638 5364
rect 19426 5352 19432 5364
rect 16632 5324 19432 5352
rect 16632 5312 16638 5324
rect 19426 5312 19432 5324
rect 19484 5312 19490 5364
rect 16022 5284 16028 5296
rect 15983 5256 16028 5284
rect 16022 5244 16028 5256
rect 16080 5244 16086 5296
rect 17037 5287 17095 5293
rect 17037 5253 17049 5287
rect 17083 5284 17095 5287
rect 19242 5284 19248 5296
rect 17083 5256 19248 5284
rect 17083 5253 17095 5256
rect 17037 5247 17095 5253
rect 19242 5244 19248 5256
rect 19300 5244 19306 5296
rect 15672 5188 15976 5216
rect 14642 5148 14648 5160
rect 14555 5120 14648 5148
rect 14642 5108 14648 5120
rect 14700 5148 14706 5160
rect 15838 5148 15844 5160
rect 14700 5120 15844 5148
rect 14700 5108 14706 5120
rect 15838 5108 15844 5120
rect 15896 5108 15902 5160
rect 14734 5080 14740 5092
rect 14016 5052 14740 5080
rect 14734 5040 14740 5052
rect 14792 5040 14798 5092
rect 14890 5083 14948 5089
rect 14890 5049 14902 5083
rect 14936 5049 14948 5083
rect 15948 5080 15976 5188
rect 16482 5176 16488 5228
rect 16540 5216 16546 5228
rect 18601 5219 18659 5225
rect 16540 5188 18460 5216
rect 16540 5176 16546 5188
rect 16850 5148 16856 5160
rect 16811 5120 16856 5148
rect 16850 5108 16856 5120
rect 16908 5108 16914 5160
rect 17954 5148 17960 5160
rect 16960 5120 17960 5148
rect 16960 5080 16988 5120
rect 17954 5108 17960 5120
rect 18012 5108 18018 5160
rect 18432 5157 18460 5188
rect 18601 5185 18613 5219
rect 18647 5216 18659 5219
rect 18782 5216 18788 5228
rect 18647 5188 18788 5216
rect 18647 5185 18659 5188
rect 18601 5179 18659 5185
rect 18782 5176 18788 5188
rect 18840 5176 18846 5228
rect 20165 5219 20223 5225
rect 20165 5216 20177 5219
rect 18892 5188 20177 5216
rect 18417 5151 18475 5157
rect 18417 5117 18429 5151
rect 18463 5117 18475 5151
rect 18417 5111 18475 5117
rect 18509 5151 18567 5157
rect 18509 5117 18521 5151
rect 18555 5148 18567 5151
rect 18690 5148 18696 5160
rect 18555 5120 18696 5148
rect 18555 5117 18567 5120
rect 18509 5111 18567 5117
rect 18690 5108 18696 5120
rect 18748 5108 18754 5160
rect 15948 5052 16988 5080
rect 14890 5043 14948 5049
rect 9030 5012 9036 5024
rect 8956 4984 9036 5012
rect 9030 4972 9036 4984
rect 9088 4972 9094 5024
rect 9861 5015 9919 5021
rect 9861 4981 9873 5015
rect 9907 5012 9919 5015
rect 10410 5012 10416 5024
rect 9907 4984 10416 5012
rect 9907 4981 9919 4984
rect 9861 4975 9919 4981
rect 10410 4972 10416 4984
rect 10468 4972 10474 5024
rect 10594 4972 10600 5024
rect 10652 5012 10658 5024
rect 12158 5012 12164 5024
rect 10652 4984 12164 5012
rect 10652 4972 10658 4984
rect 12158 4972 12164 4984
rect 12216 4972 12222 5024
rect 12360 5012 12388 5040
rect 12802 5012 12808 5024
rect 12360 4984 12808 5012
rect 12802 4972 12808 4984
rect 12860 4972 12866 5024
rect 13814 5012 13820 5024
rect 13775 4984 13820 5012
rect 13814 4972 13820 4984
rect 13872 5012 13878 5024
rect 14905 5012 14933 5043
rect 17770 5040 17776 5092
rect 17828 5080 17834 5092
rect 18892 5080 18920 5188
rect 20165 5185 20177 5188
rect 20211 5185 20223 5219
rect 20165 5179 20223 5185
rect 17828 5052 18920 5080
rect 17828 5040 17834 5052
rect 19058 5040 19064 5092
rect 19116 5080 19122 5092
rect 20073 5083 20131 5089
rect 20073 5080 20085 5083
rect 19116 5052 20085 5080
rect 19116 5040 19122 5052
rect 20073 5049 20085 5052
rect 20119 5049 20131 5083
rect 20073 5043 20131 5049
rect 13872 4984 14933 5012
rect 13872 4972 13878 4984
rect 15378 4972 15384 5024
rect 15436 5012 15442 5024
rect 17218 5012 17224 5024
rect 15436 4984 17224 5012
rect 15436 4972 15442 4984
rect 17218 4972 17224 4984
rect 17276 4972 17282 5024
rect 18046 5012 18052 5024
rect 18007 4984 18052 5012
rect 18046 4972 18052 4984
rect 18104 4972 18110 5024
rect 19610 5012 19616 5024
rect 19571 4984 19616 5012
rect 19610 4972 19616 4984
rect 19668 4972 19674 5024
rect 19978 5012 19984 5024
rect 19939 4984 19984 5012
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 3326 4808 3332 4820
rect 3287 4780 3332 4808
rect 3326 4768 3332 4780
rect 3384 4768 3390 4820
rect 3436 4780 4108 4808
rect 3237 4743 3295 4749
rect 3237 4709 3249 4743
rect 3283 4740 3295 4743
rect 3436 4740 3464 4780
rect 3283 4712 3464 4740
rect 4080 4740 4108 4780
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 5166 4808 5172 4820
rect 4212 4780 5172 4808
rect 4212 4768 4218 4780
rect 5166 4768 5172 4780
rect 5224 4768 5230 4820
rect 5350 4768 5356 4820
rect 5408 4808 5414 4820
rect 5445 4811 5503 4817
rect 5445 4808 5457 4811
rect 5408 4780 5457 4808
rect 5408 4768 5414 4780
rect 5445 4777 5457 4780
rect 5491 4777 5503 4811
rect 5994 4808 6000 4820
rect 5445 4771 5503 4777
rect 5736 4780 6000 4808
rect 5736 4740 5764 4780
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 6638 4768 6644 4820
rect 6696 4808 6702 4820
rect 6733 4811 6791 4817
rect 6733 4808 6745 4811
rect 6696 4780 6745 4808
rect 6696 4768 6702 4780
rect 6733 4777 6745 4780
rect 6779 4777 6791 4811
rect 6733 4771 6791 4777
rect 7190 4768 7196 4820
rect 7248 4808 7254 4820
rect 7466 4808 7472 4820
rect 7248 4780 7472 4808
rect 7248 4768 7254 4780
rect 7466 4768 7472 4780
rect 7524 4808 7530 4820
rect 8297 4811 8355 4817
rect 8297 4808 8309 4811
rect 7524 4780 8309 4808
rect 7524 4768 7530 4780
rect 8297 4777 8309 4780
rect 8343 4777 8355 4811
rect 8297 4771 8355 4777
rect 8665 4811 8723 4817
rect 8665 4777 8677 4811
rect 8711 4808 8723 4811
rect 8711 4780 9536 4808
rect 8711 4777 8723 4780
rect 8665 4771 8723 4777
rect 4080 4712 5764 4740
rect 3283 4709 3295 4712
rect 3237 4703 3295 4709
rect 5810 4700 5816 4752
rect 5868 4740 5874 4752
rect 5868 4712 6776 4740
rect 5868 4700 5874 4712
rect 1664 4675 1722 4681
rect 1664 4641 1676 4675
rect 1710 4672 1722 4675
rect 2682 4672 2688 4684
rect 1710 4644 2688 4672
rect 1710 4641 1722 4644
rect 1664 4635 1722 4641
rect 2682 4632 2688 4644
rect 2740 4632 2746 4684
rect 4065 4675 4123 4681
rect 4065 4641 4077 4675
rect 4111 4672 4123 4675
rect 4154 4672 4160 4684
rect 4111 4644 4160 4672
rect 4111 4641 4123 4644
rect 4065 4635 4123 4641
rect 4154 4632 4160 4644
rect 4212 4632 4218 4684
rect 4332 4675 4390 4681
rect 4332 4641 4344 4675
rect 4378 4672 4390 4675
rect 5718 4672 5724 4684
rect 4378 4644 5724 4672
rect 4378 4641 4390 4644
rect 4332 4635 4390 4641
rect 5718 4632 5724 4644
rect 5776 4632 5782 4684
rect 5905 4675 5963 4681
rect 5905 4641 5917 4675
rect 5951 4641 5963 4675
rect 5905 4635 5963 4641
rect 5997 4675 6055 4681
rect 5997 4641 6009 4675
rect 6043 4672 6055 4675
rect 6178 4672 6184 4684
rect 6043 4644 6184 4672
rect 6043 4641 6055 4644
rect 5997 4635 6055 4641
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4604 3571 4607
rect 3970 4604 3976 4616
rect 3559 4576 3976 4604
rect 3559 4573 3571 4576
rect 3513 4567 3571 4573
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 5258 4564 5264 4616
rect 5316 4604 5322 4616
rect 5316 4576 5764 4604
rect 5316 4564 5322 4576
rect 2777 4539 2835 4545
rect 2777 4505 2789 4539
rect 2823 4536 2835 4539
rect 2958 4536 2964 4548
rect 2823 4508 2964 4536
rect 2823 4505 2835 4508
rect 2777 4499 2835 4505
rect 2958 4496 2964 4508
rect 3016 4536 3022 4548
rect 3694 4536 3700 4548
rect 3016 4508 3700 4536
rect 3016 4496 3022 4508
rect 3694 4496 3700 4508
rect 3752 4496 3758 4548
rect 5626 4536 5632 4548
rect 5368 4508 5632 4536
rect 2869 4471 2927 4477
rect 2869 4437 2881 4471
rect 2915 4468 2927 4471
rect 5368 4468 5396 4508
rect 5626 4496 5632 4508
rect 5684 4496 5690 4548
rect 2915 4440 5396 4468
rect 5537 4471 5595 4477
rect 2915 4437 2927 4440
rect 2869 4431 2927 4437
rect 5537 4437 5549 4471
rect 5583 4468 5595 4471
rect 5736 4468 5764 4576
rect 5583 4440 5764 4468
rect 5583 4437 5595 4440
rect 5537 4431 5595 4437
rect 5810 4428 5816 4480
rect 5868 4468 5874 4480
rect 5920 4468 5948 4635
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 6748 4672 6776 4712
rect 6822 4700 6828 4752
rect 6880 4740 6886 4752
rect 7006 4740 7012 4752
rect 6880 4712 7012 4740
rect 6880 4700 6886 4712
rect 7006 4700 7012 4712
rect 7064 4700 7070 4752
rect 7745 4743 7803 4749
rect 7116 4712 7696 4740
rect 7116 4672 7144 4712
rect 6748 4644 7144 4672
rect 7193 4675 7251 4681
rect 7193 4641 7205 4675
rect 7239 4641 7251 4675
rect 7193 4635 7251 4641
rect 6089 4607 6147 4613
rect 6089 4573 6101 4607
rect 6135 4604 6147 4607
rect 6454 4604 6460 4616
rect 6135 4576 6460 4604
rect 6135 4573 6147 4576
rect 6089 4567 6147 4573
rect 6454 4564 6460 4576
rect 6512 4564 6518 4616
rect 6822 4604 6828 4616
rect 6783 4576 6828 4604
rect 6822 4564 6828 4576
rect 6880 4564 6886 4616
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4573 6975 4607
rect 6917 4567 6975 4573
rect 5994 4496 6000 4548
rect 6052 4536 6058 4548
rect 6730 4536 6736 4548
rect 6052 4508 6736 4536
rect 6052 4496 6058 4508
rect 6730 4496 6736 4508
rect 6788 4496 6794 4548
rect 5868 4440 5948 4468
rect 5868 4428 5874 4440
rect 6086 4428 6092 4480
rect 6144 4468 6150 4480
rect 6365 4471 6423 4477
rect 6365 4468 6377 4471
rect 6144 4440 6377 4468
rect 6144 4428 6150 4440
rect 6365 4437 6377 4440
rect 6411 4437 6423 4471
rect 6932 4468 6960 4567
rect 7199 4536 7227 4635
rect 7282 4632 7288 4684
rect 7340 4672 7346 4684
rect 7558 4672 7564 4684
rect 7340 4644 7564 4672
rect 7340 4632 7346 4644
rect 7558 4632 7564 4644
rect 7616 4632 7622 4684
rect 7668 4672 7696 4712
rect 7745 4709 7757 4743
rect 7791 4740 7803 4743
rect 7791 4712 8064 4740
rect 7791 4709 7803 4712
rect 7745 4703 7803 4709
rect 8036 4672 8064 4712
rect 8110 4700 8116 4752
rect 8168 4740 8174 4752
rect 8205 4743 8263 4749
rect 8205 4740 8217 4743
rect 8168 4712 8217 4740
rect 8168 4700 8174 4712
rect 8205 4709 8217 4712
rect 8251 4740 8263 4743
rect 9030 4740 9036 4752
rect 8251 4712 8892 4740
rect 8991 4712 9036 4740
rect 8251 4709 8263 4712
rect 8205 4703 8263 4709
rect 8864 4672 8892 4712
rect 9030 4700 9036 4712
rect 9088 4700 9094 4752
rect 9508 4740 9536 4780
rect 9674 4768 9680 4820
rect 9732 4808 9738 4820
rect 9953 4811 10011 4817
rect 9953 4808 9965 4811
rect 9732 4780 9965 4808
rect 9732 4768 9738 4780
rect 9953 4777 9965 4780
rect 9999 4777 10011 4811
rect 9953 4771 10011 4777
rect 10134 4768 10140 4820
rect 10192 4808 10198 4820
rect 10321 4811 10379 4817
rect 10321 4808 10333 4811
rect 10192 4780 10333 4808
rect 10192 4768 10198 4780
rect 10321 4777 10333 4780
rect 10367 4777 10379 4811
rect 11330 4808 11336 4820
rect 10321 4771 10379 4777
rect 10888 4780 11336 4808
rect 10226 4740 10232 4752
rect 9508 4712 10232 4740
rect 10226 4700 10232 4712
rect 10284 4700 10290 4752
rect 10413 4743 10471 4749
rect 10413 4709 10425 4743
rect 10459 4740 10471 4743
rect 10502 4740 10508 4752
rect 10459 4712 10508 4740
rect 10459 4709 10471 4712
rect 10413 4703 10471 4709
rect 10502 4700 10508 4712
rect 10560 4740 10566 4752
rect 10888 4740 10916 4780
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 13173 4811 13231 4817
rect 13173 4777 13185 4811
rect 13219 4808 13231 4811
rect 20070 4808 20076 4820
rect 13219 4780 20076 4808
rect 13219 4777 13231 4780
rect 13173 4771 13231 4777
rect 20070 4768 20076 4780
rect 20128 4768 20134 4820
rect 11054 4740 11060 4752
rect 10560 4712 10916 4740
rect 11015 4712 11060 4740
rect 10560 4700 10566 4712
rect 11054 4700 11060 4712
rect 11112 4700 11118 4752
rect 11146 4700 11152 4752
rect 11204 4740 11210 4752
rect 11977 4743 12035 4749
rect 11977 4740 11989 4743
rect 11204 4712 11989 4740
rect 11204 4700 11210 4712
rect 11977 4709 11989 4712
rect 12023 4740 12035 4743
rect 13446 4740 13452 4752
rect 12023 4712 13452 4740
rect 12023 4709 12035 4712
rect 11977 4703 12035 4709
rect 13446 4700 13452 4712
rect 13504 4700 13510 4752
rect 13630 4740 13636 4752
rect 13591 4712 13636 4740
rect 13630 4700 13636 4712
rect 13688 4700 13694 4752
rect 15194 4700 15200 4752
rect 15252 4740 15258 4752
rect 16209 4743 16267 4749
rect 16209 4740 16221 4743
rect 15252 4712 16221 4740
rect 15252 4700 15258 4712
rect 16209 4709 16221 4712
rect 16255 4709 16267 4743
rect 16209 4703 16267 4709
rect 7668 4644 7972 4672
rect 8036 4644 8340 4672
rect 8864 4644 9260 4672
rect 7469 4607 7527 4613
rect 7469 4573 7481 4607
rect 7515 4604 7527 4607
rect 7745 4607 7803 4613
rect 7745 4604 7757 4607
rect 7515 4576 7757 4604
rect 7515 4573 7527 4576
rect 7469 4567 7527 4573
rect 7745 4573 7757 4576
rect 7791 4573 7803 4607
rect 7944 4604 7972 4644
rect 7944 4576 8064 4604
rect 7745 4567 7803 4573
rect 7199 4508 7972 4536
rect 7944 4480 7972 4508
rect 7374 4468 7380 4480
rect 6932 4440 7380 4468
rect 6365 4431 6423 4437
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 7742 4428 7748 4480
rect 7800 4468 7806 4480
rect 7837 4471 7895 4477
rect 7837 4468 7849 4471
rect 7800 4440 7849 4468
rect 7800 4428 7806 4440
rect 7837 4437 7849 4440
rect 7883 4437 7895 4471
rect 7837 4431 7895 4437
rect 7926 4428 7932 4480
rect 7984 4428 7990 4480
rect 8036 4468 8064 4576
rect 8312 4548 8340 4644
rect 8478 4564 8484 4616
rect 8536 4604 8542 4616
rect 9125 4607 9183 4613
rect 8536 4576 8581 4604
rect 8536 4564 8542 4576
rect 9125 4573 9137 4607
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 8294 4496 8300 4548
rect 8352 4496 8358 4548
rect 9140 4468 9168 4567
rect 9232 4536 9260 4644
rect 9490 4632 9496 4684
rect 9548 4672 9554 4684
rect 10778 4672 10784 4684
rect 9548 4644 10640 4672
rect 10739 4644 10784 4672
rect 9548 4632 9554 4644
rect 9309 4607 9367 4613
rect 9309 4573 9321 4607
rect 9355 4604 9367 4607
rect 9674 4604 9680 4616
rect 9355 4576 9680 4604
rect 9355 4573 9367 4576
rect 9309 4567 9367 4573
rect 9674 4564 9680 4576
rect 9732 4564 9738 4616
rect 10612 4613 10640 4644
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 11606 4672 11612 4684
rect 10888 4644 11612 4672
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4604 10655 4607
rect 10888 4604 10916 4644
rect 11606 4632 11612 4644
rect 11664 4632 11670 4684
rect 11698 4632 11704 4684
rect 11756 4672 11762 4684
rect 13538 4672 13544 4684
rect 11756 4644 12296 4672
rect 13499 4644 13544 4672
rect 11756 4632 11762 4644
rect 10643 4576 10916 4604
rect 10643 4573 10655 4576
rect 10597 4567 10655 4573
rect 11054 4564 11060 4616
rect 11112 4604 11118 4616
rect 12268 4613 12296 4644
rect 13538 4632 13544 4644
rect 13596 4632 13602 4684
rect 16224 4672 16252 4703
rect 17586 4700 17592 4752
rect 17644 4749 17650 4752
rect 17644 4743 17708 4749
rect 17644 4709 17662 4743
rect 17696 4709 17708 4743
rect 17644 4703 17708 4709
rect 17644 4700 17650 4703
rect 19705 4675 19763 4681
rect 19705 4672 19717 4675
rect 16224 4644 19717 4672
rect 19705 4641 19717 4644
rect 19751 4641 19763 4675
rect 19705 4635 19763 4641
rect 12069 4607 12127 4613
rect 12069 4604 12081 4607
rect 11112 4576 12081 4604
rect 11112 4564 11118 4576
rect 12069 4573 12081 4576
rect 12115 4573 12127 4607
rect 12069 4567 12127 4573
rect 12253 4607 12311 4613
rect 12253 4573 12265 4607
rect 12299 4604 12311 4607
rect 12618 4604 12624 4616
rect 12299 4576 12624 4604
rect 12299 4573 12311 4576
rect 12253 4567 12311 4573
rect 10134 4536 10140 4548
rect 9232 4508 10140 4536
rect 10134 4496 10140 4508
rect 10192 4536 10198 4548
rect 11974 4536 11980 4548
rect 10192 4508 11980 4536
rect 10192 4496 10198 4508
rect 11974 4496 11980 4508
rect 12032 4496 12038 4548
rect 12084 4536 12112 4567
rect 12618 4564 12624 4576
rect 12676 4564 12682 4616
rect 13630 4564 13636 4616
rect 13688 4604 13694 4616
rect 13725 4607 13783 4613
rect 13725 4604 13737 4607
rect 13688 4576 13737 4604
rect 13688 4564 13694 4576
rect 13725 4573 13737 4576
rect 13771 4604 13783 4607
rect 13814 4604 13820 4616
rect 13771 4576 13820 4604
rect 13771 4573 13783 4576
rect 13725 4567 13783 4573
rect 13814 4564 13820 4576
rect 13872 4564 13878 4616
rect 14182 4564 14188 4616
rect 14240 4604 14246 4616
rect 16301 4607 16359 4613
rect 16301 4604 16313 4607
rect 14240 4576 16313 4604
rect 14240 4564 14246 4576
rect 16301 4573 16313 4576
rect 16347 4573 16359 4607
rect 16482 4604 16488 4616
rect 16443 4576 16488 4604
rect 16301 4567 16359 4573
rect 16482 4564 16488 4576
rect 16540 4564 16546 4616
rect 17402 4604 17408 4616
rect 17363 4576 17408 4604
rect 17402 4564 17408 4576
rect 17460 4564 17466 4616
rect 14090 4536 14096 4548
rect 12084 4508 14096 4536
rect 14090 4496 14096 4508
rect 14148 4496 14154 4548
rect 15838 4536 15844 4548
rect 15799 4508 15844 4536
rect 15838 4496 15844 4508
rect 15896 4496 15902 4548
rect 8036 4440 9168 4468
rect 9858 4428 9864 4480
rect 9916 4468 9922 4480
rect 11609 4471 11667 4477
rect 11609 4468 11621 4471
rect 9916 4440 11621 4468
rect 9916 4428 9922 4440
rect 11609 4437 11621 4440
rect 11655 4437 11667 4471
rect 11609 4431 11667 4437
rect 12158 4428 12164 4480
rect 12216 4468 12222 4480
rect 17586 4468 17592 4480
rect 12216 4440 17592 4468
rect 12216 4428 12222 4440
rect 17586 4428 17592 4440
rect 17644 4428 17650 4480
rect 18782 4468 18788 4480
rect 18743 4440 18788 4468
rect 18782 4428 18788 4440
rect 18840 4428 18846 4480
rect 19889 4471 19947 4477
rect 19889 4437 19901 4471
rect 19935 4468 19947 4471
rect 21266 4468 21272 4480
rect 19935 4440 21272 4468
rect 19935 4437 19947 4440
rect 19889 4431 19947 4437
rect 21266 4428 21272 4440
rect 21324 4428 21330 4480
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 2314 4224 2320 4276
rect 2372 4264 2378 4276
rect 5718 4264 5724 4276
rect 2372 4236 5580 4264
rect 5679 4236 5724 4264
rect 2372 4224 2378 4236
rect 5552 4196 5580 4236
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 5810 4224 5816 4276
rect 5868 4264 5874 4276
rect 7282 4264 7288 4276
rect 5868 4236 7288 4264
rect 5868 4224 5874 4236
rect 7282 4224 7288 4236
rect 7340 4224 7346 4276
rect 13630 4264 13636 4276
rect 7484 4236 13636 4264
rect 6086 4196 6092 4208
rect 5552 4168 6092 4196
rect 6086 4156 6092 4168
rect 6144 4156 6150 4208
rect 7098 4196 7104 4208
rect 6196 4168 7104 4196
rect 6196 4128 6224 4168
rect 7098 4156 7104 4168
rect 7156 4156 7162 4208
rect 6362 4128 6368 4140
rect 5644 4100 6224 4128
rect 6323 4100 6368 4128
rect 1486 4020 1492 4072
rect 1544 4060 1550 4072
rect 1653 4063 1711 4069
rect 1653 4060 1665 4063
rect 1544 4032 1665 4060
rect 1544 4020 1550 4032
rect 1653 4029 1665 4032
rect 1699 4029 1711 4063
rect 1653 4023 1711 4029
rect 2958 4020 2964 4072
rect 3016 4060 3022 4072
rect 3125 4063 3183 4069
rect 3125 4060 3137 4063
rect 3016 4032 3137 4060
rect 3016 4020 3022 4032
rect 3125 4029 3137 4032
rect 3171 4029 3183 4063
rect 3125 4023 3183 4029
rect 4154 4020 4160 4072
rect 4212 4060 4218 4072
rect 4341 4063 4399 4069
rect 4341 4060 4353 4063
rect 4212 4032 4353 4060
rect 4212 4020 4218 4032
rect 4341 4029 4353 4032
rect 4387 4060 4399 4063
rect 4430 4060 4436 4072
rect 4387 4032 4436 4060
rect 4387 4029 4399 4032
rect 4341 4023 4399 4029
rect 4430 4020 4436 4032
rect 4488 4020 4494 4072
rect 4608 4063 4666 4069
rect 4608 4029 4620 4063
rect 4654 4060 4666 4063
rect 5166 4060 5172 4072
rect 4654 4032 5172 4060
rect 4654 4029 4666 4032
rect 4608 4023 4666 4029
rect 5166 4020 5172 4032
rect 5224 4060 5230 4072
rect 5644 4060 5672 4100
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 7282 4128 7288 4140
rect 7243 4100 7288 4128
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 7484 4137 7512 4236
rect 13630 4224 13636 4236
rect 13688 4224 13694 4276
rect 14642 4264 14648 4276
rect 14476 4236 14648 4264
rect 9125 4199 9183 4205
rect 9125 4165 9137 4199
rect 9171 4196 9183 4199
rect 9490 4196 9496 4208
rect 9171 4168 9496 4196
rect 9171 4165 9183 4168
rect 9125 4159 9183 4165
rect 9490 4156 9496 4168
rect 9548 4156 9554 4208
rect 9674 4156 9680 4208
rect 9732 4196 9738 4208
rect 9769 4199 9827 4205
rect 9769 4196 9781 4199
rect 9732 4168 9781 4196
rect 9732 4156 9738 4168
rect 9769 4165 9781 4168
rect 9815 4165 9827 4199
rect 10686 4196 10692 4208
rect 9769 4159 9827 4165
rect 10244 4168 10692 4196
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4097 7527 4131
rect 7469 4091 7527 4097
rect 7650 4088 7656 4140
rect 7708 4128 7714 4140
rect 7745 4131 7803 4137
rect 7745 4128 7757 4131
rect 7708 4100 7757 4128
rect 7708 4088 7714 4100
rect 7745 4097 7757 4100
rect 7791 4097 7803 4131
rect 10244 4128 10272 4168
rect 10686 4156 10692 4168
rect 10744 4156 10750 4208
rect 11422 4196 11428 4208
rect 10796 4168 11428 4196
rect 7745 4091 7803 4097
rect 8772 4100 10272 4128
rect 5224 4032 5672 4060
rect 5224 4020 5230 4032
rect 5718 4020 5724 4072
rect 5776 4060 5782 4072
rect 7006 4060 7012 4072
rect 5776 4032 7012 4060
rect 5776 4020 5782 4032
rect 7006 4020 7012 4032
rect 7064 4020 7070 4072
rect 7098 4020 7104 4072
rect 7156 4060 7162 4072
rect 8001 4063 8059 4069
rect 8001 4060 8013 4063
rect 7156 4032 8013 4060
rect 7156 4020 7162 4032
rect 8001 4029 8013 4032
rect 8047 4029 8059 4063
rect 8772 4060 8800 4100
rect 10318 4088 10324 4140
rect 10376 4128 10382 4140
rect 10505 4131 10563 4137
rect 10505 4128 10517 4131
rect 10376 4100 10517 4128
rect 10376 4088 10382 4100
rect 10505 4097 10517 4100
rect 10551 4097 10563 4131
rect 10505 4091 10563 4097
rect 9214 4060 9220 4072
rect 8001 4023 8059 4029
rect 8404 4032 8800 4060
rect 9175 4032 9220 4060
rect 5074 3952 5080 4004
rect 5132 3992 5138 4004
rect 6273 3995 6331 4001
rect 6273 3992 6285 3995
rect 5132 3964 6285 3992
rect 5132 3952 5138 3964
rect 6273 3961 6285 3964
rect 6319 3961 6331 3995
rect 6273 3955 6331 3961
rect 7193 3995 7251 4001
rect 7193 3961 7205 3995
rect 7239 3992 7251 3995
rect 8404 3992 8432 4032
rect 9214 4020 9220 4032
rect 9272 4020 9278 4072
rect 9769 4063 9827 4069
rect 9769 4060 9781 4063
rect 9416 4032 9781 4060
rect 7239 3964 8432 3992
rect 7239 3961 7251 3964
rect 7193 3955 7251 3961
rect 8478 3952 8484 4004
rect 8536 3992 8542 4004
rect 9416 3992 9444 4032
rect 9769 4029 9781 4032
rect 9815 4029 9827 4063
rect 10796 4060 10824 4168
rect 11422 4156 11428 4168
rect 11480 4156 11486 4208
rect 11606 4156 11612 4208
rect 11664 4196 11670 4208
rect 11664 4168 11836 4196
rect 11664 4156 11670 4168
rect 11330 4128 11336 4140
rect 11291 4100 11336 4128
rect 11330 4088 11336 4100
rect 11388 4088 11394 4140
rect 11514 4088 11520 4140
rect 11572 4088 11578 4140
rect 11532 4060 11560 4088
rect 9769 4023 9827 4029
rect 9876 4032 10824 4060
rect 11348 4032 11560 4060
rect 11640 4063 11698 4069
rect 8536 3964 9444 3992
rect 8536 3952 8542 3964
rect 9490 3952 9496 4004
rect 9548 3992 9554 4004
rect 9548 3964 9593 3992
rect 9548 3952 9554 3964
rect 2777 3927 2835 3933
rect 2777 3893 2789 3927
rect 2823 3924 2835 3927
rect 3142 3924 3148 3936
rect 2823 3896 3148 3924
rect 2823 3893 2835 3896
rect 2777 3887 2835 3893
rect 3142 3884 3148 3896
rect 3200 3884 3206 3936
rect 3786 3884 3792 3936
rect 3844 3924 3850 3936
rect 4249 3927 4307 3933
rect 4249 3924 4261 3927
rect 3844 3896 4261 3924
rect 3844 3884 3850 3896
rect 4249 3893 4261 3896
rect 4295 3893 4307 3927
rect 4249 3887 4307 3893
rect 4338 3884 4344 3936
rect 4396 3924 4402 3936
rect 5534 3924 5540 3936
rect 4396 3896 5540 3924
rect 4396 3884 4402 3896
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 5813 3927 5871 3933
rect 5813 3893 5825 3927
rect 5859 3924 5871 3927
rect 6086 3924 6092 3936
rect 5859 3896 6092 3924
rect 5859 3893 5871 3896
rect 5813 3887 5871 3893
rect 6086 3884 6092 3896
rect 6144 3884 6150 3936
rect 6178 3884 6184 3936
rect 6236 3924 6242 3936
rect 6825 3927 6883 3933
rect 6236 3896 6281 3924
rect 6236 3884 6242 3896
rect 6825 3893 6837 3927
rect 6871 3924 6883 3927
rect 9876 3924 9904 4032
rect 10042 3952 10048 4004
rect 10100 3992 10106 4004
rect 10413 3995 10471 4001
rect 10413 3992 10425 3995
rect 10100 3964 10425 3992
rect 10100 3952 10106 3964
rect 10413 3961 10425 3964
rect 10459 3992 10471 3995
rect 11054 3992 11060 4004
rect 10459 3964 11060 3992
rect 10459 3961 10471 3964
rect 10413 3955 10471 3961
rect 11054 3952 11060 3964
rect 11112 3952 11118 4004
rect 11241 3995 11299 4001
rect 11241 3961 11253 3995
rect 11287 3992 11299 3995
rect 11348 3992 11376 4032
rect 11640 4029 11652 4063
rect 11686 4060 11698 4063
rect 11808 4060 11836 4168
rect 11974 4156 11980 4208
rect 12032 4196 12038 4208
rect 12342 4196 12348 4208
rect 12032 4168 12348 4196
rect 12032 4156 12038 4168
rect 12342 4156 12348 4168
rect 12400 4156 12406 4208
rect 12526 4156 12532 4208
rect 12584 4196 12590 4208
rect 14274 4196 14280 4208
rect 12584 4168 14280 4196
rect 12584 4156 12590 4168
rect 14274 4156 14280 4168
rect 14332 4156 14338 4208
rect 14476 4137 14504 4236
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 15841 4267 15899 4273
rect 15841 4233 15853 4267
rect 15887 4264 15899 4267
rect 16482 4264 16488 4276
rect 15887 4236 16488 4264
rect 15887 4233 15899 4236
rect 15841 4227 15899 4233
rect 16482 4224 16488 4236
rect 16540 4224 16546 4276
rect 16022 4196 16028 4208
rect 15488 4168 16028 4196
rect 14461 4131 14519 4137
rect 14461 4097 14473 4131
rect 14507 4097 14519 4131
rect 14461 4091 14519 4097
rect 11686 4032 11836 4060
rect 11885 4063 11943 4069
rect 11686 4029 11698 4032
rect 11640 4023 11698 4029
rect 11885 4029 11897 4063
rect 11931 4060 11943 4063
rect 12250 4060 12256 4072
rect 11931 4032 12256 4060
rect 11931 4029 11943 4032
rect 11885 4023 11943 4029
rect 12250 4020 12256 4032
rect 12308 4020 12314 4072
rect 12529 4063 12587 4069
rect 12529 4029 12541 4063
rect 12575 4060 12587 4063
rect 13354 4060 13360 4072
rect 12575 4032 13360 4060
rect 12575 4029 12587 4032
rect 12529 4023 12587 4029
rect 13354 4020 13360 4032
rect 13412 4020 13418 4072
rect 14090 4020 14096 4072
rect 14148 4060 14154 4072
rect 14550 4060 14556 4072
rect 14148 4032 14556 4060
rect 14148 4020 14154 4032
rect 14550 4020 14556 4032
rect 14608 4020 14614 4072
rect 14728 4063 14786 4069
rect 14728 4029 14740 4063
rect 14774 4060 14786 4063
rect 15488 4060 15516 4168
rect 16022 4156 16028 4168
rect 16080 4196 16086 4208
rect 16080 4168 20208 4196
rect 16080 4156 16086 4168
rect 16298 4088 16304 4140
rect 16356 4128 16362 4140
rect 18506 4128 18512 4140
rect 16356 4100 16804 4128
rect 18467 4100 18512 4128
rect 16356 4088 16362 4100
rect 16669 4063 16727 4069
rect 16669 4060 16681 4063
rect 14774 4032 15516 4060
rect 15580 4032 16681 4060
rect 14774 4029 14786 4032
rect 14728 4023 14786 4029
rect 11287 3964 11376 3992
rect 11287 3961 11299 3964
rect 11241 3955 11299 3961
rect 11422 3952 11428 4004
rect 11480 3992 11486 4004
rect 13906 3992 13912 4004
rect 11480 3964 13912 3992
rect 11480 3952 11486 3964
rect 13906 3952 13912 3964
rect 13964 3952 13970 4004
rect 14274 3952 14280 4004
rect 14332 3992 14338 4004
rect 15580 3992 15608 4032
rect 16669 4029 16681 4032
rect 16715 4029 16727 4063
rect 16776 4060 16804 4100
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 18690 4128 18696 4140
rect 18651 4100 18696 4128
rect 18690 4088 18696 4100
rect 18748 4088 18754 4140
rect 19058 4088 19064 4140
rect 19116 4128 19122 4140
rect 20070 4128 20076 4140
rect 19116 4100 19748 4128
rect 20031 4100 20076 4128
rect 19116 4088 19122 4100
rect 19720 4060 19748 4100
rect 20070 4088 20076 4100
rect 20128 4088 20134 4140
rect 20180 4137 20208 4168
rect 20165 4131 20223 4137
rect 20165 4097 20177 4131
rect 20211 4097 20223 4131
rect 20165 4091 20223 4097
rect 19981 4063 20039 4069
rect 19981 4060 19993 4063
rect 16776 4032 19196 4060
rect 19720 4032 19993 4060
rect 16669 4023 16727 4029
rect 14332 3964 15608 3992
rect 14332 3952 14338 3964
rect 6871 3896 9904 3924
rect 9953 3927 10011 3933
rect 6871 3893 6883 3896
rect 6825 3887 6883 3893
rect 9953 3893 9965 3927
rect 9999 3924 10011 3927
rect 10134 3924 10140 3936
rect 9999 3896 10140 3924
rect 9999 3893 10011 3896
rect 9953 3887 10011 3893
rect 10134 3884 10140 3896
rect 10192 3884 10198 3936
rect 10226 3884 10232 3936
rect 10284 3924 10290 3936
rect 10321 3927 10379 3933
rect 10321 3924 10333 3927
rect 10284 3896 10333 3924
rect 10284 3884 10290 3896
rect 10321 3893 10333 3896
rect 10367 3893 10379 3927
rect 10321 3887 10379 3893
rect 10781 3927 10839 3933
rect 10781 3893 10793 3927
rect 10827 3924 10839 3927
rect 10870 3924 10876 3936
rect 10827 3896 10876 3924
rect 10827 3893 10839 3896
rect 10781 3887 10839 3893
rect 10870 3884 10876 3896
rect 10928 3884 10934 3936
rect 11149 3927 11207 3933
rect 11149 3893 11161 3927
rect 11195 3924 11207 3927
rect 12526 3924 12532 3936
rect 11195 3896 12532 3924
rect 11195 3893 11207 3896
rect 11149 3887 11207 3893
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 12710 3924 12716 3936
rect 12671 3896 12716 3924
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 13446 3884 13452 3936
rect 13504 3924 13510 3936
rect 16853 3927 16911 3933
rect 16853 3924 16865 3927
rect 13504 3896 16865 3924
rect 13504 3884 13510 3896
rect 16853 3893 16865 3896
rect 16899 3893 16911 3927
rect 16853 3887 16911 3893
rect 18049 3927 18107 3933
rect 18049 3893 18061 3927
rect 18095 3924 18107 3927
rect 18138 3924 18144 3936
rect 18095 3896 18144 3924
rect 18095 3893 18107 3896
rect 18049 3887 18107 3893
rect 18138 3884 18144 3896
rect 18196 3884 18202 3936
rect 18230 3884 18236 3936
rect 18288 3924 18294 3936
rect 18417 3927 18475 3933
rect 18417 3924 18429 3927
rect 18288 3896 18429 3924
rect 18288 3884 18294 3896
rect 18417 3893 18429 3896
rect 18463 3893 18475 3927
rect 19168 3924 19196 4032
rect 19981 4029 19993 4032
rect 20027 4029 20039 4063
rect 19981 4023 20039 4029
rect 19613 3927 19671 3933
rect 19613 3924 19625 3927
rect 19168 3896 19625 3924
rect 18417 3887 18475 3893
rect 19613 3893 19625 3896
rect 19659 3893 19671 3927
rect 19613 3887 19671 3893
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 2590 3680 2596 3732
rect 2648 3720 2654 3732
rect 2648 3692 6488 3720
rect 2648 3680 2654 3692
rect 1118 3612 1124 3664
rect 1176 3652 1182 3664
rect 1642 3655 1700 3661
rect 1642 3652 1654 3655
rect 1176 3624 1654 3652
rect 1176 3612 1182 3624
rect 1642 3621 1654 3624
rect 1688 3621 1700 3655
rect 1642 3615 1700 3621
rect 2038 3612 2044 3664
rect 2096 3652 2102 3664
rect 4332 3655 4390 3661
rect 2096 3624 2268 3652
rect 2096 3612 2102 3624
rect 1394 3544 1400 3596
rect 1452 3584 1458 3596
rect 1946 3584 1952 3596
rect 1452 3556 1952 3584
rect 1452 3544 1458 3556
rect 1946 3544 1952 3556
rect 2004 3544 2010 3596
rect 2240 3584 2268 3624
rect 4332 3621 4344 3655
rect 4378 3652 4390 3655
rect 4522 3652 4528 3664
rect 4378 3624 4528 3652
rect 4378 3621 4390 3624
rect 4332 3615 4390 3621
rect 4522 3612 4528 3624
rect 4580 3612 4586 3664
rect 5350 3612 5356 3664
rect 5408 3652 5414 3664
rect 5718 3652 5724 3664
rect 5408 3624 5724 3652
rect 5408 3612 5414 3624
rect 5718 3612 5724 3624
rect 5776 3612 5782 3664
rect 6080 3655 6138 3661
rect 6080 3621 6092 3655
rect 6126 3652 6138 3655
rect 6362 3652 6368 3664
rect 6126 3624 6368 3652
rect 6126 3621 6138 3624
rect 6080 3615 6138 3621
rect 6362 3612 6368 3624
rect 6420 3612 6426 3664
rect 6460 3652 6488 3692
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 7193 3723 7251 3729
rect 7193 3720 7205 3723
rect 7156 3692 7205 3720
rect 7156 3680 7162 3692
rect 7193 3689 7205 3692
rect 7239 3689 7251 3723
rect 7193 3683 7251 3689
rect 7282 3680 7288 3732
rect 7340 3720 7346 3732
rect 7469 3723 7527 3729
rect 7469 3720 7481 3723
rect 7340 3692 7481 3720
rect 7340 3680 7346 3692
rect 7469 3689 7481 3692
rect 7515 3689 7527 3723
rect 7469 3683 7527 3689
rect 7653 3723 7711 3729
rect 7653 3689 7665 3723
rect 7699 3720 7711 3723
rect 7742 3720 7748 3732
rect 7699 3692 7748 3720
rect 7699 3689 7711 3692
rect 7653 3683 7711 3689
rect 7742 3680 7748 3692
rect 7800 3680 7806 3732
rect 8113 3723 8171 3729
rect 8113 3689 8125 3723
rect 8159 3720 8171 3723
rect 8386 3720 8392 3732
rect 8159 3692 8392 3720
rect 8159 3689 8171 3692
rect 8113 3683 8171 3689
rect 8386 3680 8392 3692
rect 8444 3680 8450 3732
rect 9217 3723 9275 3729
rect 9217 3689 9229 3723
rect 9263 3720 9275 3723
rect 9309 3723 9367 3729
rect 9309 3720 9321 3723
rect 9263 3692 9321 3720
rect 9263 3689 9275 3692
rect 9217 3683 9275 3689
rect 9309 3689 9321 3692
rect 9355 3720 9367 3723
rect 9582 3720 9588 3732
rect 9355 3692 9588 3720
rect 9355 3689 9367 3692
rect 9309 3683 9367 3689
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 10045 3723 10103 3729
rect 10045 3720 10057 3723
rect 10008 3692 10057 3720
rect 10008 3680 10014 3692
rect 10045 3689 10057 3692
rect 10091 3689 10103 3723
rect 11606 3720 11612 3732
rect 10045 3683 10103 3689
rect 10612 3692 11612 3720
rect 6460 3624 7246 3652
rect 2866 3584 2872 3596
rect 2240 3556 2872 3584
rect 2866 3544 2872 3556
rect 2924 3544 2930 3596
rect 3237 3587 3295 3593
rect 3237 3553 3249 3587
rect 3283 3584 3295 3587
rect 6546 3584 6552 3596
rect 3283 3556 6552 3584
rect 3283 3553 3295 3556
rect 3237 3547 3295 3553
rect 6546 3544 6552 3556
rect 6604 3544 6610 3596
rect 3326 3516 3332 3528
rect 3287 3488 3332 3516
rect 3326 3476 3332 3488
rect 3384 3476 3390 3528
rect 3418 3476 3424 3528
rect 3476 3516 3482 3528
rect 5810 3516 5816 3528
rect 3476 3488 3521 3516
rect 5771 3488 5816 3516
rect 3476 3476 3482 3488
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 2774 3448 2780 3460
rect 2735 3420 2780 3448
rect 2774 3408 2780 3420
rect 2832 3408 2838 3460
rect 5718 3448 5724 3460
rect 5368 3420 5724 3448
rect 2869 3383 2927 3389
rect 2869 3349 2881 3383
rect 2915 3380 2927 3383
rect 5368 3380 5396 3420
rect 5718 3408 5724 3420
rect 5776 3408 5782 3460
rect 2915 3352 5396 3380
rect 2915 3349 2927 3352
rect 2869 3343 2927 3349
rect 5442 3340 5448 3392
rect 5500 3380 5506 3392
rect 7218 3380 7246 3624
rect 8202 3612 8208 3664
rect 8260 3652 8266 3664
rect 10612 3652 10640 3692
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 11701 3723 11759 3729
rect 11701 3689 11713 3723
rect 11747 3720 11759 3723
rect 12250 3720 12256 3732
rect 11747 3692 12256 3720
rect 11747 3689 11759 3692
rect 11701 3683 11759 3689
rect 12250 3680 12256 3692
rect 12308 3680 12314 3732
rect 16114 3720 16120 3732
rect 12544 3692 16120 3720
rect 8260 3624 10640 3652
rect 10873 3655 10931 3661
rect 8260 3612 8266 3624
rect 10873 3621 10885 3655
rect 10919 3652 10931 3655
rect 11793 3655 11851 3661
rect 10919 3624 11744 3652
rect 10919 3621 10931 3624
rect 10873 3615 10931 3621
rect 7282 3544 7288 3596
rect 7340 3584 7346 3596
rect 8021 3587 8079 3593
rect 8021 3584 8033 3587
rect 7340 3556 8033 3584
rect 7340 3544 7346 3556
rect 8021 3553 8033 3556
rect 8067 3553 8079 3587
rect 8021 3547 8079 3553
rect 8846 3544 8852 3596
rect 8904 3584 8910 3596
rect 10226 3584 10232 3596
rect 8904 3556 10232 3584
rect 8904 3544 8910 3556
rect 10226 3544 10232 3556
rect 10284 3544 10290 3596
rect 11606 3584 11612 3596
rect 10336 3556 11612 3584
rect 7374 3476 7380 3528
rect 7432 3516 7438 3528
rect 8110 3516 8116 3528
rect 7432 3488 8116 3516
rect 7432 3476 7438 3488
rect 8110 3476 8116 3488
rect 8168 3516 8174 3528
rect 8205 3519 8263 3525
rect 8205 3516 8217 3519
rect 8168 3488 8217 3516
rect 8168 3476 8174 3488
rect 8205 3485 8217 3488
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 8662 3476 8668 3528
rect 8720 3516 8726 3528
rect 9858 3516 9864 3528
rect 8720 3488 9864 3516
rect 8720 3476 8726 3488
rect 9858 3476 9864 3488
rect 9916 3516 9922 3528
rect 10336 3525 10364 3556
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 11716 3584 11744 3624
rect 11793 3621 11805 3655
rect 11839 3652 11851 3655
rect 12544 3652 12572 3692
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 17589 3723 17647 3729
rect 17589 3689 17601 3723
rect 17635 3720 17647 3723
rect 18506 3720 18512 3732
rect 17635 3692 18512 3720
rect 17635 3689 17647 3692
rect 17589 3683 17647 3689
rect 18506 3680 18512 3692
rect 18564 3680 18570 3732
rect 15194 3652 15200 3664
rect 11839 3624 12572 3652
rect 13372 3624 15200 3652
rect 11839 3621 11851 3624
rect 11793 3615 11851 3621
rect 11974 3584 11980 3596
rect 11716 3556 11980 3584
rect 11974 3544 11980 3556
rect 12032 3544 12038 3596
rect 12158 3584 12164 3596
rect 12119 3556 12164 3584
rect 12158 3544 12164 3556
rect 12216 3544 12222 3596
rect 12526 3584 12532 3596
rect 12487 3556 12532 3584
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 12802 3544 12808 3596
rect 12860 3584 12866 3596
rect 12860 3556 12905 3584
rect 12860 3544 12866 3556
rect 10137 3519 10195 3525
rect 10137 3516 10149 3519
rect 9916 3488 10149 3516
rect 9916 3476 9922 3488
rect 10137 3485 10149 3488
rect 10183 3485 10195 3519
rect 10137 3479 10195 3485
rect 10321 3519 10379 3525
rect 10321 3485 10333 3519
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 10502 3476 10508 3528
rect 10560 3516 10566 3528
rect 10965 3519 11023 3525
rect 10965 3516 10977 3519
rect 10560 3488 10977 3516
rect 10560 3476 10566 3488
rect 10965 3485 10977 3488
rect 11011 3485 11023 3519
rect 10965 3479 11023 3485
rect 11057 3519 11115 3525
rect 11057 3485 11069 3519
rect 11103 3485 11115 3519
rect 11057 3479 11115 3485
rect 7558 3408 7564 3460
rect 7616 3448 7622 3460
rect 8938 3448 8944 3460
rect 7616 3420 8944 3448
rect 7616 3408 7622 3420
rect 8938 3408 8944 3420
rect 8996 3408 9002 3460
rect 9582 3408 9588 3460
rect 9640 3448 9646 3460
rect 9677 3451 9735 3457
rect 9677 3448 9689 3451
rect 9640 3420 9689 3448
rect 9640 3408 9646 3420
rect 9677 3417 9689 3420
rect 9723 3417 9735 3451
rect 9677 3411 9735 3417
rect 10870 3408 10876 3460
rect 10928 3448 10934 3460
rect 11072 3448 11100 3479
rect 11790 3476 11796 3528
rect 11848 3516 11854 3528
rect 11885 3519 11943 3525
rect 11885 3516 11897 3519
rect 11848 3488 11897 3516
rect 11848 3476 11854 3488
rect 11885 3485 11897 3488
rect 11931 3485 11943 3519
rect 11885 3479 11943 3485
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 12710 3516 12716 3528
rect 12400 3488 12716 3516
rect 12400 3476 12406 3488
rect 12710 3476 12716 3488
rect 12768 3476 12774 3528
rect 10928 3420 11100 3448
rect 11333 3451 11391 3457
rect 10928 3408 10934 3420
rect 11333 3417 11345 3451
rect 11379 3448 11391 3451
rect 13372 3448 13400 3624
rect 15194 3612 15200 3624
rect 15252 3612 15258 3664
rect 15378 3612 15384 3664
rect 15436 3652 15442 3664
rect 17957 3655 18015 3661
rect 17957 3652 17969 3655
rect 15436 3624 17969 3652
rect 15436 3612 15442 3624
rect 17957 3621 17969 3624
rect 18003 3621 18015 3655
rect 17957 3615 18015 3621
rect 18046 3612 18052 3664
rect 18104 3652 18110 3664
rect 19702 3652 19708 3664
rect 18104 3624 19708 3652
rect 18104 3612 18110 3624
rect 19702 3612 19708 3624
rect 19760 3612 19766 3664
rect 14090 3584 14096 3596
rect 14051 3556 14096 3584
rect 14090 3544 14096 3556
rect 14148 3544 14154 3596
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3553 15347 3587
rect 15289 3547 15347 3553
rect 16485 3587 16543 3593
rect 16485 3553 16497 3587
rect 16531 3584 16543 3587
rect 16942 3584 16948 3596
rect 16531 3556 16948 3584
rect 16531 3553 16543 3556
rect 16485 3547 16543 3553
rect 13722 3476 13728 3528
rect 13780 3516 13786 3528
rect 15304 3516 15332 3547
rect 16942 3544 16948 3556
rect 17000 3544 17006 3596
rect 19334 3544 19340 3596
rect 19392 3584 19398 3596
rect 19613 3587 19671 3593
rect 19613 3584 19625 3587
rect 19392 3556 19625 3584
rect 19392 3544 19398 3556
rect 19613 3553 19625 3556
rect 19659 3553 19671 3587
rect 19613 3547 19671 3553
rect 13780 3488 15332 3516
rect 13780 3476 13786 3488
rect 17954 3476 17960 3528
rect 18012 3516 18018 3528
rect 18049 3519 18107 3525
rect 18049 3516 18061 3519
rect 18012 3488 18061 3516
rect 18012 3476 18018 3488
rect 18049 3485 18061 3488
rect 18095 3485 18107 3519
rect 18049 3479 18107 3485
rect 18138 3476 18144 3528
rect 18196 3516 18202 3528
rect 18782 3516 18788 3528
rect 18196 3488 18788 3516
rect 18196 3476 18202 3488
rect 18782 3476 18788 3488
rect 18840 3476 18846 3528
rect 14090 3448 14096 3460
rect 11379 3420 13400 3448
rect 13924 3420 14096 3448
rect 11379 3417 11391 3420
rect 11333 3411 11391 3417
rect 8202 3380 8208 3392
rect 5500 3352 5545 3380
rect 7218 3352 8208 3380
rect 5500 3340 5506 3352
rect 8202 3340 8208 3352
rect 8260 3340 8266 3392
rect 8754 3340 8760 3392
rect 8812 3380 8818 3392
rect 9950 3380 9956 3392
rect 8812 3352 9956 3380
rect 8812 3340 8818 3352
rect 9950 3340 9956 3352
rect 10008 3340 10014 3392
rect 10505 3383 10563 3389
rect 10505 3349 10517 3383
rect 10551 3380 10563 3383
rect 12158 3380 12164 3392
rect 10551 3352 12164 3380
rect 10551 3349 10563 3352
rect 10505 3343 10563 3349
rect 12158 3340 12164 3352
rect 12216 3340 12222 3392
rect 12345 3383 12403 3389
rect 12345 3349 12357 3383
rect 12391 3380 12403 3383
rect 13924 3380 13952 3420
rect 14090 3408 14096 3420
rect 14148 3408 14154 3460
rect 12391 3352 13952 3380
rect 12391 3349 12403 3352
rect 12345 3343 12403 3349
rect 13998 3340 14004 3392
rect 14056 3380 14062 3392
rect 14277 3383 14335 3389
rect 14277 3380 14289 3383
rect 14056 3352 14289 3380
rect 14056 3340 14062 3352
rect 14277 3349 14289 3352
rect 14323 3349 14335 3383
rect 14277 3343 14335 3349
rect 15473 3383 15531 3389
rect 15473 3349 15485 3383
rect 15519 3380 15531 3383
rect 16114 3380 16120 3392
rect 15519 3352 16120 3380
rect 15519 3349 15531 3352
rect 15473 3343 15531 3349
rect 16114 3340 16120 3352
rect 16172 3340 16178 3392
rect 16669 3383 16727 3389
rect 16669 3349 16681 3383
rect 16715 3380 16727 3383
rect 17494 3380 17500 3392
rect 16715 3352 17500 3380
rect 16715 3349 16727 3352
rect 16669 3343 16727 3349
rect 17494 3340 17500 3352
rect 17552 3340 17558 3392
rect 19797 3383 19855 3389
rect 19797 3349 19809 3383
rect 19843 3380 19855 3383
rect 20346 3380 20352 3392
rect 19843 3352 20352 3380
rect 19843 3349 19855 3352
rect 19797 3343 19855 3349
rect 20346 3340 20352 3352
rect 20404 3340 20410 3392
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 3234 3136 3240 3188
rect 3292 3176 3298 3188
rect 5905 3179 5963 3185
rect 3292 3148 3924 3176
rect 3292 3136 3298 3148
rect 2498 3068 2504 3120
rect 2556 3108 2562 3120
rect 2777 3111 2835 3117
rect 2777 3108 2789 3111
rect 2556 3080 2789 3108
rect 2556 3068 2562 3080
rect 2777 3077 2789 3080
rect 2823 3077 2835 3111
rect 2777 3071 2835 3077
rect 3896 3040 3924 3148
rect 5905 3145 5917 3179
rect 5951 3176 5963 3179
rect 6086 3176 6092 3188
rect 5951 3148 6092 3176
rect 5951 3145 5963 3148
rect 5905 3139 5963 3145
rect 6086 3136 6092 3148
rect 6144 3176 6150 3188
rect 6362 3176 6368 3188
rect 6144 3148 6368 3176
rect 6144 3136 6150 3148
rect 6362 3136 6368 3148
rect 6420 3136 6426 3188
rect 7006 3136 7012 3188
rect 7064 3176 7070 3188
rect 8113 3179 8171 3185
rect 7064 3148 7246 3176
rect 7064 3136 7070 3148
rect 4249 3111 4307 3117
rect 4249 3077 4261 3111
rect 4295 3108 4307 3111
rect 4522 3108 4528 3120
rect 4295 3080 4528 3108
rect 4295 3077 4307 3080
rect 4249 3071 4307 3077
rect 4522 3068 4528 3080
rect 4580 3068 4586 3120
rect 7101 3111 7159 3117
rect 7101 3077 7113 3111
rect 7147 3077 7159 3111
rect 7101 3071 7159 3077
rect 6270 3040 6276 3052
rect 3896 3012 4651 3040
rect 1664 2975 1722 2981
rect 1664 2941 1676 2975
rect 1710 2972 1722 2975
rect 2222 2972 2228 2984
rect 1710 2944 2228 2972
rect 1710 2941 1722 2944
rect 1664 2935 1722 2941
rect 2222 2932 2228 2944
rect 2280 2932 2286 2984
rect 3136 2975 3194 2981
rect 3136 2941 3148 2975
rect 3182 2972 3194 2975
rect 3510 2972 3516 2984
rect 3182 2944 3516 2972
rect 3182 2941 3194 2944
rect 3136 2935 3194 2941
rect 3510 2932 3516 2944
rect 3568 2932 3574 2984
rect 4062 2932 4068 2984
rect 4120 2972 4126 2984
rect 4525 2975 4583 2981
rect 4525 2972 4537 2975
rect 4120 2944 4537 2972
rect 4120 2932 4126 2944
rect 4525 2941 4537 2944
rect 4571 2941 4583 2975
rect 4623 2972 4651 3012
rect 5552 3012 6276 3040
rect 5552 2972 5580 3012
rect 6270 3000 6276 3012
rect 6328 3000 6334 3052
rect 4623 2944 5580 2972
rect 6181 2975 6239 2981
rect 4525 2935 4583 2941
rect 6181 2941 6193 2975
rect 6227 2972 6239 2975
rect 7116 2972 7144 3071
rect 7218 3040 7246 3148
rect 8113 3145 8125 3179
rect 8159 3176 8171 3179
rect 8202 3176 8208 3188
rect 8159 3148 8208 3176
rect 8159 3145 8171 3148
rect 8113 3139 8171 3145
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 9582 3176 9588 3188
rect 8312 3148 9588 3176
rect 8018 3068 8024 3120
rect 8076 3108 8082 3120
rect 8312 3108 8340 3148
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 9858 3136 9864 3188
rect 9916 3176 9922 3188
rect 10042 3176 10048 3188
rect 9916 3148 10048 3176
rect 9916 3136 9922 3148
rect 10042 3136 10048 3148
rect 10100 3136 10106 3188
rect 10226 3136 10232 3188
rect 10284 3176 10290 3188
rect 11333 3179 11391 3185
rect 10284 3148 11100 3176
rect 10284 3136 10290 3148
rect 8076 3080 8340 3108
rect 8076 3068 8082 3080
rect 9306 3068 9312 3120
rect 9364 3108 9370 3120
rect 10870 3108 10876 3120
rect 9364 3080 10876 3108
rect 9364 3068 9370 3080
rect 10870 3068 10876 3080
rect 10928 3068 10934 3120
rect 11072 3108 11100 3148
rect 11333 3145 11345 3179
rect 11379 3176 11391 3179
rect 12342 3176 12348 3188
rect 11379 3148 12348 3176
rect 11379 3145 11391 3148
rect 11333 3139 11391 3145
rect 12342 3136 12348 3148
rect 12400 3136 12406 3188
rect 12437 3179 12495 3185
rect 12437 3145 12449 3179
rect 12483 3176 12495 3179
rect 13538 3176 13544 3188
rect 12483 3148 13544 3176
rect 12483 3145 12495 3148
rect 12437 3139 12495 3145
rect 13538 3136 13544 3148
rect 13596 3136 13602 3188
rect 17310 3136 17316 3188
rect 17368 3176 17374 3188
rect 17368 3148 19472 3176
rect 17368 3136 17374 3148
rect 11514 3108 11520 3120
rect 11072 3080 11520 3108
rect 11514 3068 11520 3080
rect 11572 3068 11578 3120
rect 11698 3068 11704 3120
rect 11756 3108 11762 3120
rect 11756 3080 12388 3108
rect 11756 3068 11762 3080
rect 12360 3052 12388 3080
rect 12728 3080 15608 3108
rect 7653 3043 7711 3049
rect 7653 3040 7665 3043
rect 7218 3012 7665 3040
rect 7653 3009 7665 3012
rect 7699 3009 7711 3043
rect 10226 3040 10232 3052
rect 7653 3003 7711 3009
rect 7944 3012 8432 3040
rect 6227 2944 7144 2972
rect 6227 2941 6239 2944
rect 6181 2935 6239 2941
rect 7466 2932 7472 2984
rect 7524 2972 7530 2984
rect 7944 2981 7972 3012
rect 7561 2975 7619 2981
rect 7561 2972 7573 2975
rect 7524 2944 7573 2972
rect 7524 2932 7530 2944
rect 7561 2941 7573 2944
rect 7607 2941 7619 2975
rect 7561 2935 7619 2941
rect 7929 2975 7987 2981
rect 7929 2941 7941 2975
rect 7975 2941 7987 2975
rect 7929 2935 7987 2941
rect 8018 2932 8024 2984
rect 8076 2972 8082 2984
rect 8297 2975 8355 2981
rect 8297 2972 8309 2975
rect 8076 2944 8309 2972
rect 8076 2932 8082 2944
rect 8297 2941 8309 2944
rect 8343 2941 8355 2975
rect 8404 2972 8432 3012
rect 9692 3012 10232 3040
rect 8846 2972 8852 2984
rect 8404 2944 8852 2972
rect 8297 2935 8355 2941
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 9692 2972 9720 3012
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 10318 3000 10324 3052
rect 10376 3040 10382 3052
rect 11103 3043 11161 3049
rect 11103 3040 11115 3043
rect 10376 3012 11115 3040
rect 10376 3000 10382 3012
rect 11103 3009 11115 3012
rect 11149 3009 11161 3043
rect 11882 3040 11888 3052
rect 11843 3012 11888 3040
rect 11103 3003 11161 3009
rect 11882 3000 11888 3012
rect 11940 3000 11946 3052
rect 12342 3000 12348 3052
rect 12400 3000 12406 3052
rect 8956 2944 9720 2972
rect 3418 2864 3424 2916
rect 3476 2904 3482 2916
rect 4770 2907 4828 2913
rect 4770 2904 4782 2907
rect 3476 2876 4782 2904
rect 3476 2864 3482 2876
rect 4770 2873 4782 2876
rect 4816 2904 4828 2907
rect 5258 2904 5264 2916
rect 4816 2876 5264 2904
rect 4816 2873 4828 2876
rect 4770 2867 4828 2873
rect 5258 2864 5264 2876
rect 5316 2864 5322 2916
rect 6457 2907 6515 2913
rect 6457 2873 6469 2907
rect 6503 2904 6515 2907
rect 8564 2907 8622 2913
rect 6503 2876 8524 2904
rect 6503 2873 6515 2876
rect 6457 2867 6515 2873
rect 5626 2796 5632 2848
rect 5684 2836 5690 2848
rect 7469 2839 7527 2845
rect 7469 2836 7481 2839
rect 5684 2808 7481 2836
rect 5684 2796 5690 2808
rect 7469 2805 7481 2808
rect 7515 2805 7527 2839
rect 8496 2836 8524 2876
rect 8564 2873 8576 2907
rect 8610 2904 8622 2907
rect 8754 2904 8760 2916
rect 8610 2876 8760 2904
rect 8610 2873 8622 2876
rect 8564 2867 8622 2873
rect 8754 2864 8760 2876
rect 8812 2864 8818 2916
rect 8956 2836 8984 2944
rect 9766 2932 9772 2984
rect 9824 2972 9830 2984
rect 9824 2944 9869 2972
rect 9824 2932 9830 2944
rect 10045 2907 10103 2913
rect 10045 2873 10057 2907
rect 10091 2904 10103 2907
rect 10410 2904 10416 2916
rect 10091 2876 10416 2904
rect 10091 2873 10103 2876
rect 10045 2867 10103 2873
rect 10410 2864 10416 2876
rect 10468 2864 10474 2916
rect 11164 2876 11560 2904
rect 8496 2808 8984 2836
rect 7469 2799 7527 2805
rect 9398 2796 9404 2848
rect 9456 2836 9462 2848
rect 9674 2836 9680 2848
rect 9456 2808 9680 2836
rect 9456 2796 9462 2808
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 9766 2796 9772 2848
rect 9824 2836 9830 2848
rect 10505 2839 10563 2845
rect 10505 2836 10517 2839
rect 9824 2808 10517 2836
rect 9824 2796 9830 2808
rect 10505 2805 10517 2808
rect 10551 2805 10563 2839
rect 10870 2836 10876 2848
rect 10831 2808 10876 2836
rect 10505 2799 10563 2805
rect 10870 2796 10876 2808
rect 10928 2796 10934 2848
rect 10965 2839 11023 2845
rect 10965 2805 10977 2839
rect 11011 2836 11023 2839
rect 11164 2836 11192 2876
rect 11011 2808 11192 2836
rect 11532 2836 11560 2876
rect 11606 2864 11612 2916
rect 11664 2904 11670 2916
rect 11701 2907 11759 2913
rect 11701 2904 11713 2907
rect 11664 2876 11713 2904
rect 11664 2864 11670 2876
rect 11701 2873 11713 2876
rect 11747 2873 11759 2907
rect 11701 2867 11759 2873
rect 11793 2907 11851 2913
rect 11793 2873 11805 2907
rect 11839 2904 11851 2907
rect 12434 2904 12440 2916
rect 11839 2876 12440 2904
rect 11839 2873 11851 2876
rect 11793 2867 11851 2873
rect 12434 2864 12440 2876
rect 12492 2864 12498 2916
rect 12728 2904 12756 3080
rect 13078 3040 13084 3052
rect 13039 3012 13084 3040
rect 13078 3000 13084 3012
rect 13136 3000 13142 3052
rect 14550 3040 14556 3052
rect 14511 3012 14556 3040
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 15580 3040 15608 3080
rect 15654 3068 15660 3120
rect 15712 3108 15718 3120
rect 19337 3111 19395 3117
rect 19337 3108 19349 3111
rect 15712 3080 19349 3108
rect 15712 3068 15718 3080
rect 19337 3077 19349 3080
rect 19383 3077 19395 3111
rect 19337 3071 19395 3077
rect 15930 3040 15936 3052
rect 15580 3012 15936 3040
rect 15930 3000 15936 3012
rect 15988 3000 15994 3052
rect 17126 3000 17132 3052
rect 17184 3040 17190 3052
rect 19444 3040 19472 3148
rect 20441 3043 20499 3049
rect 20441 3040 20453 3043
rect 17184 3012 18000 3040
rect 19444 3012 20453 3040
rect 17184 3000 17190 3012
rect 14366 2972 14372 2984
rect 14327 2944 14372 2972
rect 14366 2932 14372 2944
rect 14424 2932 14430 2984
rect 15562 2972 15568 2984
rect 15523 2944 15568 2972
rect 15562 2932 15568 2944
rect 15620 2932 15626 2984
rect 16666 2972 16672 2984
rect 16627 2944 16672 2972
rect 16666 2932 16672 2944
rect 16724 2932 16730 2984
rect 17972 2972 18000 3012
rect 20441 3009 20453 3012
rect 20487 3009 20499 3043
rect 20441 3003 20499 3009
rect 18037 2975 18095 2981
rect 18037 2972 18049 2975
rect 17972 2944 18049 2972
rect 18037 2941 18049 2944
rect 18083 2941 18095 2975
rect 18037 2935 18095 2941
rect 18874 2932 18880 2984
rect 18932 2972 18938 2984
rect 19153 2975 19211 2981
rect 19153 2972 19165 2975
rect 18932 2944 19165 2972
rect 18932 2932 18938 2944
rect 19153 2941 19165 2944
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 19518 2932 19524 2984
rect 19576 2972 19582 2984
rect 20257 2975 20315 2981
rect 20257 2972 20269 2975
rect 19576 2944 20269 2972
rect 19576 2932 19582 2944
rect 20257 2941 20269 2944
rect 20303 2941 20315 2975
rect 20257 2935 20315 2941
rect 12544 2876 12756 2904
rect 12805 2907 12863 2913
rect 12544 2836 12572 2876
rect 12805 2873 12817 2907
rect 12851 2904 12863 2907
rect 12851 2876 14044 2904
rect 12851 2873 12863 2876
rect 12805 2867 12863 2873
rect 11532 2808 12572 2836
rect 11011 2805 11023 2808
rect 10965 2799 11023 2805
rect 12618 2796 12624 2848
rect 12676 2836 12682 2848
rect 14016 2845 14044 2876
rect 15930 2864 15936 2916
rect 15988 2904 15994 2916
rect 19978 2904 19984 2916
rect 15988 2876 19984 2904
rect 15988 2864 15994 2876
rect 19978 2864 19984 2876
rect 20036 2904 20042 2916
rect 22646 2904 22652 2916
rect 20036 2876 22652 2904
rect 20036 2864 20042 2876
rect 22646 2864 22652 2876
rect 22704 2864 22710 2916
rect 12897 2839 12955 2845
rect 12897 2836 12909 2839
rect 12676 2808 12909 2836
rect 12676 2796 12682 2808
rect 12897 2805 12909 2808
rect 12943 2805 12955 2839
rect 12897 2799 12955 2805
rect 14001 2839 14059 2845
rect 14001 2805 14013 2839
rect 14047 2805 14059 2839
rect 14001 2799 14059 2805
rect 14458 2796 14464 2848
rect 14516 2836 14522 2848
rect 14516 2808 14561 2836
rect 14516 2796 14522 2808
rect 15194 2796 15200 2848
rect 15252 2836 15258 2848
rect 15749 2839 15807 2845
rect 15749 2836 15761 2839
rect 15252 2808 15761 2836
rect 15252 2796 15258 2808
rect 15749 2805 15761 2808
rect 15795 2805 15807 2839
rect 15749 2799 15807 2805
rect 16853 2839 16911 2845
rect 16853 2805 16865 2839
rect 16899 2836 16911 2839
rect 17034 2836 17040 2848
rect 16899 2808 17040 2836
rect 16899 2805 16911 2808
rect 16853 2799 16911 2805
rect 17034 2796 17040 2808
rect 17092 2796 17098 2848
rect 17954 2796 17960 2848
rect 18012 2836 18018 2848
rect 18233 2839 18291 2845
rect 18233 2836 18245 2839
rect 18012 2808 18245 2836
rect 18012 2796 18018 2808
rect 18233 2805 18245 2808
rect 18279 2805 18291 2839
rect 18233 2799 18291 2805
rect 20162 2796 20168 2848
rect 20220 2836 20226 2848
rect 22186 2836 22192 2848
rect 20220 2808 22192 2836
rect 20220 2796 20226 2808
rect 22186 2796 22192 2808
rect 22244 2796 22250 2848
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 2682 2592 2688 2644
rect 2740 2632 2746 2644
rect 5445 2635 5503 2641
rect 5445 2632 5457 2635
rect 2740 2604 5457 2632
rect 2740 2592 2746 2604
rect 5445 2601 5457 2604
rect 5491 2601 5503 2635
rect 5445 2595 5503 2601
rect 5537 2635 5595 2641
rect 5537 2601 5549 2635
rect 5583 2632 5595 2635
rect 5626 2632 5632 2644
rect 5583 2604 5632 2632
rect 5583 2601 5595 2604
rect 5537 2595 5595 2601
rect 1664 2567 1722 2573
rect 1664 2533 1676 2567
rect 1710 2564 1722 2567
rect 4154 2564 4160 2576
rect 1710 2536 4160 2564
rect 1710 2533 1722 2536
rect 1664 2527 1722 2533
rect 4154 2524 4160 2536
rect 4212 2524 4218 2576
rect 4332 2567 4390 2573
rect 4332 2533 4344 2567
rect 4378 2564 4390 2567
rect 4430 2564 4436 2576
rect 4378 2536 4436 2564
rect 4378 2533 4390 2536
rect 4332 2527 4390 2533
rect 4430 2524 4436 2536
rect 4488 2524 4494 2576
rect 5460 2564 5488 2595
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 5718 2592 5724 2644
rect 5776 2632 5782 2644
rect 5905 2635 5963 2641
rect 5905 2632 5917 2635
rect 5776 2604 5917 2632
rect 5776 2592 5782 2604
rect 5905 2601 5917 2604
rect 5951 2601 5963 2635
rect 5905 2595 5963 2601
rect 5994 2592 6000 2644
rect 6052 2632 6058 2644
rect 6052 2604 6097 2632
rect 7024 2604 8156 2632
rect 6052 2592 6058 2604
rect 7024 2564 7052 2604
rect 5460 2536 7052 2564
rect 7098 2524 7104 2576
rect 7156 2524 7162 2576
rect 7466 2524 7472 2576
rect 7524 2564 7530 2576
rect 7926 2564 7932 2576
rect 7524 2536 7932 2564
rect 7524 2524 7530 2536
rect 7926 2524 7932 2536
rect 7984 2524 7990 2576
rect 8128 2564 8156 2604
rect 8202 2592 8208 2644
rect 8260 2632 8266 2644
rect 8849 2635 8907 2641
rect 8849 2632 8861 2635
rect 8260 2604 8861 2632
rect 8260 2592 8266 2604
rect 8849 2601 8861 2604
rect 8895 2632 8907 2635
rect 9306 2632 9312 2644
rect 8895 2604 9312 2632
rect 8895 2601 8907 2604
rect 8849 2595 8907 2601
rect 9306 2592 9312 2604
rect 9364 2592 9370 2644
rect 9401 2635 9459 2641
rect 9401 2601 9413 2635
rect 9447 2601 9459 2635
rect 9401 2595 9459 2601
rect 8478 2564 8484 2576
rect 8128 2536 8484 2564
rect 8478 2524 8484 2536
rect 8536 2524 8542 2576
rect 8662 2564 8668 2576
rect 8579 2536 8668 2564
rect 1394 2456 1400 2508
rect 1452 2496 1458 2508
rect 3234 2496 3240 2508
rect 1452 2468 1497 2496
rect 3195 2468 3240 2496
rect 1452 2456 1458 2468
rect 3234 2456 3240 2468
rect 3292 2456 3298 2508
rect 6365 2499 6423 2505
rect 6365 2465 6377 2499
rect 6411 2496 6423 2499
rect 7116 2496 7144 2524
rect 6411 2468 7144 2496
rect 7184 2499 7242 2505
rect 6411 2465 6423 2468
rect 6365 2459 6423 2465
rect 7184 2465 7196 2499
rect 7230 2496 7242 2499
rect 8018 2496 8024 2508
rect 7230 2468 8024 2496
rect 7230 2465 7242 2468
rect 7184 2459 7242 2465
rect 8018 2456 8024 2468
rect 8076 2456 8082 2508
rect 8579 2496 8607 2536
rect 8662 2524 8668 2536
rect 8720 2564 8726 2576
rect 8757 2567 8815 2573
rect 8757 2564 8769 2567
rect 8720 2536 8769 2564
rect 8720 2524 8726 2536
rect 8757 2533 8769 2536
rect 8803 2533 8815 2567
rect 9416 2564 9444 2595
rect 9858 2592 9864 2644
rect 9916 2632 9922 2644
rect 10134 2632 10140 2644
rect 9916 2604 10140 2632
rect 9916 2592 9922 2604
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 10594 2632 10600 2644
rect 10555 2604 10600 2632
rect 10594 2592 10600 2604
rect 10652 2592 10658 2644
rect 11054 2632 11060 2644
rect 11015 2604 11060 2632
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 11146 2592 11152 2644
rect 11204 2632 11210 2644
rect 11425 2635 11483 2641
rect 11425 2632 11437 2635
rect 11204 2604 11437 2632
rect 11204 2592 11210 2604
rect 11425 2601 11437 2604
rect 11471 2601 11483 2635
rect 12618 2632 12624 2644
rect 11425 2595 11483 2601
rect 11808 2604 12112 2632
rect 12579 2604 12624 2632
rect 10410 2564 10416 2576
rect 8757 2527 8815 2533
rect 8864 2536 9352 2564
rect 9416 2536 10416 2564
rect 8864 2508 8892 2536
rect 8128 2468 8607 2496
rect 3326 2428 3332 2440
rect 3287 2400 3332 2428
rect 3326 2388 3332 2400
rect 3384 2388 3390 2440
rect 3418 2388 3424 2440
rect 3476 2428 3482 2440
rect 3694 2428 3700 2440
rect 3476 2400 3521 2428
rect 3655 2400 3700 2428
rect 3476 2388 3482 2400
rect 3694 2388 3700 2400
rect 3752 2388 3758 2440
rect 6086 2428 6092 2440
rect 6047 2400 6092 2428
rect 6086 2388 6092 2400
rect 6144 2388 6150 2440
rect 7926 2388 7932 2440
rect 7984 2428 7990 2440
rect 8128 2428 8156 2468
rect 8846 2456 8852 2508
rect 8904 2456 8910 2508
rect 9030 2456 9036 2508
rect 9088 2496 9094 2508
rect 9214 2496 9220 2508
rect 9088 2468 9220 2496
rect 9088 2456 9094 2468
rect 9214 2456 9220 2468
rect 9272 2456 9278 2508
rect 8662 2428 8668 2440
rect 7984 2400 8156 2428
rect 8220 2400 8668 2428
rect 7984 2388 7990 2400
rect 2774 2292 2780 2304
rect 2735 2264 2780 2292
rect 2774 2252 2780 2264
rect 2832 2252 2838 2304
rect 2869 2295 2927 2301
rect 2869 2261 2881 2295
rect 2915 2292 2927 2295
rect 5074 2292 5080 2304
rect 2915 2264 5080 2292
rect 2915 2261 2927 2264
rect 2869 2255 2927 2261
rect 5074 2252 5080 2264
rect 5132 2252 5138 2304
rect 6546 2292 6552 2304
rect 6507 2264 6552 2292
rect 6546 2252 6552 2264
rect 6604 2252 6610 2304
rect 7558 2252 7564 2304
rect 7616 2292 7622 2304
rect 8220 2292 8248 2400
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 8941 2431 8999 2437
rect 8941 2397 8953 2431
rect 8987 2397 8999 2431
rect 9324 2428 9352 2536
rect 10410 2524 10416 2536
rect 10468 2524 10474 2576
rect 10870 2524 10876 2576
rect 10928 2564 10934 2576
rect 11808 2564 11836 2604
rect 10928 2536 11836 2564
rect 12084 2564 12112 2604
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 12710 2592 12716 2644
rect 12768 2632 12774 2644
rect 12989 2635 13047 2641
rect 12989 2632 13001 2635
rect 12768 2604 13001 2632
rect 12768 2592 12774 2604
rect 12989 2601 13001 2604
rect 13035 2601 13047 2635
rect 12989 2595 13047 2601
rect 13814 2592 13820 2644
rect 13872 2632 13878 2644
rect 15378 2632 15384 2644
rect 13872 2604 15384 2632
rect 13872 2592 13878 2604
rect 15378 2592 15384 2604
rect 15436 2592 15442 2644
rect 15930 2632 15936 2644
rect 15891 2604 15936 2632
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 20162 2632 20168 2644
rect 20123 2604 20168 2632
rect 20162 2592 20168 2604
rect 20220 2592 20226 2644
rect 13081 2567 13139 2573
rect 13081 2564 13093 2567
rect 12084 2536 13093 2564
rect 10928 2524 10934 2536
rect 13081 2533 13093 2536
rect 13127 2533 13139 2567
rect 13081 2527 13139 2533
rect 14734 2524 14740 2576
rect 14792 2564 14798 2576
rect 15841 2567 15899 2573
rect 15841 2564 15853 2567
rect 14792 2536 15853 2564
rect 14792 2524 14798 2536
rect 15841 2533 15853 2536
rect 15887 2533 15899 2567
rect 15841 2527 15899 2533
rect 10042 2456 10048 2508
rect 10100 2496 10106 2508
rect 10137 2499 10195 2505
rect 10137 2496 10149 2499
rect 10100 2468 10149 2496
rect 10100 2456 10106 2468
rect 10137 2465 10149 2468
rect 10183 2465 10195 2499
rect 10137 2459 10195 2465
rect 10226 2456 10232 2508
rect 10284 2496 10290 2508
rect 10965 2499 11023 2505
rect 10284 2468 10329 2496
rect 10284 2456 10290 2468
rect 10965 2465 10977 2499
rect 11011 2496 11023 2499
rect 11054 2496 11060 2508
rect 11011 2468 11060 2496
rect 11011 2465 11023 2468
rect 10965 2459 11023 2465
rect 11054 2456 11060 2468
rect 11112 2456 11118 2508
rect 11790 2496 11796 2508
rect 11751 2468 11796 2496
rect 11790 2456 11796 2468
rect 11848 2456 11854 2508
rect 11885 2499 11943 2505
rect 11885 2465 11897 2499
rect 11931 2465 11943 2499
rect 11885 2459 11943 2465
rect 10318 2428 10324 2440
rect 9324 2400 10324 2428
rect 8941 2391 8999 2397
rect 8389 2363 8447 2369
rect 8389 2329 8401 2363
rect 8435 2360 8447 2363
rect 8846 2360 8852 2372
rect 8435 2332 8852 2360
rect 8435 2329 8447 2332
rect 8389 2323 8447 2329
rect 8846 2320 8852 2332
rect 8904 2320 8910 2372
rect 8956 2360 8984 2391
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 10870 2388 10876 2440
rect 10928 2428 10934 2440
rect 11149 2431 11207 2437
rect 11149 2428 11161 2431
rect 10928 2400 11161 2428
rect 10928 2388 10934 2400
rect 11149 2397 11161 2400
rect 11195 2397 11207 2431
rect 11149 2391 11207 2397
rect 11698 2388 11704 2440
rect 11756 2428 11762 2440
rect 11900 2428 11928 2459
rect 12066 2456 12072 2508
rect 12124 2496 12130 2508
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 12124 2468 14197 2496
rect 12124 2456 12130 2468
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 14185 2459 14243 2465
rect 14366 2456 14372 2508
rect 14424 2496 14430 2508
rect 17037 2499 17095 2505
rect 17037 2496 17049 2499
rect 14424 2468 17049 2496
rect 14424 2456 14430 2468
rect 17037 2465 17049 2468
rect 17083 2465 17095 2499
rect 17037 2459 17095 2465
rect 17218 2456 17224 2508
rect 17276 2496 17282 2508
rect 18877 2499 18935 2505
rect 18877 2496 18889 2499
rect 17276 2468 18889 2496
rect 17276 2456 17282 2468
rect 18877 2465 18889 2468
rect 18923 2465 18935 2499
rect 19978 2496 19984 2508
rect 19939 2468 19984 2496
rect 18877 2459 18935 2465
rect 19978 2456 19984 2468
rect 20036 2456 20042 2508
rect 11756 2400 11928 2428
rect 11756 2388 11762 2400
rect 11974 2388 11980 2440
rect 12032 2428 12038 2440
rect 12032 2400 12077 2428
rect 12032 2388 12038 2400
rect 12342 2388 12348 2440
rect 12400 2428 12406 2440
rect 13173 2431 13231 2437
rect 13173 2428 13185 2431
rect 12400 2400 13185 2428
rect 12400 2388 12406 2400
rect 13173 2397 13185 2400
rect 13219 2428 13231 2431
rect 14550 2428 14556 2440
rect 13219 2400 14556 2428
rect 13219 2397 13231 2400
rect 13173 2391 13231 2397
rect 14550 2388 14556 2400
rect 14608 2428 14614 2440
rect 16025 2431 16083 2437
rect 16025 2428 16037 2431
rect 14608 2400 16037 2428
rect 14608 2388 14614 2400
rect 16025 2397 16037 2400
rect 16071 2397 16083 2431
rect 16025 2391 16083 2397
rect 9122 2360 9128 2372
rect 8956 2332 9128 2360
rect 9122 2320 9128 2332
rect 9180 2320 9186 2372
rect 11606 2360 11612 2372
rect 9232 2332 11612 2360
rect 7616 2264 8248 2292
rect 8297 2295 8355 2301
rect 7616 2252 7622 2264
rect 8297 2261 8309 2295
rect 8343 2292 8355 2295
rect 8478 2292 8484 2304
rect 8343 2264 8484 2292
rect 8343 2261 8355 2264
rect 8297 2255 8355 2261
rect 8478 2252 8484 2264
rect 8536 2252 8542 2304
rect 8662 2252 8668 2304
rect 8720 2292 8726 2304
rect 9232 2292 9260 2332
rect 11606 2320 11612 2332
rect 11664 2320 11670 2372
rect 13722 2320 13728 2372
rect 13780 2360 13786 2372
rect 15470 2360 15476 2372
rect 13780 2332 15240 2360
rect 15431 2332 15476 2360
rect 13780 2320 13786 2332
rect 9766 2292 9772 2304
rect 8720 2264 9260 2292
rect 9727 2264 9772 2292
rect 8720 2252 8726 2264
rect 9766 2252 9772 2264
rect 9824 2252 9830 2304
rect 10134 2252 10140 2304
rect 10192 2292 10198 2304
rect 13814 2292 13820 2304
rect 10192 2264 13820 2292
rect 10192 2252 10198 2264
rect 13814 2252 13820 2264
rect 13872 2252 13878 2304
rect 14369 2295 14427 2301
rect 14369 2261 14381 2295
rect 14415 2292 14427 2295
rect 14734 2292 14740 2304
rect 14415 2264 14740 2292
rect 14415 2261 14427 2264
rect 14369 2255 14427 2261
rect 14734 2252 14740 2264
rect 14792 2252 14798 2304
rect 15212 2292 15240 2332
rect 15470 2320 15476 2332
rect 15528 2320 15534 2372
rect 17221 2295 17279 2301
rect 17221 2292 17233 2295
rect 15212 2264 17233 2292
rect 17221 2261 17233 2264
rect 17267 2261 17279 2295
rect 17221 2255 17279 2261
rect 19061 2295 19119 2301
rect 19061 2261 19073 2295
rect 19107 2292 19119 2295
rect 19886 2292 19892 2304
rect 19107 2264 19892 2292
rect 19107 2261 19119 2264
rect 19061 2255 19119 2261
rect 19886 2252 19892 2264
rect 19944 2252 19950 2304
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 3694 2048 3700 2100
rect 3752 2088 3758 2100
rect 11790 2088 11796 2100
rect 3752 2060 11796 2088
rect 3752 2048 3758 2060
rect 11790 2048 11796 2060
rect 11848 2048 11854 2100
rect 9674 2020 9680 2032
rect 6012 1992 9680 2020
rect 3234 1912 3240 1964
rect 3292 1952 3298 1964
rect 6012 1952 6040 1992
rect 9674 1980 9680 1992
rect 9732 1980 9738 2032
rect 9766 1980 9772 2032
rect 9824 2020 9830 2032
rect 12986 2020 12992 2032
rect 9824 1992 12992 2020
rect 9824 1980 9830 1992
rect 12986 1980 12992 1992
rect 13044 1980 13050 2032
rect 3292 1924 6040 1952
rect 3292 1912 3298 1924
rect 6546 1912 6552 1964
rect 6604 1952 6610 1964
rect 18414 1952 18420 1964
rect 6604 1924 18420 1952
rect 6604 1912 6610 1924
rect 18414 1912 18420 1924
rect 18472 1912 18478 1964
rect 3326 1844 3332 1896
rect 3384 1884 3390 1896
rect 9858 1884 9864 1896
rect 3384 1856 9864 1884
rect 3384 1844 3390 1856
rect 9858 1844 9864 1856
rect 9916 1844 9922 1896
rect 9950 1844 9956 1896
rect 10008 1884 10014 1896
rect 11974 1884 11980 1896
rect 10008 1856 11980 1884
rect 10008 1844 10014 1856
rect 11974 1844 11980 1856
rect 12032 1844 12038 1896
rect 12250 1844 12256 1896
rect 12308 1884 12314 1896
rect 19978 1884 19984 1896
rect 12308 1856 19984 1884
rect 12308 1844 12314 1856
rect 19978 1844 19984 1856
rect 20036 1844 20042 1896
rect 2774 1776 2780 1828
rect 2832 1816 2838 1828
rect 8754 1816 8760 1828
rect 2832 1788 8760 1816
rect 2832 1776 2838 1788
rect 8754 1776 8760 1788
rect 8812 1776 8818 1828
rect 12158 1816 12164 1828
rect 9416 1788 12164 1816
rect 1578 1708 1584 1760
rect 1636 1748 1642 1760
rect 6822 1748 6828 1760
rect 1636 1720 6828 1748
rect 1636 1708 1642 1720
rect 6822 1708 6828 1720
rect 6880 1748 6886 1760
rect 8113 1751 8171 1757
rect 8113 1748 8125 1751
rect 6880 1720 8125 1748
rect 6880 1708 6886 1720
rect 8113 1717 8125 1720
rect 8159 1717 8171 1751
rect 8113 1711 8171 1717
rect 8478 1708 8484 1760
rect 8536 1748 8542 1760
rect 9416 1748 9444 1788
rect 12158 1776 12164 1788
rect 12216 1776 12222 1828
rect 12802 1776 12808 1828
rect 12860 1816 12866 1828
rect 13262 1816 13268 1828
rect 12860 1788 13268 1816
rect 12860 1776 12866 1788
rect 13262 1776 13268 1788
rect 13320 1776 13326 1828
rect 8536 1720 9444 1748
rect 8536 1708 8542 1720
rect 9490 1708 9496 1760
rect 9548 1748 9554 1760
rect 14366 1748 14372 1760
rect 9548 1720 14372 1748
rect 9548 1708 9554 1720
rect 14366 1708 14372 1720
rect 14424 1708 14430 1760
rect 658 1640 664 1692
rect 716 1680 722 1692
rect 8202 1680 8208 1692
rect 716 1652 8208 1680
rect 716 1640 722 1652
rect 8202 1640 8208 1652
rect 8260 1640 8266 1692
rect 8846 1640 8852 1692
rect 8904 1680 8910 1692
rect 10134 1680 10140 1692
rect 8904 1652 10140 1680
rect 8904 1640 8910 1652
rect 10134 1640 10140 1652
rect 10192 1640 10198 1692
rect 10413 1683 10471 1689
rect 10413 1649 10425 1683
rect 10459 1680 10471 1683
rect 14458 1680 14464 1692
rect 10459 1652 14464 1680
rect 10459 1649 10471 1652
rect 10413 1643 10471 1649
rect 14458 1640 14464 1652
rect 14516 1640 14522 1692
rect 2314 1572 2320 1624
rect 2372 1612 2378 1624
rect 11698 1612 11704 1624
rect 2372 1584 11704 1612
rect 2372 1572 2378 1584
rect 11698 1572 11704 1584
rect 11756 1572 11762 1624
rect 13170 1612 13176 1624
rect 12728 1584 13176 1612
rect 198 1504 204 1556
rect 256 1544 262 1556
rect 8386 1544 8392 1556
rect 256 1516 8392 1544
rect 256 1504 262 1516
rect 8386 1504 8392 1516
rect 8444 1504 8450 1556
rect 8478 1504 8484 1556
rect 8536 1544 8542 1556
rect 12728 1544 12756 1584
rect 13170 1572 13176 1584
rect 13228 1572 13234 1624
rect 8536 1516 12756 1544
rect 8536 1504 8542 1516
rect 4246 1436 4252 1488
rect 4304 1476 4310 1488
rect 4982 1476 4988 1488
rect 4304 1448 4988 1476
rect 4304 1436 4310 1448
rect 4982 1436 4988 1448
rect 5040 1476 5046 1488
rect 11054 1476 11060 1488
rect 5040 1448 11060 1476
rect 5040 1436 5046 1448
rect 11054 1436 11060 1448
rect 11112 1436 11118 1488
rect 2958 1368 2964 1420
rect 3016 1408 3022 1420
rect 7374 1408 7380 1420
rect 3016 1380 7380 1408
rect 3016 1368 3022 1380
rect 7374 1368 7380 1380
rect 7432 1368 7438 1420
rect 8113 1411 8171 1417
rect 8113 1377 8125 1411
rect 8159 1408 8171 1411
rect 10226 1408 10232 1420
rect 8159 1380 10232 1408
rect 8159 1377 8171 1380
rect 8113 1371 8171 1377
rect 10226 1368 10232 1380
rect 10284 1408 10290 1420
rect 10413 1411 10471 1417
rect 10413 1408 10425 1411
rect 10284 1380 10425 1408
rect 10284 1368 10290 1380
rect 10413 1377 10425 1380
rect 10459 1377 10471 1411
rect 10413 1371 10471 1377
rect 1118 1300 1124 1352
rect 1176 1340 1182 1352
rect 6638 1340 6644 1352
rect 1176 1312 6644 1340
rect 1176 1300 1182 1312
rect 6638 1300 6644 1312
rect 6696 1300 6702 1352
rect 3418 1232 3424 1284
rect 3476 1272 3482 1284
rect 6454 1272 6460 1284
rect 3476 1244 6460 1272
rect 3476 1232 3482 1244
rect 6454 1232 6460 1244
rect 6512 1232 6518 1284
rect 10410 1232 10416 1284
rect 10468 1272 10474 1284
rect 16574 1272 16580 1284
rect 10468 1244 16580 1272
rect 10468 1232 10474 1244
rect 16574 1232 16580 1244
rect 16632 1232 16638 1284
rect 19242 552 19248 604
rect 19300 592 19306 604
rect 20806 592 20812 604
rect 19300 564 20812 592
rect 19300 552 19306 564
rect 20806 552 20812 564
rect 20864 552 20870 604
<< via1 >>
rect 7012 20748 7064 20800
rect 8116 20748 8168 20800
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 4160 20544 4212 20596
rect 12532 20544 12584 20596
rect 14096 20544 14148 20596
rect 15200 20544 15252 20596
rect 19432 20544 19484 20596
rect 21272 20544 21324 20596
rect 9680 20476 9732 20528
rect 5724 20408 5776 20460
rect 7104 20408 7156 20460
rect 3976 20340 4028 20392
rect 4160 20340 4212 20392
rect 8484 20383 8536 20392
rect 4620 20272 4672 20324
rect 8484 20349 8493 20383
rect 8493 20349 8527 20383
rect 8527 20349 8536 20383
rect 8484 20340 8536 20349
rect 10324 20451 10376 20460
rect 10324 20417 10333 20451
rect 10333 20417 10367 20451
rect 10367 20417 10376 20451
rect 10324 20408 10376 20417
rect 12900 20408 12952 20460
rect 10416 20340 10468 20392
rect 11336 20383 11388 20392
rect 11336 20349 11345 20383
rect 11345 20349 11379 20383
rect 11379 20349 11388 20383
rect 11336 20340 11388 20349
rect 12992 20340 13044 20392
rect 10968 20272 11020 20324
rect 11244 20272 11296 20324
rect 17776 20340 17828 20392
rect 19984 20383 20036 20392
rect 13544 20272 13596 20324
rect 19984 20349 19993 20383
rect 19993 20349 20027 20383
rect 20027 20349 20036 20383
rect 19984 20340 20036 20349
rect 2688 20204 2740 20256
rect 5632 20247 5684 20256
rect 5632 20213 5641 20247
rect 5641 20213 5675 20247
rect 5675 20213 5684 20247
rect 5632 20204 5684 20213
rect 6644 20204 6696 20256
rect 8668 20247 8720 20256
rect 8668 20213 8677 20247
rect 8677 20213 8711 20247
rect 8711 20213 8720 20247
rect 8668 20204 8720 20213
rect 10140 20247 10192 20256
rect 10140 20213 10149 20247
rect 10149 20213 10183 20247
rect 10183 20213 10192 20247
rect 10140 20204 10192 20213
rect 10600 20204 10652 20256
rect 11704 20204 11756 20256
rect 11796 20204 11848 20256
rect 13084 20247 13136 20256
rect 13084 20213 13093 20247
rect 13093 20213 13127 20247
rect 13127 20213 13136 20247
rect 13084 20204 13136 20213
rect 13360 20204 13412 20256
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 1952 20043 2004 20052
rect 1952 20009 1961 20043
rect 1961 20009 1995 20043
rect 1995 20009 2004 20043
rect 1952 20000 2004 20009
rect 3056 20043 3108 20052
rect 3056 20009 3065 20043
rect 3065 20009 3099 20043
rect 3099 20009 3108 20043
rect 3056 20000 3108 20009
rect 3792 20000 3844 20052
rect 7288 20000 7340 20052
rect 7380 20000 7432 20052
rect 5632 19932 5684 19984
rect 7840 19932 7892 19984
rect 9220 20000 9272 20052
rect 10324 20000 10376 20052
rect 10600 20043 10652 20052
rect 10600 20009 10609 20043
rect 10609 20009 10643 20043
rect 10643 20009 10652 20043
rect 10600 20000 10652 20009
rect 12808 20000 12860 20052
rect 14740 20000 14792 20052
rect 16120 20000 16172 20052
rect 18144 20000 18196 20052
rect 19800 20000 19852 20052
rect 20812 20000 20864 20052
rect 11244 19932 11296 19984
rect 11336 19932 11388 19984
rect 16948 19932 17000 19984
rect 1860 19864 1912 19916
rect 3516 19864 3568 19916
rect 3608 19864 3660 19916
rect 4528 19907 4580 19916
rect 4528 19873 4537 19907
rect 4537 19873 4571 19907
rect 4571 19873 4580 19907
rect 4528 19864 4580 19873
rect 7104 19864 7156 19916
rect 9864 19864 9916 19916
rect 12532 19907 12584 19916
rect 12532 19873 12541 19907
rect 12541 19873 12575 19907
rect 12575 19873 12584 19907
rect 12532 19864 12584 19873
rect 12716 19864 12768 19916
rect 4620 19839 4672 19848
rect 4620 19805 4629 19839
rect 4629 19805 4663 19839
rect 4663 19805 4672 19839
rect 4620 19796 4672 19805
rect 5540 19796 5592 19848
rect 5632 19796 5684 19848
rect 4068 19771 4120 19780
rect 4068 19737 4077 19771
rect 4077 19737 4111 19771
rect 4111 19737 4120 19771
rect 4068 19728 4120 19737
rect 8760 19796 8812 19848
rect 8852 19796 8904 19848
rect 10232 19796 10284 19848
rect 11244 19839 11296 19848
rect 11244 19805 11253 19839
rect 11253 19805 11287 19839
rect 11287 19805 11296 19839
rect 11244 19796 11296 19805
rect 11336 19796 11388 19848
rect 12808 19839 12860 19848
rect 12808 19805 12817 19839
rect 12817 19805 12851 19839
rect 12851 19805 12860 19839
rect 12808 19796 12860 19805
rect 13912 19864 13964 19916
rect 17408 19864 17460 19916
rect 7840 19728 7892 19780
rect 15200 19728 15252 19780
rect 16304 19728 16356 19780
rect 7104 19660 7156 19712
rect 7564 19660 7616 19712
rect 9772 19660 9824 19712
rect 12440 19660 12492 19712
rect 18880 19864 18932 19916
rect 17868 19796 17920 19848
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 5540 19499 5592 19508
rect 5540 19465 5549 19499
rect 5549 19465 5583 19499
rect 5583 19465 5592 19499
rect 5540 19456 5592 19465
rect 5908 19456 5960 19508
rect 9220 19456 9272 19508
rect 11980 19456 12032 19508
rect 12900 19456 12952 19508
rect 14556 19456 14608 19508
rect 14004 19388 14056 19440
rect 2136 19320 2188 19372
rect 2688 19320 2740 19372
rect 1492 19295 1544 19304
rect 1492 19261 1501 19295
rect 1501 19261 1535 19295
rect 1535 19261 1544 19295
rect 1492 19252 1544 19261
rect 3424 19252 3476 19304
rect 3976 19252 4028 19304
rect 8852 19320 8904 19372
rect 6920 19252 6972 19304
rect 7104 19295 7156 19304
rect 7104 19261 7113 19295
rect 7113 19261 7147 19295
rect 7147 19261 7156 19295
rect 7104 19252 7156 19261
rect 8208 19252 8260 19304
rect 12256 19320 12308 19372
rect 15016 19363 15068 19372
rect 15016 19329 15025 19363
rect 15025 19329 15059 19363
rect 15059 19329 15068 19363
rect 15016 19320 15068 19329
rect 12440 19295 12492 19304
rect 12440 19261 12449 19295
rect 12449 19261 12483 19295
rect 12483 19261 12492 19295
rect 12440 19252 12492 19261
rect 13084 19252 13136 19304
rect 14464 19252 14516 19304
rect 15292 19252 15344 19304
rect 2780 19184 2832 19236
rect 4252 19184 4304 19236
rect 5448 19184 5500 19236
rect 7564 19184 7616 19236
rect 2688 19116 2740 19168
rect 2964 19159 3016 19168
rect 2964 19125 2973 19159
rect 2973 19125 3007 19159
rect 3007 19125 3016 19159
rect 2964 19116 3016 19125
rect 4068 19116 4120 19168
rect 8484 19159 8536 19168
rect 8484 19125 8493 19159
rect 8493 19125 8527 19159
rect 8527 19125 8536 19159
rect 8484 19116 8536 19125
rect 9128 19184 9180 19236
rect 10232 19184 10284 19236
rect 10968 19184 11020 19236
rect 13452 19184 13504 19236
rect 17040 19252 17092 19304
rect 16396 19227 16448 19236
rect 14004 19116 14056 19168
rect 16396 19193 16405 19227
rect 16405 19193 16439 19227
rect 16439 19193 16448 19227
rect 16396 19184 16448 19193
rect 19616 19252 19668 19304
rect 15200 19116 15252 19168
rect 20352 19116 20404 19168
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 2872 18912 2924 18964
rect 6920 18912 6972 18964
rect 204 18844 256 18896
rect 1768 18819 1820 18828
rect 1768 18785 1777 18819
rect 1777 18785 1811 18819
rect 1811 18785 1820 18819
rect 1768 18776 1820 18785
rect 4252 18776 4304 18828
rect 664 18708 716 18760
rect 3792 18708 3844 18760
rect 1124 18640 1176 18692
rect 3700 18640 3752 18692
rect 7196 18844 7248 18896
rect 4712 18776 4764 18828
rect 4896 18776 4948 18828
rect 7288 18776 7340 18828
rect 7656 18912 7708 18964
rect 8208 18912 8260 18964
rect 9680 18912 9732 18964
rect 12256 18912 12308 18964
rect 22192 18912 22244 18964
rect 7840 18844 7892 18896
rect 9956 18776 10008 18828
rect 4620 18751 4672 18760
rect 4620 18717 4629 18751
rect 4629 18717 4663 18751
rect 4663 18717 4672 18751
rect 4620 18708 4672 18717
rect 4804 18708 4856 18760
rect 7104 18708 7156 18760
rect 8208 18708 8260 18760
rect 2872 18572 2924 18624
rect 4252 18572 4304 18624
rect 5264 18572 5316 18624
rect 5632 18615 5684 18624
rect 5632 18581 5641 18615
rect 5641 18581 5675 18615
rect 5675 18581 5684 18615
rect 5632 18572 5684 18581
rect 9220 18640 9272 18692
rect 8576 18615 8628 18624
rect 8576 18581 8585 18615
rect 8585 18581 8619 18615
rect 8619 18581 8628 18615
rect 8576 18572 8628 18581
rect 9312 18572 9364 18624
rect 10784 18776 10836 18828
rect 11704 18776 11756 18828
rect 15200 18844 15252 18896
rect 15476 18844 15528 18896
rect 13544 18776 13596 18828
rect 16028 18776 16080 18828
rect 17960 18844 18012 18896
rect 17224 18819 17276 18828
rect 17224 18785 17233 18819
rect 17233 18785 17267 18819
rect 17267 18785 17276 18819
rect 17224 18776 17276 18785
rect 18696 18776 18748 18828
rect 11980 18708 12032 18760
rect 12440 18708 12492 18760
rect 12624 18708 12676 18760
rect 12808 18708 12860 18760
rect 13268 18708 13320 18760
rect 13636 18708 13688 18760
rect 15292 18708 15344 18760
rect 16120 18708 16172 18760
rect 17684 18708 17736 18760
rect 12900 18572 12952 18624
rect 14004 18572 14056 18624
rect 15200 18572 15252 18624
rect 15568 18572 15620 18624
rect 18144 18572 18196 18624
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 1676 18368 1728 18420
rect 2596 18368 2648 18420
rect 12716 18368 12768 18420
rect 2504 18300 2556 18352
rect 2044 18232 2096 18284
rect 4252 18232 4304 18284
rect 7288 18300 7340 18352
rect 9220 18300 9272 18352
rect 12348 18300 12400 18352
rect 2320 18164 2372 18216
rect 3148 18164 3200 18216
rect 2596 18096 2648 18148
rect 3976 18164 4028 18216
rect 5632 18232 5684 18284
rect 7472 18232 7524 18284
rect 8208 18275 8260 18284
rect 8208 18241 8217 18275
rect 8217 18241 8251 18275
rect 8251 18241 8260 18275
rect 8208 18232 8260 18241
rect 9680 18232 9732 18284
rect 9864 18232 9916 18284
rect 10692 18232 10744 18284
rect 12900 18232 12952 18284
rect 17684 18368 17736 18420
rect 21732 18368 21784 18420
rect 15200 18300 15252 18352
rect 14740 18232 14792 18284
rect 15292 18232 15344 18284
rect 16856 18232 16908 18284
rect 17040 18232 17092 18284
rect 18972 18232 19024 18284
rect 2780 18028 2832 18080
rect 3148 18028 3200 18080
rect 3332 18071 3384 18080
rect 3332 18037 3341 18071
rect 3341 18037 3375 18071
rect 3375 18037 3384 18071
rect 3332 18028 3384 18037
rect 3884 18028 3936 18080
rect 4252 18028 4304 18080
rect 6000 18096 6052 18148
rect 8484 18139 8536 18148
rect 8484 18105 8518 18139
rect 8518 18105 8536 18139
rect 8484 18096 8536 18105
rect 8944 18164 8996 18216
rect 10876 18164 10928 18216
rect 14188 18164 14240 18216
rect 13820 18096 13872 18148
rect 15384 18096 15436 18148
rect 17684 18096 17736 18148
rect 6184 18028 6236 18080
rect 6828 18071 6880 18080
rect 6828 18037 6837 18071
rect 6837 18037 6871 18071
rect 6871 18037 6880 18071
rect 6828 18028 6880 18037
rect 9588 18071 9640 18080
rect 9588 18037 9597 18071
rect 9597 18037 9631 18071
rect 9631 18037 9640 18071
rect 9588 18028 9640 18037
rect 11152 18028 11204 18080
rect 12164 18028 12216 18080
rect 12716 18028 12768 18080
rect 14004 18028 14056 18080
rect 14372 18071 14424 18080
rect 14372 18037 14381 18071
rect 14381 18037 14415 18071
rect 14415 18037 14424 18071
rect 14372 18028 14424 18037
rect 14740 18028 14792 18080
rect 16120 18028 16172 18080
rect 16396 18028 16448 18080
rect 18052 18071 18104 18080
rect 18052 18037 18061 18071
rect 18061 18037 18095 18071
rect 18095 18037 18104 18071
rect 18052 18028 18104 18037
rect 20260 18028 20312 18080
rect 22652 18028 22704 18080
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 7656 17824 7708 17876
rect 9036 17824 9088 17876
rect 9496 17824 9548 17876
rect 9588 17824 9640 17876
rect 11704 17824 11756 17876
rect 11888 17824 11940 17876
rect 12256 17824 12308 17876
rect 4068 17756 4120 17808
rect 13360 17756 13412 17808
rect 18604 17824 18656 17876
rect 19064 17824 19116 17876
rect 4804 17688 4856 17740
rect 7196 17688 7248 17740
rect 8576 17688 8628 17740
rect 8944 17688 8996 17740
rect 11612 17688 11664 17740
rect 12348 17688 12400 17740
rect 12900 17688 12952 17740
rect 2412 17620 2464 17672
rect 2044 17552 2096 17604
rect 3976 17552 4028 17604
rect 5540 17620 5592 17672
rect 10600 17663 10652 17672
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 10968 17620 11020 17672
rect 16488 17756 16540 17808
rect 16672 17756 16724 17808
rect 20260 17756 20312 17808
rect 15384 17688 15436 17740
rect 15752 17731 15804 17740
rect 15752 17697 15761 17731
rect 15761 17697 15795 17731
rect 15795 17697 15804 17731
rect 15752 17688 15804 17697
rect 16028 17688 16080 17740
rect 18512 17688 18564 17740
rect 19892 17688 19944 17740
rect 13820 17620 13872 17672
rect 14004 17620 14056 17672
rect 14280 17620 14332 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 16396 17620 16448 17672
rect 17316 17663 17368 17672
rect 17316 17629 17325 17663
rect 17325 17629 17359 17663
rect 17359 17629 17368 17663
rect 17316 17620 17368 17629
rect 18236 17620 18288 17672
rect 2412 17484 2464 17536
rect 5448 17527 5500 17536
rect 5448 17493 5457 17527
rect 5457 17493 5491 17527
rect 5491 17493 5500 17527
rect 5448 17484 5500 17493
rect 10968 17484 11020 17536
rect 11244 17484 11296 17536
rect 11704 17484 11756 17536
rect 13084 17484 13136 17536
rect 19248 17620 19300 17672
rect 20812 17552 20864 17604
rect 16212 17484 16264 17536
rect 17132 17484 17184 17536
rect 17224 17484 17276 17536
rect 19064 17484 19116 17536
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 3332 17280 3384 17332
rect 4344 17280 4396 17332
rect 4988 17280 5040 17332
rect 5172 17280 5224 17332
rect 14280 17280 14332 17332
rect 7656 17255 7708 17264
rect 7656 17221 7665 17255
rect 7665 17221 7699 17255
rect 7699 17221 7708 17255
rect 7656 17212 7708 17221
rect 4804 17144 4856 17196
rect 5448 17144 5500 17196
rect 5724 17144 5776 17196
rect 10140 17212 10192 17264
rect 12440 17212 12492 17264
rect 12532 17212 12584 17264
rect 17592 17212 17644 17264
rect 18420 17212 18472 17264
rect 8576 17144 8628 17196
rect 2044 17076 2096 17128
rect 2504 17119 2556 17128
rect 2504 17085 2538 17119
rect 2538 17085 2556 17119
rect 2504 17076 2556 17085
rect 5356 17076 5408 17128
rect 6552 17076 6604 17128
rect 7012 17076 7064 17128
rect 7380 17076 7432 17128
rect 10784 17144 10836 17196
rect 10968 17144 11020 17196
rect 12992 17144 13044 17196
rect 14740 17144 14792 17196
rect 17316 17144 17368 17196
rect 18512 17187 18564 17196
rect 18512 17153 18521 17187
rect 18521 17153 18555 17187
rect 18555 17153 18564 17187
rect 18512 17144 18564 17153
rect 10600 17119 10652 17128
rect 2504 16940 2556 16992
rect 4988 16940 5040 16992
rect 10600 17085 10609 17119
rect 10609 17085 10643 17119
rect 10643 17085 10652 17119
rect 10600 17076 10652 17085
rect 11704 17076 11756 17128
rect 13912 17076 13964 17128
rect 15108 17076 15160 17128
rect 15292 17119 15344 17128
rect 15292 17085 15301 17119
rect 15301 17085 15335 17119
rect 15335 17085 15344 17119
rect 15292 17076 15344 17085
rect 8208 17008 8260 17060
rect 9036 17008 9088 17060
rect 8576 16940 8628 16992
rect 9128 16940 9180 16992
rect 9956 16940 10008 16992
rect 12532 17008 12584 17060
rect 19708 17076 19760 17128
rect 12348 16940 12400 16992
rect 12624 16940 12676 16992
rect 12900 16940 12952 16992
rect 14740 16940 14792 16992
rect 15660 17008 15712 17060
rect 16120 16940 16172 16992
rect 19064 16940 19116 16992
rect 19800 16940 19852 16992
rect 20076 16983 20128 16992
rect 20076 16949 20085 16983
rect 20085 16949 20119 16983
rect 20119 16949 20128 16983
rect 20076 16940 20128 16949
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 4344 16736 4396 16788
rect 5080 16736 5132 16788
rect 4160 16600 4212 16652
rect 5724 16736 5776 16788
rect 7656 16736 7708 16788
rect 7564 16668 7616 16720
rect 7012 16600 7064 16652
rect 7196 16600 7248 16652
rect 8576 16736 8628 16788
rect 11796 16736 11848 16788
rect 12348 16736 12400 16788
rect 20076 16736 20128 16788
rect 7932 16668 7984 16720
rect 12440 16668 12492 16720
rect 8024 16600 8076 16652
rect 3516 16532 3568 16584
rect 4988 16532 5040 16584
rect 8576 16600 8628 16652
rect 9864 16600 9916 16652
rect 10784 16600 10836 16652
rect 11060 16600 11112 16652
rect 11704 16600 11756 16652
rect 16120 16711 16172 16720
rect 16120 16677 16154 16711
rect 16154 16677 16172 16711
rect 16120 16668 16172 16677
rect 16212 16668 16264 16720
rect 9772 16532 9824 16584
rect 10600 16575 10652 16584
rect 10600 16541 10609 16575
rect 10609 16541 10643 16575
rect 10643 16541 10652 16575
rect 10600 16532 10652 16541
rect 2964 16396 3016 16448
rect 3516 16396 3568 16448
rect 4068 16439 4120 16448
rect 4068 16405 4077 16439
rect 4077 16405 4111 16439
rect 4111 16405 4120 16439
rect 4068 16396 4120 16405
rect 7380 16464 7432 16516
rect 10876 16532 10928 16584
rect 13084 16600 13136 16652
rect 14004 16600 14056 16652
rect 18144 16668 18196 16720
rect 18604 16668 18656 16720
rect 7288 16396 7340 16448
rect 12348 16464 12400 16516
rect 13176 16532 13228 16584
rect 13268 16532 13320 16584
rect 13636 16532 13688 16584
rect 15292 16532 15344 16584
rect 15476 16532 15528 16584
rect 13360 16464 13412 16516
rect 18144 16532 18196 16584
rect 8668 16396 8720 16448
rect 8852 16396 8904 16448
rect 12532 16396 12584 16448
rect 13176 16396 13228 16448
rect 15844 16396 15896 16448
rect 16028 16396 16080 16448
rect 17316 16396 17368 16448
rect 18420 16464 18472 16516
rect 19708 16464 19760 16516
rect 19340 16396 19392 16448
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 4160 16192 4212 16244
rect 2412 16099 2464 16108
rect 2412 16065 2421 16099
rect 2421 16065 2455 16099
rect 2455 16065 2464 16099
rect 2412 16056 2464 16065
rect 3056 15988 3108 16040
rect 3976 16124 4028 16176
rect 9772 16192 9824 16244
rect 9864 16192 9916 16244
rect 7196 16124 7248 16176
rect 7748 16124 7800 16176
rect 5356 16099 5408 16108
rect 5356 16065 5365 16099
rect 5365 16065 5399 16099
rect 5399 16065 5408 16099
rect 5356 16056 5408 16065
rect 6000 16056 6052 16108
rect 7380 15988 7432 16040
rect 8300 16056 8352 16108
rect 12716 16124 12768 16176
rect 11336 16099 11388 16108
rect 11336 16065 11345 16099
rect 11345 16065 11379 16099
rect 11379 16065 11388 16099
rect 11336 16056 11388 16065
rect 8024 15988 8076 16040
rect 10416 15988 10468 16040
rect 10600 15988 10652 16040
rect 12716 15988 12768 16040
rect 16580 16124 16632 16176
rect 15476 16056 15528 16108
rect 3700 15963 3752 15972
rect 3700 15929 3709 15963
rect 3709 15929 3743 15963
rect 3743 15929 3752 15963
rect 3700 15920 3752 15929
rect 4436 15920 4488 15972
rect 6000 15852 6052 15904
rect 7656 15852 7708 15904
rect 8668 15920 8720 15972
rect 9128 15920 9180 15972
rect 13176 15920 13228 15972
rect 13636 15920 13688 15972
rect 16120 16056 16172 16108
rect 19064 16124 19116 16176
rect 16304 15988 16356 16040
rect 16488 15920 16540 15972
rect 9864 15852 9916 15904
rect 9956 15895 10008 15904
rect 9956 15861 9965 15895
rect 9965 15861 9999 15895
rect 9999 15861 10008 15895
rect 9956 15852 10008 15861
rect 10416 15852 10468 15904
rect 13912 15852 13964 15904
rect 15292 15852 15344 15904
rect 15384 15895 15436 15904
rect 15384 15861 15393 15895
rect 15393 15861 15427 15895
rect 15427 15861 15436 15895
rect 15384 15852 15436 15861
rect 16396 15852 16448 15904
rect 18144 16056 18196 16108
rect 19340 16056 19392 16108
rect 17408 15988 17460 16040
rect 17592 15988 17644 16040
rect 20260 15988 20312 16040
rect 19524 15920 19576 15972
rect 17040 15852 17092 15904
rect 17408 15852 17460 15904
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 3608 15648 3660 15700
rect 4436 15648 4488 15700
rect 5172 15648 5224 15700
rect 5448 15648 5500 15700
rect 5540 15648 5592 15700
rect 7196 15648 7248 15700
rect 7472 15648 7524 15700
rect 8208 15648 8260 15700
rect 9220 15648 9272 15700
rect 10140 15648 10192 15700
rect 10416 15648 10468 15700
rect 10968 15648 11020 15700
rect 13636 15691 13688 15700
rect 13636 15657 13645 15691
rect 13645 15657 13679 15691
rect 13679 15657 13688 15691
rect 13636 15648 13688 15657
rect 14004 15691 14056 15700
rect 14004 15657 14013 15691
rect 14013 15657 14047 15691
rect 14047 15657 14056 15691
rect 14004 15648 14056 15657
rect 14096 15691 14148 15700
rect 14096 15657 14105 15691
rect 14105 15657 14139 15691
rect 14139 15657 14148 15691
rect 14096 15648 14148 15657
rect 16672 15648 16724 15700
rect 17592 15648 17644 15700
rect 2596 15580 2648 15632
rect 3884 15512 3936 15564
rect 9956 15580 10008 15632
rect 3056 15487 3108 15496
rect 3056 15453 3065 15487
rect 3065 15453 3099 15487
rect 3099 15453 3108 15487
rect 3056 15444 3108 15453
rect 6460 15512 6512 15564
rect 6552 15512 6604 15564
rect 1400 15376 1452 15428
rect 5632 15444 5684 15496
rect 7288 15512 7340 15564
rect 10048 15555 10100 15564
rect 10048 15521 10057 15555
rect 10057 15521 10091 15555
rect 10091 15521 10100 15555
rect 10048 15512 10100 15521
rect 9680 15444 9732 15496
rect 8300 15376 8352 15428
rect 9864 15376 9916 15428
rect 2228 15308 2280 15360
rect 7288 15308 7340 15360
rect 8208 15308 8260 15360
rect 9128 15308 9180 15360
rect 9680 15351 9732 15360
rect 9680 15317 9689 15351
rect 9689 15317 9723 15351
rect 9723 15317 9732 15351
rect 9680 15308 9732 15317
rect 10416 15512 10468 15564
rect 11612 15555 11664 15564
rect 11612 15521 11621 15555
rect 11621 15521 11655 15555
rect 11655 15521 11664 15555
rect 11612 15512 11664 15521
rect 10508 15444 10560 15496
rect 10968 15444 11020 15496
rect 14556 15580 14608 15632
rect 14924 15580 14976 15632
rect 16212 15580 16264 15632
rect 15292 15555 15344 15564
rect 15292 15521 15301 15555
rect 15301 15521 15335 15555
rect 15335 15521 15344 15555
rect 15292 15512 15344 15521
rect 17316 15512 17368 15564
rect 19156 15555 19208 15564
rect 19156 15521 19165 15555
rect 19165 15521 19199 15555
rect 19199 15521 19208 15555
rect 19156 15512 19208 15521
rect 14004 15444 14056 15496
rect 14740 15444 14792 15496
rect 15844 15444 15896 15496
rect 16488 15444 16540 15496
rect 18144 15444 18196 15496
rect 19340 15487 19392 15496
rect 12164 15376 12216 15428
rect 17592 15376 17644 15428
rect 19340 15453 19349 15487
rect 19349 15453 19383 15487
rect 19383 15453 19392 15487
rect 19340 15444 19392 15453
rect 19616 15376 19668 15428
rect 20076 15376 20128 15428
rect 10232 15308 10284 15360
rect 12716 15308 12768 15360
rect 14096 15308 14148 15360
rect 18880 15308 18932 15360
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 1952 15104 2004 15156
rect 3240 15104 3292 15156
rect 10876 15104 10928 15156
rect 15752 15104 15804 15156
rect 19524 15104 19576 15156
rect 1676 15036 1728 15088
rect 2136 15036 2188 15088
rect 5632 15036 5684 15088
rect 7472 15036 7524 15088
rect 9772 15036 9824 15088
rect 14280 15036 14332 15088
rect 14556 15036 14608 15088
rect 3516 14968 3568 15020
rect 1492 14900 1544 14952
rect 2044 14900 2096 14952
rect 3332 14832 3384 14884
rect 4988 14832 5040 14884
rect 2136 14764 2188 14816
rect 2504 14764 2556 14816
rect 5172 14807 5224 14816
rect 5172 14773 5181 14807
rect 5181 14773 5215 14807
rect 5215 14773 5224 14807
rect 5172 14764 5224 14773
rect 5356 14764 5408 14816
rect 6644 14943 6696 14952
rect 6644 14909 6653 14943
rect 6653 14909 6687 14943
rect 6687 14909 6696 14943
rect 6644 14900 6696 14909
rect 7288 14968 7340 15020
rect 7748 14968 7800 15020
rect 10232 14968 10284 15020
rect 6552 14832 6604 14884
rect 8852 14875 8904 14884
rect 8852 14841 8886 14875
rect 8886 14841 8904 14875
rect 8852 14832 8904 14841
rect 9312 14900 9364 14952
rect 11888 14968 11940 15020
rect 12532 14968 12584 15020
rect 13176 15011 13228 15020
rect 13176 14977 13185 15011
rect 13185 14977 13219 15011
rect 13219 14977 13228 15011
rect 13176 14968 13228 14977
rect 13636 14968 13688 15020
rect 17592 15036 17644 15088
rect 18420 15036 18472 15088
rect 14740 14900 14792 14952
rect 15108 14900 15160 14952
rect 16396 14968 16448 15020
rect 17316 14968 17368 15020
rect 19340 14968 19392 15020
rect 16856 14900 16908 14952
rect 17868 14900 17920 14952
rect 18144 14900 18196 14952
rect 18972 14900 19024 14952
rect 20076 14943 20128 14952
rect 20076 14909 20085 14943
rect 20085 14909 20119 14943
rect 20119 14909 20128 14943
rect 20076 14900 20128 14909
rect 11152 14875 11204 14884
rect 5632 14764 5684 14816
rect 5908 14764 5960 14816
rect 9588 14764 9640 14816
rect 9956 14807 10008 14816
rect 9956 14773 9965 14807
rect 9965 14773 9999 14807
rect 9999 14773 10008 14807
rect 9956 14764 10008 14773
rect 10784 14807 10836 14816
rect 10784 14773 10793 14807
rect 10793 14773 10827 14807
rect 10827 14773 10836 14807
rect 10784 14764 10836 14773
rect 11152 14841 11161 14875
rect 11161 14841 11195 14875
rect 11195 14841 11204 14875
rect 11152 14832 11204 14841
rect 12440 14832 12492 14884
rect 13360 14832 13412 14884
rect 14924 14832 14976 14884
rect 12716 14807 12768 14816
rect 12716 14773 12725 14807
rect 12725 14773 12759 14807
rect 12759 14773 12768 14807
rect 12716 14764 12768 14773
rect 13084 14807 13136 14816
rect 13084 14773 13093 14807
rect 13093 14773 13127 14807
rect 13127 14773 13136 14807
rect 13084 14764 13136 14773
rect 14096 14764 14148 14816
rect 14740 14764 14792 14816
rect 16396 14832 16448 14884
rect 17040 14764 17092 14816
rect 18236 14764 18288 14816
rect 18420 14807 18472 14816
rect 18420 14773 18429 14807
rect 18429 14773 18463 14807
rect 18463 14773 18472 14807
rect 18420 14764 18472 14773
rect 18604 14764 18656 14816
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 6552 14560 6604 14612
rect 6828 14603 6880 14612
rect 6828 14569 6837 14603
rect 6837 14569 6871 14603
rect 6871 14569 6880 14603
rect 6828 14560 6880 14569
rect 7012 14560 7064 14612
rect 10784 14560 10836 14612
rect 10876 14560 10928 14612
rect 12440 14560 12492 14612
rect 12532 14560 12584 14612
rect 14280 14603 14332 14612
rect 5908 14492 5960 14544
rect 6736 14492 6788 14544
rect 9680 14492 9732 14544
rect 3976 14424 4028 14476
rect 4712 14424 4764 14476
rect 5080 14424 5132 14476
rect 6368 14424 6420 14476
rect 7012 14424 7064 14476
rect 9220 14424 9272 14476
rect 11336 14492 11388 14544
rect 12992 14492 13044 14544
rect 14280 14569 14289 14603
rect 14289 14569 14323 14603
rect 14323 14569 14332 14603
rect 14280 14560 14332 14569
rect 18328 14560 18380 14612
rect 11428 14467 11480 14476
rect 1492 14356 1544 14408
rect 4988 14399 5040 14408
rect 4988 14365 4997 14399
rect 4997 14365 5031 14399
rect 5031 14365 5040 14399
rect 4988 14356 5040 14365
rect 6460 14356 6512 14408
rect 8668 14399 8720 14408
rect 6368 14288 6420 14340
rect 8668 14365 8677 14399
rect 8677 14365 8711 14399
rect 8711 14365 8720 14399
rect 8668 14356 8720 14365
rect 9680 14356 9732 14408
rect 9956 14288 10008 14340
rect 4160 14220 4212 14272
rect 6184 14220 6236 14272
rect 9312 14220 9364 14272
rect 9588 14220 9640 14272
rect 11428 14433 11437 14467
rect 11437 14433 11471 14467
rect 11471 14433 11480 14467
rect 11428 14424 11480 14433
rect 12440 14424 12492 14476
rect 14280 14424 14332 14476
rect 14464 14424 14516 14476
rect 15200 14424 15252 14476
rect 18972 14492 19024 14544
rect 18144 14424 18196 14476
rect 20260 14424 20312 14476
rect 11888 14399 11940 14408
rect 11888 14365 11897 14399
rect 11897 14365 11931 14399
rect 11931 14365 11940 14399
rect 11888 14356 11940 14365
rect 13912 14356 13964 14408
rect 17316 14399 17368 14408
rect 17316 14365 17325 14399
rect 17325 14365 17359 14399
rect 17359 14365 17368 14399
rect 17316 14356 17368 14365
rect 18880 14399 18932 14408
rect 18880 14365 18889 14399
rect 18889 14365 18923 14399
rect 18923 14365 18932 14399
rect 18880 14356 18932 14365
rect 13176 14288 13228 14340
rect 15660 14288 15712 14340
rect 17960 14288 18012 14340
rect 11152 14220 11204 14272
rect 11888 14220 11940 14272
rect 13360 14220 13412 14272
rect 15936 14220 15988 14272
rect 18144 14220 18196 14272
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 3148 14016 3200 14068
rect 9680 14059 9732 14068
rect 3792 13948 3844 14000
rect 8852 13991 8904 14000
rect 8852 13957 8861 13991
rect 8861 13957 8895 13991
rect 8895 13957 8904 13991
rect 8852 13948 8904 13957
rect 9680 14025 9689 14059
rect 9689 14025 9723 14059
rect 9723 14025 9732 14059
rect 9680 14016 9732 14025
rect 11796 14016 11848 14068
rect 20812 14059 20864 14068
rect 20812 14025 20821 14059
rect 20821 14025 20855 14059
rect 20855 14025 20864 14059
rect 20812 14016 20864 14025
rect 4068 13880 4120 13932
rect 1492 13855 1544 13864
rect 1492 13821 1501 13855
rect 1501 13821 1535 13855
rect 1535 13821 1544 13855
rect 1492 13812 1544 13821
rect 5172 13880 5224 13932
rect 13912 13948 13964 14000
rect 14096 13948 14148 14000
rect 7472 13855 7524 13864
rect 4160 13744 4212 13796
rect 2872 13719 2924 13728
rect 2872 13685 2881 13719
rect 2881 13685 2915 13719
rect 2915 13685 2924 13719
rect 2872 13676 2924 13685
rect 3240 13676 3292 13728
rect 7472 13821 7481 13855
rect 7481 13821 7515 13855
rect 7515 13821 7524 13855
rect 7472 13812 7524 13821
rect 12716 13880 12768 13932
rect 14464 13880 14516 13932
rect 15936 13948 15988 14000
rect 19340 13948 19392 14000
rect 19156 13880 19208 13932
rect 7748 13787 7800 13796
rect 7748 13753 7782 13787
rect 7782 13753 7800 13787
rect 7748 13744 7800 13753
rect 9404 13744 9456 13796
rect 13360 13812 13412 13864
rect 14096 13812 14148 13864
rect 16028 13812 16080 13864
rect 16120 13812 16172 13864
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 17040 13812 17092 13864
rect 18236 13812 18288 13864
rect 15200 13744 15252 13796
rect 8668 13676 8720 13728
rect 9772 13676 9824 13728
rect 10048 13719 10100 13728
rect 10048 13685 10057 13719
rect 10057 13685 10091 13719
rect 10091 13685 10100 13719
rect 10048 13676 10100 13685
rect 10324 13676 10376 13728
rect 10784 13676 10836 13728
rect 12624 13676 12676 13728
rect 13360 13676 13412 13728
rect 15476 13676 15528 13728
rect 17960 13744 18012 13796
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 3976 13472 4028 13524
rect 7748 13515 7800 13524
rect 2320 13447 2372 13456
rect 2320 13413 2329 13447
rect 2329 13413 2363 13447
rect 2363 13413 2372 13447
rect 2320 13404 2372 13413
rect 2412 13404 2464 13456
rect 6368 13404 6420 13456
rect 2780 13336 2832 13388
rect 4344 13336 4396 13388
rect 6460 13336 6512 13388
rect 7748 13481 7757 13515
rect 7757 13481 7791 13515
rect 7791 13481 7800 13515
rect 7748 13472 7800 13481
rect 8944 13472 8996 13524
rect 9312 13472 9364 13524
rect 11796 13472 11848 13524
rect 12348 13515 12400 13524
rect 6828 13404 6880 13456
rect 9772 13404 9824 13456
rect 9864 13404 9916 13456
rect 12348 13481 12357 13515
rect 12357 13481 12391 13515
rect 12391 13481 12400 13515
rect 12348 13472 12400 13481
rect 17316 13472 17368 13524
rect 17868 13472 17920 13524
rect 18972 13515 19024 13524
rect 18972 13481 18981 13515
rect 18981 13481 19015 13515
rect 19015 13481 19024 13515
rect 18972 13472 19024 13481
rect 19984 13472 20036 13524
rect 5172 13268 5224 13320
rect 6184 13200 6236 13252
rect 8668 13268 8720 13320
rect 9220 13268 9272 13320
rect 9312 13268 9364 13320
rect 12624 13404 12676 13456
rect 12900 13404 12952 13456
rect 13544 13404 13596 13456
rect 16856 13404 16908 13456
rect 12348 13336 12400 13388
rect 11796 13268 11848 13320
rect 15936 13336 15988 13388
rect 16488 13336 16540 13388
rect 16764 13379 16816 13388
rect 16764 13345 16773 13379
rect 16773 13345 16807 13379
rect 16807 13345 16816 13379
rect 18236 13404 18288 13456
rect 18880 13404 18932 13456
rect 16764 13336 16816 13345
rect 12808 13268 12860 13320
rect 14464 13268 14516 13320
rect 15660 13268 15712 13320
rect 12900 13200 12952 13252
rect 13268 13200 13320 13252
rect 3148 13132 3200 13184
rect 4160 13132 4212 13184
rect 5356 13132 5408 13184
rect 5724 13132 5776 13184
rect 8208 13132 8260 13184
rect 10048 13132 10100 13184
rect 11888 13132 11940 13184
rect 14004 13132 14056 13184
rect 14464 13132 14516 13184
rect 20168 13268 20220 13320
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 2780 12971 2832 12980
rect 2780 12937 2789 12971
rect 2789 12937 2823 12971
rect 2823 12937 2832 12971
rect 4344 12971 4396 12980
rect 2780 12928 2832 12937
rect 4344 12937 4353 12971
rect 4353 12937 4387 12971
rect 4387 12937 4396 12971
rect 4344 12928 4396 12937
rect 6644 12928 6696 12980
rect 6828 12971 6880 12980
rect 6828 12937 6837 12971
rect 6837 12937 6871 12971
rect 6871 12937 6880 12971
rect 6828 12928 6880 12937
rect 7196 12928 7248 12980
rect 9220 12928 9272 12980
rect 10784 12928 10836 12980
rect 11244 12928 11296 12980
rect 2872 12860 2924 12912
rect 2596 12792 2648 12844
rect 2780 12792 2832 12844
rect 3240 12835 3292 12844
rect 3240 12801 3249 12835
rect 3249 12801 3283 12835
rect 3283 12801 3292 12835
rect 3240 12792 3292 12801
rect 4436 12860 4488 12912
rect 9864 12860 9916 12912
rect 4528 12792 4580 12844
rect 4988 12792 5040 12844
rect 7288 12835 7340 12844
rect 7288 12801 7297 12835
rect 7297 12801 7331 12835
rect 7331 12801 7340 12835
rect 7288 12792 7340 12801
rect 7748 12792 7800 12844
rect 8208 12792 8260 12844
rect 9312 12792 9364 12844
rect 10140 12835 10192 12844
rect 10140 12801 10149 12835
rect 10149 12801 10183 12835
rect 10183 12801 10192 12835
rect 10140 12792 10192 12801
rect 11888 12928 11940 12980
rect 13636 12860 13688 12912
rect 16028 12903 16080 12912
rect 16028 12869 16037 12903
rect 16037 12869 16071 12903
rect 16071 12869 16080 12903
rect 16028 12860 16080 12869
rect 17040 12903 17092 12912
rect 17040 12869 17049 12903
rect 17049 12869 17083 12903
rect 17083 12869 17092 12903
rect 17040 12860 17092 12869
rect 17776 12860 17828 12912
rect 18604 12835 18656 12844
rect 3148 12767 3200 12776
rect 3148 12733 3157 12767
rect 3157 12733 3191 12767
rect 3191 12733 3200 12767
rect 3148 12724 3200 12733
rect 5356 12656 5408 12708
rect 10048 12724 10100 12776
rect 12440 12767 12492 12776
rect 12440 12733 12449 12767
rect 12449 12733 12483 12767
rect 12483 12733 12492 12767
rect 12440 12724 12492 12733
rect 18604 12801 18613 12835
rect 18613 12801 18647 12835
rect 18647 12801 18656 12835
rect 18604 12792 18656 12801
rect 2964 12588 3016 12640
rect 3148 12588 3200 12640
rect 3424 12588 3476 12640
rect 4160 12588 4212 12640
rect 4344 12588 4396 12640
rect 5172 12588 5224 12640
rect 8300 12588 8352 12640
rect 8852 12631 8904 12640
rect 8852 12597 8861 12631
rect 8861 12597 8895 12631
rect 8895 12597 8904 12631
rect 8852 12588 8904 12597
rect 9588 12656 9640 12708
rect 17960 12724 18012 12776
rect 18144 12724 18196 12776
rect 19616 12724 19668 12776
rect 9772 12588 9824 12640
rect 14740 12656 14792 12708
rect 17224 12656 17276 12708
rect 17408 12656 17460 12708
rect 17776 12656 17828 12708
rect 18972 12656 19024 12708
rect 16580 12588 16632 12640
rect 19708 12588 19760 12640
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 1308 12384 1360 12436
rect 1768 12384 1820 12436
rect 6460 12384 6512 12436
rect 8208 12384 8260 12436
rect 8300 12427 8352 12436
rect 8300 12393 8309 12427
rect 8309 12393 8343 12427
rect 8343 12393 8352 12427
rect 8300 12384 8352 12393
rect 9680 12384 9732 12436
rect 10600 12384 10652 12436
rect 10968 12384 11020 12436
rect 11612 12384 11664 12436
rect 11796 12384 11848 12436
rect 12440 12384 12492 12436
rect 14280 12384 14332 12436
rect 15476 12384 15528 12436
rect 2044 12316 2096 12368
rect 2688 12316 2740 12368
rect 4344 12316 4396 12368
rect 4804 12316 4856 12368
rect 5080 12316 5132 12368
rect 5632 12316 5684 12368
rect 5908 12316 5960 12368
rect 2136 12248 2188 12300
rect 2688 12223 2740 12232
rect 2688 12189 2697 12223
rect 2697 12189 2731 12223
rect 2731 12189 2740 12223
rect 2688 12180 2740 12189
rect 2780 12180 2832 12232
rect 3516 12180 3568 12232
rect 5264 12248 5316 12300
rect 5448 12180 5500 12232
rect 6552 12180 6604 12232
rect 7012 12248 7064 12300
rect 8392 12291 8444 12300
rect 8392 12257 8401 12291
rect 8401 12257 8435 12291
rect 8435 12257 8444 12291
rect 8392 12248 8444 12257
rect 4160 12112 4212 12164
rect 6092 12112 6144 12164
rect 7380 12180 7432 12232
rect 11980 12316 12032 12368
rect 12164 12316 12216 12368
rect 12532 12316 12584 12368
rect 13084 12316 13136 12368
rect 13636 12316 13688 12368
rect 18144 12316 18196 12368
rect 18604 12316 18656 12368
rect 19248 12384 19300 12436
rect 10784 12248 10836 12300
rect 12440 12248 12492 12300
rect 8668 12180 8720 12232
rect 9680 12180 9732 12232
rect 10324 12223 10376 12232
rect 7840 12112 7892 12164
rect 10048 12112 10100 12164
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 15108 12248 15160 12300
rect 16764 12248 16816 12300
rect 2964 12044 3016 12096
rect 3056 12044 3108 12096
rect 3424 12044 3476 12096
rect 4344 12044 4396 12096
rect 7472 12044 7524 12096
rect 11060 12044 11112 12096
rect 11704 12044 11756 12096
rect 15292 12180 15344 12232
rect 16028 12180 16080 12232
rect 13636 12044 13688 12096
rect 15660 12044 15712 12096
rect 18604 12044 18656 12096
rect 19248 12087 19300 12096
rect 19248 12053 19257 12087
rect 19257 12053 19291 12087
rect 19291 12053 19300 12087
rect 19248 12044 19300 12053
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 3056 11840 3108 11892
rect 6092 11840 6144 11892
rect 7288 11840 7340 11892
rect 7656 11840 7708 11892
rect 7932 11840 7984 11892
rect 8208 11840 8260 11892
rect 8760 11772 8812 11824
rect 1492 11636 1544 11688
rect 3516 11704 3568 11756
rect 5264 11704 5316 11756
rect 7288 11704 7340 11756
rect 7472 11747 7524 11756
rect 7472 11713 7481 11747
rect 7481 11713 7515 11747
rect 7515 11713 7524 11747
rect 7472 11704 7524 11713
rect 8024 11704 8076 11756
rect 8300 11704 8352 11756
rect 12440 11883 12492 11892
rect 12440 11849 12449 11883
rect 12449 11849 12483 11883
rect 12483 11849 12492 11883
rect 12440 11840 12492 11849
rect 17960 11840 18012 11892
rect 19064 11840 19116 11892
rect 14280 11772 14332 11824
rect 16948 11772 17000 11824
rect 12532 11704 12584 11756
rect 4896 11636 4948 11688
rect 8668 11636 8720 11688
rect 9312 11636 9364 11688
rect 9680 11679 9732 11688
rect 9680 11645 9689 11679
rect 9689 11645 9723 11679
rect 9723 11645 9732 11679
rect 9680 11636 9732 11645
rect 10324 11636 10376 11688
rect 11060 11636 11112 11688
rect 11428 11636 11480 11688
rect 2872 11568 2924 11620
rect 5264 11568 5316 11620
rect 7840 11568 7892 11620
rect 8300 11568 8352 11620
rect 4160 11500 4212 11552
rect 4804 11500 4856 11552
rect 5172 11500 5224 11552
rect 6092 11500 6144 11552
rect 11060 11543 11112 11552
rect 11060 11509 11069 11543
rect 11069 11509 11103 11543
rect 11103 11509 11112 11543
rect 11060 11500 11112 11509
rect 11796 11568 11848 11620
rect 12532 11568 12584 11620
rect 12808 11704 12860 11756
rect 13084 11704 13136 11756
rect 14464 11704 14516 11756
rect 15844 11704 15896 11756
rect 13176 11636 13228 11688
rect 14280 11636 14332 11688
rect 16304 11636 16356 11688
rect 12808 11543 12860 11552
rect 12808 11509 12817 11543
rect 12817 11509 12851 11543
rect 12851 11509 12860 11543
rect 12808 11500 12860 11509
rect 15108 11568 15160 11620
rect 16672 11568 16724 11620
rect 19064 11704 19116 11756
rect 19248 11704 19300 11756
rect 20168 11747 20220 11756
rect 20168 11713 20177 11747
rect 20177 11713 20211 11747
rect 20211 11713 20220 11747
rect 20168 11704 20220 11713
rect 15384 11543 15436 11552
rect 15384 11509 15393 11543
rect 15393 11509 15427 11543
rect 15427 11509 15436 11543
rect 15384 11500 15436 11509
rect 16028 11500 16080 11552
rect 18696 11568 18748 11620
rect 18880 11568 18932 11620
rect 17224 11500 17276 11552
rect 18236 11500 18288 11552
rect 19340 11500 19392 11552
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 1492 11228 1544 11280
rect 2044 11228 2096 11280
rect 2596 11296 2648 11348
rect 3976 11296 4028 11348
rect 4620 11296 4672 11348
rect 5908 11339 5960 11348
rect 3608 11228 3660 11280
rect 4988 11228 5040 11280
rect 3240 11160 3292 11212
rect 5908 11305 5917 11339
rect 5917 11305 5951 11339
rect 5951 11305 5960 11339
rect 5908 11296 5960 11305
rect 7472 11296 7524 11348
rect 6460 11228 6512 11280
rect 6920 11228 6972 11280
rect 11060 11228 11112 11280
rect 2044 11092 2096 11144
rect 2320 11092 2372 11144
rect 3056 11135 3108 11144
rect 3056 11101 3065 11135
rect 3065 11101 3099 11135
rect 3099 11101 3108 11135
rect 3056 11092 3108 11101
rect 4160 11092 4212 11144
rect 6276 10956 6328 11008
rect 6828 10956 6880 11008
rect 9680 11160 9732 11212
rect 10232 11160 10284 11212
rect 10692 11092 10744 11144
rect 11704 11296 11756 11348
rect 13636 11339 13688 11348
rect 13636 11305 13645 11339
rect 13645 11305 13679 11339
rect 13679 11305 13688 11339
rect 13636 11296 13688 11305
rect 14096 11339 14148 11348
rect 14096 11305 14105 11339
rect 14105 11305 14139 11339
rect 14139 11305 14148 11339
rect 14096 11296 14148 11305
rect 14464 11296 14516 11348
rect 16028 11296 16080 11348
rect 18144 11339 18196 11348
rect 18144 11305 18153 11339
rect 18153 11305 18187 11339
rect 18187 11305 18196 11339
rect 18144 11296 18196 11305
rect 18972 11339 19024 11348
rect 18972 11305 18981 11339
rect 18981 11305 19015 11339
rect 19015 11305 19024 11339
rect 18972 11296 19024 11305
rect 19340 11339 19392 11348
rect 19340 11305 19349 11339
rect 19349 11305 19383 11339
rect 19383 11305 19392 11339
rect 19340 11296 19392 11305
rect 11428 11228 11480 11280
rect 14004 11271 14056 11280
rect 14004 11237 14013 11271
rect 14013 11237 14047 11271
rect 14047 11237 14056 11271
rect 14004 11228 14056 11237
rect 15200 11228 15252 11280
rect 16764 11203 16816 11212
rect 16764 11169 16773 11203
rect 16773 11169 16807 11203
rect 16807 11169 16816 11203
rect 16764 11160 16816 11169
rect 17868 11160 17920 11212
rect 14740 11092 14792 11144
rect 15844 11092 15896 11144
rect 19432 11135 19484 11144
rect 19432 11101 19441 11135
rect 19441 11101 19475 11135
rect 19475 11101 19484 11135
rect 19432 11092 19484 11101
rect 8760 11067 8812 11076
rect 8760 11033 8769 11067
rect 8769 11033 8803 11067
rect 8803 11033 8812 11067
rect 8760 11024 8812 11033
rect 10784 11024 10836 11076
rect 8392 10956 8444 11008
rect 11152 10956 11204 11008
rect 11704 10999 11756 11008
rect 11704 10965 11713 10999
rect 11713 10965 11747 10999
rect 11747 10965 11756 10999
rect 11704 10956 11756 10965
rect 11796 10956 11848 11008
rect 13912 11024 13964 11076
rect 14832 11024 14884 11076
rect 15936 11024 15988 11076
rect 13636 10956 13688 11008
rect 18788 10956 18840 11008
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 3056 10752 3108 10804
rect 5172 10752 5224 10804
rect 6736 10752 6788 10804
rect 8392 10752 8444 10804
rect 9772 10752 9824 10804
rect 10324 10752 10376 10804
rect 11060 10752 11112 10804
rect 14096 10752 14148 10804
rect 15844 10795 15896 10804
rect 15844 10761 15853 10795
rect 15853 10761 15887 10795
rect 15887 10761 15896 10795
rect 15844 10752 15896 10761
rect 16672 10752 16724 10804
rect 19432 10752 19484 10804
rect 3976 10684 4028 10736
rect 2320 10591 2372 10600
rect 2320 10557 2354 10591
rect 2354 10557 2372 10591
rect 2320 10548 2372 10557
rect 2504 10480 2556 10532
rect 2688 10412 2740 10464
rect 11152 10684 11204 10736
rect 11888 10684 11940 10736
rect 14280 10684 14332 10736
rect 17500 10684 17552 10736
rect 3608 10548 3660 10600
rect 6828 10591 6880 10600
rect 6828 10557 6837 10591
rect 6837 10557 6871 10591
rect 6871 10557 6880 10591
rect 6828 10548 6880 10557
rect 4160 10480 4212 10532
rect 5540 10480 5592 10532
rect 6644 10480 6696 10532
rect 7104 10523 7156 10532
rect 7104 10489 7138 10523
rect 7138 10489 7156 10523
rect 7104 10480 7156 10489
rect 3608 10412 3660 10464
rect 6276 10412 6328 10464
rect 11428 10616 11480 10668
rect 15568 10616 15620 10668
rect 15844 10616 15896 10668
rect 16028 10616 16080 10668
rect 20168 10659 20220 10668
rect 20168 10625 20177 10659
rect 20177 10625 20211 10659
rect 20211 10625 20220 10659
rect 20168 10616 20220 10625
rect 11704 10548 11756 10600
rect 14464 10591 14516 10600
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 14464 10548 14516 10557
rect 9680 10480 9732 10532
rect 11152 10480 11204 10532
rect 11336 10480 11388 10532
rect 13084 10480 13136 10532
rect 16764 10548 16816 10600
rect 15660 10480 15712 10532
rect 16028 10480 16080 10532
rect 16856 10480 16908 10532
rect 17960 10480 18012 10532
rect 11060 10412 11112 10464
rect 11520 10412 11572 10464
rect 12808 10455 12860 10464
rect 12808 10421 12817 10455
rect 12817 10421 12851 10455
rect 12851 10421 12860 10455
rect 12808 10412 12860 10421
rect 14096 10412 14148 10464
rect 15936 10412 15988 10464
rect 17684 10412 17736 10464
rect 19984 10412 20036 10464
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 1860 10208 1912 10260
rect 7472 10208 7524 10260
rect 8208 10208 8260 10260
rect 8392 10208 8444 10260
rect 11336 10208 11388 10260
rect 11888 10208 11940 10260
rect 2688 10140 2740 10192
rect 4252 10140 4304 10192
rect 8300 10140 8352 10192
rect 13176 10140 13228 10192
rect 4068 10115 4120 10124
rect 4068 10081 4077 10115
rect 4077 10081 4111 10115
rect 4111 10081 4120 10115
rect 4068 10072 4120 10081
rect 5908 10072 5960 10124
rect 6092 10072 6144 10124
rect 7564 10072 7616 10124
rect 7840 10072 7892 10124
rect 7932 10072 7984 10124
rect 12348 10072 12400 10124
rect 12532 10072 12584 10124
rect 2504 10004 2556 10056
rect 6828 10004 6880 10056
rect 8024 10004 8076 10056
rect 7104 9936 7156 9988
rect 9680 10004 9732 10056
rect 11980 10004 12032 10056
rect 2872 9911 2924 9920
rect 2872 9877 2881 9911
rect 2881 9877 2915 9911
rect 2915 9877 2924 9911
rect 2872 9868 2924 9877
rect 3608 9868 3660 9920
rect 4344 9868 4396 9920
rect 6828 9868 6880 9920
rect 7656 9868 7708 9920
rect 7840 9868 7892 9920
rect 8760 9936 8812 9988
rect 9404 9936 9456 9988
rect 11428 9936 11480 9988
rect 11520 9936 11572 9988
rect 15384 10208 15436 10260
rect 15568 10208 15620 10260
rect 15660 10183 15712 10192
rect 15660 10149 15669 10183
rect 15669 10149 15703 10183
rect 15703 10149 15712 10183
rect 15660 10140 15712 10149
rect 18788 10251 18840 10260
rect 18788 10217 18797 10251
rect 18797 10217 18831 10251
rect 18831 10217 18840 10251
rect 18788 10208 18840 10217
rect 15936 10140 15988 10192
rect 13820 10004 13872 10056
rect 16120 10072 16172 10124
rect 16028 10004 16080 10056
rect 17408 10047 17460 10056
rect 17408 10013 17417 10047
rect 17417 10013 17451 10047
rect 17451 10013 17460 10047
rect 17408 10004 17460 10013
rect 18604 10004 18656 10056
rect 18788 10004 18840 10056
rect 13176 9868 13228 9920
rect 13912 9868 13964 9920
rect 14188 9868 14240 9920
rect 15292 9868 15344 9920
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 1952 9707 2004 9716
rect 1952 9673 1961 9707
rect 1961 9673 1995 9707
rect 1995 9673 2004 9707
rect 1952 9664 2004 9673
rect 5908 9664 5960 9716
rect 8392 9664 8444 9716
rect 8484 9664 8536 9716
rect 9312 9664 9364 9716
rect 9956 9664 10008 9716
rect 10232 9664 10284 9716
rect 12348 9664 12400 9716
rect 2596 9596 2648 9648
rect 3240 9596 3292 9648
rect 7012 9639 7064 9648
rect 1216 9392 1268 9444
rect 1492 9392 1544 9444
rect 2044 9460 2096 9512
rect 2688 9528 2740 9580
rect 3884 9460 3936 9512
rect 7012 9605 7021 9639
rect 7021 9605 7055 9639
rect 7055 9605 7064 9639
rect 7012 9596 7064 9605
rect 7104 9596 7156 9648
rect 2320 9392 2372 9444
rect 5540 9392 5592 9444
rect 7012 9460 7064 9512
rect 7564 9460 7616 9512
rect 7748 9460 7800 9512
rect 8024 9460 8076 9512
rect 8392 9435 8444 9444
rect 8392 9401 8401 9435
rect 8401 9401 8435 9435
rect 8435 9401 8444 9435
rect 8392 9392 8444 9401
rect 1860 9324 1912 9376
rect 2136 9367 2188 9376
rect 2136 9333 2145 9367
rect 2145 9333 2179 9367
rect 2179 9333 2188 9367
rect 2596 9367 2648 9376
rect 2136 9324 2188 9333
rect 2596 9333 2605 9367
rect 2605 9333 2639 9367
rect 2639 9333 2648 9367
rect 2596 9324 2648 9333
rect 3608 9324 3660 9376
rect 3884 9324 3936 9376
rect 4620 9324 4672 9376
rect 6460 9324 6512 9376
rect 7748 9324 7800 9376
rect 8944 9528 8996 9580
rect 9496 9528 9548 9580
rect 8576 9392 8628 9444
rect 9772 9460 9824 9512
rect 9956 9528 10008 9580
rect 10508 9571 10560 9580
rect 10508 9537 10517 9571
rect 10517 9537 10551 9571
rect 10551 9537 10560 9571
rect 10508 9528 10560 9537
rect 13084 9664 13136 9716
rect 13636 9664 13688 9716
rect 12900 9596 12952 9648
rect 13176 9571 13228 9580
rect 13176 9537 13185 9571
rect 13185 9537 13219 9571
rect 13219 9537 13228 9571
rect 13176 9528 13228 9537
rect 13912 9664 13964 9716
rect 14004 9664 14056 9716
rect 14188 9664 14240 9716
rect 16120 9707 16172 9716
rect 16120 9673 16129 9707
rect 16129 9673 16163 9707
rect 16163 9673 16172 9707
rect 16120 9664 16172 9673
rect 17500 9664 17552 9716
rect 17868 9664 17920 9716
rect 9128 9324 9180 9376
rect 9496 9367 9548 9376
rect 9496 9333 9505 9367
rect 9505 9333 9539 9367
rect 9539 9333 9548 9367
rect 9496 9324 9548 9333
rect 9864 9367 9916 9376
rect 9864 9333 9873 9367
rect 9873 9333 9907 9367
rect 9907 9333 9916 9367
rect 9864 9324 9916 9333
rect 10232 9367 10284 9376
rect 10232 9333 10241 9367
rect 10241 9333 10275 9367
rect 10275 9333 10284 9367
rect 10232 9324 10284 9333
rect 12348 9324 12400 9376
rect 17224 9596 17276 9648
rect 14464 9528 14516 9580
rect 17960 9528 18012 9580
rect 14280 9503 14332 9512
rect 14280 9469 14289 9503
rect 14289 9469 14323 9503
rect 14323 9469 14332 9503
rect 14280 9460 14332 9469
rect 15568 9460 15620 9512
rect 16212 9460 16264 9512
rect 16672 9460 16724 9512
rect 15476 9392 15528 9444
rect 15752 9392 15804 9444
rect 17040 9392 17092 9444
rect 17868 9460 17920 9512
rect 18604 9460 18656 9512
rect 18788 9392 18840 9444
rect 14004 9324 14056 9376
rect 14280 9324 14332 9376
rect 19248 9324 19300 9376
rect 19432 9367 19484 9376
rect 19432 9333 19441 9367
rect 19441 9333 19475 9367
rect 19475 9333 19484 9367
rect 19432 9324 19484 9333
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 1584 9120 1636 9172
rect 3332 9120 3384 9172
rect 3608 9120 3660 9172
rect 4160 9120 4212 9172
rect 4712 9120 4764 9172
rect 1308 9052 1360 9104
rect 2596 9052 2648 9104
rect 4620 9052 4672 9104
rect 6184 9120 6236 9172
rect 7656 9120 7708 9172
rect 9772 9120 9824 9172
rect 10232 9120 10284 9172
rect 12348 9163 12400 9172
rect 5908 9052 5960 9104
rect 1768 9027 1820 9036
rect 1768 8993 1777 9027
rect 1777 8993 1811 9027
rect 1811 8993 1820 9027
rect 1768 8984 1820 8993
rect 1860 9027 1912 9036
rect 1860 8993 1869 9027
rect 1869 8993 1903 9027
rect 1903 8993 1912 9027
rect 1860 8984 1912 8993
rect 2780 9027 2832 9036
rect 2780 8993 2789 9027
rect 2789 8993 2823 9027
rect 2823 8993 2832 9027
rect 2780 8984 2832 8993
rect 2136 8916 2188 8968
rect 2688 8916 2740 8968
rect 3608 8984 3660 9036
rect 4436 8984 4488 9036
rect 4528 8959 4580 8968
rect 1860 8848 1912 8900
rect 3976 8848 4028 8900
rect 4160 8848 4212 8900
rect 4528 8925 4537 8959
rect 4537 8925 4571 8959
rect 4571 8925 4580 8959
rect 4528 8916 4580 8925
rect 5172 8984 5224 9036
rect 5356 8916 5408 8968
rect 4988 8848 5040 8900
rect 5172 8848 5224 8900
rect 6092 8984 6144 9036
rect 6276 9052 6328 9104
rect 6552 9052 6604 9104
rect 6736 9052 6788 9104
rect 7564 9052 7616 9104
rect 7932 9052 7984 9104
rect 8576 9095 8628 9104
rect 8576 9061 8585 9095
rect 8585 9061 8619 9095
rect 8619 9061 8628 9095
rect 8576 9052 8628 9061
rect 9128 9052 9180 9104
rect 10600 9052 10652 9104
rect 8944 8984 8996 9036
rect 10232 9027 10284 9036
rect 10232 8993 10241 9027
rect 10241 8993 10275 9027
rect 10275 8993 10284 9027
rect 10232 8984 10284 8993
rect 11152 8984 11204 9036
rect 2688 8780 2740 8832
rect 6460 8848 6512 8900
rect 7840 8916 7892 8968
rect 8392 8916 8444 8968
rect 8576 8916 8628 8968
rect 9956 8916 10008 8968
rect 10600 8916 10652 8968
rect 12348 9129 12357 9163
rect 12357 9129 12391 9163
rect 12391 9129 12400 9163
rect 12348 9120 12400 9129
rect 13820 9120 13872 9172
rect 14096 9120 14148 9172
rect 14004 9052 14056 9104
rect 14464 9120 14516 9172
rect 16212 9120 16264 9172
rect 17868 9120 17920 9172
rect 18880 9163 18932 9172
rect 18880 9129 18889 9163
rect 18889 9129 18923 9163
rect 18923 9129 18932 9163
rect 18880 9120 18932 9129
rect 14740 9052 14792 9104
rect 19064 9052 19116 9104
rect 19432 9052 19484 9104
rect 6000 8780 6052 8832
rect 6092 8780 6144 8832
rect 8300 8780 8352 8832
rect 8392 8780 8444 8832
rect 9128 8780 9180 8832
rect 9680 8780 9732 8832
rect 11980 8780 12032 8832
rect 12348 8780 12400 8832
rect 12532 8848 12584 8900
rect 13820 8916 13872 8968
rect 15384 8916 15436 8968
rect 15568 8984 15620 9036
rect 16396 8984 16448 9036
rect 15844 8916 15896 8968
rect 16028 8916 16080 8968
rect 18972 8959 19024 8968
rect 18972 8925 18981 8959
rect 18981 8925 19015 8959
rect 19015 8925 19024 8959
rect 18972 8916 19024 8925
rect 16488 8848 16540 8900
rect 15752 8780 15804 8832
rect 16764 8780 16816 8832
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 1124 8576 1176 8628
rect 3608 8508 3660 8560
rect 2596 8440 2648 8492
rect 2872 8372 2924 8424
rect 3332 8372 3384 8424
rect 4988 8576 5040 8628
rect 4988 8440 5040 8492
rect 5632 8576 5684 8628
rect 6000 8576 6052 8628
rect 6552 8576 6604 8628
rect 5264 8508 5316 8560
rect 6276 8508 6328 8560
rect 7472 8508 7524 8560
rect 6368 8483 6420 8492
rect 6368 8449 6377 8483
rect 6377 8449 6411 8483
rect 6411 8449 6420 8483
rect 6368 8440 6420 8449
rect 6552 8440 6604 8492
rect 7748 8440 7800 8492
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 2504 8236 2556 8288
rect 3332 8236 3384 8288
rect 4436 8304 4488 8356
rect 5172 8304 5224 8356
rect 5908 8372 5960 8424
rect 7104 8372 7156 8424
rect 7932 8415 7984 8424
rect 7932 8381 7941 8415
rect 7941 8381 7975 8415
rect 7975 8381 7984 8415
rect 7932 8372 7984 8381
rect 9128 8576 9180 8628
rect 9772 8576 9824 8628
rect 9956 8576 10008 8628
rect 10600 8576 10652 8628
rect 14280 8576 14332 8628
rect 15476 8619 15528 8628
rect 15476 8585 15485 8619
rect 15485 8585 15519 8619
rect 15519 8585 15528 8619
rect 15476 8576 15528 8585
rect 12532 8508 12584 8560
rect 12624 8508 12676 8560
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 17960 8508 18012 8560
rect 9496 8304 9548 8356
rect 9772 8372 9824 8424
rect 16948 8483 17000 8492
rect 16948 8449 16957 8483
rect 16957 8449 16991 8483
rect 16991 8449 17000 8483
rect 16948 8440 17000 8449
rect 17868 8440 17920 8492
rect 10600 8372 10652 8424
rect 16764 8415 16816 8424
rect 11428 8304 11480 8356
rect 14280 8304 14332 8356
rect 16764 8381 16773 8415
rect 16773 8381 16807 8415
rect 16807 8381 16816 8415
rect 16764 8372 16816 8381
rect 18052 8415 18104 8424
rect 18052 8381 18061 8415
rect 18061 8381 18095 8415
rect 18095 8381 18104 8415
rect 18052 8372 18104 8381
rect 17224 8304 17276 8356
rect 18972 8304 19024 8356
rect 20260 8347 20312 8356
rect 20260 8313 20269 8347
rect 20269 8313 20303 8347
rect 20303 8313 20312 8347
rect 20260 8304 20312 8313
rect 4712 8236 4764 8288
rect 5080 8236 5132 8288
rect 6092 8236 6144 8288
rect 6828 8236 6880 8288
rect 7104 8236 7156 8288
rect 8576 8236 8628 8288
rect 15660 8236 15712 8288
rect 16764 8236 16816 8288
rect 18604 8236 18656 8288
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 1952 8032 2004 8084
rect 4344 8032 4396 8084
rect 4804 8032 4856 8084
rect 5264 8032 5316 8084
rect 6644 8075 6696 8084
rect 6644 8041 6653 8075
rect 6653 8041 6687 8075
rect 6687 8041 6696 8075
rect 6644 8032 6696 8041
rect 6736 8032 6788 8084
rect 10508 8032 10560 8084
rect 12164 8032 12216 8084
rect 12348 8032 12400 8084
rect 13084 8032 13136 8084
rect 13636 8075 13688 8084
rect 13636 8041 13645 8075
rect 13645 8041 13679 8075
rect 13679 8041 13688 8075
rect 13636 8032 13688 8041
rect 13820 8032 13872 8084
rect 14740 8032 14792 8084
rect 15384 8032 15436 8084
rect 2964 7964 3016 8016
rect 2320 7896 2372 7948
rect 2872 7828 2924 7880
rect 2504 7760 2556 7812
rect 1400 7735 1452 7744
rect 1400 7701 1409 7735
rect 1409 7701 1443 7735
rect 1443 7701 1452 7735
rect 1400 7692 1452 7701
rect 1584 7692 1636 7744
rect 2596 7692 2648 7744
rect 2964 7692 3016 7744
rect 4620 7896 4672 7948
rect 4896 7896 4948 7948
rect 5080 7896 5132 7948
rect 5816 7896 5868 7948
rect 6828 7896 6880 7948
rect 7104 7896 7156 7948
rect 7564 7939 7616 7948
rect 7564 7905 7573 7939
rect 7573 7905 7607 7939
rect 7607 7905 7616 7939
rect 7564 7896 7616 7905
rect 3332 7760 3384 7812
rect 6092 7692 6144 7744
rect 6460 7692 6512 7744
rect 9496 7896 9548 7948
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 9956 7939 10008 7948
rect 9956 7905 9990 7939
rect 9990 7905 10008 7939
rect 9956 7896 10008 7905
rect 11980 7896 12032 7948
rect 7932 7828 7984 7880
rect 8116 7760 8168 7812
rect 12532 7828 12584 7880
rect 10968 7760 11020 7812
rect 6736 7692 6788 7744
rect 8852 7692 8904 7744
rect 9864 7692 9916 7744
rect 13820 7896 13872 7948
rect 14096 7964 14148 8016
rect 16948 7964 17000 8016
rect 15660 7939 15712 7948
rect 15660 7905 15669 7939
rect 15669 7905 15703 7939
rect 15703 7905 15712 7939
rect 18052 8032 18104 8084
rect 15660 7896 15712 7905
rect 12992 7828 13044 7880
rect 14372 7828 14424 7880
rect 15476 7828 15528 7880
rect 18696 7964 18748 8016
rect 18052 7896 18104 7948
rect 18604 7896 18656 7948
rect 13084 7760 13136 7812
rect 12532 7692 12584 7744
rect 15384 7692 15436 7744
rect 16028 7692 16080 7744
rect 17040 7692 17092 7744
rect 18972 7692 19024 7744
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 1768 7488 1820 7540
rect 2136 7488 2188 7540
rect 2412 7488 2464 7540
rect 2780 7488 2832 7540
rect 5632 7488 5684 7540
rect 13084 7488 13136 7540
rect 13176 7488 13228 7540
rect 13452 7488 13504 7540
rect 15752 7488 15804 7540
rect 6460 7420 6512 7472
rect 6644 7420 6696 7472
rect 7840 7420 7892 7472
rect 8300 7420 8352 7472
rect 9496 7420 9548 7472
rect 12164 7420 12216 7472
rect 2596 7352 2648 7404
rect 4252 7352 4304 7404
rect 4344 7352 4396 7404
rect 5264 7352 5316 7404
rect 1768 7327 1820 7336
rect 1768 7293 1777 7327
rect 1777 7293 1811 7327
rect 1811 7293 1820 7327
rect 1768 7284 1820 7293
rect 1032 7216 1084 7268
rect 6000 7352 6052 7404
rect 6736 7352 6788 7404
rect 8024 7352 8076 7404
rect 6644 7284 6696 7336
rect 2412 7216 2464 7268
rect 3240 7216 3292 7268
rect 1308 7148 1360 7200
rect 1860 7191 1912 7200
rect 1860 7157 1869 7191
rect 1869 7157 1903 7191
rect 1903 7157 1912 7191
rect 1860 7148 1912 7157
rect 2044 7148 2096 7200
rect 2780 7148 2832 7200
rect 3608 7148 3660 7200
rect 5080 7216 5132 7268
rect 5724 7216 5776 7268
rect 6092 7259 6144 7268
rect 6092 7225 6101 7259
rect 6101 7225 6135 7259
rect 6135 7225 6144 7259
rect 6092 7216 6144 7225
rect 8208 7284 8260 7336
rect 7564 7216 7616 7268
rect 7932 7216 7984 7268
rect 8116 7216 8168 7268
rect 8300 7216 8352 7268
rect 8852 7216 8904 7268
rect 11428 7352 11480 7404
rect 9680 7284 9732 7336
rect 10416 7327 10468 7336
rect 10416 7293 10450 7327
rect 10450 7293 10468 7327
rect 10416 7284 10468 7293
rect 11336 7284 11388 7336
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 16120 7352 16172 7404
rect 13728 7284 13780 7336
rect 15384 7327 15436 7336
rect 15384 7293 15393 7327
rect 15393 7293 15427 7327
rect 15427 7293 15436 7327
rect 15384 7284 15436 7293
rect 18696 7420 18748 7472
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 18144 7284 18196 7336
rect 19984 7327 20036 7336
rect 19984 7293 19993 7327
rect 19993 7293 20027 7327
rect 20027 7293 20036 7327
rect 19984 7284 20036 7293
rect 11980 7216 12032 7268
rect 12164 7216 12216 7268
rect 12900 7216 12952 7268
rect 9036 7148 9088 7200
rect 9680 7148 9732 7200
rect 9864 7148 9916 7200
rect 12808 7148 12860 7200
rect 13084 7148 13136 7200
rect 15476 7191 15528 7200
rect 15476 7157 15485 7191
rect 15485 7157 15519 7191
rect 15519 7157 15528 7191
rect 15476 7148 15528 7157
rect 16672 7216 16724 7268
rect 17592 7216 17644 7268
rect 17132 7148 17184 7200
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 1308 6944 1360 6996
rect 3608 6944 3660 6996
rect 4988 6944 5040 6996
rect 5264 6987 5316 6996
rect 5264 6953 5273 6987
rect 5273 6953 5307 6987
rect 5307 6953 5316 6987
rect 5264 6944 5316 6953
rect 5632 6944 5684 6996
rect 4804 6876 4856 6928
rect 6276 6944 6328 6996
rect 6368 6944 6420 6996
rect 11428 6944 11480 6996
rect 11520 6944 11572 6996
rect 2964 6808 3016 6860
rect 3332 6808 3384 6860
rect 1308 6740 1360 6792
rect 2780 6740 2832 6792
rect 3700 6740 3752 6792
rect 1216 6604 1268 6656
rect 2780 6647 2832 6656
rect 2780 6613 2789 6647
rect 2789 6613 2823 6647
rect 2823 6613 2832 6647
rect 2780 6604 2832 6613
rect 3240 6604 3292 6656
rect 4068 6647 4120 6656
rect 4068 6613 4077 6647
rect 4077 6613 4111 6647
rect 4111 6613 4120 6647
rect 4068 6604 4120 6613
rect 4160 6604 4212 6656
rect 4988 6740 5040 6792
rect 5356 6740 5408 6792
rect 6644 6876 6696 6928
rect 7196 6876 7248 6928
rect 7472 6876 7524 6928
rect 7932 6876 7984 6928
rect 11704 6876 11756 6928
rect 10416 6851 10468 6860
rect 10416 6817 10425 6851
rect 10425 6817 10459 6851
rect 10459 6817 10468 6851
rect 10416 6808 10468 6817
rect 10968 6808 11020 6860
rect 16120 6876 16172 6928
rect 6368 6740 6420 6792
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 7748 6740 7800 6792
rect 9128 6740 9180 6792
rect 9864 6740 9916 6792
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 11336 6740 11388 6792
rect 11704 6740 11756 6792
rect 12532 6808 12584 6860
rect 14740 6808 14792 6860
rect 15844 6808 15896 6860
rect 16212 6851 16264 6860
rect 16212 6817 16221 6851
rect 16221 6817 16255 6851
rect 16255 6817 16264 6851
rect 16212 6808 16264 6817
rect 6184 6672 6236 6724
rect 11520 6672 11572 6724
rect 12164 6672 12216 6724
rect 14280 6740 14332 6792
rect 17868 6808 17920 6860
rect 17868 6672 17920 6724
rect 4804 6604 4856 6656
rect 5356 6604 5408 6656
rect 5816 6604 5868 6656
rect 7012 6604 7064 6656
rect 7656 6604 7708 6656
rect 9855 6604 9907 6656
rect 11060 6604 11112 6656
rect 15016 6604 15068 6656
rect 17592 6647 17644 6656
rect 17592 6613 17601 6647
rect 17601 6613 17635 6647
rect 17635 6613 17644 6647
rect 17592 6604 17644 6613
rect 18052 6604 18104 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 1308 6400 1360 6452
rect 3332 6400 3384 6452
rect 4804 6400 4856 6452
rect 5172 6400 5224 6452
rect 6276 6400 6328 6452
rect 6460 6400 6512 6452
rect 5540 6332 5592 6384
rect 1952 6239 2004 6248
rect 1952 6205 1961 6239
rect 1961 6205 1995 6239
rect 1995 6205 2004 6239
rect 1952 6196 2004 6205
rect 3700 6264 3752 6316
rect 4344 6196 4396 6248
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 6276 6264 6328 6316
rect 7564 6400 7616 6452
rect 8208 6400 8260 6452
rect 8392 6443 8444 6452
rect 8392 6409 8401 6443
rect 8401 6409 8435 6443
rect 8435 6409 8444 6443
rect 8392 6400 8444 6409
rect 8852 6307 8904 6316
rect 8852 6273 8861 6307
rect 8861 6273 8895 6307
rect 8895 6273 8904 6307
rect 8852 6264 8904 6273
rect 2136 6128 2188 6180
rect 2688 6128 2740 6180
rect 4620 6128 4672 6180
rect 5356 6128 5408 6180
rect 6644 6196 6696 6248
rect 8392 6128 8444 6180
rect 9772 6332 9824 6384
rect 12348 6400 12400 6452
rect 9128 6264 9180 6316
rect 9680 6264 9732 6316
rect 10416 6332 10468 6384
rect 9772 6196 9824 6248
rect 9680 6128 9732 6180
rect 3792 6060 3844 6112
rect 6184 6060 6236 6112
rect 6276 6060 6328 6112
rect 10600 6196 10652 6248
rect 11152 6264 11204 6316
rect 11428 6264 11480 6316
rect 11612 6332 11664 6384
rect 15476 6400 15528 6452
rect 16120 6400 16172 6452
rect 17500 6400 17552 6452
rect 19616 6443 19668 6452
rect 19616 6409 19625 6443
rect 19625 6409 19659 6443
rect 19659 6409 19668 6443
rect 19616 6400 19668 6409
rect 12164 6264 12216 6316
rect 12440 6307 12492 6316
rect 12440 6273 12449 6307
rect 12449 6273 12483 6307
rect 12483 6273 12492 6307
rect 12440 6264 12492 6273
rect 15568 6264 15620 6316
rect 11336 6196 11388 6248
rect 12532 6128 12584 6180
rect 12624 6128 12676 6180
rect 13084 6196 13136 6248
rect 13452 6196 13504 6248
rect 13912 6196 13964 6248
rect 15016 6239 15068 6248
rect 15016 6205 15025 6239
rect 15025 6205 15059 6239
rect 15059 6205 15068 6239
rect 15016 6196 15068 6205
rect 17040 6264 17092 6316
rect 18052 6264 18104 6316
rect 16948 6196 17000 6248
rect 17776 6196 17828 6248
rect 17960 6196 18012 6248
rect 18512 6239 18564 6248
rect 18512 6205 18521 6239
rect 18521 6205 18555 6239
rect 18555 6205 18564 6239
rect 18512 6196 18564 6205
rect 19892 6196 19944 6248
rect 12900 6128 12952 6180
rect 13728 6060 13780 6112
rect 13912 6060 13964 6112
rect 18052 6103 18104 6112
rect 18052 6069 18061 6103
rect 18061 6069 18095 6103
rect 18095 6069 18104 6103
rect 18052 6060 18104 6069
rect 20076 6103 20128 6112
rect 20076 6069 20085 6103
rect 20085 6069 20119 6103
rect 20119 6069 20128 6103
rect 20076 6060 20128 6069
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 2964 5856 3016 5908
rect 1676 5831 1728 5840
rect 1676 5797 1710 5831
rect 1710 5797 1728 5831
rect 1676 5788 1728 5797
rect 3240 5763 3292 5772
rect 3240 5729 3249 5763
rect 3249 5729 3283 5763
rect 3283 5729 3292 5763
rect 3240 5720 3292 5729
rect 3332 5695 3384 5704
rect 3332 5661 3341 5695
rect 3341 5661 3375 5695
rect 3375 5661 3384 5695
rect 3332 5652 3384 5661
rect 5356 5856 5408 5908
rect 5540 5856 5592 5908
rect 3792 5788 3844 5840
rect 5080 5788 5132 5840
rect 5172 5788 5224 5840
rect 6828 5856 6880 5908
rect 7104 5856 7156 5908
rect 7656 5856 7708 5908
rect 7748 5856 7800 5908
rect 8760 5856 8812 5908
rect 9220 5856 9272 5908
rect 9680 5856 9732 5908
rect 11152 5856 11204 5908
rect 4344 5720 4396 5772
rect 5540 5720 5592 5772
rect 7380 5788 7432 5840
rect 5632 5652 5684 5704
rect 5816 5652 5868 5704
rect 6828 5720 6880 5772
rect 9496 5788 9548 5840
rect 12900 5856 12952 5908
rect 13820 5856 13872 5908
rect 11980 5788 12032 5840
rect 12808 5788 12860 5840
rect 7196 5695 7248 5704
rect 4160 5584 4212 5636
rect 7196 5661 7205 5695
rect 7205 5661 7239 5695
rect 7239 5661 7248 5695
rect 7196 5652 7248 5661
rect 7380 5652 7432 5704
rect 7748 5652 7800 5704
rect 8024 5652 8076 5704
rect 8208 5652 8260 5704
rect 2688 5516 2740 5568
rect 5264 5516 5316 5568
rect 11704 5720 11756 5772
rect 20260 5788 20312 5840
rect 8760 5652 8812 5704
rect 9128 5652 9180 5704
rect 8668 5584 8720 5636
rect 7564 5516 7616 5568
rect 10968 5584 11020 5636
rect 11336 5652 11388 5704
rect 11612 5652 11664 5704
rect 11980 5652 12032 5704
rect 12348 5695 12400 5704
rect 12348 5661 12357 5695
rect 12357 5661 12391 5695
rect 12391 5661 12400 5695
rect 12348 5652 12400 5661
rect 15844 5763 15896 5772
rect 15844 5729 15853 5763
rect 15853 5729 15887 5763
rect 15887 5729 15896 5763
rect 15844 5720 15896 5729
rect 16396 5720 16448 5772
rect 17868 5720 17920 5772
rect 18604 5763 18656 5772
rect 18604 5729 18638 5763
rect 18638 5729 18656 5763
rect 18604 5720 18656 5729
rect 13912 5652 13964 5704
rect 17408 5652 17460 5704
rect 14464 5584 14516 5636
rect 19432 5584 19484 5636
rect 11888 5559 11940 5568
rect 11888 5525 11897 5559
rect 11897 5525 11931 5559
rect 11931 5525 11940 5559
rect 11888 5516 11940 5525
rect 12164 5516 12216 5568
rect 13544 5516 13596 5568
rect 16580 5516 16632 5568
rect 17224 5559 17276 5568
rect 17224 5525 17233 5559
rect 17233 5525 17267 5559
rect 17267 5525 17276 5559
rect 17224 5516 17276 5525
rect 17776 5516 17828 5568
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 2412 5312 2464 5364
rect 4068 5244 4120 5296
rect 4160 5244 4212 5296
rect 2780 5176 2832 5228
rect 6368 5219 6420 5228
rect 2872 5151 2924 5160
rect 2872 5117 2881 5151
rect 2881 5117 2915 5151
rect 2915 5117 2924 5151
rect 2872 5108 2924 5117
rect 4068 5108 4120 5160
rect 1676 5083 1728 5092
rect 1676 5049 1710 5083
rect 1710 5049 1728 5083
rect 1676 5040 1728 5049
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 6368 5176 6420 5185
rect 5356 5108 5408 5160
rect 6276 5108 6328 5160
rect 7840 5312 7892 5364
rect 6736 5176 6788 5228
rect 6920 5176 6972 5228
rect 7380 5176 7432 5228
rect 8300 5244 8352 5296
rect 8668 5287 8720 5296
rect 8668 5253 8677 5287
rect 8677 5253 8711 5287
rect 8711 5253 8720 5287
rect 8668 5244 8720 5253
rect 9036 5244 9088 5296
rect 8392 5219 8444 5228
rect 5172 5040 5224 5092
rect 4252 4972 4304 5024
rect 4436 4972 4488 5024
rect 5908 5040 5960 5092
rect 6460 5040 6512 5092
rect 7104 5108 7156 5160
rect 8392 5185 8401 5219
rect 8401 5185 8435 5219
rect 8435 5185 8444 5219
rect 8392 5176 8444 5185
rect 9680 5244 9732 5296
rect 11888 5312 11940 5364
rect 7288 5040 7340 5092
rect 7932 5108 7984 5160
rect 8208 5151 8260 5160
rect 8208 5117 8217 5151
rect 8217 5117 8251 5151
rect 8251 5117 8260 5151
rect 8208 5108 8260 5117
rect 8668 5108 8720 5160
rect 9956 5108 10008 5160
rect 8484 5040 8536 5092
rect 11336 5244 11388 5296
rect 10692 5176 10744 5228
rect 12164 5176 12216 5228
rect 12440 5219 12492 5228
rect 12440 5185 12449 5219
rect 12449 5185 12483 5219
rect 12483 5185 12492 5219
rect 12440 5176 12492 5185
rect 10508 5108 10560 5160
rect 10600 5108 10652 5160
rect 10968 5108 11020 5160
rect 11980 5108 12032 5160
rect 13084 5108 13136 5160
rect 13912 5108 13964 5160
rect 5632 4972 5684 5024
rect 5816 5015 5868 5024
rect 5816 4981 5825 5015
rect 5825 4981 5859 5015
rect 5859 4981 5868 5015
rect 6276 5015 6328 5024
rect 5816 4972 5868 4981
rect 6276 4981 6285 5015
rect 6285 4981 6319 5015
rect 6319 4981 6328 5015
rect 6276 4972 6328 4981
rect 6552 4972 6604 5024
rect 7380 4972 7432 5024
rect 7564 4972 7616 5024
rect 8760 4972 8812 5024
rect 11888 5040 11940 5092
rect 12348 5040 12400 5092
rect 14556 5312 14608 5364
rect 16580 5312 16632 5364
rect 19432 5312 19484 5364
rect 16028 5287 16080 5296
rect 16028 5253 16037 5287
rect 16037 5253 16071 5287
rect 16071 5253 16080 5287
rect 16028 5244 16080 5253
rect 19248 5244 19300 5296
rect 14648 5151 14700 5160
rect 14648 5117 14657 5151
rect 14657 5117 14691 5151
rect 14691 5117 14700 5151
rect 14648 5108 14700 5117
rect 15844 5108 15896 5160
rect 14740 5040 14792 5092
rect 16488 5176 16540 5228
rect 16856 5151 16908 5160
rect 16856 5117 16865 5151
rect 16865 5117 16899 5151
rect 16899 5117 16908 5151
rect 16856 5108 16908 5117
rect 17960 5108 18012 5160
rect 18788 5176 18840 5228
rect 18696 5108 18748 5160
rect 9036 4972 9088 5024
rect 10416 4972 10468 5024
rect 10600 4972 10652 5024
rect 12164 4972 12216 5024
rect 12808 4972 12860 5024
rect 13820 5015 13872 5024
rect 13820 4981 13829 5015
rect 13829 4981 13863 5015
rect 13863 4981 13872 5015
rect 17776 5040 17828 5092
rect 19064 5040 19116 5092
rect 13820 4972 13872 4981
rect 15384 4972 15436 5024
rect 17224 4972 17276 5024
rect 18052 5015 18104 5024
rect 18052 4981 18061 5015
rect 18061 4981 18095 5015
rect 18095 4981 18104 5015
rect 18052 4972 18104 4981
rect 19616 5015 19668 5024
rect 19616 4981 19625 5015
rect 19625 4981 19659 5015
rect 19659 4981 19668 5015
rect 19616 4972 19668 4981
rect 19984 5015 20036 5024
rect 19984 4981 19993 5015
rect 19993 4981 20027 5015
rect 20027 4981 20036 5015
rect 19984 4972 20036 4981
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 3332 4811 3384 4820
rect 3332 4777 3341 4811
rect 3341 4777 3375 4811
rect 3375 4777 3384 4811
rect 3332 4768 3384 4777
rect 4160 4768 4212 4820
rect 5172 4768 5224 4820
rect 5356 4768 5408 4820
rect 6000 4768 6052 4820
rect 6644 4768 6696 4820
rect 7196 4768 7248 4820
rect 7472 4768 7524 4820
rect 5816 4700 5868 4752
rect 2688 4632 2740 4684
rect 4160 4632 4212 4684
rect 5724 4632 5776 4684
rect 3976 4564 4028 4616
rect 5264 4564 5316 4616
rect 2964 4496 3016 4548
rect 3700 4496 3752 4548
rect 5632 4496 5684 4548
rect 5816 4428 5868 4480
rect 6184 4632 6236 4684
rect 6828 4700 6880 4752
rect 7012 4700 7064 4752
rect 6460 4564 6512 4616
rect 6828 4607 6880 4616
rect 6828 4573 6837 4607
rect 6837 4573 6871 4607
rect 6871 4573 6880 4607
rect 6828 4564 6880 4573
rect 6000 4496 6052 4548
rect 6736 4496 6788 4548
rect 6092 4428 6144 4480
rect 7288 4632 7340 4684
rect 7564 4632 7616 4684
rect 8116 4700 8168 4752
rect 9036 4743 9088 4752
rect 9036 4709 9045 4743
rect 9045 4709 9079 4743
rect 9079 4709 9088 4743
rect 9036 4700 9088 4709
rect 9680 4768 9732 4820
rect 10140 4768 10192 4820
rect 10232 4700 10284 4752
rect 10508 4700 10560 4752
rect 11336 4768 11388 4820
rect 20076 4768 20128 4820
rect 11060 4743 11112 4752
rect 11060 4709 11069 4743
rect 11069 4709 11103 4743
rect 11103 4709 11112 4743
rect 11060 4700 11112 4709
rect 11152 4700 11204 4752
rect 13452 4700 13504 4752
rect 13636 4743 13688 4752
rect 13636 4709 13645 4743
rect 13645 4709 13679 4743
rect 13679 4709 13688 4743
rect 13636 4700 13688 4709
rect 15200 4700 15252 4752
rect 7380 4428 7432 4480
rect 7748 4428 7800 4480
rect 7932 4428 7984 4480
rect 8484 4607 8536 4616
rect 8484 4573 8493 4607
rect 8493 4573 8527 4607
rect 8527 4573 8536 4607
rect 8484 4564 8536 4573
rect 8300 4496 8352 4548
rect 9496 4632 9548 4684
rect 10784 4675 10836 4684
rect 9680 4564 9732 4616
rect 10784 4641 10793 4675
rect 10793 4641 10827 4675
rect 10827 4641 10836 4675
rect 10784 4632 10836 4641
rect 11612 4632 11664 4684
rect 11704 4632 11756 4684
rect 13544 4675 13596 4684
rect 11060 4564 11112 4616
rect 13544 4641 13553 4675
rect 13553 4641 13587 4675
rect 13587 4641 13596 4675
rect 13544 4632 13596 4641
rect 17592 4700 17644 4752
rect 10140 4496 10192 4548
rect 11980 4496 12032 4548
rect 12624 4564 12676 4616
rect 13636 4564 13688 4616
rect 13820 4564 13872 4616
rect 14188 4564 14240 4616
rect 16488 4607 16540 4616
rect 16488 4573 16497 4607
rect 16497 4573 16531 4607
rect 16531 4573 16540 4607
rect 16488 4564 16540 4573
rect 17408 4607 17460 4616
rect 17408 4573 17417 4607
rect 17417 4573 17451 4607
rect 17451 4573 17460 4607
rect 17408 4564 17460 4573
rect 14096 4496 14148 4548
rect 15844 4539 15896 4548
rect 15844 4505 15853 4539
rect 15853 4505 15887 4539
rect 15887 4505 15896 4539
rect 15844 4496 15896 4505
rect 9864 4428 9916 4480
rect 12164 4428 12216 4480
rect 17592 4428 17644 4480
rect 18788 4471 18840 4480
rect 18788 4437 18797 4471
rect 18797 4437 18831 4471
rect 18831 4437 18840 4471
rect 18788 4428 18840 4437
rect 21272 4428 21324 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 2320 4224 2372 4276
rect 5724 4267 5776 4276
rect 5724 4233 5733 4267
rect 5733 4233 5767 4267
rect 5767 4233 5776 4267
rect 5724 4224 5776 4233
rect 5816 4224 5868 4276
rect 7288 4224 7340 4276
rect 6092 4156 6144 4208
rect 7104 4156 7156 4208
rect 6368 4131 6420 4140
rect 1492 4020 1544 4072
rect 2964 4020 3016 4072
rect 4160 4020 4212 4072
rect 4436 4020 4488 4072
rect 5172 4020 5224 4072
rect 6368 4097 6377 4131
rect 6377 4097 6411 4131
rect 6411 4097 6420 4131
rect 6368 4088 6420 4097
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 13636 4224 13688 4276
rect 9496 4156 9548 4208
rect 9680 4156 9732 4208
rect 7656 4088 7708 4140
rect 10692 4156 10744 4208
rect 5724 4020 5776 4072
rect 7012 4020 7064 4072
rect 7104 4020 7156 4072
rect 10324 4088 10376 4140
rect 9220 4063 9272 4072
rect 5080 3952 5132 4004
rect 9220 4029 9229 4063
rect 9229 4029 9263 4063
rect 9263 4029 9272 4063
rect 9220 4020 9272 4029
rect 8484 3952 8536 4004
rect 11428 4156 11480 4208
rect 11612 4156 11664 4208
rect 11336 4131 11388 4140
rect 11336 4097 11345 4131
rect 11345 4097 11379 4131
rect 11379 4097 11388 4131
rect 11336 4088 11388 4097
rect 11520 4088 11572 4140
rect 9496 3995 9548 4004
rect 9496 3961 9505 3995
rect 9505 3961 9539 3995
rect 9539 3961 9548 3995
rect 9496 3952 9548 3961
rect 3148 3884 3200 3936
rect 3792 3884 3844 3936
rect 4344 3884 4396 3936
rect 5540 3884 5592 3936
rect 6092 3884 6144 3936
rect 6184 3927 6236 3936
rect 6184 3893 6193 3927
rect 6193 3893 6227 3927
rect 6227 3893 6236 3927
rect 6184 3884 6236 3893
rect 10048 3952 10100 4004
rect 11060 3952 11112 4004
rect 11980 4156 12032 4208
rect 12348 4156 12400 4208
rect 12532 4156 12584 4208
rect 14280 4156 14332 4208
rect 14648 4224 14700 4276
rect 16488 4224 16540 4276
rect 12256 4020 12308 4072
rect 13360 4020 13412 4072
rect 14096 4020 14148 4072
rect 14556 4020 14608 4072
rect 16028 4156 16080 4208
rect 16304 4088 16356 4140
rect 18512 4131 18564 4140
rect 11428 3952 11480 4004
rect 13912 3952 13964 4004
rect 14280 3952 14332 4004
rect 18512 4097 18521 4131
rect 18521 4097 18555 4131
rect 18555 4097 18564 4131
rect 18512 4088 18564 4097
rect 18696 4131 18748 4140
rect 18696 4097 18705 4131
rect 18705 4097 18739 4131
rect 18739 4097 18748 4131
rect 18696 4088 18748 4097
rect 19064 4088 19116 4140
rect 20076 4131 20128 4140
rect 20076 4097 20085 4131
rect 20085 4097 20119 4131
rect 20119 4097 20128 4131
rect 20076 4088 20128 4097
rect 10140 3884 10192 3936
rect 10232 3884 10284 3936
rect 10876 3884 10928 3936
rect 12532 3884 12584 3936
rect 12716 3927 12768 3936
rect 12716 3893 12725 3927
rect 12725 3893 12759 3927
rect 12759 3893 12768 3927
rect 12716 3884 12768 3893
rect 13452 3884 13504 3936
rect 18144 3884 18196 3936
rect 18236 3884 18288 3936
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 2596 3680 2648 3732
rect 1124 3612 1176 3664
rect 2044 3612 2096 3664
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 1952 3544 2004 3596
rect 4528 3612 4580 3664
rect 5356 3612 5408 3664
rect 5724 3612 5776 3664
rect 6368 3612 6420 3664
rect 7104 3680 7156 3732
rect 7288 3680 7340 3732
rect 7748 3680 7800 3732
rect 8392 3680 8444 3732
rect 9588 3680 9640 3732
rect 9956 3680 10008 3732
rect 2872 3544 2924 3596
rect 6552 3544 6604 3596
rect 3332 3519 3384 3528
rect 3332 3485 3341 3519
rect 3341 3485 3375 3519
rect 3375 3485 3384 3519
rect 3332 3476 3384 3485
rect 3424 3519 3476 3528
rect 3424 3485 3433 3519
rect 3433 3485 3467 3519
rect 3467 3485 3476 3519
rect 5816 3519 5868 3528
rect 3424 3476 3476 3485
rect 5816 3485 5825 3519
rect 5825 3485 5859 3519
rect 5859 3485 5868 3519
rect 5816 3476 5868 3485
rect 2780 3451 2832 3460
rect 2780 3417 2789 3451
rect 2789 3417 2823 3451
rect 2823 3417 2832 3451
rect 2780 3408 2832 3417
rect 5724 3408 5776 3460
rect 5448 3383 5500 3392
rect 5448 3349 5457 3383
rect 5457 3349 5491 3383
rect 5491 3349 5500 3383
rect 8208 3612 8260 3664
rect 11612 3680 11664 3732
rect 12256 3680 12308 3732
rect 7288 3544 7340 3596
rect 8852 3544 8904 3596
rect 10232 3544 10284 3596
rect 7380 3476 7432 3528
rect 8116 3476 8168 3528
rect 8668 3476 8720 3528
rect 9864 3476 9916 3528
rect 11612 3544 11664 3596
rect 16120 3680 16172 3732
rect 18512 3680 18564 3732
rect 11980 3544 12032 3596
rect 12164 3587 12216 3596
rect 12164 3553 12173 3587
rect 12173 3553 12207 3587
rect 12207 3553 12216 3587
rect 12164 3544 12216 3553
rect 12532 3587 12584 3596
rect 12532 3553 12541 3587
rect 12541 3553 12575 3587
rect 12575 3553 12584 3587
rect 12532 3544 12584 3553
rect 12808 3587 12860 3596
rect 12808 3553 12817 3587
rect 12817 3553 12851 3587
rect 12851 3553 12860 3587
rect 12808 3544 12860 3553
rect 10508 3476 10560 3528
rect 7564 3408 7616 3460
rect 8944 3408 8996 3460
rect 9588 3408 9640 3460
rect 10876 3408 10928 3460
rect 11796 3476 11848 3528
rect 12348 3476 12400 3528
rect 12716 3476 12768 3528
rect 15200 3612 15252 3664
rect 15384 3612 15436 3664
rect 18052 3612 18104 3664
rect 19708 3612 19760 3664
rect 14096 3587 14148 3596
rect 14096 3553 14105 3587
rect 14105 3553 14139 3587
rect 14139 3553 14148 3587
rect 14096 3544 14148 3553
rect 13728 3476 13780 3528
rect 16948 3544 17000 3596
rect 19340 3544 19392 3596
rect 17960 3476 18012 3528
rect 18144 3519 18196 3528
rect 18144 3485 18153 3519
rect 18153 3485 18187 3519
rect 18187 3485 18196 3519
rect 18144 3476 18196 3485
rect 18788 3476 18840 3528
rect 5448 3340 5500 3349
rect 8208 3340 8260 3392
rect 8760 3340 8812 3392
rect 9956 3340 10008 3392
rect 12164 3340 12216 3392
rect 14096 3408 14148 3460
rect 14004 3340 14056 3392
rect 16120 3340 16172 3392
rect 17500 3340 17552 3392
rect 20352 3340 20404 3392
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 3240 3136 3292 3188
rect 2504 3068 2556 3120
rect 6092 3136 6144 3188
rect 6368 3136 6420 3188
rect 7012 3136 7064 3188
rect 4528 3068 4580 3120
rect 2228 2932 2280 2984
rect 3516 2932 3568 2984
rect 4068 2932 4120 2984
rect 6276 3000 6328 3052
rect 8208 3136 8260 3188
rect 8024 3068 8076 3120
rect 9588 3136 9640 3188
rect 9864 3136 9916 3188
rect 10048 3136 10100 3188
rect 10232 3136 10284 3188
rect 9312 3068 9364 3120
rect 10876 3068 10928 3120
rect 12348 3136 12400 3188
rect 13544 3136 13596 3188
rect 17316 3136 17368 3188
rect 11520 3068 11572 3120
rect 11704 3068 11756 3120
rect 7472 2932 7524 2984
rect 8024 2932 8076 2984
rect 8852 2932 8904 2984
rect 10232 3000 10284 3052
rect 10324 3000 10376 3052
rect 11888 3043 11940 3052
rect 11888 3009 11897 3043
rect 11897 3009 11931 3043
rect 11931 3009 11940 3043
rect 11888 3000 11940 3009
rect 12348 3000 12400 3052
rect 3424 2864 3476 2916
rect 5264 2864 5316 2916
rect 5632 2796 5684 2848
rect 8760 2864 8812 2916
rect 9772 2975 9824 2984
rect 9772 2941 9781 2975
rect 9781 2941 9815 2975
rect 9815 2941 9824 2975
rect 9772 2932 9824 2941
rect 10416 2864 10468 2916
rect 9404 2796 9456 2848
rect 9680 2839 9732 2848
rect 9680 2805 9689 2839
rect 9689 2805 9723 2839
rect 9723 2805 9732 2839
rect 9680 2796 9732 2805
rect 9772 2796 9824 2848
rect 10876 2839 10928 2848
rect 10876 2805 10885 2839
rect 10885 2805 10919 2839
rect 10919 2805 10928 2839
rect 10876 2796 10928 2805
rect 11612 2864 11664 2916
rect 12440 2864 12492 2916
rect 13084 3043 13136 3052
rect 13084 3009 13093 3043
rect 13093 3009 13127 3043
rect 13127 3009 13136 3043
rect 13084 3000 13136 3009
rect 14556 3043 14608 3052
rect 14556 3009 14565 3043
rect 14565 3009 14599 3043
rect 14599 3009 14608 3043
rect 14556 3000 14608 3009
rect 15660 3068 15712 3120
rect 15936 3000 15988 3052
rect 17132 3000 17184 3052
rect 14372 2975 14424 2984
rect 14372 2941 14381 2975
rect 14381 2941 14415 2975
rect 14415 2941 14424 2975
rect 14372 2932 14424 2941
rect 15568 2975 15620 2984
rect 15568 2941 15577 2975
rect 15577 2941 15611 2975
rect 15611 2941 15620 2975
rect 15568 2932 15620 2941
rect 16672 2975 16724 2984
rect 16672 2941 16681 2975
rect 16681 2941 16715 2975
rect 16715 2941 16724 2975
rect 16672 2932 16724 2941
rect 18880 2932 18932 2984
rect 19524 2932 19576 2984
rect 12624 2796 12676 2848
rect 15936 2864 15988 2916
rect 19984 2864 20036 2916
rect 22652 2864 22704 2916
rect 14464 2839 14516 2848
rect 14464 2805 14473 2839
rect 14473 2805 14507 2839
rect 14507 2805 14516 2839
rect 14464 2796 14516 2805
rect 15200 2796 15252 2848
rect 17040 2796 17092 2848
rect 17960 2796 18012 2848
rect 20168 2796 20220 2848
rect 22192 2796 22244 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 2688 2592 2740 2644
rect 4160 2524 4212 2576
rect 4436 2524 4488 2576
rect 5632 2592 5684 2644
rect 5724 2592 5776 2644
rect 6000 2635 6052 2644
rect 6000 2601 6009 2635
rect 6009 2601 6043 2635
rect 6043 2601 6052 2635
rect 6000 2592 6052 2601
rect 7104 2524 7156 2576
rect 7472 2524 7524 2576
rect 7932 2524 7984 2576
rect 8208 2592 8260 2644
rect 9312 2592 9364 2644
rect 8484 2524 8536 2576
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 3240 2499 3292 2508
rect 1400 2456 1452 2465
rect 3240 2465 3249 2499
rect 3249 2465 3283 2499
rect 3283 2465 3292 2499
rect 3240 2456 3292 2465
rect 8024 2456 8076 2508
rect 8668 2524 8720 2576
rect 9864 2592 9916 2644
rect 10140 2592 10192 2644
rect 10600 2635 10652 2644
rect 10600 2601 10609 2635
rect 10609 2601 10643 2635
rect 10643 2601 10652 2635
rect 10600 2592 10652 2601
rect 11060 2635 11112 2644
rect 11060 2601 11069 2635
rect 11069 2601 11103 2635
rect 11103 2601 11112 2635
rect 11060 2592 11112 2601
rect 11152 2592 11204 2644
rect 12624 2635 12676 2644
rect 3332 2431 3384 2440
rect 3332 2397 3341 2431
rect 3341 2397 3375 2431
rect 3375 2397 3384 2431
rect 3332 2388 3384 2397
rect 3424 2431 3476 2440
rect 3424 2397 3433 2431
rect 3433 2397 3467 2431
rect 3467 2397 3476 2431
rect 3700 2431 3752 2440
rect 3424 2388 3476 2397
rect 3700 2397 3709 2431
rect 3709 2397 3743 2431
rect 3743 2397 3752 2431
rect 3700 2388 3752 2397
rect 6092 2431 6144 2440
rect 6092 2397 6101 2431
rect 6101 2397 6135 2431
rect 6135 2397 6144 2431
rect 6092 2388 6144 2397
rect 7932 2388 7984 2440
rect 8852 2456 8904 2508
rect 9036 2456 9088 2508
rect 9220 2499 9272 2508
rect 9220 2465 9229 2499
rect 9229 2465 9263 2499
rect 9263 2465 9272 2499
rect 9220 2456 9272 2465
rect 2780 2295 2832 2304
rect 2780 2261 2789 2295
rect 2789 2261 2823 2295
rect 2823 2261 2832 2295
rect 2780 2252 2832 2261
rect 5080 2252 5132 2304
rect 6552 2295 6604 2304
rect 6552 2261 6561 2295
rect 6561 2261 6595 2295
rect 6595 2261 6604 2295
rect 6552 2252 6604 2261
rect 7564 2252 7616 2304
rect 8668 2388 8720 2440
rect 10416 2524 10468 2576
rect 10876 2524 10928 2576
rect 12624 2601 12633 2635
rect 12633 2601 12667 2635
rect 12667 2601 12676 2635
rect 12624 2592 12676 2601
rect 12716 2592 12768 2644
rect 13820 2592 13872 2644
rect 15384 2592 15436 2644
rect 15936 2635 15988 2644
rect 15936 2601 15945 2635
rect 15945 2601 15979 2635
rect 15979 2601 15988 2635
rect 15936 2592 15988 2601
rect 20168 2635 20220 2644
rect 20168 2601 20177 2635
rect 20177 2601 20211 2635
rect 20211 2601 20220 2635
rect 20168 2592 20220 2601
rect 14740 2524 14792 2576
rect 10048 2456 10100 2508
rect 10232 2499 10284 2508
rect 10232 2465 10241 2499
rect 10241 2465 10275 2499
rect 10275 2465 10284 2499
rect 10232 2456 10284 2465
rect 11060 2456 11112 2508
rect 11796 2499 11848 2508
rect 11796 2465 11805 2499
rect 11805 2465 11839 2499
rect 11839 2465 11848 2499
rect 11796 2456 11848 2465
rect 10324 2431 10376 2440
rect 8852 2320 8904 2372
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 10876 2388 10928 2440
rect 11704 2388 11756 2440
rect 12072 2456 12124 2508
rect 14372 2456 14424 2508
rect 17224 2456 17276 2508
rect 19984 2499 20036 2508
rect 19984 2465 19993 2499
rect 19993 2465 20027 2499
rect 20027 2465 20036 2499
rect 19984 2456 20036 2465
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 12348 2388 12400 2440
rect 14556 2388 14608 2440
rect 9128 2320 9180 2372
rect 8484 2252 8536 2304
rect 8668 2252 8720 2304
rect 11612 2320 11664 2372
rect 13728 2320 13780 2372
rect 15476 2363 15528 2372
rect 9772 2295 9824 2304
rect 9772 2261 9781 2295
rect 9781 2261 9815 2295
rect 9815 2261 9824 2295
rect 9772 2252 9824 2261
rect 10140 2252 10192 2304
rect 13820 2252 13872 2304
rect 14740 2252 14792 2304
rect 15476 2329 15485 2363
rect 15485 2329 15519 2363
rect 15519 2329 15528 2363
rect 15476 2320 15528 2329
rect 19892 2252 19944 2304
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 3700 2048 3752 2100
rect 11796 2048 11848 2100
rect 3240 1912 3292 1964
rect 9680 1980 9732 2032
rect 9772 1980 9824 2032
rect 12992 1980 13044 2032
rect 6552 1912 6604 1964
rect 18420 1912 18472 1964
rect 3332 1844 3384 1896
rect 9864 1844 9916 1896
rect 9956 1844 10008 1896
rect 11980 1844 12032 1896
rect 12256 1844 12308 1896
rect 19984 1844 20036 1896
rect 2780 1776 2832 1828
rect 8760 1776 8812 1828
rect 1584 1708 1636 1760
rect 6828 1708 6880 1760
rect 8484 1708 8536 1760
rect 12164 1776 12216 1828
rect 12808 1776 12860 1828
rect 13268 1776 13320 1828
rect 9496 1708 9548 1760
rect 14372 1708 14424 1760
rect 664 1640 716 1692
rect 8208 1640 8260 1692
rect 8852 1640 8904 1692
rect 10140 1640 10192 1692
rect 14464 1640 14516 1692
rect 2320 1572 2372 1624
rect 11704 1572 11756 1624
rect 204 1504 256 1556
rect 8392 1504 8444 1556
rect 8484 1504 8536 1556
rect 13176 1572 13228 1624
rect 4252 1436 4304 1488
rect 4988 1436 5040 1488
rect 11060 1436 11112 1488
rect 2964 1368 3016 1420
rect 7380 1368 7432 1420
rect 10232 1368 10284 1420
rect 1124 1300 1176 1352
rect 6644 1300 6696 1352
rect 3424 1232 3476 1284
rect 6460 1232 6512 1284
rect 10416 1232 10468 1284
rect 16580 1232 16632 1284
rect 19248 552 19300 604
rect 20812 552 20864 604
<< metal2 >>
rect 202 22520 258 23000
rect 662 22520 718 23000
rect 1122 22520 1178 23000
rect 1582 22520 1638 23000
rect 2042 22520 2098 23000
rect 2502 22520 2558 23000
rect 2962 22522 3018 23000
rect 2962 22520 3280 22522
rect 3422 22520 3478 23000
rect 3882 22520 3938 23000
rect 4066 22672 4122 22681
rect 4122 22630 4200 22658
rect 4066 22607 4122 22616
rect 216 18902 244 22520
rect 204 18896 256 18902
rect 204 18838 256 18844
rect 676 18766 704 22520
rect 664 18760 716 18766
rect 664 18702 716 18708
rect 1136 18698 1164 22520
rect 1492 19304 1544 19310
rect 1492 19246 1544 19252
rect 1124 18692 1176 18698
rect 1124 18634 1176 18640
rect 1504 18057 1532 19246
rect 1596 19145 1624 22520
rect 1950 20768 2006 20777
rect 1950 20703 2006 20712
rect 1964 20058 1992 20703
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 1860 19916 1912 19922
rect 1860 19858 1912 19864
rect 1582 19136 1638 19145
rect 1582 19071 1638 19080
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 1676 18420 1728 18426
rect 1676 18362 1728 18368
rect 1490 18048 1546 18057
rect 1490 17983 1546 17992
rect 1400 15428 1452 15434
rect 1400 15370 1452 15376
rect 1308 12436 1360 12442
rect 1308 12378 1360 12384
rect 1216 9444 1268 9450
rect 1216 9386 1268 9392
rect 1124 8628 1176 8634
rect 1124 8570 1176 8576
rect 1032 7268 1084 7274
rect 1032 7210 1084 7216
rect 1044 2553 1072 7210
rect 1136 3670 1164 8570
rect 1228 6662 1256 9386
rect 1320 9110 1348 12378
rect 1412 9330 1440 15370
rect 1688 15314 1716 18362
rect 1596 15286 1716 15314
rect 1492 14952 1544 14958
rect 1492 14894 1544 14900
rect 1504 14414 1532 14894
rect 1492 14408 1544 14414
rect 1492 14350 1544 14356
rect 1504 13870 1532 14350
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 1504 11694 1532 13806
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 1492 11280 1544 11286
rect 1492 11222 1544 11228
rect 1504 9450 1532 11222
rect 1492 9444 1544 9450
rect 1492 9386 1544 9392
rect 1412 9302 1532 9330
rect 1308 9104 1360 9110
rect 1308 9046 1360 9052
rect 1400 7744 1452 7750
rect 1400 7686 1452 7692
rect 1308 7200 1360 7206
rect 1308 7142 1360 7148
rect 1320 7002 1348 7142
rect 1308 6996 1360 7002
rect 1308 6938 1360 6944
rect 1308 6792 1360 6798
rect 1308 6734 1360 6740
rect 1216 6656 1268 6662
rect 1216 6598 1268 6604
rect 1320 6458 1348 6734
rect 1308 6452 1360 6458
rect 1308 6394 1360 6400
rect 1412 5681 1440 7686
rect 1398 5672 1454 5681
rect 1398 5607 1454 5616
rect 1504 4078 1532 9302
rect 1596 9178 1624 15286
rect 1676 15088 1728 15094
rect 1676 15030 1728 15036
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1124 3664 1176 3670
rect 1124 3606 1176 3612
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 1030 2544 1086 2553
rect 1412 2514 1440 3538
rect 1596 3097 1624 7686
rect 1688 5846 1716 15030
rect 1780 12442 1808 18770
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 1872 10418 1900 19858
rect 2056 18290 2084 22520
rect 2136 19372 2188 19378
rect 2136 19314 2188 19320
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 2044 17604 2096 17610
rect 2044 17546 2096 17552
rect 2056 17134 2084 17546
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 1952 15156 2004 15162
rect 1952 15098 2004 15104
rect 1780 10390 1900 10418
rect 1780 9897 1808 10390
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 1766 9888 1822 9897
rect 1766 9823 1822 9832
rect 1872 9602 1900 10202
rect 1964 9722 1992 15098
rect 2056 14958 2084 17070
rect 2148 15094 2176 19314
rect 2516 18358 2544 22520
rect 2976 22494 3280 22520
rect 2870 22128 2926 22137
rect 2870 22063 2926 22072
rect 2778 21720 2834 21729
rect 2778 21655 2834 21664
rect 2688 20256 2740 20262
rect 2688 20198 2740 20204
rect 2700 19378 2728 20198
rect 2688 19372 2740 19378
rect 2688 19314 2740 19320
rect 2792 19242 2820 21655
rect 2780 19236 2832 19242
rect 2780 19178 2832 19184
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 2504 18352 2556 18358
rect 2504 18294 2556 18300
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2228 15360 2280 15366
rect 2228 15302 2280 15308
rect 2136 15088 2188 15094
rect 2136 15030 2188 15036
rect 2044 14952 2096 14958
rect 2044 14894 2096 14900
rect 2136 14816 2188 14822
rect 2136 14758 2188 14764
rect 2148 12481 2176 14758
rect 2134 12472 2190 12481
rect 2134 12407 2190 12416
rect 2044 12368 2096 12374
rect 2044 12310 2096 12316
rect 2056 11286 2084 12310
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2044 11280 2096 11286
rect 2044 11222 2096 11228
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 1952 9716 2004 9722
rect 1952 9658 2004 9664
rect 1872 9574 1992 9602
rect 1858 9480 1914 9489
rect 1858 9415 1914 9424
rect 1872 9382 1900 9415
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1858 9072 1914 9081
rect 1768 9036 1820 9042
rect 1858 9007 1860 9016
rect 1768 8978 1820 8984
rect 1912 9007 1914 9016
rect 1860 8978 1912 8984
rect 1780 7546 1808 8978
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1872 7857 1900 8842
rect 1964 8090 1992 9574
rect 2056 9518 2084 11086
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 2148 9382 2176 12242
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 2148 8673 2176 8910
rect 2134 8664 2190 8673
rect 2134 8599 2190 8608
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1858 7848 1914 7857
rect 1858 7783 1914 7792
rect 2042 7848 2098 7857
rect 2042 7783 2098 7792
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1766 7440 1822 7449
rect 1766 7375 1822 7384
rect 1780 7342 1808 7375
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 2056 7206 2084 7783
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 1860 7200 1912 7206
rect 1860 7142 1912 7148
rect 2044 7200 2096 7206
rect 2148 7177 2176 7482
rect 2044 7142 2096 7148
rect 2134 7168 2190 7177
rect 1872 6497 1900 7142
rect 2134 7103 2190 7112
rect 1858 6488 1914 6497
rect 1858 6423 1914 6432
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 1676 5840 1728 5846
rect 1676 5782 1728 5788
rect 1676 5092 1728 5098
rect 1676 5034 1728 5040
rect 1688 4729 1716 5034
rect 1674 4720 1730 4729
rect 1674 4655 1730 4664
rect 1964 3602 1992 6190
rect 2136 6180 2188 6186
rect 2136 6122 2188 6128
rect 2148 4593 2176 6122
rect 2134 4584 2190 4593
rect 2134 4519 2190 4528
rect 2044 3664 2096 3670
rect 2044 3606 2096 3612
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1582 3088 1638 3097
rect 1582 3023 1638 3032
rect 1030 2479 1086 2488
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1584 1760 1636 1766
rect 1584 1702 1636 1708
rect 664 1692 716 1698
rect 664 1634 716 1640
rect 204 1556 256 1562
rect 204 1498 256 1504
rect 216 480 244 1498
rect 676 480 704 1634
rect 1124 1352 1176 1358
rect 1124 1294 1176 1300
rect 1136 480 1164 1294
rect 1596 480 1624 1702
rect 2056 480 2084 3606
rect 2240 3074 2268 15302
rect 2332 13462 2360 18158
rect 2608 18154 2636 18362
rect 2596 18148 2648 18154
rect 2596 18090 2648 18096
rect 2502 18048 2558 18057
rect 2502 17983 2558 17992
rect 2412 17672 2464 17678
rect 2410 17640 2412 17649
rect 2464 17640 2466 17649
rect 2410 17575 2466 17584
rect 2412 17536 2464 17542
rect 2412 17478 2464 17484
rect 2424 16114 2452 17478
rect 2516 17134 2544 17983
rect 2504 17128 2556 17134
rect 2504 17070 2556 17076
rect 2504 16992 2556 16998
rect 2504 16934 2556 16940
rect 2412 16108 2464 16114
rect 2412 16050 2464 16056
rect 2516 14822 2544 16934
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 2504 14816 2556 14822
rect 2502 14784 2504 14793
rect 2556 14784 2558 14793
rect 2502 14719 2558 14728
rect 2320 13456 2372 13462
rect 2320 13398 2372 13404
rect 2412 13456 2464 13462
rect 2412 13398 2464 13404
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2332 10606 2360 11086
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 2332 10033 2360 10542
rect 2318 10024 2374 10033
rect 2318 9959 2374 9968
rect 2318 9480 2374 9489
rect 2318 9415 2320 9424
rect 2372 9415 2374 9424
rect 2320 9386 2372 9392
rect 2318 9208 2374 9217
rect 2318 9143 2374 9152
rect 2332 8537 2360 9143
rect 2318 8528 2374 8537
rect 2318 8463 2374 8472
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2332 4282 2360 7890
rect 2424 7546 2452 13398
rect 2608 12850 2636 15574
rect 2596 12844 2648 12850
rect 2596 12786 2648 12792
rect 2700 12374 2728 19110
rect 2884 18970 2912 22063
rect 3054 21176 3110 21185
rect 3054 21111 3110 21120
rect 3068 20058 3096 21111
rect 3146 20224 3202 20233
rect 3146 20159 3202 20168
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 2872 18964 2924 18970
rect 2872 18906 2924 18912
rect 2872 18624 2924 18630
rect 2872 18566 2924 18572
rect 2780 18080 2832 18086
rect 2780 18022 2832 18028
rect 2792 13569 2820 18022
rect 2884 14521 2912 18566
rect 2976 16454 3004 19110
rect 3160 18222 3188 20159
rect 3252 19009 3280 22494
rect 3436 19310 3464 22520
rect 3792 20052 3844 20058
rect 3792 19994 3844 20000
rect 3516 19916 3568 19922
rect 3516 19858 3568 19864
rect 3608 19916 3660 19922
rect 3608 19858 3660 19864
rect 3424 19304 3476 19310
rect 3330 19272 3386 19281
rect 3424 19246 3476 19252
rect 3330 19207 3386 19216
rect 3344 19156 3372 19207
rect 3344 19128 3464 19156
rect 3238 19000 3294 19009
rect 3238 18935 3294 18944
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 3148 18080 3200 18086
rect 3148 18022 3200 18028
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 3068 15609 3096 15982
rect 3054 15600 3110 15609
rect 3054 15535 3110 15544
rect 3056 15496 3108 15502
rect 2962 15464 3018 15473
rect 3056 15438 3108 15444
rect 2962 15399 3018 15408
rect 2870 14512 2926 14521
rect 2870 14447 2926 14456
rect 2872 13728 2924 13734
rect 2872 13670 2924 13676
rect 2778 13560 2834 13569
rect 2778 13495 2834 13504
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2792 12986 2820 13330
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 2884 12918 2912 13670
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2780 12844 2832 12850
rect 2780 12786 2832 12792
rect 2688 12368 2740 12374
rect 2792 12345 2820 12786
rect 2688 12310 2740 12316
rect 2778 12336 2834 12345
rect 2778 12271 2834 12280
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 2780 12232 2832 12238
rect 2780 12174 2832 12180
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2504 10532 2556 10538
rect 2504 10474 2556 10480
rect 2516 10062 2544 10474
rect 2608 10305 2636 11290
rect 2700 10470 2728 12174
rect 2688 10464 2740 10470
rect 2688 10406 2740 10412
rect 2594 10296 2650 10305
rect 2594 10231 2650 10240
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2516 8294 2544 9998
rect 2608 9654 2636 10231
rect 2700 10198 2728 10406
rect 2688 10192 2740 10198
rect 2688 10134 2740 10140
rect 2686 10024 2742 10033
rect 2686 9959 2742 9968
rect 2596 9648 2648 9654
rect 2596 9590 2648 9596
rect 2700 9586 2728 9959
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2608 9217 2636 9318
rect 2594 9208 2650 9217
rect 2792 9160 2820 12174
rect 2884 11626 2912 12854
rect 2976 12646 3004 15399
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 3068 12102 3096 15438
rect 3160 14249 3188 18022
rect 3344 17338 3372 18022
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3238 17096 3294 17105
rect 3238 17031 3294 17040
rect 3252 15162 3280 17031
rect 3436 16946 3464 19128
rect 3344 16918 3464 16946
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 3344 15042 3372 16918
rect 3528 16590 3556 19858
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3516 16448 3568 16454
rect 3516 16390 3568 16396
rect 3528 16153 3556 16390
rect 3514 16144 3570 16153
rect 3514 16079 3570 16088
rect 3422 15872 3478 15881
rect 3422 15807 3478 15816
rect 3252 15014 3372 15042
rect 3146 14240 3202 14249
rect 3146 14175 3202 14184
rect 3146 14104 3202 14113
rect 3146 14039 3148 14048
rect 3200 14039 3202 14048
rect 3148 14010 3200 14016
rect 3252 13841 3280 15014
rect 3332 14884 3384 14890
rect 3332 14826 3384 14832
rect 3238 13832 3294 13841
rect 3238 13767 3294 13776
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3160 12782 3188 13126
rect 3252 12850 3280 13670
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 2872 11620 2924 11626
rect 2872 11562 2924 11568
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2594 9143 2650 9152
rect 2700 9132 2820 9160
rect 2596 9104 2648 9110
rect 2596 9046 2648 9052
rect 2608 8498 2636 9046
rect 2700 8974 2728 9132
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2594 8392 2650 8401
rect 2594 8327 2650 8336
rect 2504 8288 2556 8294
rect 2504 8230 2556 8236
rect 2504 7812 2556 7818
rect 2504 7754 2556 7760
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2412 7268 2464 7274
rect 2412 7210 2464 7216
rect 2424 5370 2452 7210
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2320 4276 2372 4282
rect 2320 4218 2372 4224
rect 2318 3496 2374 3505
rect 2318 3431 2374 3440
rect 2148 3046 2268 3074
rect 2148 2417 2176 3046
rect 2228 2984 2280 2990
rect 2226 2952 2228 2961
rect 2280 2952 2282 2961
rect 2226 2887 2282 2896
rect 2134 2408 2190 2417
rect 2134 2343 2190 2352
rect 2332 1630 2360 3431
rect 2320 1624 2372 1630
rect 2320 1566 2372 1572
rect 2424 649 2452 5306
rect 2516 5137 2544 7754
rect 2608 7750 2636 8327
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 2608 7410 2636 7686
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2700 7154 2728 8774
rect 2792 7546 2820 8978
rect 2884 8430 2912 9862
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2884 7886 2912 8366
rect 2976 8022 3004 12038
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 3068 11150 3096 11834
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 2964 8016 3016 8022
rect 2964 7958 3016 7964
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2870 7576 2926 7585
rect 2780 7540 2832 7546
rect 2870 7511 2926 7520
rect 2780 7482 2832 7488
rect 2608 7126 2728 7154
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2502 5128 2558 5137
rect 2502 5063 2558 5072
rect 2608 3738 2636 7126
rect 2792 7018 2820 7142
rect 2700 6990 2820 7018
rect 2700 6186 2728 6990
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2792 6662 2820 6734
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2688 6180 2740 6186
rect 2688 6122 2740 6128
rect 2700 5574 2728 6122
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 2792 5234 2820 6598
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2884 5166 2912 7511
rect 2976 6866 3004 7686
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2962 6760 3018 6769
rect 2962 6695 3018 6704
rect 2976 5914 3004 6695
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2504 3120 2556 3126
rect 2502 3088 2504 3097
rect 2556 3088 2558 3097
rect 2502 3023 2558 3032
rect 2700 2650 2728 4626
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2870 4176 2926 4185
rect 2870 4111 2926 4120
rect 2884 3602 2912 4111
rect 2976 4078 3004 4490
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2778 3496 2834 3505
rect 2778 3431 2780 3440
rect 2832 3431 2834 3440
rect 2780 3402 2832 3408
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 2792 1834 2820 2246
rect 2780 1828 2832 1834
rect 2780 1770 2832 1776
rect 2502 1456 2558 1465
rect 2502 1391 2558 1400
rect 2964 1420 3016 1426
rect 2410 640 2466 649
rect 2410 575 2466 584
rect 2516 480 2544 1391
rect 2964 1362 3016 1368
rect 2976 480 3004 1362
rect 3068 1193 3096 10746
rect 3160 3942 3188 12582
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 3252 9654 3280 11154
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 3252 7274 3280 9590
rect 3344 9178 3372 14826
rect 3436 12646 3464 15807
rect 3528 15586 3556 16079
rect 3620 15706 3648 19858
rect 3804 19825 3832 19994
rect 3790 19816 3846 19825
rect 3790 19751 3846 19760
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 3700 18692 3752 18698
rect 3700 18634 3752 18640
rect 3712 17785 3740 18634
rect 3698 17776 3754 17785
rect 3698 17711 3754 17720
rect 3804 16697 3832 18702
rect 3896 18086 3924 22520
rect 4172 20602 4200 22630
rect 4342 22520 4398 23000
rect 4894 22520 4950 23000
rect 5354 22520 5410 23000
rect 5814 22520 5870 23000
rect 6274 22520 6330 23000
rect 6734 22520 6790 23000
rect 7194 22520 7250 23000
rect 7654 22520 7710 23000
rect 8114 22520 8170 23000
rect 8574 22520 8630 23000
rect 9034 22520 9090 23000
rect 9586 22520 9642 23000
rect 10046 22520 10102 23000
rect 10506 22520 10562 23000
rect 10966 22520 11022 23000
rect 11426 22520 11482 23000
rect 11886 22520 11942 23000
rect 12346 22520 12402 23000
rect 12806 22520 12862 23000
rect 13266 22520 13322 23000
rect 13726 22520 13782 23000
rect 14278 22520 14334 23000
rect 14738 22520 14794 23000
rect 15198 22520 15254 23000
rect 15658 22520 15714 23000
rect 16118 22520 16174 23000
rect 16578 22520 16634 23000
rect 17038 22520 17094 23000
rect 17498 22520 17554 23000
rect 17958 22520 18014 23000
rect 18418 22520 18474 23000
rect 18970 22520 19026 23000
rect 19430 22520 19486 23000
rect 19890 22520 19946 23000
rect 20350 22520 20406 23000
rect 20810 22520 20866 23000
rect 21270 22520 21326 23000
rect 21730 22520 21786 23000
rect 22190 22520 22246 23000
rect 22650 22520 22706 23000
rect 4160 20596 4212 20602
rect 4160 20538 4212 20544
rect 3976 20392 4028 20398
rect 3976 20334 4028 20340
rect 4160 20392 4212 20398
rect 4160 20334 4212 20340
rect 3988 19310 4016 20334
rect 4066 19816 4122 19825
rect 4066 19751 4068 19760
rect 4120 19751 4122 19760
rect 4068 19722 4120 19728
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3988 18222 4016 19246
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 4080 18329 4108 19110
rect 4066 18320 4122 18329
rect 4066 18255 4122 18264
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 3884 18080 3936 18086
rect 3884 18022 3936 18028
rect 3988 17610 4016 18158
rect 4066 17912 4122 17921
rect 4066 17847 4122 17856
rect 4080 17814 4108 17847
rect 4068 17808 4120 17814
rect 4068 17750 4120 17756
rect 3976 17604 4028 17610
rect 3976 17546 4028 17552
rect 4066 17368 4122 17377
rect 4066 17303 4122 17312
rect 4080 16833 4108 17303
rect 4066 16824 4122 16833
rect 4066 16759 4122 16768
rect 4172 16776 4200 20334
rect 4356 19938 4384 22520
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 4620 20324 4672 20330
rect 4620 20266 4672 20272
rect 4264 19910 4384 19938
rect 4528 19916 4580 19922
rect 4264 19242 4292 19910
rect 4528 19858 4580 19864
rect 4540 19700 4568 19858
rect 4632 19854 4660 20266
rect 4620 19848 4672 19854
rect 4620 19790 4672 19796
rect 4356 19672 4568 19700
rect 4252 19236 4304 19242
rect 4252 19178 4304 19184
rect 4252 18828 4304 18834
rect 4252 18770 4304 18776
rect 4264 18737 4292 18770
rect 4250 18728 4306 18737
rect 4250 18663 4306 18672
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 4264 18290 4292 18566
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 4264 16946 4292 18022
rect 4356 17338 4384 19672
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4618 19272 4674 19281
rect 4618 19207 4674 19216
rect 4632 18766 4660 19207
rect 4908 19122 4936 22520
rect 5170 19544 5226 19553
rect 5170 19479 5226 19488
rect 4908 19094 5120 19122
rect 4724 18924 5028 18952
rect 4724 18834 4752 18924
rect 4712 18828 4764 18834
rect 4712 18770 4764 18776
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4816 17746 4844 18702
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4816 17202 4844 17682
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 4264 16918 4384 16946
rect 4356 16794 4384 16918
rect 4344 16788 4396 16794
rect 4172 16748 4292 16776
rect 3790 16688 3846 16697
rect 3790 16623 3846 16632
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 3976 16176 4028 16182
rect 3976 16118 4028 16124
rect 3988 16017 4016 16118
rect 3974 16008 4030 16017
rect 3700 15972 3752 15978
rect 3974 15943 4030 15952
rect 3700 15914 3752 15920
rect 3608 15700 3660 15706
rect 3608 15642 3660 15648
rect 3528 15558 3648 15586
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 3528 12238 3556 14962
rect 3620 14906 3648 15558
rect 3712 15473 3740 15914
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 3698 15464 3754 15473
rect 3698 15399 3754 15408
rect 3790 15056 3846 15065
rect 3790 14991 3846 15000
rect 3620 14878 3740 14906
rect 3606 14784 3662 14793
rect 3606 14719 3662 14728
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3344 8294 3372 8366
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3344 7818 3372 8230
rect 3332 7812 3384 7818
rect 3332 7754 3384 7760
rect 3344 7585 3372 7754
rect 3330 7576 3386 7585
rect 3330 7511 3386 7520
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3252 6089 3280 6598
rect 3344 6458 3372 6802
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3238 6080 3294 6089
rect 3238 6015 3294 6024
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 3252 3194 3280 5714
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3344 5545 3372 5646
rect 3330 5536 3386 5545
rect 3330 5471 3386 5480
rect 3330 4856 3386 4865
rect 3330 4791 3332 4800
rect 3384 4791 3386 4800
rect 3332 4762 3384 4768
rect 3436 3534 3464 12038
rect 3528 11762 3556 12174
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3620 11642 3648 14719
rect 3528 11614 3648 11642
rect 3332 3528 3384 3534
rect 3330 3496 3332 3505
rect 3424 3528 3476 3534
rect 3384 3496 3386 3505
rect 3424 3470 3476 3476
rect 3330 3431 3386 3440
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3436 2922 3464 3470
rect 3528 2990 3556 11614
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3620 10606 3648 11222
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3620 9926 3648 10406
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3620 9178 3648 9318
rect 3712 9217 3740 14878
rect 3804 14006 3832 14991
rect 3792 14000 3844 14006
rect 3792 13942 3844 13948
rect 3790 13696 3846 13705
rect 3790 13631 3846 13640
rect 3698 9208 3754 9217
rect 3608 9172 3660 9178
rect 3698 9143 3754 9152
rect 3608 9114 3660 9120
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 3620 8566 3648 8978
rect 3608 8560 3660 8566
rect 3608 8502 3660 8508
rect 3698 8528 3754 8537
rect 3620 7206 3648 8502
rect 3698 8463 3754 8472
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3606 7032 3662 7041
rect 3606 6967 3608 6976
rect 3660 6967 3662 6976
rect 3608 6938 3660 6944
rect 3712 6905 3740 8463
rect 3698 6896 3754 6905
rect 3698 6831 3754 6840
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3712 6322 3740 6734
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3804 6202 3832 13631
rect 3896 10044 3924 15506
rect 3976 14476 4028 14482
rect 3976 14418 4028 14424
rect 3988 14249 4016 14418
rect 3974 14240 4030 14249
rect 3974 14175 4030 14184
rect 4080 13938 4108 16390
rect 4172 16250 4200 16594
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 4172 13802 4200 14214
rect 4160 13796 4212 13802
rect 4160 13738 4212 13744
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 3988 11354 4016 13466
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4172 12646 4200 13126
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 4172 11558 4200 12106
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 4172 11150 4200 11494
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 3988 10169 4016 10678
rect 4160 10532 4212 10538
rect 4160 10474 4212 10480
rect 3974 10160 4030 10169
rect 3974 10095 4030 10104
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 3896 10016 4016 10044
rect 3882 9888 3938 9897
rect 3882 9823 3938 9832
rect 3896 9518 3924 9823
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3712 6174 3832 6202
rect 3606 5400 3662 5409
rect 3606 5335 3662 5344
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3424 2916 3476 2922
rect 3424 2858 3476 2864
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 3252 1970 3280 2450
rect 3436 2446 3464 2858
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 3424 2440 3476 2446
rect 3424 2382 3476 2388
rect 3240 1964 3292 1970
rect 3240 1906 3292 1912
rect 3344 1902 3372 2382
rect 3620 2009 3648 5335
rect 3712 4554 3740 6174
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3804 5846 3832 6054
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3790 4720 3846 4729
rect 3790 4655 3846 4664
rect 3700 4548 3752 4554
rect 3700 4490 3752 4496
rect 3804 3942 3832 4655
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3700 2440 3752 2446
rect 3700 2382 3752 2388
rect 3712 2106 3740 2382
rect 3700 2100 3752 2106
rect 3700 2042 3752 2048
rect 3606 2000 3662 2009
rect 3606 1935 3662 1944
rect 3332 1896 3384 1902
rect 3332 1838 3384 1844
rect 3424 1284 3476 1290
rect 3424 1226 3476 1232
rect 3054 1184 3110 1193
rect 3054 1119 3110 1128
rect 3436 480 3464 1226
rect 3896 480 3924 9318
rect 3988 8906 4016 10016
rect 3976 8900 4028 8906
rect 3976 8842 4028 8848
rect 3974 7984 4030 7993
rect 3974 7919 4030 7928
rect 3988 6361 4016 7919
rect 4080 6662 4108 10066
rect 4172 9178 4200 10474
rect 4264 10198 4292 16748
rect 4344 16730 4396 16736
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4436 15972 4488 15978
rect 4436 15914 4488 15920
rect 4448 15706 4476 15914
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4710 14512 4766 14521
rect 4710 14447 4712 14456
rect 4764 14447 4766 14456
rect 4712 14418 4764 14424
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4344 13388 4396 13394
rect 4344 13330 4396 13336
rect 4356 12986 4384 13330
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 4344 12640 4396 12646
rect 4448 12617 4476 12854
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4344 12582 4396 12588
rect 4434 12608 4490 12617
rect 4356 12374 4384 12582
rect 4434 12543 4490 12552
rect 4344 12368 4396 12374
rect 4344 12310 4396 12316
rect 4344 12096 4396 12102
rect 4540 12084 4568 12786
rect 4804 12368 4856 12374
rect 4804 12310 4856 12316
rect 4396 12056 4568 12084
rect 4344 12038 4396 12044
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4356 10044 4384 12038
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4816 11665 4844 12310
rect 4908 11694 4936 18770
rect 5000 17338 5028 18924
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 4988 16992 5040 16998
rect 4986 16960 4988 16969
rect 5040 16960 5042 16969
rect 4986 16895 5042 16904
rect 5092 16794 5120 19094
rect 5184 18193 5212 19479
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 5170 18184 5226 18193
rect 5170 18119 5226 18128
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 5000 14890 5028 16526
rect 5184 15706 5212 17274
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 4988 14884 5040 14890
rect 4988 14826 5040 14832
rect 5000 14414 5028 14826
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 5000 12850 5028 14350
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4986 12472 5042 12481
rect 4986 12407 5042 12416
rect 4896 11688 4948 11694
rect 4618 11656 4674 11665
rect 4618 11591 4674 11600
rect 4802 11656 4858 11665
rect 4896 11630 4948 11636
rect 4802 11591 4858 11600
rect 4632 11354 4660 11591
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4264 10016 4384 10044
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4158 8936 4214 8945
rect 4158 8871 4160 8880
rect 4212 8871 4214 8880
rect 4160 8842 4212 8848
rect 4158 8800 4214 8809
rect 4158 8735 4214 8744
rect 4172 6746 4200 8735
rect 4264 7410 4292 10016
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4356 8090 4384 9862
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4526 9480 4582 9489
rect 4526 9415 4582 9424
rect 4434 9344 4490 9353
rect 4434 9279 4490 9288
rect 4448 9042 4476 9279
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4540 8974 4568 9415
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4632 9110 4660 9318
rect 4710 9208 4766 9217
rect 4710 9143 4712 9152
rect 4764 9143 4766 9152
rect 4712 9114 4764 9120
rect 4620 9104 4672 9110
rect 4620 9046 4672 9052
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4448 7857 4476 8298
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4632 7857 4660 7890
rect 4434 7848 4490 7857
rect 4356 7806 4434 7834
rect 4356 7410 4384 7806
rect 4434 7783 4490 7792
rect 4618 7848 4674 7857
rect 4618 7783 4674 7792
rect 4724 7732 4752 8230
rect 4816 8090 4844 11494
rect 5000 11370 5028 12407
rect 5092 12374 5120 14418
rect 5184 13938 5212 14758
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 5184 13326 5212 13874
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5080 12368 5132 12374
rect 5080 12310 5132 12316
rect 5184 11558 5212 12582
rect 5276 12481 5304 18566
rect 5368 17134 5396 22520
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 5632 20256 5684 20262
rect 5632 20198 5684 20204
rect 5644 19990 5672 20198
rect 5632 19984 5684 19990
rect 5632 19926 5684 19932
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 5552 19514 5580 19790
rect 5540 19508 5592 19514
rect 5540 19450 5592 19456
rect 5644 19417 5672 19790
rect 5630 19408 5686 19417
rect 5630 19343 5686 19352
rect 5736 19281 5764 20402
rect 5722 19272 5778 19281
rect 5448 19236 5500 19242
rect 5722 19207 5778 19216
rect 5448 19178 5500 19184
rect 5460 17542 5488 19178
rect 5538 18864 5594 18873
rect 5538 18799 5594 18808
rect 5552 18170 5580 18799
rect 5722 18728 5778 18737
rect 5722 18663 5778 18672
rect 5632 18624 5684 18630
rect 5632 18566 5684 18572
rect 5644 18290 5672 18566
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5552 18142 5672 18170
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5460 17202 5488 17478
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5356 17128 5408 17134
rect 5356 17070 5408 17076
rect 5354 16824 5410 16833
rect 5354 16759 5410 16768
rect 5368 16289 5396 16759
rect 5354 16280 5410 16289
rect 5354 16215 5410 16224
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5368 15881 5396 16050
rect 5354 15872 5410 15881
rect 5354 15807 5410 15816
rect 5552 15706 5580 17614
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5368 13190 5396 14758
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 5262 12472 5318 12481
rect 5262 12407 5318 12416
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 5276 11762 5304 12242
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5262 11656 5318 11665
rect 5262 11591 5264 11600
rect 5316 11591 5318 11600
rect 5264 11562 5316 11568
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 4908 11342 5028 11370
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4908 7954 4936 11342
rect 4988 11280 5040 11286
rect 4988 11222 5040 11228
rect 5000 8906 5028 11222
rect 5184 10810 5212 11494
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5172 9036 5224 9042
rect 5092 8996 5172 9024
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 5000 8634 5028 8842
rect 5092 8809 5120 8996
rect 5172 8978 5224 8984
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5078 8800 5134 8809
rect 5078 8735 5134 8744
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 5000 7834 5028 8434
rect 5184 8362 5212 8842
rect 5276 8786 5304 11562
rect 5368 8974 5396 12650
rect 5460 12238 5488 15642
rect 5644 15586 5672 18142
rect 5736 17377 5764 18663
rect 5722 17368 5778 17377
rect 5722 17303 5778 17312
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 5736 16794 5764 17138
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 5552 15558 5672 15586
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5460 12073 5488 12174
rect 5446 12064 5502 12073
rect 5446 11999 5502 12008
rect 5446 11248 5502 11257
rect 5446 11183 5502 11192
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5276 8758 5396 8786
rect 5264 8560 5316 8566
rect 5264 8502 5316 8508
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 8072 5120 8230
rect 5276 8090 5304 8502
rect 5264 8084 5316 8090
rect 5092 8044 5212 8072
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 4908 7806 5028 7834
rect 4724 7704 4844 7732
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 4816 6934 4844 7704
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 4172 6718 4292 6746
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4160 6656 4212 6662
rect 4264 6633 4292 6718
rect 4804 6656 4856 6662
rect 4160 6598 4212 6604
rect 4250 6624 4306 6633
rect 4066 6488 4122 6497
rect 4066 6423 4122 6432
rect 3974 6352 4030 6361
rect 3974 6287 4030 6296
rect 3974 5944 4030 5953
rect 3974 5879 4030 5888
rect 3988 4622 4016 5879
rect 4080 5302 4108 6423
rect 4172 5642 4200 6598
rect 4804 6598 4856 6604
rect 4250 6559 4306 6568
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4816 6458 4844 6598
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4344 6248 4396 6254
rect 4396 6225 4476 6236
rect 4396 6216 4490 6225
rect 4396 6208 4434 6216
rect 4344 6190 4396 6196
rect 4434 6151 4490 6160
rect 4344 5772 4396 5778
rect 4540 5760 4568 6258
rect 4620 6180 4672 6186
rect 4672 6140 4844 6168
rect 4620 6122 4672 6128
rect 4396 5732 4568 5760
rect 4344 5714 4396 5720
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 4250 5264 4306 5273
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 4080 2990 4108 5102
rect 4172 4826 4200 5238
rect 4250 5199 4306 5208
rect 4264 5030 4292 5199
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4160 4684 4212 4690
rect 4356 4672 4384 5714
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4212 4644 4384 4672
rect 4160 4626 4212 4632
rect 4172 4078 4200 4626
rect 4448 4604 4476 4966
rect 4264 4576 4476 4604
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 4160 2576 4212 2582
rect 4264 2564 4292 4576
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4816 4321 4844 6140
rect 4802 4312 4858 4321
rect 4802 4247 4858 4256
rect 4436 4072 4488 4078
rect 4436 4014 4488 4020
rect 4526 4040 4582 4049
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4212 2536 4292 2564
rect 4160 2518 4212 2524
rect 4250 2136 4306 2145
rect 4250 2071 4306 2080
rect 4264 1494 4292 2071
rect 4252 1488 4304 1494
rect 4252 1430 4304 1436
rect 4356 480 4384 3878
rect 4448 3641 4476 4014
rect 4526 3975 4582 3984
rect 4540 3670 4568 3975
rect 4710 3768 4766 3777
rect 4710 3703 4766 3712
rect 4528 3664 4580 3670
rect 4434 3632 4490 3641
rect 4528 3606 4580 3612
rect 4434 3567 4490 3576
rect 4724 3380 4752 3703
rect 4724 3352 4844 3380
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4528 3120 4580 3126
rect 4816 3108 4844 3352
rect 4580 3080 4844 3108
rect 4528 3062 4580 3068
rect 4434 2680 4490 2689
rect 4434 2615 4490 2624
rect 4448 2582 4476 2615
rect 4436 2576 4488 2582
rect 4436 2518 4488 2524
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4908 480 4936 7806
rect 4986 7576 5042 7585
rect 4986 7511 5042 7520
rect 5092 7528 5120 7890
rect 5184 7698 5212 8044
rect 5264 8026 5316 8032
rect 5184 7670 5304 7698
rect 5000 7002 5028 7511
rect 5092 7500 5212 7528
rect 5078 7440 5134 7449
rect 5078 7375 5134 7384
rect 5092 7274 5120 7375
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 4988 6996 5040 7002
rect 4988 6938 5040 6944
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 5000 6633 5028 6734
rect 4986 6624 5042 6633
rect 4986 6559 5042 6568
rect 5184 6458 5212 7500
rect 5276 7410 5304 7670
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5262 7304 5318 7313
rect 5262 7239 5318 7248
rect 5276 7002 5304 7239
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5368 6882 5396 8758
rect 5276 6854 5396 6882
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5276 6168 5304 6854
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5368 6662 5396 6734
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5354 6488 5410 6497
rect 5354 6423 5410 6432
rect 5368 6186 5396 6423
rect 5000 6140 5304 6168
rect 5356 6180 5408 6186
rect 5000 1494 5028 6140
rect 5356 6122 5408 6128
rect 5368 6066 5396 6122
rect 5276 6038 5396 6066
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 5172 5840 5224 5846
rect 5172 5782 5224 5788
rect 5092 4457 5120 5782
rect 5184 5098 5212 5782
rect 5276 5574 5304 6038
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 5368 5409 5396 5850
rect 5354 5400 5410 5409
rect 5354 5335 5410 5344
rect 5262 5264 5318 5273
rect 5262 5199 5318 5208
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5078 4448 5134 4457
rect 5078 4383 5134 4392
rect 5184 4078 5212 4762
rect 5276 4622 5304 5199
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5368 4865 5396 5102
rect 5354 4856 5410 4865
rect 5354 4791 5356 4800
rect 5408 4791 5410 4800
rect 5356 4762 5408 4768
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5080 4004 5132 4010
rect 5080 3946 5132 3952
rect 5092 2310 5120 3946
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5264 2916 5316 2922
rect 5264 2858 5316 2864
rect 5080 2304 5132 2310
rect 5276 2281 5304 2858
rect 5080 2246 5132 2252
rect 5262 2272 5318 2281
rect 5262 2207 5318 2216
rect 4988 1488 5040 1494
rect 4988 1430 5040 1436
rect 5368 480 5396 3606
rect 5460 3398 5488 11183
rect 5552 10538 5580 15558
rect 5632 15496 5684 15502
rect 5632 15438 5684 15444
rect 5644 15094 5672 15438
rect 5632 15088 5684 15094
rect 5632 15030 5684 15036
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5644 13705 5672 14758
rect 5630 13696 5686 13705
rect 5630 13631 5686 13640
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 5632 12368 5684 12374
rect 5632 12310 5684 12316
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5538 10160 5594 10169
rect 5538 10095 5594 10104
rect 5552 9450 5580 10095
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5644 9364 5672 12310
rect 5624 9336 5672 9364
rect 5624 9194 5652 9336
rect 5624 9166 5672 9194
rect 5644 8634 5672 9166
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5736 7732 5764 13126
rect 5828 10169 5856 22520
rect 5908 19508 5960 19514
rect 5908 19450 5960 19456
rect 5920 14822 5948 19450
rect 6090 19408 6146 19417
rect 6090 19343 6146 19352
rect 6000 18148 6052 18154
rect 6000 18090 6052 18096
rect 6012 16114 6040 18090
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 5908 14544 5960 14550
rect 5908 14486 5960 14492
rect 5920 12374 5948 14486
rect 5908 12368 5960 12374
rect 5908 12310 5960 12316
rect 5920 11354 5948 12310
rect 5908 11348 5960 11354
rect 5908 11290 5960 11296
rect 5906 10976 5962 10985
rect 5906 10911 5962 10920
rect 5814 10160 5870 10169
rect 5920 10130 5948 10911
rect 5814 10095 5870 10104
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 6012 10010 6040 15846
rect 6104 12345 6132 19343
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6196 14278 6224 18022
rect 6184 14272 6236 14278
rect 6184 14214 6236 14220
rect 6184 13252 6236 13258
rect 6184 13194 6236 13200
rect 6196 12628 6224 13194
rect 6288 12696 6316 22520
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 6366 17232 6422 17241
rect 6366 17167 6422 17176
rect 6380 14482 6408 17167
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6564 15570 6592 17070
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 6472 14414 6500 15506
rect 6656 15314 6684 20198
rect 6564 15286 6684 15314
rect 6564 15042 6592 15286
rect 6748 15201 6776 22520
rect 7012 20800 7064 20806
rect 7012 20742 7064 20748
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 6932 18970 6960 19246
rect 6920 18964 6972 18970
rect 6920 18906 6972 18912
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 6734 15192 6790 15201
rect 6734 15127 6790 15136
rect 6564 15014 6776 15042
rect 6644 14952 6696 14958
rect 6644 14894 6696 14900
rect 6552 14884 6604 14890
rect 6552 14826 6604 14832
rect 6564 14618 6592 14826
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 6368 14340 6420 14346
rect 6368 14282 6420 14288
rect 6380 13462 6408 14282
rect 6368 13456 6420 13462
rect 6656 13410 6684 14894
rect 6748 14550 6776 15014
rect 6840 14618 6868 18022
rect 7024 17218 7052 20742
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7116 19922 7144 20402
rect 7104 19916 7156 19922
rect 7104 19858 7156 19864
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7116 19310 7144 19654
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 7116 18766 7144 19246
rect 7208 18902 7236 22520
rect 7300 20182 7512 20210
rect 7300 20058 7328 20182
rect 7288 20052 7340 20058
rect 7288 19994 7340 20000
rect 7380 20052 7432 20058
rect 7380 19994 7432 20000
rect 7196 18896 7248 18902
rect 7196 18838 7248 18844
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7116 18306 7144 18702
rect 7300 18358 7328 18770
rect 7288 18352 7340 18358
rect 7116 18278 7236 18306
rect 7288 18294 7340 18300
rect 7208 17746 7236 18278
rect 7196 17740 7248 17746
rect 7196 17682 7248 17688
rect 6932 17190 7052 17218
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6736 14544 6788 14550
rect 6736 14486 6788 14492
rect 6368 13398 6420 13404
rect 6380 12832 6408 13398
rect 6472 13394 6684 13410
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 6460 13388 6684 13394
rect 6512 13382 6684 13388
rect 6460 13330 6512 13336
rect 6656 12986 6684 13382
rect 6840 12986 6868 13398
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6380 12804 6500 12832
rect 6288 12668 6408 12696
rect 6196 12600 6316 12628
rect 6090 12336 6146 12345
rect 6090 12271 6146 12280
rect 6092 12164 6144 12170
rect 6092 12106 6144 12112
rect 6104 11898 6132 12106
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 6092 11552 6144 11558
rect 6090 11520 6092 11529
rect 6144 11520 6146 11529
rect 6090 11455 6146 11464
rect 6182 11112 6238 11121
rect 6182 11047 6238 11056
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 5828 9982 6040 10010
rect 5828 8786 5856 9982
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 5920 9110 5948 9658
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 6104 9042 6132 10066
rect 6196 9178 6224 11047
rect 6288 11014 6316 12600
rect 6276 11008 6328 11014
rect 6276 10950 6328 10956
rect 6276 10464 6328 10470
rect 6380 10441 6408 12668
rect 6472 12442 6500 12804
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6460 11280 6512 11286
rect 6460 11222 6512 11228
rect 6276 10406 6328 10412
rect 6366 10432 6422 10441
rect 6288 10282 6316 10406
rect 6366 10367 6422 10376
rect 6472 10305 6500 11222
rect 6458 10296 6514 10305
rect 6288 10254 6408 10282
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6276 9104 6328 9110
rect 6196 9052 6276 9058
rect 6196 9046 6328 9052
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6196 9030 6316 9046
rect 6000 8832 6052 8838
rect 5828 8758 5948 8786
rect 6000 8774 6052 8780
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 5814 8664 5870 8673
rect 5814 8599 5870 8608
rect 5828 7954 5856 8599
rect 5920 8514 5948 8758
rect 6012 8634 6040 8774
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5920 8486 6040 8514
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5814 7848 5870 7857
rect 5814 7783 5870 7792
rect 5644 7704 5764 7732
rect 5644 7546 5672 7704
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5724 7268 5776 7274
rect 5828 7256 5856 7783
rect 5776 7228 5856 7256
rect 5724 7210 5776 7216
rect 5538 7032 5594 7041
rect 5538 6967 5594 6976
rect 5632 6996 5684 7002
rect 5552 6390 5580 6967
rect 5632 6938 5684 6944
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5644 6066 5672 6938
rect 5736 6361 5764 7210
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5722 6352 5778 6361
rect 5722 6287 5778 6296
rect 5552 6038 5672 6066
rect 5552 5914 5580 6038
rect 5828 5930 5856 6598
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5644 5902 5856 5930
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5552 3942 5580 5714
rect 5644 5710 5672 5902
rect 5632 5704 5684 5710
rect 5816 5704 5868 5710
rect 5632 5646 5684 5652
rect 5814 5672 5816 5681
rect 5868 5672 5870 5681
rect 5644 5030 5672 5646
rect 5814 5607 5870 5616
rect 5920 5098 5948 8366
rect 6012 7410 6040 8486
rect 6104 8294 6132 8774
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6196 7857 6224 9030
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 6182 7848 6238 7857
rect 6182 7783 6238 7792
rect 6288 7800 6316 8502
rect 6380 8498 6408 10254
rect 6458 10231 6514 10240
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6472 8906 6500 9318
rect 6564 9110 6592 12174
rect 6932 11286 6960 17190
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 7024 16658 7052 17070
rect 7208 16658 7236 17682
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 7208 16182 7236 16594
rect 7300 16454 7328 18294
rect 7392 17134 7420 19994
rect 7484 18465 7512 20182
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7576 19242 7604 19654
rect 7564 19236 7616 19242
rect 7564 19178 7616 19184
rect 7576 18850 7604 19178
rect 7668 18970 7696 22520
rect 8128 20806 8156 22520
rect 8116 20800 8168 20806
rect 8116 20742 8168 20748
rect 8484 20392 8536 20398
rect 8484 20334 8536 20340
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 7840 19984 7892 19990
rect 7840 19926 7892 19932
rect 7852 19786 7880 19926
rect 7840 19780 7892 19786
rect 7840 19722 7892 19728
rect 8496 19417 8524 20334
rect 8482 19408 8538 19417
rect 8482 19343 8538 19352
rect 8208 19304 8260 19310
rect 8588 19258 8616 22520
rect 8668 20256 8720 20262
rect 8668 20198 8720 20204
rect 8208 19246 8260 19252
rect 8220 19122 8248 19246
rect 8404 19230 8616 19258
rect 8220 19094 8340 19122
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 7840 18896 7892 18902
rect 7576 18844 7840 18850
rect 7576 18838 7892 18844
rect 7576 18822 7880 18838
rect 8220 18766 8248 18906
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8312 18578 8340 19094
rect 8220 18550 8340 18578
rect 7470 18456 7526 18465
rect 7470 18391 7526 18400
rect 8220 18290 8248 18550
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7380 16516 7432 16522
rect 7380 16458 7432 16464
rect 7288 16448 7340 16454
rect 7392 16425 7420 16458
rect 7288 16390 7340 16396
rect 7378 16416 7434 16425
rect 7196 16176 7248 16182
rect 7196 16118 7248 16124
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7010 15600 7066 15609
rect 7010 15535 7066 15544
rect 7024 14618 7052 15535
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 7024 12306 7052 14418
rect 7208 12986 7236 15642
rect 7300 15570 7328 16390
rect 7378 16351 7434 16360
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7300 15026 7328 15302
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7300 14793 7328 14962
rect 7286 14784 7342 14793
rect 7286 14719 7342 14728
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7010 12064 7066 12073
rect 7010 11999 7066 12008
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 6918 11112 6974 11121
rect 6918 11047 6974 11056
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6644 10532 6696 10538
rect 6644 10474 6696 10480
rect 6552 9104 6604 9110
rect 6552 9046 6604 9052
rect 6460 8900 6512 8906
rect 6460 8842 6512 8848
rect 6550 8664 6606 8673
rect 6550 8599 6552 8608
rect 6604 8599 6606 8608
rect 6552 8570 6604 8576
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6288 7772 6408 7800
rect 6092 7744 6144 7750
rect 6380 7732 6408 7772
rect 6460 7744 6512 7750
rect 6144 7704 6316 7732
rect 6380 7704 6460 7732
rect 6092 7686 6144 7692
rect 6090 7440 6146 7449
rect 6000 7404 6052 7410
rect 6090 7375 6146 7384
rect 6000 7346 6052 7352
rect 6104 7274 6132 7375
rect 6092 7268 6144 7274
rect 6092 7210 6144 7216
rect 6288 7002 6316 7704
rect 6460 7686 6512 7692
rect 6460 7472 6512 7478
rect 6460 7414 6512 7420
rect 6472 7177 6500 7414
rect 6458 7168 6514 7177
rect 6458 7103 6514 7112
rect 6366 7032 6422 7041
rect 6276 6996 6328 7002
rect 6366 6967 6368 6976
rect 6276 6938 6328 6944
rect 6420 6967 6422 6976
rect 6368 6938 6420 6944
rect 6564 6882 6592 8434
rect 6656 8090 6684 10474
rect 6748 9353 6776 10746
rect 6840 10606 6868 10950
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6826 10296 6882 10305
rect 6826 10231 6882 10240
rect 6840 10062 6868 10231
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6734 9344 6790 9353
rect 6734 9279 6790 9288
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 6748 8090 6776 9046
rect 6840 8294 6868 9862
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6828 7948 6880 7954
rect 6828 7890 6880 7896
rect 6642 7848 6698 7857
rect 6642 7783 6698 7792
rect 6656 7478 6684 7783
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6748 7410 6776 7686
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6656 6934 6684 7278
rect 6012 6854 6592 6882
rect 6644 6928 6696 6934
rect 6644 6870 6696 6876
rect 5908 5092 5960 5098
rect 5908 5034 5960 5040
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5828 4758 5856 4966
rect 6012 4826 6040 6854
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6184 6724 6236 6730
rect 6184 6666 6236 6672
rect 6196 6118 6224 6666
rect 6274 6488 6330 6497
rect 6274 6423 6276 6432
rect 6328 6423 6330 6432
rect 6276 6394 6328 6400
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6288 6118 6316 6258
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 6380 5953 6408 6734
rect 6458 6488 6514 6497
rect 6458 6423 6460 6432
rect 6512 6423 6514 6432
rect 6460 6394 6512 6400
rect 6366 5944 6422 5953
rect 6366 5879 6422 5888
rect 6366 5264 6422 5273
rect 6564 5216 6592 6734
rect 6840 6610 6868 7890
rect 6748 6582 6868 6610
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6656 6089 6684 6190
rect 6642 6080 6698 6089
rect 6642 6015 6698 6024
rect 6748 5681 6776 6582
rect 6826 6488 6882 6497
rect 6826 6423 6882 6432
rect 6840 5914 6868 6423
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6734 5672 6790 5681
rect 6734 5607 6790 5616
rect 6366 5199 6368 5208
rect 6420 5199 6422 5208
rect 6368 5170 6420 5176
rect 6472 5188 6592 5216
rect 6736 5228 6788 5234
rect 6276 5160 6328 5166
rect 6328 5108 6408 5114
rect 6276 5102 6408 5108
rect 6288 5086 6408 5102
rect 6472 5098 6500 5188
rect 6736 5170 6788 5176
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 5816 4752 5868 4758
rect 5630 4720 5686 4729
rect 5816 4694 5868 4700
rect 5630 4655 5686 4664
rect 5724 4684 5776 4690
rect 5644 4554 5672 4655
rect 5724 4626 5776 4632
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 5736 4570 5764 4626
rect 5736 4554 6040 4570
rect 5632 4548 5684 4554
rect 5632 4490 5684 4496
rect 5736 4548 6052 4554
rect 5736 4542 6000 4548
rect 5630 4448 5686 4457
rect 5630 4383 5686 4392
rect 5644 4162 5672 4383
rect 5736 4282 5764 4542
rect 6000 4490 6052 4496
rect 5816 4480 5868 4486
rect 5814 4448 5816 4457
rect 6092 4480 6144 4486
rect 5868 4448 5870 4457
rect 6196 4457 6224 4626
rect 6092 4422 6144 4428
rect 6182 4448 6238 4457
rect 5814 4383 5870 4392
rect 5998 4312 6054 4321
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5816 4276 5868 4282
rect 5998 4247 6054 4256
rect 5816 4218 5868 4224
rect 5828 4162 5856 4218
rect 5644 4134 5856 4162
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5736 3670 5764 4014
rect 5724 3664 5776 3670
rect 6012 3641 6040 4247
rect 6104 4214 6132 4422
rect 6182 4383 6238 4392
rect 6092 4208 6144 4214
rect 6092 4150 6144 4156
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 5724 3606 5776 3612
rect 5998 3632 6054 3641
rect 5998 3567 6054 3576
rect 5816 3528 5868 3534
rect 5814 3496 5816 3505
rect 5868 3496 5870 3505
rect 5724 3460 5776 3466
rect 5814 3431 5870 3440
rect 5724 3402 5776 3408
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5538 3224 5594 3233
rect 5538 3159 5594 3168
rect 5552 2825 5580 3159
rect 5632 2848 5684 2854
rect 5538 2816 5594 2825
rect 5632 2790 5684 2796
rect 5538 2751 5594 2760
rect 5644 2650 5672 2790
rect 5736 2650 5764 3402
rect 6104 3369 6132 3878
rect 6090 3360 6146 3369
rect 6090 3295 6146 3304
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 6012 2417 6040 2586
rect 6104 2446 6132 3130
rect 6092 2440 6144 2446
rect 5998 2408 6054 2417
rect 6092 2382 6144 2388
rect 5998 2343 6054 2352
rect 6196 2009 6224 3878
rect 6288 3074 6316 4966
rect 6380 4321 6408 5086
rect 6460 5092 6512 5098
rect 6460 5034 6512 5040
rect 6552 5024 6604 5030
rect 6458 4992 6514 5001
rect 6552 4966 6604 4972
rect 6458 4927 6514 4936
rect 6472 4622 6500 4927
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6458 4448 6514 4457
rect 6458 4383 6514 4392
rect 6366 4312 6422 4321
rect 6366 4247 6422 4256
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6380 3670 6408 4082
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 6380 3194 6408 3606
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6288 3058 6408 3074
rect 6276 3052 6408 3058
rect 6328 3046 6408 3052
rect 6276 2994 6328 3000
rect 6288 2963 6316 2994
rect 6274 2816 6330 2825
rect 6274 2751 6330 2760
rect 6182 2000 6238 2009
rect 6182 1935 6238 1944
rect 5814 1728 5870 1737
rect 5814 1663 5870 1672
rect 5828 480 5856 1663
rect 6288 480 6316 2751
rect 6380 2417 6408 3046
rect 6366 2408 6422 2417
rect 6366 2343 6422 2352
rect 6472 1290 6500 4383
rect 6564 3602 6592 4966
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6656 4457 6684 4762
rect 6748 4554 6776 5170
rect 6840 4758 6868 5714
rect 6932 5234 6960 11047
rect 7024 9654 7052 11999
rect 7300 11898 7328 12786
rect 7392 12345 7420 15982
rect 7484 15706 7512 18226
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 8298 17912 8354 17921
rect 7656 17876 7708 17882
rect 8298 17847 8354 17856
rect 7656 17818 7708 17824
rect 7668 17270 7696 17818
rect 8312 17649 8340 17847
rect 8298 17640 8354 17649
rect 8298 17575 8354 17584
rect 7656 17264 7708 17270
rect 7656 17206 7708 17212
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 7564 16720 7616 16726
rect 7564 16662 7616 16668
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7472 15088 7524 15094
rect 7472 15030 7524 15036
rect 7484 13870 7512 15030
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7378 12336 7434 12345
rect 7378 12271 7434 12280
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7288 11756 7340 11762
rect 7288 11698 7340 11704
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 7116 9994 7144 10474
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7102 9888 7158 9897
rect 7102 9823 7158 9832
rect 7116 9738 7144 9823
rect 7116 9710 7227 9738
rect 7012 9648 7064 9654
rect 7012 9590 7064 9596
rect 7104 9648 7156 9654
rect 7104 9590 7156 9596
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 7024 6662 7052 9454
rect 7116 8430 7144 9590
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7104 8288 7156 8294
rect 7104 8230 7156 8236
rect 7116 7954 7144 8230
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7199 7188 7227 9710
rect 7116 7160 7227 7188
rect 7300 7177 7328 11698
rect 7286 7168 7342 7177
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7116 5914 7144 7160
rect 7286 7103 7342 7112
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7116 5250 7144 5850
rect 7208 5710 7236 6870
rect 7392 6440 7420 12174
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7484 11762 7512 12038
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7484 10266 7512 11290
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7576 10130 7604 16662
rect 7668 16017 7696 16730
rect 7932 16720 7984 16726
rect 7932 16662 7984 16668
rect 7944 16289 7972 16662
rect 8024 16652 8076 16658
rect 8024 16594 8076 16600
rect 7930 16280 7986 16289
rect 7930 16215 7986 16224
rect 7748 16176 7800 16182
rect 7748 16118 7800 16124
rect 7654 16008 7710 16017
rect 7654 15943 7710 15952
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 7668 12288 7696 15846
rect 7760 15026 7788 16118
rect 8036 16046 8064 16594
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 8220 15706 8248 17002
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8312 15434 8340 16050
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 7748 13796 7800 13802
rect 7748 13738 7800 13744
rect 7760 13530 7788 13738
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7760 12850 7788 13466
rect 8220 13190 8248 15302
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 8220 12442 8248 12786
rect 8298 12744 8354 12753
rect 8298 12679 8354 12688
rect 8312 12646 8340 12679
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 8298 12472 8354 12481
rect 8208 12436 8260 12442
rect 8036 12396 8208 12424
rect 7930 12336 7986 12345
rect 7668 12260 7788 12288
rect 7930 12271 7986 12280
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7668 10010 7696 11834
rect 7576 9982 7696 10010
rect 7470 9888 7526 9897
rect 7470 9823 7526 9832
rect 7484 8786 7512 9823
rect 7576 9518 7604 9982
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7668 9330 7696 9862
rect 7760 9518 7788 12260
rect 7840 12164 7892 12170
rect 7840 12106 7892 12112
rect 7852 11626 7880 12106
rect 7944 11898 7972 12271
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 8036 11762 8064 12396
rect 8298 12407 8300 12416
rect 8208 12378 8260 12384
rect 8352 12407 8354 12416
rect 8300 12378 8352 12384
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 7840 11620 7892 11626
rect 7840 11562 7892 11568
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 8220 10266 8248 11834
rect 8312 11762 8340 12378
rect 8404 12306 8432 19230
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8496 18154 8524 19110
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8484 18148 8536 18154
rect 8484 18090 8536 18096
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8300 11620 8352 11626
rect 8300 11562 8352 11568
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8312 10198 8340 11562
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8404 10810 8432 10950
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 7852 9926 7880 10066
rect 7944 10033 7972 10066
rect 8024 10056 8076 10062
rect 7930 10024 7986 10033
rect 8076 10016 8248 10044
rect 8024 9998 8076 10004
rect 7930 9959 7986 9968
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 8022 9752 8078 9761
rect 8022 9687 8078 9696
rect 8036 9518 8064 9687
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 7576 9302 7696 9330
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7576 9110 7604 9302
rect 7654 9208 7710 9217
rect 7654 9143 7656 9152
rect 7708 9143 7710 9152
rect 7656 9114 7708 9120
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7484 8758 7696 8786
rect 7562 8664 7618 8673
rect 7562 8599 7618 8608
rect 7472 8560 7524 8566
rect 7472 8502 7524 8508
rect 7484 6934 7512 8502
rect 7576 7954 7604 8599
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 7472 6928 7524 6934
rect 7472 6870 7524 6876
rect 7576 6458 7604 7210
rect 7668 6662 7696 8758
rect 7760 8498 7788 9318
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7852 8378 7880 8910
rect 7944 8430 7972 9046
rect 8220 8650 8248 10016
rect 8298 10024 8354 10033
rect 8298 9959 8354 9968
rect 8312 8838 8340 9959
rect 8404 9722 8432 10202
rect 8496 9722 8524 18090
rect 8588 17746 8616 18566
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8588 17202 8616 17682
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8588 16794 8616 16934
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8588 9568 8616 16594
rect 8680 16561 8708 20198
rect 8760 19848 8812 19854
rect 8760 19790 8812 19796
rect 8852 19848 8904 19854
rect 8852 19790 8904 19796
rect 8666 16552 8722 16561
rect 8666 16487 8722 16496
rect 8668 16448 8720 16454
rect 8668 16390 8720 16396
rect 8680 15978 8708 16390
rect 8668 15972 8720 15978
rect 8668 15914 8720 15920
rect 8680 14414 8708 15914
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8666 13968 8722 13977
rect 8666 13903 8722 13912
rect 8680 13734 8708 13903
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8680 12345 8708 13262
rect 8666 12336 8722 12345
rect 8666 12271 8722 12280
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8680 11801 8708 12174
rect 8772 11937 8800 19790
rect 8864 19553 8892 19790
rect 8850 19544 8906 19553
rect 8850 19479 8906 19488
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 8864 16833 8892 19314
rect 8942 19272 8998 19281
rect 8942 19207 8998 19216
rect 8956 18222 8984 19207
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 9048 17882 9076 22520
rect 9220 20052 9272 20058
rect 9220 19994 9272 20000
rect 9232 19514 9260 19994
rect 9600 19666 9628 22520
rect 9680 20528 9732 20534
rect 9680 20470 9732 20476
rect 9416 19638 9628 19666
rect 9220 19508 9272 19514
rect 9220 19450 9272 19456
rect 9128 19236 9180 19242
rect 9128 19178 9180 19184
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 8850 16824 8906 16833
rect 8850 16759 8906 16768
rect 8850 16688 8906 16697
rect 8850 16623 8906 16632
rect 8864 16454 8892 16623
rect 8852 16448 8904 16454
rect 8852 16390 8904 16396
rect 8852 14884 8904 14890
rect 8852 14826 8904 14832
rect 8864 14006 8892 14826
rect 8852 14000 8904 14006
rect 8852 13942 8904 13948
rect 8956 13530 8984 17682
rect 9140 17105 9168 19178
rect 9220 18692 9272 18698
rect 9220 18634 9272 18640
rect 9232 18358 9260 18634
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9220 18352 9272 18358
rect 9220 18294 9272 18300
rect 9126 17096 9182 17105
rect 9036 17060 9088 17066
rect 9126 17031 9182 17040
rect 9036 17002 9088 17008
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 9048 13410 9076 17002
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 9140 16674 9168 16934
rect 9140 16646 9260 16674
rect 9128 15972 9180 15978
rect 9128 15914 9180 15920
rect 9140 15366 9168 15914
rect 9232 15706 9260 16646
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 9128 15360 9180 15366
rect 9128 15302 9180 15308
rect 9324 15042 9352 18566
rect 9416 16969 9444 19638
rect 9692 18970 9720 20470
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9588 18080 9640 18086
rect 9586 18048 9588 18057
rect 9640 18048 9642 18057
rect 9586 17983 9642 17992
rect 9586 17912 9642 17921
rect 9496 17876 9548 17882
rect 9586 17847 9588 17856
rect 9496 17818 9548 17824
rect 9640 17847 9642 17856
rect 9588 17818 9640 17824
rect 9402 16960 9458 16969
rect 9402 16895 9458 16904
rect 9402 16688 9458 16697
rect 9402 16623 9458 16632
rect 8956 13382 9076 13410
rect 9140 15014 9352 15042
rect 8850 12744 8906 12753
rect 8850 12679 8906 12688
rect 8864 12646 8892 12679
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8850 12472 8906 12481
rect 8850 12407 8906 12416
rect 8758 11928 8814 11937
rect 8758 11863 8814 11872
rect 8760 11824 8812 11830
rect 8666 11792 8722 11801
rect 8760 11766 8812 11772
rect 8666 11727 8722 11736
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8496 9540 8616 9568
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8404 8974 8432 9386
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8220 8622 8340 8650
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 7760 8350 7880 8378
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7760 7857 7788 8350
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 7932 7880 7984 7886
rect 7746 7848 7802 7857
rect 7932 7822 7984 7828
rect 8022 7848 8078 7857
rect 7746 7783 7802 7792
rect 7840 7472 7892 7478
rect 7760 7432 7840 7460
rect 7760 7177 7788 7432
rect 7840 7414 7892 7420
rect 7944 7274 7972 7822
rect 8022 7783 8078 7792
rect 8116 7812 8168 7818
rect 8036 7410 8064 7783
rect 8116 7754 8168 7760
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 8128 7274 8156 7754
rect 8220 7342 8248 8434
rect 8312 7478 8340 8622
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 7932 7268 7984 7274
rect 7932 7210 7984 7216
rect 8116 7268 8168 7274
rect 8116 7210 8168 7216
rect 7746 7168 7802 7177
rect 7746 7103 7802 7112
rect 7760 6798 7788 7103
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 7932 6928 7984 6934
rect 7932 6870 7984 6876
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7564 6452 7616 6458
rect 7392 6412 7512 6440
rect 7378 6352 7434 6361
rect 7378 6287 7434 6296
rect 7286 5944 7342 5953
rect 7286 5879 7342 5888
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 6920 5228 6972 5234
rect 7116 5222 7236 5250
rect 6920 5170 6972 5176
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6736 4548 6788 4554
rect 6736 4490 6788 4496
rect 6642 4448 6698 4457
rect 6642 4383 6698 4392
rect 6734 4312 6790 4321
rect 6734 4247 6790 4256
rect 6642 4040 6698 4049
rect 6642 3975 6698 3984
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6564 1970 6592 2246
rect 6552 1964 6604 1970
rect 6552 1906 6604 1912
rect 6656 1358 6684 3975
rect 6748 1737 6776 4247
rect 6840 1766 6868 4558
rect 6828 1760 6880 1766
rect 6734 1728 6790 1737
rect 6828 1702 6880 1708
rect 6734 1663 6790 1672
rect 6932 1612 6960 5170
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 7024 4078 7052 4694
rect 7116 4214 7144 5102
rect 7208 4978 7236 5222
rect 7300 5098 7328 5879
rect 7392 5846 7420 6287
rect 7380 5840 7432 5846
rect 7380 5782 7432 5788
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7392 5234 7420 5646
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7288 5092 7340 5098
rect 7288 5034 7340 5040
rect 7380 5024 7432 5030
rect 7208 4950 7328 4978
rect 7380 4966 7432 4972
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7104 4208 7156 4214
rect 7104 4150 7156 4156
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7116 3738 7144 4014
rect 7104 3732 7156 3738
rect 7024 3692 7104 3720
rect 7024 3194 7052 3692
rect 7104 3674 7156 3680
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7104 2576 7156 2582
rect 7208 2564 7236 4762
rect 7300 4690 7328 4950
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7392 4570 7420 4966
rect 7484 4826 7512 6412
rect 7564 6394 7616 6400
rect 7576 5574 7604 6394
rect 7944 6304 7972 6870
rect 8220 6458 8248 7278
rect 8312 7274 8340 7414
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 8404 6458 8432 8774
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 7760 6276 7972 6304
rect 7760 6168 7788 6276
rect 7668 6140 7788 6168
rect 7668 5914 7696 6140
rect 7746 6080 7802 6089
rect 7746 6015 7802 6024
rect 7760 5914 7788 6015
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 8220 5710 8248 6394
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 8404 6089 8432 6122
rect 8390 6080 8446 6089
rect 8390 6015 8446 6024
rect 8298 5944 8354 5953
rect 8298 5879 8354 5888
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 7564 5568 7616 5574
rect 7760 5556 7788 5646
rect 7616 5528 7696 5556
rect 7564 5510 7616 5516
rect 7564 5024 7616 5030
rect 7562 4992 7564 5001
rect 7616 4992 7618 5001
rect 7562 4927 7618 4936
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7392 4542 7512 4570
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7300 4146 7328 4218
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7286 3904 7342 3913
rect 7286 3839 7342 3848
rect 7300 3738 7328 3839
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7300 3602 7328 3674
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7392 3534 7420 4422
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7378 3360 7434 3369
rect 7378 3295 7434 3304
rect 7156 2536 7236 2564
rect 7104 2518 7156 2524
rect 6748 1584 6960 1612
rect 6644 1352 6696 1358
rect 6644 1294 6696 1300
rect 6460 1284 6512 1290
rect 6460 1226 6512 1232
rect 6748 480 6776 1584
rect 7194 1456 7250 1465
rect 7392 1426 7420 3295
rect 7484 3074 7512 4542
rect 7576 3466 7604 4626
rect 7668 4146 7696 5528
rect 7751 5528 7788 5556
rect 7751 4486 7779 5528
rect 7840 5364 7892 5370
rect 8036 5352 8064 5646
rect 7892 5324 8064 5352
rect 7840 5306 7892 5312
rect 8312 5302 8340 5879
rect 8300 5296 8352 5302
rect 7930 5264 7986 5273
rect 7930 5199 7986 5208
rect 8206 5264 8262 5273
rect 8300 5238 8352 5244
rect 8206 5199 8262 5208
rect 7944 5166 7972 5199
rect 8220 5166 8248 5199
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 8116 4752 8168 4758
rect 8036 4712 8116 4740
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7746 4312 7802 4321
rect 7746 4247 7802 4256
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7668 3505 7696 4082
rect 7760 3738 7788 4247
rect 7944 3924 7972 4422
rect 8036 4049 8064 4712
rect 8116 4694 8168 4700
rect 8312 4672 8340 5238
rect 8404 5234 8432 6015
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8404 5001 8432 5170
rect 8496 5098 8524 9540
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 8588 9110 8616 9386
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8588 8294 8616 8910
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8680 7936 8708 11630
rect 8772 11082 8800 11766
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8772 10985 8800 11018
rect 8758 10976 8814 10985
rect 8758 10911 8814 10920
rect 8760 9988 8812 9994
rect 8760 9930 8812 9936
rect 8588 7908 8708 7936
rect 8484 5092 8536 5098
rect 8588 5080 8616 7908
rect 8666 7848 8722 7857
rect 8666 7783 8722 7792
rect 8680 5642 8708 7783
rect 8772 6168 8800 9930
rect 8864 7750 8892 12407
rect 8956 10713 8984 13382
rect 9034 11520 9090 11529
rect 9034 11455 9090 11464
rect 8942 10704 8998 10713
rect 8942 10639 8998 10648
rect 8956 9761 8984 10639
rect 8942 9752 8998 9761
rect 8942 9687 8998 9696
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8956 9217 8984 9522
rect 8942 9208 8998 9217
rect 8942 9143 8998 9152
rect 8944 9036 8996 9042
rect 8944 8978 8996 8984
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8852 7268 8904 7274
rect 8852 7210 8904 7216
rect 8864 6322 8892 7210
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8772 6140 8892 6168
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8772 5710 8800 5850
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 8758 5536 8814 5545
rect 8758 5471 8814 5480
rect 8668 5296 8720 5302
rect 8666 5264 8668 5273
rect 8720 5264 8722 5273
rect 8666 5199 8722 5208
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8484 5034 8536 5040
rect 8579 5052 8616 5080
rect 8390 4992 8446 5001
rect 8446 4950 8524 4978
rect 8390 4927 8446 4936
rect 8312 4644 8432 4672
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8022 4040 8078 4049
rect 8022 3975 8078 3984
rect 8206 4040 8262 4049
rect 8206 3975 8262 3984
rect 8220 3924 8248 3975
rect 7944 3896 8248 3924
rect 8312 3913 8340 4490
rect 8298 3904 8354 3913
rect 7886 3836 8182 3856
rect 8298 3839 8354 3848
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 8404 3738 8432 4644
rect 8496 4622 8524 4950
rect 8579 4672 8607 5052
rect 8680 4842 8708 5102
rect 8772 5030 8800 5471
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8680 4814 8800 4842
rect 8579 4644 8616 4672
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8208 3664 8260 3670
rect 8022 3632 8078 3641
rect 8208 3606 8260 3612
rect 8390 3632 8446 3641
rect 8022 3567 8078 3576
rect 7654 3496 7710 3505
rect 7564 3460 7616 3466
rect 7654 3431 7710 3440
rect 7564 3402 7616 3408
rect 7484 3046 7604 3074
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7484 2825 7512 2926
rect 7470 2816 7526 2825
rect 7470 2751 7526 2760
rect 7472 2576 7524 2582
rect 7472 2518 7524 2524
rect 7484 1601 7512 2518
rect 7576 2310 7604 3046
rect 7668 2972 7696 3431
rect 8036 3126 8064 3567
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 8128 3074 8156 3470
rect 8220 3398 8248 3606
rect 8390 3567 8446 3576
rect 8298 3496 8354 3505
rect 8298 3431 8354 3440
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 8312 3210 8340 3431
rect 8220 3194 8340 3210
rect 8208 3188 8340 3194
rect 8260 3182 8340 3188
rect 8208 3130 8260 3136
rect 8128 3046 8340 3074
rect 8024 2984 8076 2990
rect 7668 2944 8024 2972
rect 8024 2926 8076 2932
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 7932 2576 7984 2582
rect 7654 2544 7710 2553
rect 7932 2518 7984 2524
rect 8114 2544 8170 2553
rect 7654 2479 7710 2488
rect 7564 2304 7616 2310
rect 7564 2246 7616 2252
rect 7470 1592 7526 1601
rect 7470 1527 7526 1536
rect 7194 1391 7250 1400
rect 7380 1420 7432 1426
rect 7208 480 7236 1391
rect 7380 1362 7432 1368
rect 7668 480 7696 2479
rect 7944 2446 7972 2518
rect 8024 2508 8076 2514
rect 8114 2479 8170 2488
rect 8024 2450 8076 2456
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 8036 1601 8064 2450
rect 8022 1592 8078 1601
rect 8022 1527 8078 1536
rect 8128 480 8156 2479
rect 8220 1698 8248 2586
rect 8312 1737 8340 3046
rect 8298 1728 8354 1737
rect 8208 1692 8260 1698
rect 8298 1663 8354 1672
rect 8208 1634 8260 1640
rect 8404 1562 8432 3567
rect 8496 2582 8524 3946
rect 8484 2576 8536 2582
rect 8484 2518 8536 2524
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 8496 1766 8524 2246
rect 8484 1760 8536 1766
rect 8484 1702 8536 1708
rect 8482 1592 8538 1601
rect 8392 1556 8444 1562
rect 8482 1527 8484 1536
rect 8392 1498 8444 1504
rect 8536 1527 8538 1536
rect 8484 1498 8536 1504
rect 8588 480 8616 4644
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8680 2582 8708 3470
rect 8772 3398 8800 4814
rect 8864 3602 8892 6140
rect 8956 4604 8984 8978
rect 9048 7585 9076 11455
rect 9140 9382 9168 15014
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 9324 14521 9352 14894
rect 9310 14512 9366 14521
rect 9220 14476 9272 14482
rect 9310 14447 9366 14456
rect 9220 14418 9272 14424
rect 9232 13326 9260 14418
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9324 13530 9352 14214
rect 9416 13802 9444 16623
rect 9404 13796 9456 13802
rect 9404 13738 9456 13744
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 9140 8838 9168 9046
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9034 7576 9090 7585
rect 9034 7511 9090 7520
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9048 5302 9076 7142
rect 9140 6905 9168 8570
rect 9126 6896 9182 6905
rect 9126 6831 9182 6840
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9140 6474 9168 6734
rect 9232 6610 9260 12922
rect 9324 12850 9352 13262
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9324 11694 9352 12786
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9416 9994 9444 13738
rect 9404 9988 9456 9994
rect 9404 9930 9456 9936
rect 9508 9874 9536 17818
rect 9586 16552 9642 16561
rect 9692 16538 9720 18226
rect 9784 16590 9812 19654
rect 9876 18290 9904 19858
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9968 18737 9996 18770
rect 9954 18728 10010 18737
rect 9954 18663 10010 18672
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9862 17776 9918 17785
rect 9862 17711 9918 17720
rect 9876 16833 9904 17711
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9862 16824 9918 16833
rect 9862 16759 9918 16768
rect 9862 16688 9918 16697
rect 9862 16623 9864 16632
rect 9916 16623 9918 16632
rect 9864 16594 9916 16600
rect 9642 16510 9720 16538
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9586 16487 9642 16496
rect 9862 16416 9918 16425
rect 9862 16351 9918 16360
rect 9876 16250 9904 16351
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9678 16008 9734 16017
rect 9678 15943 9734 15952
rect 9692 15502 9720 15943
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9600 14278 9628 14758
rect 9692 14550 9720 15302
rect 9784 15094 9812 16186
rect 9968 16153 9996 16934
rect 9954 16144 10010 16153
rect 9954 16079 10010 16088
rect 10060 16096 10088 22520
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10140 20256 10192 20262
rect 10140 20198 10192 20204
rect 10152 19961 10180 20198
rect 10336 20058 10364 20402
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10324 20052 10376 20058
rect 10324 19994 10376 20000
rect 10138 19952 10194 19961
rect 10138 19887 10194 19896
rect 10232 19848 10284 19854
rect 10230 19816 10232 19825
rect 10284 19816 10286 19825
rect 10230 19751 10286 19760
rect 10230 19272 10286 19281
rect 10230 19207 10232 19216
rect 10284 19207 10286 19216
rect 10232 19178 10284 19184
rect 10322 19000 10378 19009
rect 10322 18935 10378 18944
rect 10140 17264 10192 17270
rect 10192 17224 10272 17252
rect 10140 17206 10192 17212
rect 10060 16068 10180 16096
rect 9864 15904 9916 15910
rect 9862 15872 9864 15881
rect 9956 15904 10008 15910
rect 9916 15872 9918 15881
rect 9956 15846 10008 15852
rect 9862 15807 9918 15816
rect 9968 15638 9996 15846
rect 10152 15706 10180 16068
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 9956 15632 10008 15638
rect 9956 15574 10008 15580
rect 10046 15600 10102 15609
rect 10244 15586 10272 17224
rect 10046 15535 10048 15544
rect 10100 15535 10102 15544
rect 10152 15558 10272 15586
rect 10048 15506 10100 15512
rect 9864 15428 9916 15434
rect 9864 15370 9916 15376
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 9876 14793 9904 15370
rect 10152 14906 10180 15558
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10244 15026 10272 15302
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 10152 14878 10272 14906
rect 9956 14816 10008 14822
rect 9862 14784 9918 14793
rect 9956 14758 10008 14764
rect 9862 14719 9918 14728
rect 9770 14648 9826 14657
rect 9770 14583 9826 14592
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9588 14272 9640 14278
rect 9588 14214 9640 14220
rect 9692 14074 9720 14350
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9784 13734 9812 14583
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9876 13462 9904 14719
rect 9968 14346 9996 14758
rect 9956 14340 10008 14346
rect 9956 14282 10008 14288
rect 10048 13728 10100 13734
rect 10046 13696 10048 13705
rect 10100 13696 10102 13705
rect 10046 13631 10102 13640
rect 9772 13456 9824 13462
rect 9772 13398 9824 13404
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9784 13002 9812 13398
rect 9876 13161 9904 13398
rect 10138 13288 10194 13297
rect 10138 13223 10194 13232
rect 10048 13184 10100 13190
rect 9862 13152 9918 13161
rect 10048 13126 10100 13132
rect 9862 13087 9918 13096
rect 9784 12974 9996 13002
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9876 12753 9904 12854
rect 9862 12744 9918 12753
rect 9588 12708 9640 12714
rect 9862 12679 9918 12688
rect 9588 12650 9640 12656
rect 9416 9846 9536 9874
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 9324 6905 9352 9658
rect 9310 6896 9366 6905
rect 9310 6831 9366 6840
rect 9232 6582 9352 6610
rect 9140 6446 9260 6474
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9140 5710 9168 6258
rect 9232 5914 9260 6446
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9324 5794 9352 6582
rect 9232 5766 9352 5794
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9126 5400 9182 5409
rect 9126 5335 9182 5344
rect 9036 5296 9088 5302
rect 9036 5238 9088 5244
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 9048 4758 9076 4966
rect 9036 4752 9088 4758
rect 9036 4694 9088 4700
rect 8956 4576 9076 4604
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8864 2990 8892 3538
rect 8944 3460 8996 3466
rect 8944 3402 8996 3408
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 8772 2496 8800 2858
rect 8852 2508 8904 2514
rect 8772 2468 8852 2496
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 8680 2310 8708 2382
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 8666 2000 8722 2009
rect 8666 1935 8722 1944
rect 8680 1601 8708 1935
rect 8772 1834 8800 2468
rect 8956 2496 8984 3402
rect 9048 2689 9076 4576
rect 9140 4321 9168 5335
rect 9126 4312 9182 4321
rect 9126 4247 9182 4256
rect 9034 2680 9090 2689
rect 9034 2615 9090 2624
rect 9036 2508 9088 2514
rect 8956 2468 9036 2496
rect 8852 2450 8904 2456
rect 9036 2450 9088 2456
rect 9140 2378 9168 4247
rect 9232 4078 9260 5766
rect 9416 5522 9444 9846
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9508 9489 9536 9522
rect 9494 9480 9550 9489
rect 9494 9415 9550 9424
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9508 8362 9536 9318
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9508 7954 9536 8298
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9508 7177 9536 7414
rect 9494 7168 9550 7177
rect 9494 7103 9550 7112
rect 9496 5840 9548 5846
rect 9496 5782 9548 5788
rect 9324 5494 9444 5522
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9324 3210 9352 5494
rect 9402 5400 9458 5409
rect 9402 5335 9458 5344
rect 9416 4049 9444 5335
rect 9508 4865 9536 5782
rect 9494 4856 9550 4865
rect 9494 4791 9550 4800
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9508 4214 9536 4626
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9402 4040 9458 4049
rect 9402 3975 9458 3984
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 9402 3768 9458 3777
rect 9402 3703 9458 3712
rect 9232 3182 9352 3210
rect 9232 2689 9260 3182
rect 9312 3120 9364 3126
rect 9312 3062 9364 3068
rect 9218 2680 9274 2689
rect 9324 2650 9352 3062
rect 9416 2938 9444 3703
rect 9508 3233 9536 3946
rect 9600 3738 9628 12650
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9692 12238 9720 12378
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9692 11218 9720 11630
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9784 10810 9812 12582
rect 9968 11529 9996 12974
rect 10060 12782 10088 13126
rect 10152 12850 10180 13223
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10048 12776 10100 12782
rect 10244 12730 10272 14878
rect 10336 13734 10364 18935
rect 10428 16046 10456 20334
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10428 15706 10456 15846
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10416 15564 10468 15570
rect 10416 15506 10468 15512
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 10048 12718 10100 12724
rect 10060 12481 10088 12718
rect 10152 12702 10272 12730
rect 10046 12472 10102 12481
rect 10046 12407 10102 12416
rect 10048 12164 10100 12170
rect 10048 12106 10100 12112
rect 9954 11520 10010 11529
rect 9954 11455 10010 11464
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9692 10062 9720 10474
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9692 8838 9720 9998
rect 9784 9518 9812 10746
rect 9954 10568 10010 10577
rect 9954 10503 10010 10512
rect 9862 10296 9918 10305
rect 9862 10231 9918 10240
rect 9876 9897 9904 10231
rect 9862 9888 9918 9897
rect 9862 9823 9918 9832
rect 9968 9722 9996 10503
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9770 9208 9826 9217
rect 9770 9143 9772 9152
rect 9824 9143 9826 9152
rect 9772 9114 9824 9120
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9692 7954 9720 8774
rect 9876 8673 9904 9318
rect 9968 8974 9996 9522
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9862 8664 9918 8673
rect 9772 8628 9824 8634
rect 9862 8599 9918 8608
rect 9956 8628 10008 8634
rect 9772 8570 9824 8576
rect 9956 8570 10008 8576
rect 9784 8430 9812 8570
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9968 7954 9996 8570
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9692 7342 9720 7890
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9770 7576 9826 7585
rect 9770 7511 9826 7520
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 6322 9720 7142
rect 9784 6390 9812 7511
rect 9876 7206 9904 7686
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9862 7032 9918 7041
rect 9862 6967 9918 6976
rect 9876 6798 9904 6967
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9855 6656 9907 6662
rect 9855 6598 9907 6604
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9680 6180 9732 6186
rect 9680 6122 9732 6128
rect 9692 5914 9720 6122
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9692 4826 9720 5238
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9692 4214 9720 4558
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9678 4040 9734 4049
rect 9678 3975 9734 3984
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9494 3224 9550 3233
rect 9600 3194 9628 3402
rect 9494 3159 9550 3168
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9416 2910 9536 2938
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9218 2615 9274 2624
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 8852 2372 8904 2378
rect 8852 2314 8904 2320
rect 9128 2372 9180 2378
rect 9128 2314 9180 2320
rect 8760 1828 8812 1834
rect 8760 1770 8812 1776
rect 8864 1698 8892 2314
rect 9232 2009 9260 2450
rect 9416 2281 9444 2790
rect 9402 2272 9458 2281
rect 9402 2207 9458 2216
rect 9034 2000 9090 2009
rect 9034 1935 9090 1944
rect 9218 2000 9274 2009
rect 9218 1935 9274 1944
rect 8852 1692 8904 1698
rect 8852 1634 8904 1640
rect 8666 1592 8722 1601
rect 8666 1527 8722 1536
rect 9048 480 9076 1935
rect 9508 1766 9536 2910
rect 9692 2854 9720 3975
rect 9784 3618 9812 6190
rect 9876 4486 9904 6598
rect 9968 5545 9996 7890
rect 10060 6089 10088 12106
rect 10046 6080 10102 6089
rect 10046 6015 10102 6024
rect 9954 5536 10010 5545
rect 9954 5471 10010 5480
rect 10152 5386 10180 12702
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10336 11694 10364 12174
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10244 9722 10272 11154
rect 10336 10810 10364 11630
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10322 9480 10378 9489
rect 10322 9415 10378 9424
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10244 9178 10272 9318
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 10244 8498 10272 8978
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10336 7528 10364 9415
rect 10060 5358 10180 5386
rect 10244 7500 10364 7528
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 9968 3890 9996 5102
rect 10060 4010 10088 5358
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10152 4554 10180 4762
rect 10244 4758 10272 7500
rect 10428 7426 10456 15506
rect 10520 15502 10548 22520
rect 10980 20330 11008 22520
rect 11440 20890 11468 22520
rect 11072 20862 11468 20890
rect 10968 20324 11020 20330
rect 10968 20266 11020 20272
rect 10600 20256 10652 20262
rect 10600 20198 10652 20204
rect 10612 20058 10640 20198
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 10968 19236 11020 19242
rect 10968 19178 11020 19184
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10612 17134 10640 17614
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10600 16584 10652 16590
rect 10598 16552 10600 16561
rect 10652 16552 10654 16561
rect 10598 16487 10654 16496
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10612 15348 10640 15982
rect 10520 15320 10640 15348
rect 10520 9897 10548 15320
rect 10704 15178 10732 18226
rect 10796 17202 10824 18770
rect 10876 18216 10928 18222
rect 10876 18158 10928 18164
rect 10784 17196 10836 17202
rect 10784 17138 10836 17144
rect 10782 17096 10838 17105
rect 10782 17031 10838 17040
rect 10796 16658 10824 17031
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10888 16590 10916 18158
rect 10980 17678 11008 19178
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 10980 17542 11008 17614
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10980 17202 11008 17478
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 11072 16776 11100 20862
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 11336 20392 11388 20398
rect 11336 20334 11388 20340
rect 11244 20324 11296 20330
rect 11244 20266 11296 20272
rect 11256 19990 11284 20266
rect 11348 19990 11376 20334
rect 11704 20256 11756 20262
rect 11704 20198 11756 20204
rect 11796 20256 11848 20262
rect 11796 20198 11848 20204
rect 11244 19984 11296 19990
rect 11244 19926 11296 19932
rect 11336 19984 11388 19990
rect 11336 19926 11388 19932
rect 11244 19848 11296 19854
rect 11242 19816 11244 19825
rect 11336 19848 11388 19854
rect 11296 19816 11298 19825
rect 11336 19790 11388 19796
rect 11242 19751 11298 19760
rect 11348 19700 11376 19790
rect 11256 19672 11376 19700
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 10980 16748 11100 16776
rect 10876 16584 10928 16590
rect 10980 16561 11008 16748
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 10876 16526 10928 16532
rect 10966 16552 11022 16561
rect 10966 16487 11022 16496
rect 10966 15872 11022 15881
rect 10966 15807 11022 15816
rect 10980 15706 11008 15807
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10612 15150 10732 15178
rect 10876 15156 10928 15162
rect 10612 14396 10640 15150
rect 10876 15098 10928 15104
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10796 14618 10824 14758
rect 10888 14618 10916 15098
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10612 14368 10732 14396
rect 10704 13852 10732 14368
rect 10612 13824 10732 13852
rect 10612 12442 10640 13824
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 10796 12986 10824 13670
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10980 12617 11008 15438
rect 11072 12764 11100 16594
rect 11164 14890 11192 18022
rect 11256 17542 11284 19672
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 11716 18834 11744 20198
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11704 17876 11756 17882
rect 11704 17818 11756 17824
rect 11610 17776 11666 17785
rect 11610 17711 11612 17720
rect 11664 17711 11666 17720
rect 11612 17682 11664 17688
rect 11716 17542 11744 17818
rect 11244 17536 11296 17542
rect 11244 17478 11296 17484
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11702 17232 11758 17241
rect 11702 17167 11758 17176
rect 11716 17134 11744 17167
rect 11704 17128 11756 17134
rect 11704 17070 11756 17076
rect 11808 16794 11836 20198
rect 11900 17882 11928 22520
rect 11978 19816 12034 19825
rect 11978 19751 12034 19760
rect 11992 19514 12020 19751
rect 11980 19508 12032 19514
rect 11980 19450 12032 19456
rect 12254 19408 12310 19417
rect 12254 19343 12256 19352
rect 12308 19343 12310 19352
rect 12256 19314 12308 19320
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 12268 18873 12296 18906
rect 12254 18864 12310 18873
rect 12254 18799 12310 18808
rect 11980 18760 12032 18766
rect 11980 18702 12032 18708
rect 11888 17876 11940 17882
rect 11888 17818 11940 17824
rect 11886 17368 11942 17377
rect 11886 17303 11942 17312
rect 11796 16788 11848 16794
rect 11796 16730 11848 16736
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11336 16108 11388 16114
rect 11256 16068 11336 16096
rect 11152 14884 11204 14890
rect 11152 14826 11204 14832
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11164 12889 11192 14214
rect 11256 12986 11284 16068
rect 11336 16050 11388 16056
rect 11612 15564 11664 15570
rect 11612 15506 11664 15512
rect 11624 15473 11652 15506
rect 11610 15464 11666 15473
rect 11610 15399 11666 15408
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11426 14920 11482 14929
rect 11426 14855 11482 14864
rect 11336 14544 11388 14550
rect 11334 14512 11336 14521
rect 11388 14512 11390 14521
rect 11440 14482 11468 14855
rect 11334 14447 11390 14456
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11150 12880 11206 12889
rect 11150 12815 11206 12824
rect 11072 12736 11284 12764
rect 10966 12608 11022 12617
rect 10966 12543 11022 12552
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10796 11200 10824 12242
rect 10796 11172 10916 11200
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10506 9888 10562 9897
rect 10704 9874 10732 11086
rect 10784 11076 10836 11082
rect 10784 11018 10836 11024
rect 10506 9823 10562 9832
rect 10612 9846 10732 9874
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10520 8090 10548 9522
rect 10612 9110 10640 9846
rect 10690 9752 10746 9761
rect 10690 9687 10746 9696
rect 10600 9104 10652 9110
rect 10600 9046 10652 9052
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10612 8634 10640 8910
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10336 7398 10456 7426
rect 10232 4752 10284 4758
rect 10232 4694 10284 4700
rect 10140 4548 10192 4554
rect 10336 4536 10364 7398
rect 10416 7336 10468 7342
rect 10520 7324 10548 8026
rect 10612 7585 10640 8366
rect 10598 7576 10654 7585
rect 10598 7511 10654 7520
rect 10468 7296 10548 7324
rect 10416 7278 10468 7284
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10428 6390 10456 6802
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 10520 6168 10548 6734
rect 10598 6488 10654 6497
rect 10598 6423 10654 6432
rect 10612 6254 10640 6423
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10428 6140 10548 6168
rect 10428 5030 10456 6140
rect 10704 6089 10732 9687
rect 10506 6080 10562 6089
rect 10690 6080 10746 6089
rect 10562 6038 10640 6066
rect 10506 6015 10562 6024
rect 10506 5536 10562 5545
rect 10506 5471 10562 5480
rect 10520 5166 10548 5471
rect 10612 5166 10640 6038
rect 10690 6015 10746 6024
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10508 4752 10560 4758
rect 10508 4694 10560 4700
rect 10336 4508 10456 4536
rect 10140 4490 10192 4496
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 10140 3936 10192 3942
rect 9968 3862 10088 3890
rect 10140 3878 10192 3884
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 9968 3618 9996 3674
rect 9784 3590 9996 3618
rect 9784 3369 9812 3590
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9770 3360 9826 3369
rect 9770 3295 9826 3304
rect 9876 3194 9904 3470
rect 9956 3392 10008 3398
rect 10060 3369 10088 3862
rect 9956 3334 10008 3340
rect 10046 3360 10102 3369
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9772 2984 9824 2990
rect 9824 2944 9904 2972
rect 9772 2926 9824 2932
rect 9680 2848 9732 2854
rect 9586 2816 9642 2825
rect 9680 2790 9732 2796
rect 9772 2848 9824 2854
rect 9876 2825 9904 2944
rect 9772 2790 9824 2796
rect 9862 2816 9918 2825
rect 9586 2751 9642 2760
rect 9496 1760 9548 1766
rect 9496 1702 9548 1708
rect 9600 480 9628 2751
rect 9784 2394 9812 2790
rect 9862 2751 9918 2760
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 9692 2366 9812 2394
rect 9692 2038 9720 2366
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9784 2038 9812 2246
rect 9680 2032 9732 2038
rect 9680 1974 9732 1980
rect 9772 2032 9824 2038
rect 9772 1974 9824 1980
rect 9876 1902 9904 2586
rect 9968 1902 9996 3334
rect 10046 3295 10102 3304
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 10060 2514 10088 3130
rect 10152 2650 10180 3878
rect 10244 3602 10272 3878
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10244 3058 10272 3130
rect 10336 3058 10364 4082
rect 10428 3108 10456 4508
rect 10520 3641 10548 4694
rect 10612 4321 10640 4966
rect 10598 4312 10654 4321
rect 10598 4247 10654 4256
rect 10704 4214 10732 5170
rect 10796 4690 10824 11018
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10782 4312 10838 4321
rect 10782 4247 10838 4256
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 10506 3632 10562 3641
rect 10506 3567 10562 3576
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10520 3233 10548 3470
rect 10506 3224 10562 3233
rect 10506 3159 10562 3168
rect 10428 3080 10548 3108
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 10140 2304 10192 2310
rect 10046 2272 10102 2281
rect 10140 2246 10192 2252
rect 10046 2207 10102 2216
rect 9864 1896 9916 1902
rect 9864 1838 9916 1844
rect 9956 1896 10008 1902
rect 9956 1838 10008 1844
rect 10060 480 10088 2207
rect 10152 1698 10180 2246
rect 10140 1692 10192 1698
rect 10140 1634 10192 1640
rect 10244 1426 10272 2450
rect 10336 2446 10364 2994
rect 10416 2916 10468 2922
rect 10416 2858 10468 2864
rect 10428 2825 10456 2858
rect 10414 2816 10470 2825
rect 10414 2751 10470 2760
rect 10416 2576 10468 2582
rect 10416 2518 10468 2524
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10232 1420 10284 1426
rect 10232 1362 10284 1368
rect 10428 1290 10456 2518
rect 10416 1284 10468 1290
rect 10416 1226 10468 1232
rect 10520 480 10548 3080
rect 10598 2816 10654 2825
rect 10598 2751 10654 2760
rect 10612 2650 10640 2751
rect 10600 2644 10652 2650
rect 10796 2632 10824 4247
rect 10888 3942 10916 11172
rect 10980 10033 11008 12378
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 11072 11694 11100 12038
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 11072 11286 11100 11494
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11072 10470 11100 10746
rect 11164 10742 11192 10950
rect 11152 10736 11204 10742
rect 11152 10678 11204 10684
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 11164 10033 11192 10474
rect 10966 10024 11022 10033
rect 11150 10024 11206 10033
rect 10966 9959 11022 9968
rect 11072 9982 11150 10010
rect 11072 8673 11100 9982
rect 11150 9959 11206 9968
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11058 8664 11114 8673
rect 11058 8599 11114 8608
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 10980 7585 11008 7754
rect 10966 7576 11022 7585
rect 10966 7511 11022 7520
rect 10966 7440 11022 7449
rect 10966 7375 11022 7384
rect 10980 6866 11008 7375
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10980 5545 11008 5578
rect 10966 5536 11022 5545
rect 10966 5471 11022 5480
rect 11072 5409 11100 6598
rect 11164 6322 11192 8978
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11058 5400 11114 5409
rect 11058 5335 11114 5344
rect 11164 5284 11192 5850
rect 11072 5256 11192 5284
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10874 3768 10930 3777
rect 10874 3703 10930 3712
rect 10888 3466 10916 3703
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 10876 3120 10928 3126
rect 10876 3062 10928 3068
rect 10888 2854 10916 3062
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 10600 2586 10652 2592
rect 10704 2604 10824 2632
rect 10704 2145 10732 2604
rect 10888 2582 10916 2790
rect 10876 2576 10928 2582
rect 10782 2544 10838 2553
rect 10876 2518 10928 2524
rect 10782 2479 10838 2488
rect 10796 2394 10824 2479
rect 10876 2440 10928 2446
rect 10796 2388 10876 2394
rect 10796 2382 10928 2388
rect 10796 2366 10916 2382
rect 10690 2136 10746 2145
rect 10690 2071 10746 2080
rect 10980 480 11008 5102
rect 11072 4758 11100 5256
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 11152 4752 11204 4758
rect 11152 4694 11204 4700
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11072 4457 11100 4558
rect 11058 4448 11114 4457
rect 11058 4383 11114 4392
rect 11164 4321 11192 4694
rect 11150 4312 11206 4321
rect 11150 4247 11206 4256
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 11072 2825 11100 3946
rect 11150 3360 11206 3369
rect 11150 3295 11206 3304
rect 11058 2816 11114 2825
rect 11058 2751 11114 2760
rect 11058 2680 11114 2689
rect 11164 2650 11192 3295
rect 11058 2615 11060 2624
rect 11112 2615 11114 2624
rect 11152 2644 11204 2650
rect 11060 2586 11112 2592
rect 11152 2586 11204 2592
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 11072 1494 11100 2450
rect 11256 2088 11284 12736
rect 11612 12436 11664 12442
rect 11716 12424 11744 16594
rect 11900 15026 11928 17303
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11900 14278 11928 14350
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11808 13841 11836 14010
rect 11794 13832 11850 13841
rect 11794 13767 11850 13776
rect 11794 13560 11850 13569
rect 11794 13495 11796 13504
rect 11848 13495 11850 13504
rect 11796 13466 11848 13472
rect 11796 13320 11848 13326
rect 11900 13297 11928 14214
rect 11796 13262 11848 13268
rect 11886 13288 11942 13297
rect 11808 12442 11836 13262
rect 11886 13223 11942 13232
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11900 12986 11928 13126
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11992 12481 12020 18702
rect 12360 18578 12388 22520
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 12544 20346 12572 20538
rect 12544 20318 12756 20346
rect 12728 19922 12756 20318
rect 12820 20058 12848 22520
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12808 20052 12860 20058
rect 12808 19994 12860 20000
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12452 19417 12480 19654
rect 12438 19408 12494 19417
rect 12438 19343 12494 19352
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 12452 18766 12480 19246
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12084 18550 12388 18578
rect 11978 12472 12034 12481
rect 11664 12396 11744 12424
rect 11796 12436 11848 12442
rect 11612 12378 11664 12384
rect 11978 12407 12034 12416
rect 11796 12378 11848 12384
rect 11980 12368 12032 12374
rect 11980 12310 12032 12316
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11440 11286 11468 11630
rect 11716 11354 11744 12038
rect 11794 11928 11850 11937
rect 11794 11863 11850 11872
rect 11808 11626 11836 11863
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11428 11280 11480 11286
rect 11428 11222 11480 11228
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11610 10704 11666 10713
rect 11428 10668 11480 10674
rect 11610 10639 11666 10648
rect 11428 10610 11480 10616
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11348 10266 11376 10474
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11440 9994 11468 10610
rect 11518 10568 11574 10577
rect 11518 10503 11574 10512
rect 11532 10470 11560 10503
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11518 10024 11574 10033
rect 11428 9988 11480 9994
rect 11624 10010 11652 10639
rect 11716 10606 11744 10950
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11574 9982 11652 10010
rect 11702 10024 11758 10033
rect 11518 9959 11520 9968
rect 11428 9930 11480 9936
rect 11572 9959 11574 9968
rect 11702 9959 11758 9968
rect 11520 9930 11572 9936
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11428 8356 11480 8362
rect 11428 8298 11480 8304
rect 11440 7993 11468 8298
rect 11426 7984 11482 7993
rect 11426 7919 11482 7928
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11348 6798 11376 7278
rect 11440 7002 11468 7346
rect 11716 7041 11744 9959
rect 11702 7032 11758 7041
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11520 6996 11572 7002
rect 11702 6967 11758 6976
rect 11520 6938 11572 6944
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11532 6730 11560 6938
rect 11704 6928 11756 6934
rect 11704 6870 11756 6876
rect 11716 6798 11744 6870
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11612 6384 11664 6390
rect 11612 6326 11664 6332
rect 11428 6316 11480 6322
rect 11428 6258 11480 6264
rect 11336 6248 11388 6254
rect 11336 6190 11388 6196
rect 11348 5710 11376 6190
rect 11440 6089 11468 6258
rect 11426 6080 11482 6089
rect 11426 6015 11482 6024
rect 11624 5710 11652 6326
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11336 5296 11388 5302
rect 11336 5238 11388 5244
rect 11348 4826 11376 5238
rect 11336 4820 11388 4826
rect 11716 4808 11744 5714
rect 11336 4762 11388 4768
rect 11624 4780 11744 4808
rect 11624 4690 11652 4780
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11428 4208 11480 4214
rect 11428 4150 11480 4156
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11348 3641 11376 4082
rect 11440 4010 11468 4150
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11428 4004 11480 4010
rect 11428 3946 11480 3952
rect 11532 3777 11560 4082
rect 11518 3768 11574 3777
rect 11624 3738 11652 4150
rect 11518 3703 11574 3712
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11334 3632 11390 3641
rect 11334 3567 11390 3576
rect 11612 3596 11664 3602
rect 11716 3584 11744 4626
rect 11664 3556 11744 3584
rect 11612 3538 11664 3544
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11716 3126 11744 3556
rect 11808 3534 11836 10950
rect 11888 10736 11940 10742
rect 11888 10678 11940 10684
rect 11900 10266 11928 10678
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11992 10146 12020 12310
rect 11900 10118 12020 10146
rect 11900 6338 11928 10118
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11992 8838 12020 9998
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11992 7274 12020 7890
rect 11980 7268 12032 7274
rect 11980 7210 12032 7216
rect 11900 6310 12020 6338
rect 11992 5846 12020 6310
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11900 5370 11928 5510
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11992 5166 12020 5646
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 11888 5092 11940 5098
rect 11888 5034 11940 5040
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11520 3120 11572 3126
rect 11520 3062 11572 3068
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 11532 2689 11560 3062
rect 11612 2916 11664 2922
rect 11808 2904 11836 3470
rect 11900 3058 11928 5034
rect 11980 4548 12032 4554
rect 11980 4490 12032 4496
rect 11992 4214 12020 4490
rect 11980 4208 12032 4214
rect 11980 4150 12032 4156
rect 11978 3632 12034 3641
rect 11978 3567 11980 3576
rect 12032 3567 12034 3576
rect 11980 3538 12032 3544
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 12084 2972 12112 18550
rect 12346 18456 12402 18465
rect 12346 18391 12402 18400
rect 12360 18358 12388 18391
rect 12348 18352 12400 18358
rect 12544 18306 12572 19858
rect 12808 19848 12860 19854
rect 12806 19816 12808 19825
rect 12860 19816 12862 19825
rect 12806 19751 12862 19760
rect 12912 19514 12940 20402
rect 12992 20392 13044 20398
rect 13044 20352 13216 20380
rect 12992 20334 13044 20340
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 13096 19417 13124 20198
rect 13082 19408 13138 19417
rect 13082 19343 13138 19352
rect 13084 19304 13136 19310
rect 13084 19246 13136 19252
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12348 18294 12400 18300
rect 12452 18278 12572 18306
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 12176 16697 12204 18022
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 12162 16688 12218 16697
rect 12162 16623 12218 16632
rect 12164 15428 12216 15434
rect 12164 15370 12216 15376
rect 12176 12374 12204 15370
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 12268 10418 12296 17818
rect 12348 17740 12400 17746
rect 12348 17682 12400 17688
rect 12360 17649 12388 17682
rect 12346 17640 12402 17649
rect 12346 17575 12402 17584
rect 12452 17270 12480 18278
rect 12530 17776 12586 17785
rect 12530 17711 12586 17720
rect 12544 17270 12572 17711
rect 12440 17264 12492 17270
rect 12440 17206 12492 17212
rect 12532 17264 12584 17270
rect 12532 17206 12584 17212
rect 12636 17082 12664 18702
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12728 18193 12756 18362
rect 12714 18184 12770 18193
rect 12714 18119 12770 18128
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12728 17377 12756 18022
rect 12714 17368 12770 17377
rect 12714 17303 12770 17312
rect 12532 17060 12584 17066
rect 12636 17054 12756 17082
rect 12532 17002 12584 17008
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12360 16794 12388 16934
rect 12544 16810 12572 17002
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12452 16782 12572 16810
rect 12452 16726 12480 16782
rect 12440 16720 12492 16726
rect 12440 16662 12492 16668
rect 12348 16516 12400 16522
rect 12348 16458 12400 16464
rect 12360 13530 12388 16458
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12544 15026 12572 16390
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12440 14884 12492 14890
rect 12440 14826 12492 14832
rect 12452 14618 12480 14826
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12544 14521 12572 14554
rect 12530 14512 12586 14521
rect 12440 14476 12492 14482
rect 12530 14447 12586 14456
rect 12440 14418 12492 14424
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12346 13424 12402 13433
rect 12346 13359 12348 13368
rect 12400 13359 12402 13368
rect 12348 13330 12400 13336
rect 12452 13274 12480 14418
rect 12636 13734 12664 16934
rect 12728 16182 12756 17054
rect 12716 16176 12768 16182
rect 12716 16118 12768 16124
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12728 15366 12756 15982
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12728 13938 12756 14758
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12820 13818 12848 18702
rect 12900 18624 12952 18630
rect 12898 18592 12900 18601
rect 12952 18592 12954 18601
rect 12898 18527 12954 18536
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 12912 17746 12940 18226
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 13096 17542 13124 19246
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12728 13790 12848 13818
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12624 13456 12676 13462
rect 12624 13398 12676 13404
rect 12176 10390 12296 10418
rect 12360 13246 12480 13274
rect 12176 8090 12204 10390
rect 12360 10282 12388 13246
rect 12438 13152 12494 13161
rect 12438 13087 12494 13096
rect 12452 12782 12480 13087
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12452 12442 12480 12718
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12532 12368 12584 12374
rect 12532 12310 12584 12316
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12452 11898 12480 12242
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12544 11762 12572 12310
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12544 10713 12572 11562
rect 12530 10704 12586 10713
rect 12530 10639 12586 10648
rect 12268 10254 12388 10282
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12164 7472 12216 7478
rect 12164 7414 12216 7420
rect 12176 7274 12204 7414
rect 12164 7268 12216 7274
rect 12164 7210 12216 7216
rect 12176 6730 12204 7210
rect 12164 6724 12216 6730
rect 12164 6666 12216 6672
rect 12162 6488 12218 6497
rect 12162 6423 12218 6432
rect 12176 6322 12204 6423
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 12176 5234 12204 5510
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 12176 4486 12204 4966
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12162 4312 12218 4321
rect 12162 4247 12218 4256
rect 12176 3602 12204 4247
rect 12268 4078 12296 10254
rect 12346 10160 12402 10169
rect 12346 10095 12348 10104
rect 12400 10095 12402 10104
rect 12532 10124 12584 10130
rect 12348 10066 12400 10072
rect 12532 10066 12584 10072
rect 12346 9752 12402 9761
rect 12346 9687 12348 9696
rect 12400 9687 12402 9696
rect 12348 9658 12400 9664
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12360 9178 12388 9318
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12544 8906 12572 10066
rect 12636 9353 12664 13398
rect 12622 9344 12678 9353
rect 12622 9279 12678 9288
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 12348 8832 12400 8838
rect 12400 8792 12480 8820
rect 12348 8774 12400 8780
rect 12452 8786 12480 8792
rect 12452 8758 12664 8786
rect 12530 8664 12586 8673
rect 12530 8599 12586 8608
rect 12544 8566 12572 8599
rect 12636 8566 12664 8758
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12360 6458 12388 8026
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12544 7750 12572 7822
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12440 7336 12492 7342
rect 12636 7324 12664 8502
rect 12492 7296 12664 7324
rect 12440 7278 12492 7284
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12452 6322 12480 7278
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12346 6080 12402 6089
rect 12346 6015 12402 6024
rect 12360 5710 12388 6015
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12360 5098 12388 5646
rect 12452 5234 12480 6258
rect 12544 6186 12572 6802
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12348 5092 12400 5098
rect 12348 5034 12400 5040
rect 12544 4978 12572 6122
rect 12360 4950 12572 4978
rect 12360 4457 12388 4950
rect 12438 4856 12494 4865
rect 12438 4791 12494 4800
rect 12346 4448 12402 4457
rect 12346 4383 12402 4392
rect 12348 4208 12400 4214
rect 12348 4150 12400 4156
rect 12256 4072 12308 4078
rect 12256 4014 12308 4020
rect 12254 3768 12310 3777
rect 12254 3703 12256 3712
rect 12308 3703 12310 3712
rect 12256 3674 12308 3680
rect 12164 3596 12216 3602
rect 12164 3538 12216 3544
rect 12360 3534 12388 4150
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12164 3392 12216 3398
rect 12162 3360 12164 3369
rect 12216 3360 12218 3369
rect 12162 3295 12218 3304
rect 12346 3224 12402 3233
rect 12346 3159 12348 3168
rect 12400 3159 12402 3168
rect 12348 3130 12400 3136
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12084 2944 12296 2972
rect 11808 2876 12204 2904
rect 11612 2858 11664 2864
rect 11518 2680 11574 2689
rect 11518 2615 11574 2624
rect 11624 2378 11652 2858
rect 12070 2816 12126 2825
rect 12070 2751 12126 2760
rect 11886 2544 11942 2553
rect 11796 2508 11848 2514
rect 12084 2514 12112 2751
rect 11886 2479 11942 2488
rect 12072 2508 12124 2514
rect 11796 2450 11848 2456
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11256 2060 11468 2088
rect 11060 1488 11112 1494
rect 11060 1430 11112 1436
rect 11440 480 11468 2060
rect 11716 1630 11744 2382
rect 11808 2106 11836 2450
rect 11796 2100 11848 2106
rect 11796 2042 11848 2048
rect 11704 1624 11756 1630
rect 11704 1566 11756 1572
rect 11900 480 11928 2479
rect 12072 2450 12124 2456
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 11992 1902 12020 2382
rect 11980 1896 12032 1902
rect 11980 1838 12032 1844
rect 12176 1834 12204 2876
rect 12268 2417 12296 2944
rect 12360 2446 12388 2994
rect 12452 2922 12480 4791
rect 12544 4214 12572 4950
rect 12636 4622 12664 6122
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12622 4448 12678 4457
rect 12622 4383 12678 4392
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12532 3936 12584 3942
rect 12636 3924 12664 4383
rect 12728 3942 12756 13790
rect 12912 13462 12940 16934
rect 13004 14550 13032 17138
rect 13188 16697 13216 20352
rect 13280 18766 13308 22520
rect 13544 20324 13596 20330
rect 13544 20266 13596 20272
rect 13360 20256 13412 20262
rect 13360 20198 13412 20204
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 13372 17814 13400 20198
rect 13452 19236 13504 19242
rect 13452 19178 13504 19184
rect 13360 17808 13412 17814
rect 13360 17750 13412 17756
rect 13358 17232 13414 17241
rect 13358 17167 13414 17176
rect 13372 16833 13400 17167
rect 13358 16824 13414 16833
rect 13358 16759 13414 16768
rect 13174 16688 13230 16697
rect 13084 16652 13136 16658
rect 13174 16623 13230 16632
rect 13084 16594 13136 16600
rect 13096 14822 13124 16594
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 13188 16454 13216 16526
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 13188 15978 13216 16390
rect 13176 15972 13228 15978
rect 13176 15914 13228 15920
rect 13174 15056 13230 15065
rect 13174 14991 13176 15000
rect 13228 14991 13230 15000
rect 13176 14962 13228 14968
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13174 14784 13230 14793
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 12900 13456 12952 13462
rect 12900 13398 12952 13404
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12820 11762 12848 13262
rect 12900 13252 12952 13258
rect 12900 13194 12952 13200
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12820 11393 12848 11494
rect 12806 11384 12862 11393
rect 12806 11319 12862 11328
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12820 7206 12848 10406
rect 12912 9654 12940 13194
rect 13096 12374 13124 14758
rect 13174 14719 13230 14728
rect 13188 14346 13216 14719
rect 13176 14340 13228 14346
rect 13176 14282 13228 14288
rect 13174 13696 13230 13705
rect 13174 13631 13230 13640
rect 13084 12368 13136 12374
rect 13084 12310 13136 12316
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 12990 11520 13046 11529
rect 12990 11455 13046 11464
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 13004 7993 13032 11455
rect 13096 11121 13124 11698
rect 13188 11694 13216 13631
rect 13280 13258 13308 16526
rect 13372 16522 13400 16759
rect 13360 16516 13412 16522
rect 13360 16458 13412 16464
rect 13360 14884 13412 14890
rect 13360 14826 13412 14832
rect 13372 14278 13400 14826
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13372 13734 13400 13806
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13266 12880 13322 12889
rect 13464 12866 13492 19178
rect 13556 19009 13584 20266
rect 13542 19000 13598 19009
rect 13542 18935 13598 18944
rect 13544 18828 13596 18834
rect 13544 18770 13596 18776
rect 13556 13705 13584 18770
rect 13636 18760 13688 18766
rect 13636 18702 13688 18708
rect 13648 16590 13676 18702
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13636 15972 13688 15978
rect 13636 15914 13688 15920
rect 13648 15706 13676 15914
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13636 15020 13688 15026
rect 13636 14962 13688 14968
rect 13542 13696 13598 13705
rect 13542 13631 13598 13640
rect 13542 13560 13598 13569
rect 13542 13495 13598 13504
rect 13556 13462 13584 13495
rect 13544 13456 13596 13462
rect 13544 13398 13596 13404
rect 13648 12918 13676 14962
rect 13636 12912 13688 12918
rect 13464 12838 13584 12866
rect 13636 12854 13688 12860
rect 13266 12815 13322 12824
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13082 11112 13138 11121
rect 13082 11047 13138 11056
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 13096 10305 13124 10474
rect 13188 10441 13216 11630
rect 13174 10432 13230 10441
rect 13174 10367 13230 10376
rect 13082 10296 13138 10305
rect 13082 10231 13138 10240
rect 13176 10192 13228 10198
rect 13176 10134 13228 10140
rect 13188 9926 13216 10134
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13096 8090 13124 9658
rect 13188 9586 13216 9862
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 12990 7984 13046 7993
rect 12990 7919 13046 7928
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 12808 7200 12860 7206
rect 12912 7177 12940 7210
rect 12808 7142 12860 7148
rect 12898 7168 12954 7177
rect 12898 7103 12954 7112
rect 12900 6180 12952 6186
rect 12900 6122 12952 6128
rect 12912 5914 12940 6122
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 12820 5545 12848 5782
rect 12806 5536 12862 5545
rect 12806 5471 12862 5480
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12820 4593 12848 4966
rect 12806 4584 12862 4593
rect 12806 4519 12862 4528
rect 12584 3896 12664 3924
rect 12716 3936 12768 3942
rect 12532 3878 12584 3884
rect 12716 3878 12768 3884
rect 12806 3904 12862 3913
rect 12806 3839 12862 3848
rect 12530 3768 12586 3777
rect 12530 3703 12586 3712
rect 12544 3602 12572 3703
rect 12820 3602 12848 3839
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12440 2916 12492 2922
rect 12440 2858 12492 2864
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12636 2650 12664 2790
rect 12728 2650 12756 3470
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12348 2440 12400 2446
rect 12254 2408 12310 2417
rect 12348 2382 12400 2388
rect 12254 2343 12310 2352
rect 12268 1902 12296 2343
rect 13004 2038 13032 7822
rect 13084 7812 13136 7818
rect 13084 7754 13136 7760
rect 13096 7546 13124 7754
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13096 7206 13124 7482
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 13096 6254 13124 7142
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 13096 3058 13124 5102
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 12992 2032 13044 2038
rect 12992 1974 13044 1980
rect 12256 1896 12308 1902
rect 12256 1838 12308 1844
rect 12164 1828 12216 1834
rect 12164 1770 12216 1776
rect 12808 1828 12860 1834
rect 12808 1770 12860 1776
rect 12346 1456 12402 1465
rect 12346 1391 12402 1400
rect 12360 480 12388 1391
rect 12820 480 12848 1770
rect 13188 1630 13216 7482
rect 13280 1834 13308 12815
rect 13556 12322 13584 12838
rect 13648 12374 13676 12854
rect 13372 12294 13584 12322
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 13372 4078 13400 12294
rect 13636 12096 13688 12102
rect 13450 12064 13506 12073
rect 13636 12038 13688 12044
rect 13450 11999 13506 12008
rect 13464 7546 13492 11999
rect 13648 11354 13676 12038
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13542 9888 13598 9897
rect 13542 9823 13598 9832
rect 13556 8537 13584 9823
rect 13648 9722 13676 10950
rect 13740 10418 13768 22520
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 14002 19952 14058 19961
rect 13912 19916 13964 19922
rect 14002 19887 14058 19896
rect 13912 19858 13964 19864
rect 13820 18148 13872 18154
rect 13820 18090 13872 18096
rect 13832 17678 13860 18090
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13924 17134 13952 19858
rect 14016 19446 14044 19887
rect 14004 19440 14056 19446
rect 14004 19382 14056 19388
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 14016 18630 14044 19110
rect 14004 18624 14056 18630
rect 14004 18566 14056 18572
rect 14004 18080 14056 18086
rect 14004 18022 14056 18028
rect 14016 17785 14044 18022
rect 14002 17776 14058 17785
rect 14002 17711 14058 17720
rect 14004 17672 14056 17678
rect 14002 17640 14004 17649
rect 14056 17640 14058 17649
rect 14002 17575 14058 17584
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 13910 16688 13966 16697
rect 13910 16623 13966 16632
rect 14004 16652 14056 16658
rect 13924 15910 13952 16623
rect 14004 16594 14056 16600
rect 13912 15904 13964 15910
rect 13910 15872 13912 15881
rect 13964 15872 13966 15881
rect 13910 15807 13966 15816
rect 14016 15706 14044 16594
rect 14108 15706 14136 20538
rect 14292 19281 14320 22520
rect 14752 20058 14780 22520
rect 15212 20602 15240 22520
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 15382 19816 15438 19825
rect 15200 19780 15252 19786
rect 15382 19751 15438 19760
rect 15200 19722 15252 19728
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14464 19304 14516 19310
rect 14278 19272 14334 19281
rect 14464 19246 14516 19252
rect 14278 19207 14334 19216
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14004 15496 14056 15502
rect 14004 15438 14056 15444
rect 13818 14920 13874 14929
rect 13818 14855 13874 14864
rect 13832 11937 13860 14855
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 13924 14006 13952 14350
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 14016 13852 14044 15438
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 14108 14822 14136 15302
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14108 14006 14136 14758
rect 14096 14000 14148 14006
rect 14094 13968 14096 13977
rect 14148 13968 14150 13977
rect 14094 13903 14150 13912
rect 13924 13824 14044 13852
rect 14096 13864 14148 13870
rect 13818 11928 13874 11937
rect 13818 11863 13874 11872
rect 13924 11082 13952 13824
rect 14096 13806 14148 13812
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 14016 11286 14044 13126
rect 14108 11354 14136 13806
rect 14200 12345 14228 18158
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14292 17338 14320 17614
rect 14280 17332 14332 17338
rect 14280 17274 14332 17280
rect 14280 15088 14332 15094
rect 14280 15030 14332 15036
rect 14292 14618 14320 15030
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14292 12442 14320 14418
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14186 12336 14242 12345
rect 14186 12271 14242 12280
rect 14186 12200 14242 12209
rect 14186 12135 14242 12144
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14004 11280 14056 11286
rect 14004 11222 14056 11228
rect 13912 11076 13964 11082
rect 13912 11018 13964 11024
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14108 10577 14136 10746
rect 14094 10568 14150 10577
rect 14094 10503 14150 10512
rect 14096 10464 14148 10470
rect 13740 10390 14044 10418
rect 14096 10406 14148 10412
rect 13820 10056 13872 10062
rect 13726 10024 13782 10033
rect 13820 9998 13872 10004
rect 13726 9959 13782 9968
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13542 8528 13598 8537
rect 13542 8463 13598 8472
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13648 7721 13676 8026
rect 13634 7712 13690 7721
rect 13634 7647 13690 7656
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13740 7342 13768 9959
rect 13832 9178 13860 9998
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13924 9722 13952 9862
rect 14016 9722 14044 10390
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 14108 9466 14136 10406
rect 14200 9926 14228 12135
rect 14278 11928 14334 11937
rect 14278 11863 14334 11872
rect 14292 11830 14320 11863
rect 14280 11824 14332 11830
rect 14280 11766 14332 11772
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14292 10742 14320 11630
rect 14384 10849 14412 18022
rect 14476 14482 14504 19246
rect 14568 15638 14596 19450
rect 15016 19372 15068 19378
rect 14660 19332 15016 19360
rect 14556 15632 14608 15638
rect 14556 15574 14608 15580
rect 14556 15088 14608 15094
rect 14556 15030 14608 15036
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14476 13326 14504 13874
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14464 13184 14516 13190
rect 14462 13152 14464 13161
rect 14516 13152 14518 13161
rect 14462 13087 14518 13096
rect 14476 11762 14504 13087
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14370 10840 14426 10849
rect 14370 10775 14426 10784
rect 14280 10736 14332 10742
rect 14476 10690 14504 11290
rect 14280 10678 14332 10684
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 13924 9438 14136 9466
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13832 8090 13860 8910
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13452 6248 13504 6254
rect 13452 6190 13504 6196
rect 13464 4758 13492 6190
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13634 5808 13690 5817
rect 13634 5743 13690 5752
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13556 5001 13584 5510
rect 13542 4992 13598 5001
rect 13542 4927 13598 4936
rect 13648 4758 13676 5743
rect 13452 4752 13504 4758
rect 13452 4694 13504 4700
rect 13636 4752 13688 4758
rect 13636 4694 13688 4700
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13268 1828 13320 1834
rect 13268 1770 13320 1776
rect 13176 1624 13228 1630
rect 13176 1566 13228 1572
rect 13464 1442 13492 3878
rect 13556 3194 13584 4626
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13648 4282 13676 4558
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13740 3534 13768 6054
rect 13832 5914 13860 7890
rect 13924 6254 13952 9438
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 14016 9110 14044 9318
rect 14094 9208 14150 9217
rect 14094 9143 14096 9152
rect 14148 9143 14150 9152
rect 14096 9114 14148 9120
rect 14004 9104 14056 9110
rect 14004 9046 14056 9052
rect 14200 8956 14228 9658
rect 14292 9518 14320 10678
rect 14384 10662 14504 10690
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14016 8928 14228 8956
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13924 5710 13952 6054
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13924 5166 13952 5646
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13832 4622 13860 4966
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13910 4040 13966 4049
rect 13910 3975 13912 3984
rect 13964 3975 13966 3984
rect 13912 3946 13964 3952
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 14016 3398 14044 8928
rect 14292 8634 14320 9318
rect 14384 8809 14412 10662
rect 14464 10600 14516 10606
rect 14464 10542 14516 10548
rect 14476 9586 14504 10542
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14476 9217 14504 9522
rect 14462 9208 14518 9217
rect 14462 9143 14464 9152
rect 14516 9143 14518 9152
rect 14464 9114 14516 9120
rect 14476 9083 14504 9114
rect 14370 8800 14426 8809
rect 14370 8735 14426 8744
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14278 8528 14334 8537
rect 14278 8463 14334 8472
rect 14292 8362 14320 8463
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 14096 8016 14148 8022
rect 14096 7958 14148 7964
rect 14108 4554 14136 7958
rect 14292 6798 14320 8298
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14096 4548 14148 4554
rect 14096 4490 14148 4496
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 14108 3602 14136 4014
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 14096 3460 14148 3466
rect 14096 3402 14148 3408
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 13728 2372 13780 2378
rect 13728 2314 13780 2320
rect 13280 1414 13492 1442
rect 13280 480 13308 1414
rect 13740 480 13768 2314
rect 13832 2310 13860 2586
rect 13820 2304 13872 2310
rect 13820 2246 13872 2252
rect 14108 1714 14136 3402
rect 14200 2009 14228 4558
rect 14384 4321 14412 7822
rect 14462 7576 14518 7585
rect 14462 7511 14518 7520
rect 14476 5642 14504 7511
rect 14568 7041 14596 15030
rect 14554 7032 14610 7041
rect 14554 6967 14610 6976
rect 14554 6760 14610 6769
rect 14554 6695 14610 6704
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 14568 5370 14596 6695
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14660 5250 14688 19332
rect 15016 19314 15068 19320
rect 15212 19174 15240 19722
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 15198 19000 15254 19009
rect 15198 18935 15254 18944
rect 15212 18902 15240 18935
rect 15200 18896 15252 18902
rect 15200 18838 15252 18844
rect 15304 18766 15332 19246
rect 15292 18760 15344 18766
rect 15198 18728 15254 18737
rect 15292 18702 15344 18708
rect 15198 18663 15254 18672
rect 15212 18630 15240 18663
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 15200 18352 15252 18358
rect 14738 18320 14794 18329
rect 15200 18294 15252 18300
rect 14738 18255 14740 18264
rect 14792 18255 14794 18264
rect 14740 18226 14792 18232
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14752 17202 14780 18022
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 14922 17640 14978 17649
rect 14922 17575 14978 17584
rect 14936 17377 14964 17575
rect 14922 17368 14978 17377
rect 14922 17303 14978 17312
rect 15106 17368 15162 17377
rect 15106 17303 15162 17312
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 15120 17134 15148 17303
rect 15108 17128 15160 17134
rect 15108 17070 15160 17076
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14752 15502 14780 16934
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 14924 15632 14976 15638
rect 14924 15574 14976 15580
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 14740 14952 14792 14958
rect 14738 14920 14740 14929
rect 14792 14920 14794 14929
rect 14936 14890 14964 15574
rect 15106 15192 15162 15201
rect 15106 15127 15162 15136
rect 15120 14958 15148 15127
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 14738 14855 14794 14864
rect 14924 14884 14976 14890
rect 14924 14826 14976 14832
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14752 12889 14780 14758
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 15212 14482 15240 18294
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15304 17134 15332 18226
rect 15396 18154 15424 19751
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15672 18850 15700 22520
rect 16132 20058 16160 22520
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16304 19780 16356 19786
rect 16304 19722 16356 19728
rect 15488 18193 15516 18838
rect 15672 18822 15976 18850
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15474 18184 15530 18193
rect 15384 18148 15436 18154
rect 15474 18119 15530 18128
rect 15384 18090 15436 18096
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15304 16590 15332 17070
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15396 15994 15424 17682
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 15488 16114 15516 16526
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15396 15966 15516 15994
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15304 15570 15332 15846
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 14738 12880 14794 12889
rect 14738 12815 14794 12824
rect 14740 12708 14792 12714
rect 14740 12650 14792 12656
rect 14752 11150 14780 12650
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 15120 11626 15148 12242
rect 15108 11620 15160 11626
rect 15108 11562 15160 11568
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 15212 11286 15240 13738
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15200 11280 15252 11286
rect 15200 11222 15252 11228
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14844 10452 14872 11018
rect 15198 10976 15254 10985
rect 15198 10911 15254 10920
rect 14752 10424 14872 10452
rect 14752 9489 14780 10424
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 14738 9480 14794 9489
rect 14738 9415 14794 9424
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 14740 9104 14792 9110
rect 14740 9046 14792 9052
rect 14752 8090 14780 9046
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14568 5222 14688 5250
rect 14370 4312 14426 4321
rect 14370 4247 14426 4256
rect 14280 4208 14332 4214
rect 14332 4168 14412 4196
rect 14280 4150 14332 4156
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14292 2689 14320 3946
rect 14384 2990 14412 4168
rect 14568 4078 14596 5222
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14660 4282 14688 5102
rect 14752 5098 14780 6802
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 15028 6254 15056 6598
rect 15016 6248 15068 6254
rect 15016 6190 15068 6196
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 14740 5092 14792 5098
rect 14740 5034 14792 5040
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14556 4072 14608 4078
rect 14556 4014 14608 4020
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 14278 2680 14334 2689
rect 14278 2615 14334 2624
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14186 2000 14242 2009
rect 14186 1935 14242 1944
rect 14384 1766 14412 2450
rect 14372 1760 14424 1766
rect 14108 1686 14320 1714
rect 14372 1702 14424 1708
rect 14476 1698 14504 2790
rect 14568 2446 14596 2994
rect 14752 2582 14780 5034
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 15212 4758 15240 10911
rect 15304 9926 15332 12174
rect 15396 11642 15424 15846
rect 15488 13734 15516 15966
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 12442 15516 13670
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15396 11614 15516 11642
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15396 10266 15424 11494
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15488 9738 15516 11614
rect 15580 10674 15608 18566
rect 15750 18184 15806 18193
rect 15750 18119 15806 18128
rect 15764 17746 15792 18119
rect 15752 17740 15804 17746
rect 15752 17682 15804 17688
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 15672 14346 15700 17002
rect 15764 15162 15792 17682
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15856 16454 15884 17614
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15672 12102 15700 13262
rect 15856 12594 15884 15438
rect 15948 14385 15976 18822
rect 16028 18828 16080 18834
rect 16028 18770 16080 18776
rect 16040 18737 16068 18770
rect 16120 18760 16172 18766
rect 16026 18728 16082 18737
rect 16120 18702 16172 18708
rect 16026 18663 16082 18672
rect 16132 18086 16160 18702
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 16132 17921 16160 18022
rect 16118 17912 16174 17921
rect 16118 17847 16174 17856
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 16040 17241 16068 17682
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 16026 17232 16082 17241
rect 16026 17167 16082 17176
rect 16120 16992 16172 16998
rect 16120 16934 16172 16940
rect 16132 16726 16160 16934
rect 16224 16726 16252 17478
rect 16120 16720 16172 16726
rect 16120 16662 16172 16668
rect 16212 16720 16264 16726
rect 16212 16662 16264 16668
rect 16028 16448 16080 16454
rect 16028 16390 16080 16396
rect 15934 14376 15990 14385
rect 15934 14311 15990 14320
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 15948 14006 15976 14214
rect 15936 14000 15988 14006
rect 15936 13942 15988 13948
rect 16040 13954 16068 16390
rect 16132 16114 16160 16662
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16316 16046 16344 19722
rect 16396 19236 16448 19242
rect 16396 19178 16448 19184
rect 16408 19009 16436 19178
rect 16394 19000 16450 19009
rect 16394 18935 16450 18944
rect 16396 18080 16448 18086
rect 16592 18034 16620 22520
rect 16948 19984 17000 19990
rect 16948 19926 17000 19932
rect 16854 18592 16910 18601
rect 16854 18527 16910 18536
rect 16868 18290 16896 18527
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 16396 18022 16448 18028
rect 16408 17678 16436 18022
rect 16500 18006 16620 18034
rect 16500 17814 16528 18006
rect 16488 17808 16540 17814
rect 16488 17750 16540 17756
rect 16672 17808 16724 17814
rect 16672 17750 16724 17756
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 16684 17377 16712 17750
rect 16670 17368 16726 17377
rect 16670 17303 16726 17312
rect 16580 16176 16632 16182
rect 16580 16118 16632 16124
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 16488 15972 16540 15978
rect 16488 15914 16540 15920
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16212 15632 16264 15638
rect 16212 15574 16264 15580
rect 16040 13926 16160 13954
rect 16132 13870 16160 13926
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 15936 13388 15988 13394
rect 15936 13330 15988 13336
rect 15764 12566 15884 12594
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15672 10538 15700 12038
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15566 10296 15622 10305
rect 15566 10231 15568 10240
rect 15620 10231 15622 10240
rect 15568 10202 15620 10208
rect 15660 10192 15712 10198
rect 15566 10160 15622 10169
rect 15660 10134 15712 10140
rect 15566 10095 15622 10104
rect 15304 9710 15516 9738
rect 15200 4752 15252 4758
rect 15200 4694 15252 4700
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 15200 3664 15252 3670
rect 15304 3652 15332 9710
rect 15580 9518 15608 10095
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15396 8090 15424 8910
rect 15488 8634 15516 9386
rect 15580 9042 15608 9454
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15488 7886 15516 8570
rect 15672 8294 15700 10134
rect 15764 9625 15792 12566
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 15856 11150 15884 11698
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15856 10810 15884 11086
rect 15948 11082 15976 13330
rect 16040 12918 16068 13806
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 16040 12238 16068 12854
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 16040 11354 16068 11494
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 15936 11076 15988 11082
rect 15936 11018 15988 11024
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 15856 9908 15884 10610
rect 16040 10538 16068 10610
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 15948 10198 15976 10406
rect 15936 10192 15988 10198
rect 15936 10134 15988 10140
rect 16040 10062 16068 10474
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 16028 10056 16080 10062
rect 16132 10033 16160 10066
rect 16028 9998 16080 10004
rect 16118 10024 16174 10033
rect 16118 9959 16174 9968
rect 15856 9880 16068 9908
rect 15750 9616 15806 9625
rect 16040 9602 16068 9880
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 15750 9551 15806 9560
rect 15948 9574 16068 9602
rect 15752 9444 15804 9450
rect 15752 9386 15804 9392
rect 15764 8838 15792 9386
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15672 8106 15700 8230
rect 15672 8078 15792 8106
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15476 7880 15528 7886
rect 15528 7840 15608 7868
rect 15476 7822 15528 7828
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15396 7342 15424 7686
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15488 6458 15516 7142
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15580 6322 15608 7840
rect 15568 6316 15620 6322
rect 15568 6258 15620 6264
rect 15382 5536 15438 5545
rect 15382 5471 15438 5480
rect 15396 5030 15424 5471
rect 15566 5400 15622 5409
rect 15672 5386 15700 7890
rect 15764 7546 15792 8078
rect 15856 7993 15884 8910
rect 15842 7984 15898 7993
rect 15842 7919 15898 7928
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 15750 6488 15806 6497
rect 15750 6423 15806 6432
rect 15764 5545 15792 6423
rect 15856 5778 15884 6802
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15750 5536 15806 5545
rect 15750 5471 15806 5480
rect 15622 5358 15700 5386
rect 15566 5335 15622 5344
rect 15856 5166 15884 5714
rect 15948 5545 15976 9574
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 16040 8537 16068 8910
rect 16026 8528 16082 8537
rect 16026 8463 16082 8472
rect 16040 7750 16068 8463
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 16132 7410 16160 9658
rect 16224 9518 16252 15574
rect 16408 15026 16436 15846
rect 16500 15502 16528 15914
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 16396 15020 16448 15026
rect 16396 14962 16448 14968
rect 16396 14884 16448 14890
rect 16396 14826 16448 14832
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16132 6934 16160 7346
rect 16120 6928 16172 6934
rect 16120 6870 16172 6876
rect 16224 6866 16252 9114
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16120 6452 16172 6458
rect 16120 6394 16172 6400
rect 16132 5624 16160 6394
rect 16123 5596 16160 5624
rect 16123 5556 16151 5596
rect 15934 5536 15990 5545
rect 16123 5528 16160 5556
rect 15934 5471 15990 5480
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15566 4720 15622 4729
rect 15566 4655 15622 4664
rect 15842 4720 15898 4729
rect 15842 4655 15898 4664
rect 15252 3624 15332 3652
rect 15384 3664 15436 3670
rect 15200 3606 15252 3612
rect 15384 3606 15436 3612
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 14740 2576 14792 2582
rect 14740 2518 14792 2524
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14292 480 14320 1686
rect 14464 1692 14516 1698
rect 14464 1634 14516 1640
rect 14752 480 14780 2246
rect 15212 480 15240 2790
rect 15396 2650 15424 3606
rect 15580 2990 15608 4655
rect 15856 4554 15884 4655
rect 15844 4548 15896 4554
rect 15844 4490 15896 4496
rect 16040 4214 16068 5238
rect 16028 4208 16080 4214
rect 16028 4150 16080 4156
rect 16132 3738 16160 5528
rect 16316 4146 16344 11630
rect 16408 9042 16436 14826
rect 16500 13977 16528 15438
rect 16486 13968 16542 13977
rect 16486 13903 16542 13912
rect 16500 13394 16528 13903
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16592 12646 16620 16118
rect 16672 15700 16724 15706
rect 16672 15642 16724 15648
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16684 12458 16712 15642
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16868 13954 16896 14894
rect 16960 14113 16988 19926
rect 17052 19310 17080 22520
rect 17408 19916 17460 19922
rect 17408 19858 17460 19864
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 17222 18864 17278 18873
rect 17222 18799 17224 18808
rect 17276 18799 17278 18808
rect 17224 18770 17276 18776
rect 17314 18456 17370 18465
rect 17314 18391 17370 18400
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 17052 15910 17080 18226
rect 17328 17678 17356 18391
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 17040 14816 17092 14822
rect 17040 14758 17092 14764
rect 16946 14104 17002 14113
rect 16946 14039 17002 14048
rect 16868 13926 16988 13954
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16868 13462 16896 13806
rect 16856 13456 16908 13462
rect 16856 13398 16908 13404
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 16592 12430 16712 12458
rect 16592 10690 16620 12430
rect 16776 12306 16804 13330
rect 16960 12322 16988 13926
rect 17052 13870 17080 14758
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 17038 13424 17094 13433
rect 17038 13359 17094 13368
rect 17052 12918 17080 13359
rect 17040 12912 17092 12918
rect 17040 12854 17092 12860
rect 16764 12300 16816 12306
rect 16960 12294 17080 12322
rect 16764 12242 16816 12248
rect 16672 11620 16724 11626
rect 16672 11562 16724 11568
rect 16684 10810 16712 11562
rect 16776 11218 16804 12242
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 16764 11212 16816 11218
rect 16764 11154 16816 11160
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16592 10662 16712 10690
rect 16684 9636 16712 10662
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16776 9897 16804 10542
rect 16856 10532 16908 10538
rect 16856 10474 16908 10480
rect 16762 9888 16818 9897
rect 16762 9823 16818 9832
rect 16592 9608 16712 9636
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 16408 5114 16436 5714
rect 16500 5234 16528 8842
rect 16592 5681 16620 9608
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16684 7585 16712 9454
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16776 8430 16804 8774
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16670 7576 16726 7585
rect 16670 7511 16726 7520
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16578 5672 16634 5681
rect 16578 5607 16634 5616
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 16592 5370 16620 5510
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16408 5086 16528 5114
rect 16500 4622 16528 5086
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 16500 4282 16528 4558
rect 16488 4276 16540 4282
rect 16488 4218 16540 4224
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 15660 3120 15712 3126
rect 15660 3062 15712 3068
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 15488 1873 15516 2314
rect 15474 1864 15530 1873
rect 15474 1799 15530 1808
rect 15672 480 15700 3062
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 15948 2922 15976 2994
rect 15936 2916 15988 2922
rect 15936 2858 15988 2864
rect 15948 2650 15976 2858
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 16132 480 16160 3334
rect 16684 2990 16712 7210
rect 16776 4457 16804 8230
rect 16868 5166 16896 10474
rect 16960 8673 16988 11766
rect 17052 9450 17080 12294
rect 17040 9444 17092 9450
rect 17040 9386 17092 9392
rect 16946 8664 17002 8673
rect 16946 8599 17002 8608
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16960 8022 16988 8434
rect 17144 8401 17172 17478
rect 17236 12714 17264 17478
rect 17328 17202 17356 17614
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 17316 16448 17368 16454
rect 17316 16390 17368 16396
rect 17328 15570 17356 16390
rect 17420 16046 17448 19858
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17316 15564 17368 15570
rect 17316 15506 17368 15512
rect 17328 15026 17356 15506
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17328 13530 17356 14350
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17314 13424 17370 13433
rect 17314 13359 17370 13368
rect 17224 12708 17276 12714
rect 17224 12650 17276 12656
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 17236 9654 17264 11494
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 17130 8392 17186 8401
rect 17130 8327 17186 8336
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 16948 8016 17000 8022
rect 16948 7958 17000 7964
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 17052 6322 17080 7686
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16762 4448 16818 4457
rect 16762 4383 16818 4392
rect 16960 3602 16988 6190
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 17144 3058 17172 7142
rect 17236 5574 17264 8298
rect 17224 5568 17276 5574
rect 17224 5510 17276 5516
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 16580 1284 16632 1290
rect 16580 1226 16632 1232
rect 16592 480 16620 1226
rect 17052 480 17080 2790
rect 17236 2514 17264 4966
rect 17328 3194 17356 13359
rect 17420 12714 17448 15846
rect 17408 12708 17460 12714
rect 17408 12650 17460 12656
rect 17512 11257 17540 22520
rect 17776 20392 17828 20398
rect 17776 20334 17828 20340
rect 17590 19408 17646 19417
rect 17590 19343 17646 19352
rect 17604 17270 17632 19343
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 17696 18426 17724 18702
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 17684 18148 17736 18154
rect 17684 18090 17736 18096
rect 17592 17264 17644 17270
rect 17592 17206 17644 17212
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17604 15706 17632 15982
rect 17592 15700 17644 15706
rect 17592 15642 17644 15648
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 17604 15094 17632 15370
rect 17592 15088 17644 15094
rect 17592 15030 17644 15036
rect 17696 11801 17724 18090
rect 17788 12918 17816 20334
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17880 14958 17908 19790
rect 17972 18902 18000 22520
rect 18432 20890 18460 22520
rect 18156 20862 18460 20890
rect 18156 20058 18184 20862
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18880 19916 18932 19922
rect 18880 19858 18932 19864
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18786 19136 18842 19145
rect 18786 19071 18842 19080
rect 17960 18896 18012 18902
rect 17960 18838 18012 18844
rect 18696 18828 18748 18834
rect 18696 18770 18748 18776
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 17958 17776 18014 17785
rect 17958 17711 18014 17720
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17972 14346 18000 17711
rect 17960 14340 18012 14346
rect 17960 14282 18012 14288
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17776 12912 17828 12918
rect 17776 12854 17828 12860
rect 17776 12708 17828 12714
rect 17776 12650 17828 12656
rect 17682 11792 17738 11801
rect 17682 11727 17738 11736
rect 17498 11248 17554 11257
rect 17498 11183 17554 11192
rect 17500 10736 17552 10742
rect 17406 10704 17462 10713
rect 17500 10678 17552 10684
rect 17406 10639 17462 10648
rect 17420 10062 17448 10639
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17512 9874 17540 10678
rect 17682 10568 17738 10577
rect 17682 10503 17738 10512
rect 17696 10470 17724 10503
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17420 9846 17540 9874
rect 17420 5817 17448 9846
rect 17590 9752 17646 9761
rect 17500 9716 17552 9722
rect 17590 9687 17646 9696
rect 17500 9658 17552 9664
rect 17512 6458 17540 9658
rect 17604 7834 17632 9687
rect 17604 7806 17724 7834
rect 17592 7268 17644 7274
rect 17592 7210 17644 7216
rect 17604 6662 17632 7210
rect 17592 6656 17644 6662
rect 17592 6598 17644 6604
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17406 5808 17462 5817
rect 17406 5743 17462 5752
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17420 4622 17448 5646
rect 17604 4758 17632 6598
rect 17592 4752 17644 4758
rect 17592 4694 17644 4700
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17604 4486 17632 4694
rect 17592 4480 17644 4486
rect 17592 4422 17644 4428
rect 17696 3913 17724 7806
rect 17788 6254 17816 12650
rect 17880 11218 17908 13466
rect 17972 12782 18000 13738
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17972 10656 18000 11834
rect 17880 10628 18000 10656
rect 17880 9722 17908 10628
rect 17960 10532 18012 10538
rect 17960 10474 18012 10480
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17972 9586 18000 10474
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17880 9178 17908 9454
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17880 8650 17908 9114
rect 18064 9081 18092 18022
rect 18156 16726 18184 18566
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18234 17912 18290 17921
rect 18234 17847 18290 17856
rect 18604 17876 18656 17882
rect 18248 17678 18276 17847
rect 18604 17818 18656 17824
rect 18512 17740 18564 17746
rect 18512 17682 18564 17688
rect 18236 17672 18288 17678
rect 18524 17649 18552 17682
rect 18236 17614 18288 17620
rect 18510 17640 18566 17649
rect 18510 17575 18566 17584
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 18420 17264 18472 17270
rect 18420 17206 18472 17212
rect 18144 16720 18196 16726
rect 18144 16662 18196 16668
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 18156 16114 18184 16526
rect 18432 16522 18460 17206
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 18420 16516 18472 16522
rect 18420 16458 18472 16464
rect 18524 16436 18552 17138
rect 18616 16726 18644 17818
rect 18604 16720 18656 16726
rect 18604 16662 18656 16668
rect 18524 16408 18644 16436
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18144 16108 18196 16114
rect 18144 16050 18196 16056
rect 18144 15496 18196 15502
rect 18142 15464 18144 15473
rect 18196 15464 18198 15473
rect 18142 15399 18198 15408
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 18420 15088 18472 15094
rect 18420 15030 18472 15036
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 18156 14482 18184 14894
rect 18432 14822 18460 15030
rect 18616 14822 18644 16408
rect 18236 14816 18288 14822
rect 18236 14758 18288 14764
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18248 14634 18276 14758
rect 18248 14618 18368 14634
rect 18248 14612 18380 14618
rect 18248 14606 18328 14612
rect 18328 14554 18380 14560
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 18156 12782 18184 14214
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 18248 13462 18276 13806
rect 18236 13456 18288 13462
rect 18236 13398 18288 13404
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 18616 12374 18644 12786
rect 18144 12368 18196 12374
rect 18144 12310 18196 12316
rect 18604 12368 18656 12374
rect 18604 12310 18656 12316
rect 18156 11354 18184 12310
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18248 10996 18276 11494
rect 18156 10968 18276 10996
rect 18050 9072 18106 9081
rect 18050 9007 18106 9016
rect 17880 8622 18092 8650
rect 17960 8560 18012 8566
rect 17960 8502 18012 8508
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17880 6866 17908 8434
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 17880 5778 17908 6666
rect 17972 6254 18000 8502
rect 18064 8430 18092 8622
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 18064 8090 18092 8366
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 18064 6662 18092 7890
rect 18156 7857 18184 10968
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18616 10062 18644 12038
rect 18708 11626 18736 18770
rect 18696 11620 18748 11626
rect 18696 11562 18748 11568
rect 18800 11098 18828 19071
rect 18892 15609 18920 19858
rect 18984 19281 19012 22520
rect 19444 20602 19472 22520
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19904 20074 19932 22520
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 19812 20058 19932 20074
rect 19800 20052 19932 20058
rect 19852 20046 19932 20052
rect 19800 19994 19852 20000
rect 19616 19304 19668 19310
rect 18970 19272 19026 19281
rect 19616 19246 19668 19252
rect 18970 19207 19026 19216
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18878 15600 18934 15609
rect 18878 15535 18934 15544
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18892 14414 18920 15302
rect 18984 14958 19012 18226
rect 19064 17876 19116 17882
rect 19064 17818 19116 17824
rect 19076 17542 19104 17818
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 19064 16992 19116 16998
rect 19062 16960 19064 16969
rect 19116 16960 19118 16969
rect 19062 16895 19118 16904
rect 19064 16176 19116 16182
rect 19064 16118 19116 16124
rect 18972 14952 19024 14958
rect 18972 14894 19024 14900
rect 18972 14544 19024 14550
rect 18972 14486 19024 14492
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 18892 13462 18920 14350
rect 18984 13530 19012 14486
rect 18972 13524 19024 13530
rect 18972 13466 19024 13472
rect 18880 13456 18932 13462
rect 18880 13398 18932 13404
rect 18878 12744 18934 12753
rect 18878 12679 18934 12688
rect 18972 12708 19024 12714
rect 18892 11626 18920 12679
rect 18972 12650 19024 12656
rect 18880 11620 18932 11626
rect 18880 11562 18932 11568
rect 18708 11070 18828 11098
rect 18604 10056 18656 10062
rect 18604 9998 18656 10004
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18604 9512 18656 9518
rect 18604 9454 18656 9460
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18616 8294 18644 9454
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18708 8022 18736 11070
rect 18788 11008 18840 11014
rect 18788 10950 18840 10956
rect 18800 10266 18828 10950
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18800 9450 18828 9998
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 18892 9178 18920 11562
rect 18984 11354 19012 12650
rect 19076 11898 19104 16118
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 19168 14521 19196 15506
rect 19154 14512 19210 14521
rect 19154 14447 19210 14456
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 19064 11756 19116 11762
rect 19064 11698 19116 11704
rect 18972 11348 19024 11354
rect 18972 11290 19024 11296
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 19076 9110 19104 11698
rect 19168 11529 19196 13874
rect 19260 12594 19288 17614
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19352 16114 19380 16390
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19352 15502 19380 16050
rect 19524 15972 19576 15978
rect 19524 15914 19576 15920
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19352 15026 19380 15438
rect 19536 15162 19564 15914
rect 19628 15434 19656 19246
rect 19892 17740 19944 17746
rect 19892 17682 19944 17688
rect 19708 17128 19760 17134
rect 19708 17070 19760 17076
rect 19720 16522 19748 17070
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 19708 16516 19760 16522
rect 19708 16458 19760 16464
rect 19616 15428 19668 15434
rect 19616 15370 19668 15376
rect 19524 15156 19576 15162
rect 19524 15098 19576 15104
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19340 14000 19392 14006
rect 19392 13960 19564 13988
rect 19340 13942 19392 13948
rect 19260 12566 19380 12594
rect 19246 12472 19302 12481
rect 19246 12407 19248 12416
rect 19300 12407 19302 12416
rect 19248 12378 19300 12384
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19260 11762 19288 12038
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19352 11642 19380 12566
rect 19260 11614 19380 11642
rect 19154 11520 19210 11529
rect 19154 11455 19210 11464
rect 19260 9382 19288 11614
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19352 11354 19380 11494
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19444 10810 19472 11086
rect 19432 10804 19484 10810
rect 19432 10746 19484 10752
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19444 9110 19472 9318
rect 19064 9104 19116 9110
rect 19064 9046 19116 9052
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 18984 8362 19012 8910
rect 18972 8356 19024 8362
rect 18972 8298 19024 8304
rect 18696 8016 18748 8022
rect 18696 7958 18748 7964
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18142 7848 18198 7857
rect 18142 7783 18198 7792
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18616 7410 18644 7890
rect 18972 7744 19024 7750
rect 18972 7686 19024 7692
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 18064 6322 18092 6598
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 18050 6216 18106 6225
rect 18050 6151 18106 6160
rect 18064 6118 18092 6151
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17788 5098 17816 5510
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 17776 5092 17828 5098
rect 17776 5034 17828 5040
rect 17682 3904 17738 3913
rect 17682 3839 17738 3848
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 17512 480 17540 3334
rect 17788 1737 17816 5034
rect 17972 3534 18000 5102
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 18064 3754 18092 4966
rect 18156 3942 18184 7278
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18510 6352 18566 6361
rect 18510 6287 18566 6296
rect 18524 6254 18552 6287
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18604 5772 18656 5778
rect 18604 5714 18656 5720
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18512 4140 18564 4146
rect 18616 4128 18644 5714
rect 18708 5166 18736 7414
rect 18788 5228 18840 5234
rect 18788 5170 18840 5176
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18800 4486 18828 5170
rect 18878 4584 18934 4593
rect 18878 4519 18934 4528
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18696 4140 18748 4146
rect 18616 4100 18696 4128
rect 18512 4082 18564 4088
rect 18696 4082 18748 4088
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18248 3754 18276 3878
rect 18064 3726 18276 3754
rect 18524 3738 18552 4082
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 18052 3664 18104 3670
rect 18052 3606 18104 3612
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 18064 3369 18092 3606
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 18050 3360 18106 3369
rect 18050 3295 18106 3304
rect 18156 2961 18184 3470
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18708 3097 18736 4082
rect 18800 3534 18828 4422
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 18694 3088 18750 3097
rect 18694 3023 18750 3032
rect 18892 2990 18920 4519
rect 18880 2984 18932 2990
rect 18142 2952 18198 2961
rect 18880 2926 18932 2932
rect 18142 2887 18198 2896
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 17774 1728 17830 1737
rect 17774 1663 17830 1672
rect 17972 480 18000 2790
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 18420 1964 18472 1970
rect 18420 1906 18472 1912
rect 18432 480 18460 1906
rect 18984 480 19012 7686
rect 19338 7440 19394 7449
rect 19338 7375 19394 7384
rect 19248 5296 19300 5302
rect 19248 5238 19300 5244
rect 19064 5092 19116 5098
rect 19064 5034 19116 5040
rect 19076 4729 19104 5034
rect 19062 4720 19118 4729
rect 19062 4655 19118 4664
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 19076 4049 19104 4082
rect 19062 4040 19118 4049
rect 19062 3975 19118 3984
rect 19260 610 19288 5238
rect 19352 3602 19380 7375
rect 19432 5636 19484 5642
rect 19432 5578 19484 5584
rect 19444 5370 19472 5578
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 19430 3496 19486 3505
rect 19430 3431 19486 3440
rect 19248 604 19300 610
rect 19248 546 19300 552
rect 19444 480 19472 3431
rect 19536 2990 19564 13960
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19628 6984 19656 12718
rect 19708 12640 19760 12646
rect 19708 12582 19760 12588
rect 19720 8945 19748 12582
rect 19706 8936 19762 8945
rect 19706 8871 19762 8880
rect 19812 7313 19840 16934
rect 19798 7304 19854 7313
rect 19798 7239 19854 7248
rect 19628 6956 19748 6984
rect 19614 6896 19670 6905
rect 19614 6831 19670 6840
rect 19628 6458 19656 6831
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19614 5128 19670 5137
rect 19614 5063 19670 5072
rect 19628 5030 19656 5063
rect 19616 5024 19668 5030
rect 19616 4966 19668 4972
rect 19720 3670 19748 6956
rect 19904 6254 19932 17682
rect 19996 17105 20024 20334
rect 20364 19174 20392 22520
rect 20824 20058 20852 22520
rect 21284 20602 21312 22520
rect 21272 20596 21324 20602
rect 21272 20538 21324 20544
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20352 19168 20404 19174
rect 20352 19110 20404 19116
rect 21744 18426 21772 22520
rect 22204 18970 22232 22520
rect 22192 18964 22244 18970
rect 22192 18906 22244 18912
rect 21732 18420 21784 18426
rect 21732 18362 21784 18368
rect 22664 18086 22692 22520
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 22652 18080 22704 18086
rect 22652 18022 22704 18028
rect 20272 17814 20300 18022
rect 20260 17808 20312 17814
rect 20260 17750 20312 17756
rect 19982 17096 20038 17105
rect 19982 17031 20038 17040
rect 19996 13530 20024 17031
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 20088 16794 20116 16934
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 20272 16046 20300 17750
rect 20812 17604 20864 17610
rect 20812 17546 20864 17552
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 20076 15428 20128 15434
rect 20076 15370 20128 15376
rect 20088 14958 20116 15370
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 20272 14482 20300 15982
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20824 14074 20852 17546
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 20180 11762 20208 13262
rect 20168 11756 20220 11762
rect 20168 11698 20220 11704
rect 20180 10674 20208 11698
rect 20168 10668 20220 10674
rect 20168 10610 20220 10616
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19996 7342 20024 10406
rect 20260 8356 20312 8362
rect 20260 8298 20312 8304
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 19892 6248 19944 6254
rect 19892 6190 19944 6196
rect 20076 6112 20128 6118
rect 20076 6054 20128 6060
rect 20088 5681 20116 6054
rect 20272 5846 20300 8298
rect 20260 5840 20312 5846
rect 20260 5782 20312 5788
rect 20074 5672 20130 5681
rect 20074 5607 20130 5616
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19708 3664 19760 3670
rect 19708 3606 19760 3612
rect 19524 2984 19576 2990
rect 19524 2926 19576 2932
rect 19996 2922 20024 4966
rect 20076 4820 20128 4826
rect 20076 4762 20128 4768
rect 20088 4146 20116 4762
rect 21272 4480 21324 4486
rect 21272 4422 21324 4428
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 20352 3392 20404 3398
rect 20352 3334 20404 3340
rect 19984 2916 20036 2922
rect 19984 2858 20036 2864
rect 20168 2848 20220 2854
rect 20168 2790 20220 2796
rect 20180 2650 20208 2790
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 19892 2304 19944 2310
rect 19892 2246 19944 2252
rect 19904 480 19932 2246
rect 19996 1902 20024 2450
rect 19984 1896 20036 1902
rect 19984 1838 20036 1844
rect 20364 480 20392 3334
rect 20812 604 20864 610
rect 20812 546 20864 552
rect 20824 480 20852 546
rect 21284 480 21312 4422
rect 22652 2916 22704 2922
rect 22652 2858 22704 2864
rect 22192 2848 22244 2854
rect 21730 2816 21786 2825
rect 22192 2790 22244 2796
rect 21730 2751 21786 2760
rect 21744 480 21772 2751
rect 22204 480 22232 2790
rect 22664 480 22692 2858
rect 202 0 258 480
rect 662 0 718 480
rect 1122 0 1178 480
rect 1582 0 1638 480
rect 2042 0 2098 480
rect 2502 0 2558 480
rect 2962 0 3018 480
rect 3422 0 3478 480
rect 3882 0 3938 480
rect 4342 0 4398 480
rect 4894 0 4950 480
rect 5354 0 5410 480
rect 5814 0 5870 480
rect 6274 0 6330 480
rect 6734 0 6790 480
rect 7194 0 7250 480
rect 7654 0 7710 480
rect 8114 0 8170 480
rect 8574 0 8630 480
rect 9034 0 9090 480
rect 9586 0 9642 480
rect 10046 0 10102 480
rect 10506 0 10562 480
rect 10966 0 11022 480
rect 11426 0 11482 480
rect 11886 0 11942 480
rect 12346 0 12402 480
rect 12806 0 12862 480
rect 13266 0 13322 480
rect 13726 0 13782 480
rect 14278 0 14334 480
rect 14738 0 14794 480
rect 15198 0 15254 480
rect 15658 0 15714 480
rect 16118 0 16174 480
rect 16578 0 16634 480
rect 17038 0 17094 480
rect 17498 0 17554 480
rect 17958 0 18014 480
rect 18418 0 18474 480
rect 18970 0 19026 480
rect 19430 0 19486 480
rect 19890 0 19946 480
rect 20350 0 20406 480
rect 20810 0 20866 480
rect 21270 0 21326 480
rect 21730 0 21786 480
rect 22190 0 22246 480
rect 22650 0 22706 480
<< via2 >>
rect 4066 22616 4122 22672
rect 1950 20712 2006 20768
rect 1582 19080 1638 19136
rect 1490 17992 1546 18048
rect 1398 5616 1454 5672
rect 1030 2488 1086 2544
rect 1766 9832 1822 9888
rect 2870 22072 2926 22128
rect 2778 21664 2834 21720
rect 2134 12416 2190 12472
rect 1858 9424 1914 9480
rect 1858 9036 1914 9072
rect 1858 9016 1860 9036
rect 1860 9016 1912 9036
rect 1912 9016 1914 9036
rect 2134 8608 2190 8664
rect 1858 7792 1914 7848
rect 2042 7792 2098 7848
rect 1766 7384 1822 7440
rect 2134 7112 2190 7168
rect 1858 6432 1914 6488
rect 1674 4664 1730 4720
rect 2134 4528 2190 4584
rect 1582 3032 1638 3088
rect 2502 17992 2558 18048
rect 2410 17620 2412 17640
rect 2412 17620 2464 17640
rect 2464 17620 2466 17640
rect 2410 17584 2466 17620
rect 2502 14764 2504 14784
rect 2504 14764 2556 14784
rect 2556 14764 2558 14784
rect 2502 14728 2558 14764
rect 2318 9968 2374 10024
rect 2318 9444 2374 9480
rect 2318 9424 2320 9444
rect 2320 9424 2372 9444
rect 2372 9424 2374 9444
rect 2318 9152 2374 9208
rect 2318 8472 2374 8528
rect 3054 21120 3110 21176
rect 3146 20168 3202 20224
rect 3330 19216 3386 19272
rect 3238 18944 3294 19000
rect 3054 15544 3110 15600
rect 2962 15408 3018 15464
rect 2870 14456 2926 14512
rect 2778 13504 2834 13560
rect 2778 12280 2834 12336
rect 2594 10240 2650 10296
rect 2686 9968 2742 10024
rect 2594 9152 2650 9208
rect 3238 17040 3294 17096
rect 3514 16088 3570 16144
rect 3422 15816 3478 15872
rect 3146 14184 3202 14240
rect 3146 14068 3202 14104
rect 3146 14048 3148 14068
rect 3148 14048 3200 14068
rect 3200 14048 3202 14068
rect 3238 13776 3294 13832
rect 2594 8336 2650 8392
rect 2318 3440 2374 3496
rect 2226 2932 2228 2952
rect 2228 2932 2280 2952
rect 2280 2932 2282 2952
rect 2226 2896 2282 2932
rect 2134 2352 2190 2408
rect 2870 7520 2926 7576
rect 2502 5072 2558 5128
rect 2962 6704 3018 6760
rect 2502 3068 2504 3088
rect 2504 3068 2556 3088
rect 2556 3068 2558 3088
rect 2502 3032 2558 3068
rect 2870 4120 2926 4176
rect 2778 3460 2834 3496
rect 2778 3440 2780 3460
rect 2780 3440 2832 3460
rect 2832 3440 2834 3460
rect 2502 1400 2558 1456
rect 2410 584 2466 640
rect 3790 19760 3846 19816
rect 3698 17720 3754 17776
rect 4066 19780 4122 19816
rect 4066 19760 4068 19780
rect 4068 19760 4120 19780
rect 4120 19760 4122 19780
rect 4066 18264 4122 18320
rect 4066 17856 4122 17912
rect 4066 17312 4122 17368
rect 4066 16768 4122 16824
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 4250 18672 4306 18728
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 4618 19216 4674 19272
rect 5170 19488 5226 19544
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 3790 16632 3846 16688
rect 3974 15952 4030 16008
rect 3698 15408 3754 15464
rect 3790 15000 3846 15056
rect 3606 14728 3662 14784
rect 3330 7520 3386 7576
rect 3238 6024 3294 6080
rect 3330 5480 3386 5536
rect 3330 4820 3386 4856
rect 3330 4800 3332 4820
rect 3332 4800 3384 4820
rect 3384 4800 3386 4820
rect 3330 3476 3332 3496
rect 3332 3476 3384 3496
rect 3384 3476 3386 3496
rect 3330 3440 3386 3476
rect 3790 13640 3846 13696
rect 3698 9152 3754 9208
rect 3698 8472 3754 8528
rect 3606 6996 3662 7032
rect 3606 6976 3608 6996
rect 3608 6976 3660 6996
rect 3660 6976 3662 6996
rect 3698 6840 3754 6896
rect 3974 14184 4030 14240
rect 3974 10104 4030 10160
rect 3882 9832 3938 9888
rect 3606 5344 3662 5400
rect 3790 4664 3846 4720
rect 3606 1944 3662 2000
rect 3054 1128 3110 1184
rect 3974 7928 4030 7984
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4710 14476 4766 14512
rect 4710 14456 4712 14476
rect 4712 14456 4764 14476
rect 4764 14456 4766 14476
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 4434 12552 4490 12608
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4986 16940 4988 16960
rect 4988 16940 5040 16960
rect 5040 16940 5042 16960
rect 4986 16904 5042 16940
rect 5170 18128 5226 18184
rect 4986 12416 5042 12472
rect 4618 11600 4674 11656
rect 4802 11600 4858 11656
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4158 8900 4214 8936
rect 4158 8880 4160 8900
rect 4160 8880 4212 8900
rect 4212 8880 4214 8900
rect 4158 8744 4214 8800
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4526 9424 4582 9480
rect 4434 9288 4490 9344
rect 4710 9172 4766 9208
rect 4710 9152 4712 9172
rect 4712 9152 4764 9172
rect 4764 9152 4766 9172
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4434 7792 4490 7848
rect 4618 7792 4674 7848
rect 5630 19352 5686 19408
rect 5722 19216 5778 19272
rect 5538 18808 5594 18864
rect 5722 18672 5778 18728
rect 5354 16768 5410 16824
rect 5354 16224 5410 16280
rect 5354 15816 5410 15872
rect 5262 12416 5318 12472
rect 5262 11620 5318 11656
rect 5262 11600 5264 11620
rect 5264 11600 5316 11620
rect 5316 11600 5318 11620
rect 5078 8744 5134 8800
rect 5722 17312 5778 17368
rect 5446 12008 5502 12064
rect 5446 11192 5502 11248
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4066 6432 4122 6488
rect 3974 6296 4030 6352
rect 3974 5888 4030 5944
rect 4250 6568 4306 6624
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4434 6160 4490 6216
rect 4250 5208 4306 5264
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4802 4256 4858 4312
rect 4250 2080 4306 2136
rect 4526 3984 4582 4040
rect 4710 3712 4766 3768
rect 4434 3576 4490 3632
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 4434 2624 4490 2680
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 4986 7520 5042 7576
rect 5078 7384 5134 7440
rect 4986 6568 5042 6624
rect 5262 7248 5318 7304
rect 5354 6432 5410 6488
rect 5354 5344 5410 5400
rect 5262 5208 5318 5264
rect 5078 4392 5134 4448
rect 5354 4820 5410 4856
rect 5354 4800 5356 4820
rect 5356 4800 5408 4820
rect 5408 4800 5410 4820
rect 5262 2216 5318 2272
rect 5630 13640 5686 13696
rect 5538 10104 5594 10160
rect 6090 19352 6146 19408
rect 5906 10920 5962 10976
rect 5814 10104 5870 10160
rect 6366 17176 6422 17232
rect 6734 15136 6790 15192
rect 6090 12280 6146 12336
rect 6090 11500 6092 11520
rect 6092 11500 6144 11520
rect 6144 11500 6146 11520
rect 6090 11464 6146 11500
rect 6182 11056 6238 11112
rect 6366 10376 6422 10432
rect 5814 8608 5870 8664
rect 5814 7792 5870 7848
rect 5538 6976 5594 7032
rect 5722 6296 5778 6352
rect 5814 5652 5816 5672
rect 5816 5652 5868 5672
rect 5868 5652 5870 5672
rect 5814 5616 5870 5652
rect 6182 7792 6238 7848
rect 6458 10240 6514 10296
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 8482 19352 8538 19408
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7470 18400 7526 18456
rect 7010 15544 7066 15600
rect 7378 16360 7434 16416
rect 7286 14728 7342 14784
rect 7010 12008 7066 12064
rect 6918 11056 6974 11112
rect 6550 8628 6606 8664
rect 6550 8608 6552 8628
rect 6552 8608 6604 8628
rect 6604 8608 6606 8628
rect 6090 7384 6146 7440
rect 6458 7112 6514 7168
rect 6366 6996 6422 7032
rect 6366 6976 6368 6996
rect 6368 6976 6420 6996
rect 6420 6976 6422 6996
rect 6826 10240 6882 10296
rect 6734 9288 6790 9344
rect 6642 7792 6698 7848
rect 6274 6452 6330 6488
rect 6274 6432 6276 6452
rect 6276 6432 6328 6452
rect 6328 6432 6330 6452
rect 6458 6452 6514 6488
rect 6458 6432 6460 6452
rect 6460 6432 6512 6452
rect 6512 6432 6514 6452
rect 6366 5888 6422 5944
rect 6366 5228 6422 5264
rect 6366 5208 6368 5228
rect 6368 5208 6420 5228
rect 6420 5208 6422 5228
rect 6642 6024 6698 6080
rect 6826 6432 6882 6488
rect 6734 5616 6790 5672
rect 5630 4664 5686 4720
rect 5630 4392 5686 4448
rect 5814 4428 5816 4448
rect 5816 4428 5868 4448
rect 5868 4428 5870 4448
rect 5814 4392 5870 4428
rect 5998 4256 6054 4312
rect 6182 4392 6238 4448
rect 5998 3576 6054 3632
rect 5814 3476 5816 3496
rect 5816 3476 5868 3496
rect 5868 3476 5870 3496
rect 5814 3440 5870 3476
rect 5538 3168 5594 3224
rect 5538 2760 5594 2816
rect 6090 3304 6146 3360
rect 5998 2352 6054 2408
rect 6458 4936 6514 4992
rect 6458 4392 6514 4448
rect 6366 4256 6422 4312
rect 6274 2760 6330 2816
rect 6182 1944 6238 2000
rect 5814 1672 5870 1728
rect 6366 2352 6422 2408
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 8298 17856 8354 17912
rect 8298 17584 8354 17640
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7378 12280 7434 12336
rect 7102 9832 7158 9888
rect 7286 7112 7342 7168
rect 7930 16224 7986 16280
rect 7654 15952 7710 16008
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 8298 12688 8354 12744
rect 7930 12280 7986 12336
rect 7470 9832 7526 9888
rect 8298 12436 8354 12472
rect 8298 12416 8300 12436
rect 8300 12416 8352 12436
rect 8352 12416 8354 12436
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 7930 9968 7986 10024
rect 8022 9696 8078 9752
rect 7654 9172 7710 9208
rect 7654 9152 7656 9172
rect 7656 9152 7708 9172
rect 7708 9152 7710 9172
rect 7562 8608 7618 8664
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 8298 9968 8354 10024
rect 8666 16496 8722 16552
rect 8666 13912 8722 13968
rect 8666 12280 8722 12336
rect 8850 19488 8906 19544
rect 8942 19216 8998 19272
rect 8850 16768 8906 16824
rect 8850 16632 8906 16688
rect 9126 17040 9182 17096
rect 9586 18028 9588 18048
rect 9588 18028 9640 18048
rect 9640 18028 9642 18048
rect 9586 17992 9642 18028
rect 9586 17876 9642 17912
rect 9586 17856 9588 17876
rect 9588 17856 9640 17876
rect 9640 17856 9642 17876
rect 9402 16904 9458 16960
rect 9402 16632 9458 16688
rect 8850 12688 8906 12744
rect 8850 12416 8906 12472
rect 8758 11872 8814 11928
rect 8666 11736 8722 11792
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7746 7792 7802 7848
rect 8022 7792 8078 7848
rect 7746 7112 7802 7168
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 7378 6296 7434 6352
rect 7286 5888 7342 5944
rect 6642 4392 6698 4448
rect 6734 4256 6790 4312
rect 6642 3984 6698 4040
rect 6734 1672 6790 1728
rect 7746 6024 7802 6080
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 8390 6024 8446 6080
rect 8298 5888 8354 5944
rect 7562 4972 7564 4992
rect 7564 4972 7616 4992
rect 7616 4972 7618 4992
rect 7562 4936 7618 4972
rect 7286 3848 7342 3904
rect 7378 3304 7434 3360
rect 7194 1400 7250 1456
rect 7930 5208 7986 5264
rect 8206 5208 8262 5264
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 7746 4256 7802 4312
rect 8758 10920 8814 10976
rect 8666 7792 8722 7848
rect 9034 11464 9090 11520
rect 8942 10648 8998 10704
rect 8942 9696 8998 9752
rect 8942 9152 8998 9208
rect 8758 5480 8814 5536
rect 8666 5244 8668 5264
rect 8668 5244 8720 5264
rect 8720 5244 8722 5264
rect 8666 5208 8722 5244
rect 8390 4936 8446 4992
rect 8022 3984 8078 4040
rect 8206 3984 8262 4040
rect 8298 3848 8354 3904
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 8022 3576 8078 3632
rect 7654 3440 7710 3496
rect 7470 2760 7526 2816
rect 8390 3576 8446 3632
rect 8298 3440 8354 3496
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 7654 2488 7710 2544
rect 7470 1536 7526 1592
rect 8114 2488 8170 2544
rect 8022 1536 8078 1592
rect 8298 1672 8354 1728
rect 8482 1556 8538 1592
rect 8482 1536 8484 1556
rect 8484 1536 8536 1556
rect 8536 1536 8538 1556
rect 9310 14456 9366 14512
rect 9034 7520 9090 7576
rect 9126 6840 9182 6896
rect 9586 16496 9642 16552
rect 9954 18672 10010 18728
rect 9862 17720 9918 17776
rect 9862 16768 9918 16824
rect 9862 16652 9918 16688
rect 9862 16632 9864 16652
rect 9864 16632 9916 16652
rect 9916 16632 9918 16652
rect 9862 16360 9918 16416
rect 9678 15952 9734 16008
rect 9954 16088 10010 16144
rect 10138 19896 10194 19952
rect 10230 19796 10232 19816
rect 10232 19796 10284 19816
rect 10284 19796 10286 19816
rect 10230 19760 10286 19796
rect 10230 19236 10286 19272
rect 10230 19216 10232 19236
rect 10232 19216 10284 19236
rect 10284 19216 10286 19236
rect 10322 18944 10378 19000
rect 9862 15852 9864 15872
rect 9864 15852 9916 15872
rect 9916 15852 9918 15872
rect 9862 15816 9918 15852
rect 10046 15564 10102 15600
rect 10046 15544 10048 15564
rect 10048 15544 10100 15564
rect 10100 15544 10102 15564
rect 9862 14728 9918 14784
rect 9770 14592 9826 14648
rect 10046 13676 10048 13696
rect 10048 13676 10100 13696
rect 10100 13676 10102 13696
rect 10046 13640 10102 13676
rect 10138 13232 10194 13288
rect 9862 13096 9918 13152
rect 9862 12688 9918 12744
rect 9310 6840 9366 6896
rect 9126 5344 9182 5400
rect 8666 1944 8722 2000
rect 9126 4256 9182 4312
rect 9034 2624 9090 2680
rect 9494 9424 9550 9480
rect 9494 7112 9550 7168
rect 9402 5344 9458 5400
rect 9494 4800 9550 4856
rect 9402 3984 9458 4040
rect 9402 3712 9458 3768
rect 9218 2624 9274 2680
rect 10046 12416 10102 12472
rect 9954 11464 10010 11520
rect 9954 10512 10010 10568
rect 9862 10240 9918 10296
rect 9862 9832 9918 9888
rect 9770 9172 9826 9208
rect 9770 9152 9772 9172
rect 9772 9152 9824 9172
rect 9824 9152 9826 9172
rect 9862 8608 9918 8664
rect 9770 7520 9826 7576
rect 9862 6976 9918 7032
rect 9678 3984 9734 4040
rect 9494 3168 9550 3224
rect 9402 2216 9458 2272
rect 9034 1944 9090 2000
rect 9218 1944 9274 2000
rect 8666 1536 8722 1592
rect 10046 6024 10102 6080
rect 9954 5480 10010 5536
rect 10322 9424 10378 9480
rect 10598 16532 10600 16552
rect 10600 16532 10652 16552
rect 10652 16532 10654 16552
rect 10598 16496 10654 16532
rect 10782 17040 10838 17096
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11242 19796 11244 19816
rect 11244 19796 11296 19816
rect 11296 19796 11298 19816
rect 11242 19760 11298 19796
rect 10966 16496 11022 16552
rect 10966 15816 11022 15872
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11610 17740 11666 17776
rect 11610 17720 11612 17740
rect 11612 17720 11664 17740
rect 11664 17720 11666 17740
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11702 17176 11758 17232
rect 11978 19760 12034 19816
rect 12254 19372 12310 19408
rect 12254 19352 12256 19372
rect 12256 19352 12308 19372
rect 12308 19352 12310 19372
rect 12254 18808 12310 18864
rect 11886 17312 11942 17368
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11610 15408 11666 15464
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11426 14864 11482 14920
rect 11334 14492 11336 14512
rect 11336 14492 11388 14512
rect 11388 14492 11390 14512
rect 11334 14456 11390 14492
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11150 12824 11206 12880
rect 10966 12552 11022 12608
rect 10506 9832 10562 9888
rect 10690 9696 10746 9752
rect 10598 7520 10654 7576
rect 10598 6432 10654 6488
rect 10506 6024 10562 6080
rect 10506 5480 10562 5536
rect 10690 6024 10746 6080
rect 9770 3304 9826 3360
rect 9586 2760 9642 2816
rect 9862 2760 9918 2816
rect 10046 3304 10102 3360
rect 10598 4256 10654 4312
rect 10782 4256 10838 4312
rect 10506 3576 10562 3632
rect 10506 3168 10562 3224
rect 10046 2216 10102 2272
rect 10414 2760 10470 2816
rect 10598 2760 10654 2816
rect 10966 9968 11022 10024
rect 11150 9968 11206 10024
rect 11058 8608 11114 8664
rect 10966 7520 11022 7576
rect 10966 7384 11022 7440
rect 10966 5480 11022 5536
rect 11058 5344 11114 5400
rect 10874 3712 10930 3768
rect 10782 2488 10838 2544
rect 10690 2080 10746 2136
rect 11058 4392 11114 4448
rect 11150 4256 11206 4312
rect 11150 3304 11206 3360
rect 11058 2760 11114 2816
rect 11058 2644 11114 2680
rect 11058 2624 11060 2644
rect 11060 2624 11112 2644
rect 11112 2624 11114 2644
rect 11794 13776 11850 13832
rect 11794 13524 11850 13560
rect 11794 13504 11796 13524
rect 11796 13504 11848 13524
rect 11848 13504 11850 13524
rect 11886 13232 11942 13288
rect 12438 19352 12494 19408
rect 11978 12416 12034 12472
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11794 11872 11850 11928
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11610 10648 11666 10704
rect 11518 10512 11574 10568
rect 11518 9988 11574 10024
rect 11518 9968 11520 9988
rect 11520 9968 11572 9988
rect 11572 9968 11574 9988
rect 11702 9968 11758 10024
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11426 7928 11482 7984
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11702 6976 11758 7032
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11426 6024 11482 6080
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11518 3712 11574 3768
rect 11334 3576 11390 3632
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11978 3596 12034 3632
rect 11978 3576 11980 3596
rect 11980 3576 12032 3596
rect 12032 3576 12034 3596
rect 12346 18400 12402 18456
rect 12806 19796 12808 19816
rect 12808 19796 12860 19816
rect 12860 19796 12862 19816
rect 12806 19760 12862 19796
rect 13082 19352 13138 19408
rect 12162 16632 12218 16688
rect 12346 17584 12402 17640
rect 12530 17720 12586 17776
rect 12714 18128 12770 18184
rect 12714 17312 12770 17368
rect 12530 14456 12586 14512
rect 12346 13388 12402 13424
rect 12346 13368 12348 13388
rect 12348 13368 12400 13388
rect 12400 13368 12402 13388
rect 12898 18572 12900 18592
rect 12900 18572 12952 18592
rect 12952 18572 12954 18592
rect 12898 18536 12954 18572
rect 12438 13096 12494 13152
rect 12530 10648 12586 10704
rect 12162 6432 12218 6488
rect 12162 4256 12218 4312
rect 12346 10124 12402 10160
rect 12346 10104 12348 10124
rect 12348 10104 12400 10124
rect 12400 10104 12402 10124
rect 12346 9716 12402 9752
rect 12346 9696 12348 9716
rect 12348 9696 12400 9716
rect 12400 9696 12402 9716
rect 12622 9288 12678 9344
rect 12530 8608 12586 8664
rect 12346 6024 12402 6080
rect 12438 4800 12494 4856
rect 12346 4392 12402 4448
rect 12254 3732 12310 3768
rect 12254 3712 12256 3732
rect 12256 3712 12308 3732
rect 12308 3712 12310 3732
rect 12162 3340 12164 3360
rect 12164 3340 12216 3360
rect 12216 3340 12218 3360
rect 12162 3304 12218 3340
rect 12346 3188 12402 3224
rect 12346 3168 12348 3188
rect 12348 3168 12400 3188
rect 12400 3168 12402 3188
rect 11518 2624 11574 2680
rect 12070 2760 12126 2816
rect 11886 2488 11942 2544
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12622 4392 12678 4448
rect 13358 17176 13414 17232
rect 13358 16768 13414 16824
rect 13174 16632 13230 16688
rect 13174 15020 13230 15056
rect 13174 15000 13176 15020
rect 13176 15000 13228 15020
rect 13228 15000 13230 15020
rect 12806 11328 12862 11384
rect 13174 14728 13230 14784
rect 13174 13640 13230 13696
rect 12990 11464 13046 11520
rect 13266 12824 13322 12880
rect 13542 18944 13598 19000
rect 13542 13640 13598 13696
rect 13542 13504 13598 13560
rect 13082 11056 13138 11112
rect 13174 10376 13230 10432
rect 13082 10240 13138 10296
rect 12990 7928 13046 7984
rect 12898 7112 12954 7168
rect 12806 5480 12862 5536
rect 12806 4528 12862 4584
rect 12806 3848 12862 3904
rect 12530 3712 12586 3768
rect 12254 2352 12310 2408
rect 12346 1400 12402 1456
rect 13450 12008 13506 12064
rect 13542 9832 13598 9888
rect 14002 19896 14058 19952
rect 14002 17720 14058 17776
rect 14002 17620 14004 17640
rect 14004 17620 14056 17640
rect 14056 17620 14058 17640
rect 14002 17584 14058 17620
rect 13910 16632 13966 16688
rect 13910 15852 13912 15872
rect 13912 15852 13964 15872
rect 13964 15852 13966 15872
rect 13910 15816 13966 15852
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 15382 19760 15438 19816
rect 14278 19216 14334 19272
rect 13818 14864 13874 14920
rect 14094 13948 14096 13968
rect 14096 13948 14148 13968
rect 14148 13948 14150 13968
rect 14094 13912 14150 13948
rect 13818 11872 13874 11928
rect 14186 12280 14242 12336
rect 14186 12144 14242 12200
rect 14094 10512 14150 10568
rect 13726 9968 13782 10024
rect 13542 8472 13598 8528
rect 13634 7656 13690 7712
rect 14278 11872 14334 11928
rect 14462 13132 14464 13152
rect 14464 13132 14516 13152
rect 14516 13132 14518 13152
rect 14462 13096 14518 13132
rect 14370 10784 14426 10840
rect 13634 5752 13690 5808
rect 13542 4936 13598 4992
rect 14094 9172 14150 9208
rect 14094 9152 14096 9172
rect 14096 9152 14148 9172
rect 14148 9152 14150 9172
rect 13910 4004 13966 4040
rect 13910 3984 13912 4004
rect 13912 3984 13964 4004
rect 13964 3984 13966 4004
rect 14462 9172 14518 9208
rect 14462 9152 14464 9172
rect 14464 9152 14516 9172
rect 14516 9152 14518 9172
rect 14370 8744 14426 8800
rect 14278 8472 14334 8528
rect 14462 7520 14518 7576
rect 14554 6976 14610 7032
rect 14554 6704 14610 6760
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 15198 18944 15254 19000
rect 15198 18672 15254 18728
rect 14738 18284 14794 18320
rect 14738 18264 14740 18284
rect 14740 18264 14792 18284
rect 14792 18264 14794 18284
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 14922 17584 14978 17640
rect 14922 17312 14978 17368
rect 15106 17312 15162 17368
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14738 14900 14740 14920
rect 14740 14900 14792 14920
rect 14792 14900 14794 14920
rect 14738 14864 14794 14900
rect 15106 15136 15162 15192
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 15474 18128 15530 18184
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 14738 12824 14794 12880
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 15198 10920 15254 10976
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 14738 9424 14794 9480
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 14370 4256 14426 4312
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 14278 2624 14334 2680
rect 14186 1944 14242 2000
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 15750 18128 15806 18184
rect 16026 18672 16082 18728
rect 16118 17856 16174 17912
rect 16026 17176 16082 17232
rect 15934 14320 15990 14376
rect 16394 18944 16450 19000
rect 16854 18536 16910 18592
rect 16670 17312 16726 17368
rect 15566 10260 15622 10296
rect 15566 10240 15568 10260
rect 15568 10240 15620 10260
rect 15620 10240 15622 10260
rect 15566 10104 15622 10160
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 16118 9968 16174 10024
rect 15750 9560 15806 9616
rect 15382 5480 15438 5536
rect 15566 5344 15622 5400
rect 15842 7928 15898 7984
rect 15750 6432 15806 6488
rect 15750 5480 15806 5536
rect 16026 8472 16082 8528
rect 15934 5480 15990 5536
rect 15566 4664 15622 4720
rect 15842 4664 15898 4720
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 16486 13912 16542 13968
rect 17222 18828 17278 18864
rect 17222 18808 17224 18828
rect 17224 18808 17276 18828
rect 17276 18808 17278 18828
rect 17314 18400 17370 18456
rect 16946 14048 17002 14104
rect 17038 13368 17094 13424
rect 16762 9832 16818 9888
rect 16670 7520 16726 7576
rect 16578 5616 16634 5672
rect 15474 1808 15530 1864
rect 16946 8608 17002 8664
rect 17314 13368 17370 13424
rect 17130 8336 17186 8392
rect 16762 4392 16818 4448
rect 17590 19352 17646 19408
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 18786 19080 18842 19136
rect 17958 17720 18014 17776
rect 17682 11736 17738 11792
rect 17498 11192 17554 11248
rect 17406 10648 17462 10704
rect 17682 10512 17738 10568
rect 17590 9696 17646 9752
rect 17406 5752 17462 5808
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18234 17856 18290 17912
rect 18510 17584 18566 17640
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 18142 15444 18144 15464
rect 18144 15444 18196 15464
rect 18196 15444 18198 15464
rect 18142 15408 18198 15444
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18050 9016 18106 9072
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 18970 19216 19026 19272
rect 18878 15544 18934 15600
rect 19062 16940 19064 16960
rect 19064 16940 19116 16960
rect 19116 16940 19118 16960
rect 19062 16904 19118 16940
rect 18878 12688 18934 12744
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 19154 14456 19210 14512
rect 19246 12436 19302 12472
rect 19246 12416 19248 12436
rect 19248 12416 19300 12436
rect 19300 12416 19302 12436
rect 19154 11464 19210 11520
rect 18142 7792 18198 7848
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18050 6160 18106 6216
rect 17682 3848 17738 3904
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18510 6296 18566 6352
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 18878 4528 18934 4584
rect 18050 3304 18106 3360
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 18694 3032 18750 3088
rect 18142 2896 18198 2952
rect 17774 1672 17830 1728
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 19338 7384 19394 7440
rect 19062 4664 19118 4720
rect 19062 3984 19118 4040
rect 19430 3440 19486 3496
rect 19706 8880 19762 8936
rect 19798 7248 19854 7304
rect 19614 6840 19670 6896
rect 19614 5072 19670 5128
rect 19982 17040 20038 17096
rect 20074 5616 20130 5672
rect 21730 2760 21786 2816
<< metal3 >>
rect 0 22674 480 22704
rect 4061 22674 4127 22677
rect 0 22672 4127 22674
rect 0 22616 4066 22672
rect 4122 22616 4127 22672
rect 0 22614 4127 22616
rect 0 22584 480 22614
rect 4061 22611 4127 22614
rect 0 22130 480 22160
rect 2865 22130 2931 22133
rect 0 22128 2931 22130
rect 0 22072 2870 22128
rect 2926 22072 2931 22128
rect 0 22070 2931 22072
rect 0 22040 480 22070
rect 2865 22067 2931 22070
rect 0 21722 480 21752
rect 2773 21722 2839 21725
rect 0 21720 2839 21722
rect 0 21664 2778 21720
rect 2834 21664 2839 21720
rect 0 21662 2839 21664
rect 0 21632 480 21662
rect 2773 21659 2839 21662
rect 0 21178 480 21208
rect 3049 21178 3115 21181
rect 0 21176 3115 21178
rect 0 21120 3054 21176
rect 3110 21120 3115 21176
rect 0 21118 3115 21120
rect 0 21088 480 21118
rect 3049 21115 3115 21118
rect 0 20770 480 20800
rect 1945 20770 2011 20773
rect 0 20768 2011 20770
rect 0 20712 1950 20768
rect 2006 20712 2011 20768
rect 0 20710 2011 20712
rect 0 20680 480 20710
rect 1945 20707 2011 20710
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 20639 18590 20640
rect 0 20226 480 20256
rect 3141 20226 3207 20229
rect 0 20224 3207 20226
rect 0 20168 3146 20224
rect 3202 20168 3207 20224
rect 0 20166 3207 20168
rect 0 20136 480 20166
rect 3141 20163 3207 20166
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 10133 19954 10199 19957
rect 13997 19954 14063 19957
rect 10133 19952 14063 19954
rect 10133 19896 10138 19952
rect 10194 19896 14002 19952
rect 14058 19896 14063 19952
rect 10133 19894 14063 19896
rect 10133 19891 10199 19894
rect 13997 19891 14063 19894
rect 0 19818 480 19848
rect 3785 19818 3851 19821
rect 0 19816 3851 19818
rect 0 19760 3790 19816
rect 3846 19760 3851 19816
rect 0 19758 3851 19760
rect 0 19728 480 19758
rect 3785 19755 3851 19758
rect 4061 19818 4127 19821
rect 9806 19818 9812 19820
rect 4061 19816 9812 19818
rect 4061 19760 4066 19816
rect 4122 19760 9812 19816
rect 4061 19758 9812 19760
rect 4061 19755 4127 19758
rect 9806 19756 9812 19758
rect 9876 19756 9882 19820
rect 10225 19818 10291 19821
rect 11237 19818 11303 19821
rect 10225 19816 11303 19818
rect 10225 19760 10230 19816
rect 10286 19760 11242 19816
rect 11298 19760 11303 19816
rect 10225 19758 11303 19760
rect 10225 19755 10291 19758
rect 11237 19755 11303 19758
rect 11973 19818 12039 19821
rect 12801 19818 12867 19821
rect 15377 19818 15443 19821
rect 11973 19816 15443 19818
rect 11973 19760 11978 19816
rect 12034 19760 12806 19816
rect 12862 19760 15382 19816
rect 15438 19760 15443 19816
rect 11973 19758 15443 19760
rect 11973 19755 12039 19758
rect 12801 19755 12867 19758
rect 15377 19755 15443 19758
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 5165 19546 5231 19549
rect 8845 19546 8911 19549
rect 5165 19544 8911 19546
rect 5165 19488 5170 19544
rect 5226 19488 8850 19544
rect 8906 19488 8911 19544
rect 5165 19486 8911 19488
rect 5165 19483 5231 19486
rect 8845 19483 8911 19486
rect 5625 19410 5691 19413
rect 6085 19410 6151 19413
rect 5625 19408 6151 19410
rect 5625 19352 5630 19408
rect 5686 19352 6090 19408
rect 6146 19352 6151 19408
rect 5625 19350 6151 19352
rect 5625 19347 5691 19350
rect 6085 19347 6151 19350
rect 8477 19412 8543 19413
rect 8477 19408 8524 19412
rect 8588 19410 8594 19412
rect 12249 19410 12315 19413
rect 12433 19410 12499 19413
rect 8477 19352 8482 19408
rect 8477 19348 8524 19352
rect 8588 19350 8634 19410
rect 12249 19408 12499 19410
rect 12249 19352 12254 19408
rect 12310 19352 12438 19408
rect 12494 19352 12499 19408
rect 12249 19350 12499 19352
rect 8588 19348 8594 19350
rect 8477 19347 8543 19348
rect 12249 19347 12315 19350
rect 12433 19347 12499 19350
rect 13077 19410 13143 19413
rect 17585 19410 17651 19413
rect 13077 19408 17651 19410
rect 13077 19352 13082 19408
rect 13138 19352 17590 19408
rect 17646 19352 17651 19408
rect 13077 19350 17651 19352
rect 13077 19347 13143 19350
rect 17585 19347 17651 19350
rect 0 19274 480 19304
rect 3325 19274 3391 19277
rect 0 19272 3391 19274
rect 0 19216 3330 19272
rect 3386 19216 3391 19272
rect 0 19214 3391 19216
rect 0 19184 480 19214
rect 3325 19211 3391 19214
rect 4613 19274 4679 19277
rect 5022 19274 5028 19276
rect 4613 19272 5028 19274
rect 4613 19216 4618 19272
rect 4674 19216 5028 19272
rect 4613 19214 5028 19216
rect 4613 19211 4679 19214
rect 5022 19212 5028 19214
rect 5092 19212 5098 19276
rect 5574 19212 5580 19276
rect 5644 19274 5650 19276
rect 5717 19274 5783 19277
rect 8937 19274 9003 19277
rect 5644 19272 5783 19274
rect 5644 19216 5722 19272
rect 5778 19216 5783 19272
rect 5644 19214 5783 19216
rect 5644 19212 5650 19214
rect 5717 19211 5783 19214
rect 5904 19272 9003 19274
rect 5904 19216 8942 19272
rect 8998 19216 9003 19272
rect 5904 19214 9003 19216
rect 1577 19138 1643 19141
rect 5904 19138 5964 19214
rect 8937 19211 9003 19214
rect 10225 19274 10291 19277
rect 14273 19274 14339 19277
rect 18965 19274 19031 19277
rect 10225 19272 14339 19274
rect 10225 19216 10230 19272
rect 10286 19216 14278 19272
rect 14334 19216 14339 19272
rect 10225 19214 14339 19216
rect 10225 19211 10291 19214
rect 14273 19211 14339 19214
rect 14414 19272 19031 19274
rect 14414 19216 18970 19272
rect 19026 19216 19031 19272
rect 14414 19214 19031 19216
rect 1577 19136 5964 19138
rect 1577 19080 1582 19136
rect 1638 19080 5964 19136
rect 1577 19078 5964 19080
rect 1577 19075 1643 19078
rect 12014 19076 12020 19140
rect 12084 19138 12090 19140
rect 14414 19138 14474 19214
rect 18965 19211 19031 19214
rect 12084 19078 14474 19138
rect 18781 19138 18847 19141
rect 22520 19138 23000 19168
rect 18781 19136 23000 19138
rect 18781 19080 18786 19136
rect 18842 19080 23000 19136
rect 18781 19078 23000 19080
rect 12084 19076 12090 19078
rect 18781 19075 18847 19078
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 22520 19048 23000 19078
rect 14805 19007 15125 19008
rect 3233 19002 3299 19005
rect 10317 19002 10383 19005
rect 13537 19002 13603 19005
rect 3233 19000 5780 19002
rect 3233 18944 3238 19000
rect 3294 18944 5780 19000
rect 3233 18942 5780 18944
rect 3233 18939 3299 18942
rect 0 18866 480 18896
rect 5533 18866 5599 18869
rect 0 18864 5599 18866
rect 0 18808 5538 18864
rect 5594 18808 5599 18864
rect 0 18806 5599 18808
rect 5720 18866 5780 18942
rect 10317 19000 13603 19002
rect 10317 18944 10322 19000
rect 10378 18944 13542 19000
rect 13598 18944 13603 19000
rect 10317 18942 13603 18944
rect 10317 18939 10383 18942
rect 13537 18939 13603 18942
rect 15193 19002 15259 19005
rect 16389 19002 16455 19005
rect 15193 19000 16455 19002
rect 15193 18944 15198 19000
rect 15254 18944 16394 19000
rect 16450 18944 16455 19000
rect 15193 18942 16455 18944
rect 15193 18939 15259 18942
rect 16389 18939 16455 18942
rect 12249 18868 12315 18869
rect 12198 18866 12204 18868
rect 5720 18806 12204 18866
rect 12268 18864 12315 18868
rect 13486 18866 13492 18868
rect 12310 18808 12315 18864
rect 0 18776 480 18806
rect 5533 18803 5599 18806
rect 12198 18804 12204 18806
rect 12268 18804 12315 18808
rect 12249 18803 12315 18804
rect 12528 18806 13492 18866
rect 4245 18730 4311 18733
rect 5717 18730 5783 18733
rect 4245 18728 5783 18730
rect 4245 18672 4250 18728
rect 4306 18672 5722 18728
rect 5778 18672 5783 18728
rect 4245 18670 5783 18672
rect 4245 18667 4311 18670
rect 5717 18667 5783 18670
rect 9949 18730 10015 18733
rect 12528 18730 12588 18806
rect 13486 18804 13492 18806
rect 13556 18866 13562 18868
rect 17217 18866 17283 18869
rect 13556 18864 17283 18866
rect 13556 18808 17222 18864
rect 17278 18808 17283 18864
rect 13556 18806 17283 18808
rect 13556 18804 13562 18806
rect 17217 18803 17283 18806
rect 9949 18728 12588 18730
rect 9949 18672 9954 18728
rect 10010 18672 12588 18728
rect 9949 18670 12588 18672
rect 15193 18730 15259 18733
rect 16021 18730 16087 18733
rect 15193 18728 16087 18730
rect 15193 18672 15198 18728
rect 15254 18672 16026 18728
rect 16082 18672 16087 18728
rect 15193 18670 16087 18672
rect 9949 18667 10015 18670
rect 15193 18667 15259 18670
rect 16021 18667 16087 18670
rect 12893 18594 12959 18597
rect 16849 18594 16915 18597
rect 12893 18592 16915 18594
rect 12893 18536 12898 18592
rect 12954 18536 16854 18592
rect 16910 18536 16915 18592
rect 12893 18534 16915 18536
rect 12893 18531 12959 18534
rect 16849 18531 16915 18534
rect 4409 18528 4729 18529
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 7046 18396 7052 18460
rect 7116 18458 7122 18460
rect 7465 18458 7531 18461
rect 7116 18456 7531 18458
rect 7116 18400 7470 18456
rect 7526 18400 7531 18456
rect 7116 18398 7531 18400
rect 7116 18396 7122 18398
rect 7465 18395 7531 18398
rect 12341 18458 12407 18461
rect 17309 18458 17375 18461
rect 12341 18456 17375 18458
rect 12341 18400 12346 18456
rect 12402 18400 17314 18456
rect 17370 18400 17375 18456
rect 12341 18398 17375 18400
rect 12341 18395 12407 18398
rect 17309 18395 17375 18398
rect 0 18322 480 18352
rect 4061 18322 4127 18325
rect 0 18320 4127 18322
rect 0 18264 4066 18320
rect 4122 18264 4127 18320
rect 0 18262 4127 18264
rect 0 18232 480 18262
rect 4061 18259 4127 18262
rect 6494 18260 6500 18324
rect 6564 18322 6570 18324
rect 14733 18322 14799 18325
rect 6564 18320 14799 18322
rect 6564 18264 14738 18320
rect 14794 18264 14799 18320
rect 6564 18262 14799 18264
rect 6564 18260 6570 18262
rect 14733 18259 14799 18262
rect 4102 18124 4108 18188
rect 4172 18186 4178 18188
rect 5165 18186 5231 18189
rect 4172 18184 5231 18186
rect 4172 18128 5170 18184
rect 5226 18128 5231 18184
rect 4172 18126 5231 18128
rect 4172 18124 4178 18126
rect 5165 18123 5231 18126
rect 5574 18124 5580 18188
rect 5644 18186 5650 18188
rect 12709 18186 12775 18189
rect 15469 18186 15535 18189
rect 15745 18186 15811 18189
rect 5644 18126 9506 18186
rect 5644 18124 5650 18126
rect 1485 18052 1551 18053
rect 1485 18048 1532 18052
rect 1596 18050 1602 18052
rect 2497 18050 2563 18053
rect 5022 18050 5028 18052
rect 1485 17992 1490 18048
rect 1485 17988 1532 17992
rect 1596 17990 1642 18050
rect 2497 18048 5028 18050
rect 2497 17992 2502 18048
rect 2558 17992 5028 18048
rect 2497 17990 5028 17992
rect 1596 17988 1602 17990
rect 1485 17987 1551 17988
rect 2497 17987 2563 17990
rect 5022 17988 5028 17990
rect 5092 17988 5098 18052
rect 9446 18050 9506 18126
rect 12709 18184 15811 18186
rect 12709 18128 12714 18184
rect 12770 18128 15474 18184
rect 15530 18128 15750 18184
rect 15806 18128 15811 18184
rect 12709 18126 15811 18128
rect 12709 18123 12775 18126
rect 15469 18123 15535 18126
rect 15745 18123 15811 18126
rect 9581 18050 9647 18053
rect 9446 18048 9647 18050
rect 9446 17992 9586 18048
rect 9642 17992 9647 18048
rect 9446 17990 9647 17992
rect 9581 17987 9647 17990
rect 7874 17984 8194 17985
rect 0 17914 480 17944
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 17919 15125 17920
rect 4061 17914 4127 17917
rect 0 17912 4127 17914
rect 0 17856 4066 17912
rect 4122 17856 4127 17912
rect 0 17854 4127 17856
rect 0 17824 480 17854
rect 4061 17851 4127 17854
rect 8293 17914 8359 17917
rect 9581 17914 9647 17917
rect 8293 17912 9647 17914
rect 8293 17856 8298 17912
rect 8354 17856 9586 17912
rect 9642 17856 9647 17912
rect 8293 17854 9647 17856
rect 8293 17851 8359 17854
rect 9581 17851 9647 17854
rect 16113 17914 16179 17917
rect 18229 17914 18295 17917
rect 16113 17912 18295 17914
rect 16113 17856 16118 17912
rect 16174 17856 18234 17912
rect 18290 17856 18295 17912
rect 16113 17854 18295 17856
rect 16113 17851 16179 17854
rect 18229 17851 18295 17854
rect 3693 17778 3759 17781
rect 9857 17778 9923 17781
rect 3693 17776 9923 17778
rect 3693 17720 3698 17776
rect 3754 17720 9862 17776
rect 9918 17720 9923 17776
rect 3693 17718 9923 17720
rect 3693 17715 3759 17718
rect 9857 17715 9923 17718
rect 11605 17778 11671 17781
rect 12525 17778 12591 17781
rect 11605 17776 12591 17778
rect 11605 17720 11610 17776
rect 11666 17720 12530 17776
rect 12586 17720 12591 17776
rect 11605 17718 12591 17720
rect 11605 17715 11671 17718
rect 12525 17715 12591 17718
rect 13997 17778 14063 17781
rect 17953 17778 18019 17781
rect 13997 17776 18019 17778
rect 13997 17720 14002 17776
rect 14058 17720 17958 17776
rect 18014 17720 18019 17776
rect 13997 17718 18019 17720
rect 13997 17715 14063 17718
rect 17953 17715 18019 17718
rect 2405 17642 2471 17645
rect 8293 17642 8359 17645
rect 12341 17644 12407 17645
rect 13997 17644 14063 17645
rect 12341 17642 12388 17644
rect 2405 17640 8359 17642
rect 2405 17584 2410 17640
rect 2466 17584 8298 17640
rect 8354 17584 8359 17640
rect 2405 17582 8359 17584
rect 12296 17640 12388 17642
rect 12296 17584 12346 17640
rect 12296 17582 12388 17584
rect 2405 17579 2471 17582
rect 8293 17579 8359 17582
rect 12341 17580 12388 17582
rect 12452 17580 12458 17644
rect 13997 17642 14044 17644
rect 13952 17640 14044 17642
rect 13952 17584 14002 17640
rect 13952 17582 14044 17584
rect 13997 17580 14044 17582
rect 14108 17580 14114 17644
rect 14917 17642 14983 17645
rect 18505 17642 18571 17645
rect 14917 17640 18571 17642
rect 14917 17584 14922 17640
rect 14978 17584 18510 17640
rect 18566 17584 18571 17640
rect 14917 17582 18571 17584
rect 12341 17579 12407 17580
rect 13997 17579 14063 17580
rect 14917 17579 14983 17582
rect 18505 17579 18571 17582
rect 4409 17440 4729 17441
rect 0 17370 480 17400
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 17375 18590 17376
rect 4061 17370 4127 17373
rect 0 17368 4127 17370
rect 0 17312 4066 17368
rect 4122 17312 4127 17368
rect 0 17310 4127 17312
rect 0 17280 480 17310
rect 4061 17307 4127 17310
rect 5717 17370 5783 17373
rect 10174 17370 10180 17372
rect 5717 17368 10180 17370
rect 5717 17312 5722 17368
rect 5778 17312 10180 17368
rect 5717 17310 10180 17312
rect 5717 17307 5783 17310
rect 10174 17308 10180 17310
rect 10244 17308 10250 17372
rect 11881 17370 11947 17373
rect 12709 17370 12775 17373
rect 14917 17370 14983 17373
rect 11881 17368 14983 17370
rect 11881 17312 11886 17368
rect 11942 17312 12714 17368
rect 12770 17312 14922 17368
rect 14978 17312 14983 17368
rect 11881 17310 14983 17312
rect 11881 17307 11947 17310
rect 12709 17307 12775 17310
rect 14917 17307 14983 17310
rect 15101 17370 15167 17373
rect 16665 17370 16731 17373
rect 15101 17368 16731 17370
rect 15101 17312 15106 17368
rect 15162 17312 16670 17368
rect 16726 17312 16731 17368
rect 15101 17310 16731 17312
rect 15101 17307 15167 17310
rect 16665 17307 16731 17310
rect 6361 17234 6427 17237
rect 11697 17234 11763 17237
rect 6361 17232 11763 17234
rect 6361 17176 6366 17232
rect 6422 17176 11702 17232
rect 11758 17176 11763 17232
rect 6361 17174 11763 17176
rect 6361 17171 6427 17174
rect 11697 17171 11763 17174
rect 13353 17234 13419 17237
rect 16021 17234 16087 17237
rect 13353 17232 16087 17234
rect 13353 17176 13358 17232
rect 13414 17176 16026 17232
rect 16082 17176 16087 17232
rect 13353 17174 16087 17176
rect 13353 17171 13419 17174
rect 16021 17171 16087 17174
rect 3233 17098 3299 17101
rect 9121 17098 9187 17101
rect 3233 17096 9187 17098
rect 3233 17040 3238 17096
rect 3294 17040 9126 17096
rect 9182 17040 9187 17096
rect 3233 17038 9187 17040
rect 3233 17035 3299 17038
rect 9121 17035 9187 17038
rect 10777 17098 10843 17101
rect 19977 17098 20043 17101
rect 10777 17096 20043 17098
rect 10777 17040 10782 17096
rect 10838 17040 19982 17096
rect 20038 17040 20043 17096
rect 10777 17038 20043 17040
rect 10777 17035 10843 17038
rect 19977 17035 20043 17038
rect 0 16962 480 16992
rect 4981 16962 5047 16965
rect 9397 16962 9463 16965
rect 0 16960 5047 16962
rect 0 16904 4986 16960
rect 5042 16904 5047 16960
rect 0 16902 5047 16904
rect 0 16872 480 16902
rect 4981 16899 5047 16902
rect 9262 16960 9463 16962
rect 9262 16904 9402 16960
rect 9458 16904 9463 16960
rect 9262 16902 9463 16904
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 4061 16826 4127 16829
rect 5349 16826 5415 16829
rect 4061 16824 5415 16826
rect 4061 16768 4066 16824
rect 4122 16768 5354 16824
rect 5410 16768 5415 16824
rect 4061 16766 5415 16768
rect 4061 16763 4127 16766
rect 5349 16763 5415 16766
rect 8334 16764 8340 16828
rect 8404 16826 8410 16828
rect 8845 16826 8911 16829
rect 8404 16824 8911 16826
rect 8404 16768 8850 16824
rect 8906 16768 8911 16824
rect 8404 16766 8911 16768
rect 8404 16764 8410 16766
rect 8845 16763 8911 16766
rect 3785 16690 3851 16693
rect 8845 16690 8911 16693
rect 3785 16688 8911 16690
rect 3785 16632 3790 16688
rect 3846 16632 8850 16688
rect 8906 16632 8911 16688
rect 3785 16630 8911 16632
rect 9262 16690 9322 16902
rect 9397 16899 9463 16902
rect 19057 16962 19123 16965
rect 19190 16962 19196 16964
rect 19057 16960 19196 16962
rect 19057 16904 19062 16960
rect 19118 16904 19196 16960
rect 19057 16902 19196 16904
rect 19057 16899 19123 16902
rect 19190 16900 19196 16902
rect 19260 16900 19266 16964
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 9857 16826 9923 16829
rect 13353 16826 13419 16829
rect 9857 16824 13419 16826
rect 9857 16768 9862 16824
rect 9918 16768 13358 16824
rect 13414 16768 13419 16824
rect 9857 16766 13419 16768
rect 9857 16763 9923 16766
rect 13353 16763 13419 16766
rect 9397 16690 9463 16693
rect 9262 16688 9463 16690
rect 9262 16632 9402 16688
rect 9458 16632 9463 16688
rect 9262 16630 9463 16632
rect 3785 16627 3851 16630
rect 8845 16627 8911 16630
rect 9397 16627 9463 16630
rect 9857 16690 9923 16693
rect 12157 16690 12223 16693
rect 9857 16688 12223 16690
rect 9857 16632 9862 16688
rect 9918 16632 12162 16688
rect 12218 16632 12223 16688
rect 9857 16630 12223 16632
rect 9857 16627 9923 16630
rect 12157 16627 12223 16630
rect 13169 16690 13235 16693
rect 13905 16690 13971 16693
rect 13169 16688 13971 16690
rect 13169 16632 13174 16688
rect 13230 16632 13910 16688
rect 13966 16632 13971 16688
rect 13169 16630 13971 16632
rect 13169 16627 13235 16630
rect 13905 16627 13971 16630
rect 8661 16554 8727 16557
rect 4248 16552 8727 16554
rect 4248 16496 8666 16552
rect 8722 16496 8727 16552
rect 4248 16494 8727 16496
rect 0 16418 480 16448
rect 4248 16418 4308 16494
rect 8661 16491 8727 16494
rect 8886 16492 8892 16556
rect 8956 16554 8962 16556
rect 9581 16554 9647 16557
rect 8956 16552 9647 16554
rect 8956 16496 9586 16552
rect 9642 16496 9647 16552
rect 8956 16494 9647 16496
rect 8956 16492 8962 16494
rect 9581 16491 9647 16494
rect 10593 16554 10659 16557
rect 10961 16554 11027 16557
rect 12566 16554 12572 16556
rect 10593 16552 12572 16554
rect 10593 16496 10598 16552
rect 10654 16496 10966 16552
rect 11022 16496 12572 16552
rect 10593 16494 12572 16496
rect 10593 16491 10659 16494
rect 10961 16491 11027 16494
rect 12566 16492 12572 16494
rect 12636 16492 12642 16556
rect 0 16358 4308 16418
rect 7373 16418 7439 16421
rect 9857 16418 9923 16421
rect 7373 16416 9923 16418
rect 7373 16360 7378 16416
rect 7434 16360 9862 16416
rect 9918 16360 9923 16416
rect 7373 16358 9923 16360
rect 0 16328 480 16358
rect 7373 16355 7439 16358
rect 9857 16355 9923 16358
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 5349 16282 5415 16285
rect 7925 16282 7991 16285
rect 5349 16280 7991 16282
rect 5349 16224 5354 16280
rect 5410 16224 7930 16280
rect 7986 16224 7991 16280
rect 5349 16222 7991 16224
rect 5349 16219 5415 16222
rect 7925 16219 7991 16222
rect 3509 16146 3575 16149
rect 9949 16146 10015 16149
rect 3509 16144 10015 16146
rect 3509 16088 3514 16144
rect 3570 16088 9954 16144
rect 10010 16088 10015 16144
rect 3509 16086 10015 16088
rect 3509 16083 3575 16086
rect 9949 16083 10015 16086
rect 0 16010 480 16040
rect 3969 16010 4035 16013
rect 7649 16012 7715 16013
rect 7598 16010 7604 16012
rect 0 16008 4035 16010
rect 0 15952 3974 16008
rect 4030 15952 4035 16008
rect 0 15950 4035 15952
rect 7522 15950 7604 16010
rect 7668 16010 7715 16012
rect 9673 16010 9739 16013
rect 7668 16008 9739 16010
rect 7710 15952 9678 16008
rect 9734 15952 9739 16008
rect 0 15920 480 15950
rect 3969 15947 4035 15950
rect 7598 15948 7604 15950
rect 7668 15950 9739 15952
rect 7668 15948 7715 15950
rect 7649 15947 7715 15948
rect 9673 15947 9739 15950
rect 3417 15874 3483 15877
rect 5349 15874 5415 15877
rect 3417 15872 5415 15874
rect 3417 15816 3422 15872
rect 3478 15816 5354 15872
rect 5410 15816 5415 15872
rect 3417 15814 5415 15816
rect 3417 15811 3483 15814
rect 5349 15811 5415 15814
rect 9857 15874 9923 15877
rect 10961 15874 11027 15877
rect 13905 15876 13971 15877
rect 9857 15872 11027 15874
rect 9857 15816 9862 15872
rect 9918 15816 10966 15872
rect 11022 15816 11027 15872
rect 9857 15814 11027 15816
rect 9857 15811 9923 15814
rect 10961 15811 11027 15814
rect 13854 15812 13860 15876
rect 13924 15874 13971 15876
rect 13924 15872 14016 15874
rect 13966 15816 14016 15872
rect 13924 15814 14016 15816
rect 13924 15812 13971 15814
rect 13905 15811 13971 15812
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 3049 15602 3115 15605
rect 7005 15602 7071 15605
rect 10041 15604 10107 15605
rect 9990 15602 9996 15604
rect 3049 15600 7071 15602
rect 3049 15544 3054 15600
rect 3110 15544 7010 15600
rect 7066 15544 7071 15600
rect 3049 15542 7071 15544
rect 9914 15542 9996 15602
rect 10060 15602 10107 15604
rect 15694 15602 15700 15604
rect 10060 15600 15700 15602
rect 10102 15544 15700 15600
rect 3049 15539 3115 15542
rect 7005 15539 7071 15542
rect 9990 15540 9996 15542
rect 10060 15542 15700 15544
rect 10060 15540 10107 15542
rect 15694 15540 15700 15542
rect 15764 15602 15770 15604
rect 18873 15602 18939 15605
rect 15764 15600 18939 15602
rect 15764 15544 18878 15600
rect 18934 15544 18939 15600
rect 15764 15542 18939 15544
rect 15764 15540 15770 15542
rect 10041 15539 10107 15540
rect 18873 15539 18939 15542
rect 0 15466 480 15496
rect 2957 15466 3023 15469
rect 0 15464 3023 15466
rect 0 15408 2962 15464
rect 3018 15408 3023 15464
rect 0 15406 3023 15408
rect 0 15376 480 15406
rect 2957 15403 3023 15406
rect 3693 15466 3759 15469
rect 5758 15466 5764 15468
rect 3693 15464 5764 15466
rect 3693 15408 3698 15464
rect 3754 15408 5764 15464
rect 3693 15406 5764 15408
rect 3693 15403 3759 15406
rect 5758 15404 5764 15406
rect 5828 15404 5834 15468
rect 11605 15466 11671 15469
rect 18137 15466 18203 15469
rect 11605 15464 18203 15466
rect 11605 15408 11610 15464
rect 11666 15408 18142 15464
rect 18198 15408 18203 15464
rect 11605 15406 18203 15408
rect 11605 15403 11671 15406
rect 18137 15403 18203 15406
rect 4409 15264 4729 15265
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 6126 15132 6132 15196
rect 6196 15194 6202 15196
rect 6729 15194 6795 15197
rect 6196 15192 6795 15194
rect 6196 15136 6734 15192
rect 6790 15136 6795 15192
rect 6196 15134 6795 15136
rect 6196 15132 6202 15134
rect 6729 15131 6795 15134
rect 13854 15132 13860 15196
rect 13924 15194 13930 15196
rect 15101 15194 15167 15197
rect 13924 15192 15167 15194
rect 13924 15136 15106 15192
rect 15162 15136 15167 15192
rect 13924 15134 15167 15136
rect 13924 15132 13930 15134
rect 15101 15131 15167 15134
rect 0 15058 480 15088
rect 3785 15058 3851 15061
rect 0 15056 3851 15058
rect 0 15000 3790 15056
rect 3846 15000 3851 15056
rect 0 14998 3851 15000
rect 0 14968 480 14998
rect 3785 14995 3851 14998
rect 13169 15058 13235 15061
rect 19190 15058 19196 15060
rect 13169 15056 19196 15058
rect 13169 15000 13174 15056
rect 13230 15000 19196 15056
rect 13169 14998 19196 15000
rect 13169 14995 13235 14998
rect 19190 14996 19196 14998
rect 19260 14996 19266 15060
rect 11421 14922 11487 14925
rect 13813 14922 13879 14925
rect 14733 14922 14799 14925
rect 11421 14920 14799 14922
rect 11421 14864 11426 14920
rect 11482 14864 13818 14920
rect 13874 14864 14738 14920
rect 14794 14864 14799 14920
rect 11421 14862 14799 14864
rect 11421 14859 11487 14862
rect 13813 14859 13879 14862
rect 14733 14859 14799 14862
rect 2497 14786 2563 14789
rect 2630 14786 2636 14788
rect 2497 14784 2636 14786
rect 2497 14728 2502 14784
rect 2558 14728 2636 14784
rect 2497 14726 2636 14728
rect 2497 14723 2563 14726
rect 2630 14724 2636 14726
rect 2700 14724 2706 14788
rect 3601 14786 3667 14789
rect 7281 14786 7347 14789
rect 3601 14784 7347 14786
rect 3601 14728 3606 14784
rect 3662 14728 7286 14784
rect 7342 14728 7347 14784
rect 3601 14726 7347 14728
rect 3601 14723 3667 14726
rect 7281 14723 7347 14726
rect 9857 14786 9923 14789
rect 13169 14786 13235 14789
rect 9857 14784 13235 14786
rect 9857 14728 9862 14784
rect 9918 14728 13174 14784
rect 13230 14728 13235 14784
rect 9857 14726 13235 14728
rect 9857 14723 9923 14726
rect 13169 14723 13235 14726
rect 7874 14720 8194 14721
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 9765 14650 9831 14653
rect 9765 14648 12772 14650
rect 9765 14592 9770 14648
rect 9826 14592 12772 14648
rect 9765 14590 12772 14592
rect 9765 14587 9831 14590
rect 0 14514 480 14544
rect 2865 14514 2931 14517
rect 0 14512 2931 14514
rect 0 14456 2870 14512
rect 2926 14456 2931 14512
rect 0 14454 2931 14456
rect 0 14424 480 14454
rect 2865 14451 2931 14454
rect 4705 14514 4771 14517
rect 9305 14514 9371 14517
rect 4705 14512 9371 14514
rect 4705 14456 4710 14512
rect 4766 14456 9310 14512
rect 9366 14456 9371 14512
rect 4705 14454 9371 14456
rect 4705 14451 4771 14454
rect 9305 14451 9371 14454
rect 11329 14514 11395 14517
rect 12525 14514 12591 14517
rect 11329 14512 12591 14514
rect 11329 14456 11334 14512
rect 11390 14456 12530 14512
rect 12586 14456 12591 14512
rect 11329 14454 12591 14456
rect 12712 14514 12772 14590
rect 19149 14514 19215 14517
rect 12712 14512 19215 14514
rect 12712 14456 19154 14512
rect 19210 14456 19215 14512
rect 12712 14454 19215 14456
rect 11329 14451 11395 14454
rect 12525 14451 12591 14454
rect 19149 14451 19215 14454
rect 2078 14316 2084 14380
rect 2148 14378 2154 14380
rect 15929 14378 15995 14381
rect 2148 14376 15995 14378
rect 2148 14320 15934 14376
rect 15990 14320 15995 14376
rect 2148 14318 15995 14320
rect 2148 14316 2154 14318
rect 15929 14315 15995 14318
rect 3141 14244 3207 14245
rect 3141 14242 3188 14244
rect 3096 14240 3188 14242
rect 3096 14184 3146 14240
rect 3096 14182 3188 14184
rect 3141 14180 3188 14182
rect 3252 14180 3258 14244
rect 3734 14180 3740 14244
rect 3804 14242 3810 14244
rect 3969 14242 4035 14245
rect 3804 14240 4035 14242
rect 3804 14184 3974 14240
rect 4030 14184 4035 14240
rect 3804 14182 4035 14184
rect 3804 14180 3810 14182
rect 3141 14179 3207 14180
rect 3969 14179 4035 14182
rect 4409 14176 4729 14177
rect 0 14106 480 14136
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 14111 18590 14112
rect 3141 14106 3207 14109
rect 0 14104 3207 14106
rect 0 14048 3146 14104
rect 3202 14048 3207 14104
rect 0 14046 3207 14048
rect 0 14016 480 14046
rect 3141 14043 3207 14046
rect 16941 14106 17007 14109
rect 16941 14104 17234 14106
rect 16941 14048 16946 14104
rect 17002 14048 17234 14104
rect 16941 14046 17234 14048
rect 16941 14043 17007 14046
rect 4838 13908 4844 13972
rect 4908 13970 4914 13972
rect 8661 13970 8727 13973
rect 4908 13968 8727 13970
rect 4908 13912 8666 13968
rect 8722 13912 8727 13968
rect 4908 13910 8727 13912
rect 4908 13908 4914 13910
rect 8661 13907 8727 13910
rect 14089 13970 14155 13973
rect 16481 13970 16547 13973
rect 14089 13968 16547 13970
rect 14089 13912 14094 13968
rect 14150 13912 16486 13968
rect 16542 13912 16547 13968
rect 14089 13910 16547 13912
rect 14089 13907 14155 13910
rect 16481 13907 16547 13910
rect 3233 13834 3299 13837
rect 11789 13834 11855 13837
rect 3233 13832 11855 13834
rect 3233 13776 3238 13832
rect 3294 13776 11794 13832
rect 11850 13776 11855 13832
rect 3233 13774 11855 13776
rect 3233 13771 3299 13774
rect 11789 13771 11855 13774
rect 3785 13698 3851 13701
rect 4102 13698 4108 13700
rect 3785 13696 4108 13698
rect 3785 13640 3790 13696
rect 3846 13640 4108 13696
rect 3785 13638 4108 13640
rect 3785 13635 3851 13638
rect 4102 13636 4108 13638
rect 4172 13636 4178 13700
rect 5390 13636 5396 13700
rect 5460 13698 5466 13700
rect 5625 13698 5691 13701
rect 5460 13696 5691 13698
rect 5460 13640 5630 13696
rect 5686 13640 5691 13696
rect 5460 13638 5691 13640
rect 5460 13636 5466 13638
rect 5625 13635 5691 13638
rect 9622 13636 9628 13700
rect 9692 13698 9698 13700
rect 10041 13698 10107 13701
rect 9692 13696 10107 13698
rect 9692 13640 10046 13696
rect 10102 13640 10107 13696
rect 9692 13638 10107 13640
rect 9692 13636 9698 13638
rect 10041 13635 10107 13638
rect 13169 13698 13235 13701
rect 13537 13698 13603 13701
rect 13169 13696 13603 13698
rect 13169 13640 13174 13696
rect 13230 13640 13542 13696
rect 13598 13640 13603 13696
rect 13169 13638 13603 13640
rect 13169 13635 13235 13638
rect 13537 13635 13603 13638
rect 7874 13632 8194 13633
rect 0 13562 480 13592
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 2773 13562 2839 13565
rect 0 13560 2839 13562
rect 0 13504 2778 13560
rect 2834 13504 2839 13560
rect 0 13502 2839 13504
rect 0 13472 480 13502
rect 2773 13499 2839 13502
rect 11789 13562 11855 13565
rect 13537 13564 13603 13565
rect 11789 13560 12588 13562
rect 11789 13504 11794 13560
rect 11850 13504 12588 13560
rect 11789 13502 12588 13504
rect 11789 13499 11855 13502
rect 6310 13364 6316 13428
rect 6380 13426 6386 13428
rect 12014 13426 12020 13428
rect 6380 13366 12020 13426
rect 6380 13364 6386 13366
rect 12014 13364 12020 13366
rect 12084 13364 12090 13428
rect 12198 13364 12204 13428
rect 12268 13426 12274 13428
rect 12341 13426 12407 13429
rect 12268 13424 12407 13426
rect 12268 13368 12346 13424
rect 12402 13368 12407 13424
rect 12268 13366 12407 13368
rect 12528 13426 12588 13502
rect 13486 13500 13492 13564
rect 13556 13562 13603 13564
rect 13556 13560 13648 13562
rect 13598 13504 13648 13560
rect 13556 13502 13648 13504
rect 13556 13500 13603 13502
rect 13537 13499 13603 13500
rect 17033 13426 17099 13429
rect 12528 13424 17099 13426
rect 12528 13368 17038 13424
rect 17094 13368 17099 13424
rect 12528 13366 17099 13368
rect 17174 13426 17234 14046
rect 17309 13426 17375 13429
rect 17174 13424 17375 13426
rect 17174 13368 17314 13424
rect 17370 13368 17375 13424
rect 17174 13366 17375 13368
rect 12268 13364 12274 13366
rect 12341 13363 12407 13366
rect 17033 13363 17099 13366
rect 17309 13363 17375 13366
rect 4838 13290 4844 13292
rect 4248 13230 4844 13290
rect 0 13154 480 13184
rect 3550 13154 3556 13156
rect 0 13094 3556 13154
rect 0 13064 480 13094
rect 3550 13092 3556 13094
rect 3620 13154 3626 13156
rect 4248 13154 4308 13230
rect 4838 13228 4844 13230
rect 4908 13228 4914 13292
rect 10133 13290 10199 13293
rect 11881 13290 11947 13293
rect 10133 13288 11947 13290
rect 10133 13232 10138 13288
rect 10194 13232 11886 13288
rect 11942 13232 11947 13288
rect 10133 13230 11947 13232
rect 10133 13227 10199 13230
rect 11881 13227 11947 13230
rect 3620 13094 4308 13154
rect 9857 13154 9923 13157
rect 10358 13154 10364 13156
rect 9857 13152 10364 13154
rect 9857 13096 9862 13152
rect 9918 13096 10364 13152
rect 9857 13094 10364 13096
rect 3620 13092 3626 13094
rect 9857 13091 9923 13094
rect 10358 13092 10364 13094
rect 10428 13092 10434 13156
rect 11884 13154 11944 13227
rect 12433 13154 12499 13157
rect 11884 13152 12499 13154
rect 11884 13096 12438 13152
rect 12494 13096 12499 13152
rect 11884 13094 12499 13096
rect 12433 13091 12499 13094
rect 14038 13092 14044 13156
rect 14108 13154 14114 13156
rect 14457 13154 14523 13157
rect 14108 13152 14523 13154
rect 14108 13096 14462 13152
rect 14518 13096 14523 13152
rect 14108 13094 14523 13096
rect 14108 13092 14114 13094
rect 14457 13091 14523 13094
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 11145 12882 11211 12885
rect 13261 12882 13327 12885
rect 11145 12880 13327 12882
rect 11145 12824 11150 12880
rect 11206 12824 13266 12880
rect 13322 12824 13327 12880
rect 11145 12822 13327 12824
rect 11145 12819 11211 12822
rect 13261 12819 13327 12822
rect 14222 12820 14228 12884
rect 14292 12882 14298 12884
rect 14733 12882 14799 12885
rect 14292 12880 14799 12882
rect 14292 12824 14738 12880
rect 14794 12824 14799 12880
rect 14292 12822 14799 12824
rect 14292 12820 14298 12822
rect 14733 12819 14799 12822
rect 8293 12746 8359 12749
rect 8845 12748 8911 12749
rect 8845 12746 8892 12748
rect 8293 12744 8892 12746
rect 8293 12688 8298 12744
rect 8354 12688 8850 12744
rect 8293 12686 8892 12688
rect 8293 12683 8359 12686
rect 8845 12684 8892 12686
rect 8956 12684 8962 12748
rect 9857 12746 9923 12749
rect 18873 12746 18939 12749
rect 9857 12744 18939 12746
rect 9857 12688 9862 12744
rect 9918 12688 18878 12744
rect 18934 12688 18939 12744
rect 9857 12686 18939 12688
rect 8845 12683 8911 12684
rect 9857 12683 9923 12686
rect 18873 12683 18939 12686
rect 0 12610 480 12640
rect 4429 12610 4495 12613
rect 0 12608 4495 12610
rect 0 12552 4434 12608
rect 4490 12552 4495 12608
rect 0 12550 4495 12552
rect 0 12520 480 12550
rect 4429 12547 4495 12550
rect 10961 12610 11027 12613
rect 11830 12610 11836 12612
rect 10961 12608 11836 12610
rect 10961 12552 10966 12608
rect 11022 12552 11836 12608
rect 10961 12550 11836 12552
rect 10961 12547 11027 12550
rect 11830 12548 11836 12550
rect 11900 12548 11906 12612
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 2129 12474 2195 12477
rect 4838 12474 4844 12476
rect 2129 12472 4844 12474
rect 2129 12416 2134 12472
rect 2190 12416 4844 12472
rect 2129 12414 4844 12416
rect 2129 12411 2195 12414
rect 4838 12412 4844 12414
rect 4908 12412 4914 12476
rect 4981 12474 5047 12477
rect 5257 12474 5323 12477
rect 4981 12472 5323 12474
rect 4981 12416 4986 12472
rect 5042 12416 5262 12472
rect 5318 12416 5323 12472
rect 4981 12414 5323 12416
rect 4981 12411 5047 12414
rect 5257 12411 5323 12414
rect 8293 12476 8359 12477
rect 8293 12472 8340 12476
rect 8404 12474 8410 12476
rect 8845 12474 8911 12477
rect 10041 12474 10107 12477
rect 8293 12416 8298 12472
rect 8293 12412 8340 12416
rect 8404 12414 8450 12474
rect 8845 12472 10107 12474
rect 8845 12416 8850 12472
rect 8906 12416 10046 12472
rect 10102 12416 10107 12472
rect 8845 12414 10107 12416
rect 8404 12412 8410 12414
rect 8293 12411 8359 12412
rect 8845 12411 8911 12414
rect 10041 12411 10107 12414
rect 11973 12476 12039 12477
rect 19241 12476 19307 12477
rect 11973 12472 12020 12476
rect 12084 12474 12090 12476
rect 19190 12474 19196 12476
rect 11973 12416 11978 12472
rect 11973 12412 12020 12416
rect 12084 12414 12130 12474
rect 19150 12414 19196 12474
rect 19260 12472 19307 12476
rect 19302 12416 19307 12472
rect 12084 12412 12090 12414
rect 19190 12412 19196 12414
rect 19260 12412 19307 12416
rect 11973 12411 12039 12412
rect 19241 12411 19307 12412
rect 2773 12340 2839 12341
rect 2773 12336 2820 12340
rect 2884 12338 2890 12340
rect 2773 12280 2778 12336
rect 2773 12276 2820 12280
rect 2884 12278 2930 12338
rect 2884 12276 2890 12278
rect 4102 12276 4108 12340
rect 4172 12338 4178 12340
rect 6085 12338 6151 12341
rect 4172 12336 6151 12338
rect 4172 12280 6090 12336
rect 6146 12280 6151 12336
rect 4172 12278 6151 12280
rect 4172 12276 4178 12278
rect 2773 12275 2839 12276
rect 6085 12275 6151 12278
rect 6862 12276 6868 12340
rect 6932 12338 6938 12340
rect 7373 12338 7439 12341
rect 6932 12336 7439 12338
rect 6932 12280 7378 12336
rect 7434 12280 7439 12336
rect 6932 12278 7439 12280
rect 6932 12276 6938 12278
rect 7373 12275 7439 12278
rect 7925 12338 7991 12341
rect 8661 12338 8727 12341
rect 7925 12336 8727 12338
rect 7925 12280 7930 12336
rect 7986 12280 8666 12336
rect 8722 12280 8727 12336
rect 7925 12278 8727 12280
rect 7925 12275 7991 12278
rect 8661 12275 8727 12278
rect 12750 12276 12756 12340
rect 12820 12338 12826 12340
rect 14181 12338 14247 12341
rect 12820 12336 14247 12338
rect 12820 12280 14186 12336
rect 14242 12280 14247 12336
rect 12820 12278 14247 12280
rect 12820 12276 12826 12278
rect 14181 12275 14247 12278
rect 0 12202 480 12232
rect 14181 12204 14247 12205
rect 14181 12202 14228 12204
rect 0 12142 4860 12202
rect 14136 12200 14228 12202
rect 14136 12144 14186 12200
rect 14136 12142 14228 12144
rect 0 12112 480 12142
rect 4409 12000 4729 12001
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 4800 11794 4860 12142
rect 14181 12140 14228 12142
rect 14292 12140 14298 12204
rect 14181 12139 14247 12140
rect 5206 12004 5212 12068
rect 5276 12066 5282 12068
rect 5441 12066 5507 12069
rect 7005 12068 7071 12069
rect 7005 12066 7052 12068
rect 5276 12064 5507 12066
rect 5276 12008 5446 12064
rect 5502 12008 5507 12064
rect 5276 12006 5507 12008
rect 6960 12064 7052 12066
rect 6960 12008 7010 12064
rect 6960 12006 7052 12008
rect 5276 12004 5282 12006
rect 5441 12003 5507 12006
rect 7005 12004 7052 12006
rect 7116 12004 7122 12068
rect 7230 12004 7236 12068
rect 7300 12066 7306 12068
rect 13445 12066 13511 12069
rect 13854 12066 13860 12068
rect 7300 12006 9138 12066
rect 7300 12004 7306 12006
rect 7005 12003 7071 12004
rect 8753 11930 8819 11933
rect 8753 11928 8954 11930
rect 8753 11872 8758 11928
rect 8814 11872 8954 11928
rect 8753 11870 8954 11872
rect 8753 11867 8819 11870
rect 8334 11794 8340 11796
rect 4800 11734 8340 11794
rect 8334 11732 8340 11734
rect 8404 11732 8410 11796
rect 8661 11792 8727 11797
rect 8661 11736 8666 11792
rect 8722 11736 8727 11792
rect 8661 11731 8727 11736
rect 0 11658 480 11688
rect 4613 11658 4679 11661
rect 0 11656 4679 11658
rect 0 11600 4618 11656
rect 4674 11600 4679 11656
rect 0 11598 4679 11600
rect 0 11568 480 11598
rect 4613 11595 4679 11598
rect 4797 11658 4863 11661
rect 5257 11658 5323 11661
rect 4797 11656 5323 11658
rect 4797 11600 4802 11656
rect 4858 11600 5262 11656
rect 5318 11600 5323 11656
rect 4797 11598 5323 11600
rect 4797 11595 4863 11598
rect 5257 11595 5323 11598
rect 7414 11596 7420 11660
rect 7484 11658 7490 11660
rect 8664 11658 8724 11731
rect 7484 11598 8724 11658
rect 7484 11596 7490 11598
rect 2814 11460 2820 11524
rect 2884 11522 2890 11524
rect 6085 11522 6151 11525
rect 2884 11520 6151 11522
rect 2884 11464 6090 11520
rect 6146 11464 6151 11520
rect 2884 11462 6151 11464
rect 8894 11522 8954 11870
rect 9078 11794 9138 12006
rect 13445 12064 13860 12066
rect 13445 12008 13450 12064
rect 13506 12008 13860 12064
rect 13445 12006 13860 12008
rect 13445 12003 13511 12006
rect 13854 12004 13860 12006
rect 13924 12004 13930 12068
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 11789 11930 11855 11933
rect 13486 11930 13492 11932
rect 11789 11928 13492 11930
rect 11789 11872 11794 11928
rect 11850 11872 13492 11928
rect 11789 11870 13492 11872
rect 11789 11867 11855 11870
rect 13486 11868 13492 11870
rect 13556 11868 13562 11932
rect 13813 11930 13879 11933
rect 14273 11930 14339 11933
rect 13813 11928 14339 11930
rect 13813 11872 13818 11928
rect 13874 11872 14278 11928
rect 14334 11872 14339 11928
rect 13813 11870 14339 11872
rect 13813 11867 13879 11870
rect 14273 11867 14339 11870
rect 17677 11794 17743 11797
rect 9078 11792 17743 11794
rect 9078 11736 17682 11792
rect 17738 11736 17743 11792
rect 9078 11734 17743 11736
rect 17677 11731 17743 11734
rect 9029 11522 9095 11525
rect 8894 11520 9095 11522
rect 8894 11464 9034 11520
rect 9090 11464 9095 11520
rect 8894 11462 9095 11464
rect 2884 11460 2890 11462
rect 6085 11459 6151 11462
rect 9029 11459 9095 11462
rect 9949 11522 10015 11525
rect 12985 11522 13051 11525
rect 9949 11520 13051 11522
rect 9949 11464 9954 11520
rect 10010 11464 12990 11520
rect 13046 11464 13051 11520
rect 9949 11462 13051 11464
rect 9949 11459 10015 11462
rect 12985 11459 13051 11462
rect 19149 11522 19215 11525
rect 22520 11522 23000 11552
rect 19149 11520 23000 11522
rect 19149 11464 19154 11520
rect 19210 11464 23000 11520
rect 19149 11462 23000 11464
rect 19149 11459 19215 11462
rect 7874 11456 8194 11457
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 22520 11432 23000 11462
rect 14805 11391 15125 11392
rect 9438 11324 9444 11388
rect 9508 11386 9514 11388
rect 12801 11386 12867 11389
rect 9508 11384 12867 11386
rect 9508 11328 12806 11384
rect 12862 11328 12867 11384
rect 9508 11326 12867 11328
rect 9508 11324 9514 11326
rect 12801 11323 12867 11326
rect 5022 11188 5028 11252
rect 5092 11250 5098 11252
rect 5441 11250 5507 11253
rect 5092 11248 5507 11250
rect 5092 11192 5446 11248
rect 5502 11192 5507 11248
rect 5092 11190 5507 11192
rect 5092 11188 5098 11190
rect 5441 11187 5507 11190
rect 6678 11188 6684 11252
rect 6748 11250 6754 11252
rect 17493 11250 17559 11253
rect 6748 11248 17559 11250
rect 6748 11192 17498 11248
rect 17554 11192 17559 11248
rect 6748 11190 17559 11192
rect 6748 11188 6754 11190
rect 17493 11187 17559 11190
rect 0 11114 480 11144
rect 5022 11114 5028 11116
rect 0 11054 5028 11114
rect 0 11024 480 11054
rect 5022 11052 5028 11054
rect 5092 11114 5098 11116
rect 6177 11114 6243 11117
rect 5092 11112 6243 11114
rect 5092 11056 6182 11112
rect 6238 11056 6243 11112
rect 5092 11054 6243 11056
rect 5092 11052 5098 11054
rect 6177 11051 6243 11054
rect 6913 11114 6979 11117
rect 13077 11114 13143 11117
rect 6913 11112 13143 11114
rect 6913 11056 6918 11112
rect 6974 11056 13082 11112
rect 13138 11056 13143 11112
rect 6913 11054 13143 11056
rect 6913 11051 6979 11054
rect 13077 11051 13143 11054
rect 5901 10978 5967 10981
rect 8753 10978 8819 10981
rect 5901 10976 8819 10978
rect 5901 10920 5906 10976
rect 5962 10920 8758 10976
rect 8814 10920 8819 10976
rect 5901 10918 8819 10920
rect 5901 10915 5967 10918
rect 8753 10915 8819 10918
rect 12566 10916 12572 10980
rect 12636 10978 12642 10980
rect 15193 10978 15259 10981
rect 12636 10976 15259 10978
rect 12636 10920 15198 10976
rect 15254 10920 15259 10976
rect 12636 10918 15259 10920
rect 12636 10916 12642 10918
rect 15193 10915 15259 10918
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 12566 10780 12572 10844
rect 12636 10842 12642 10844
rect 14365 10842 14431 10845
rect 12636 10840 14431 10842
rect 12636 10784 14370 10840
rect 14426 10784 14431 10840
rect 12636 10782 14431 10784
rect 12636 10780 12642 10782
rect 14365 10779 14431 10782
rect 0 10706 480 10736
rect 8937 10706 9003 10709
rect 0 10704 9003 10706
rect 0 10648 8942 10704
rect 8998 10648 9003 10704
rect 0 10646 9003 10648
rect 0 10616 480 10646
rect 8937 10643 9003 10646
rect 11605 10706 11671 10709
rect 12525 10706 12591 10709
rect 17401 10706 17467 10709
rect 11605 10704 17467 10706
rect 11605 10648 11610 10704
rect 11666 10648 12530 10704
rect 12586 10648 17406 10704
rect 17462 10648 17467 10704
rect 11605 10646 17467 10648
rect 11605 10643 11671 10646
rect 12525 10643 12591 10646
rect 17401 10643 17467 10646
rect 9949 10570 10015 10573
rect 11513 10570 11579 10573
rect 9949 10568 11579 10570
rect 9949 10512 9954 10568
rect 10010 10512 11518 10568
rect 11574 10512 11579 10568
rect 9949 10510 11579 10512
rect 9949 10507 10015 10510
rect 11513 10507 11579 10510
rect 14089 10570 14155 10573
rect 17677 10570 17743 10573
rect 14089 10568 17743 10570
rect 14089 10512 14094 10568
rect 14150 10512 17682 10568
rect 17738 10512 17743 10568
rect 14089 10510 17743 10512
rect 14089 10507 14155 10510
rect 17677 10507 17743 10510
rect 6361 10434 6427 10437
rect 7046 10434 7052 10436
rect 6361 10432 7052 10434
rect 6361 10376 6366 10432
rect 6422 10376 7052 10432
rect 6361 10374 7052 10376
rect 6361 10371 6427 10374
rect 7046 10372 7052 10374
rect 7116 10372 7122 10436
rect 8702 10372 8708 10436
rect 8772 10434 8778 10436
rect 13169 10434 13235 10437
rect 8772 10432 13235 10434
rect 8772 10376 13174 10432
rect 13230 10376 13235 10432
rect 8772 10374 13235 10376
rect 8772 10372 8778 10374
rect 13169 10371 13235 10374
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 10303 15125 10304
rect 2262 10236 2268 10300
rect 2332 10298 2338 10300
rect 2589 10298 2655 10301
rect 2332 10296 2655 10298
rect 2332 10240 2594 10296
rect 2650 10240 2655 10296
rect 2332 10238 2655 10240
rect 2332 10236 2338 10238
rect 2589 10235 2655 10238
rect 3918 10236 3924 10300
rect 3988 10298 3994 10300
rect 6453 10298 6519 10301
rect 6821 10298 6887 10301
rect 3988 10296 6887 10298
rect 3988 10240 6458 10296
rect 6514 10240 6826 10296
rect 6882 10240 6887 10296
rect 3988 10238 6887 10240
rect 3988 10236 3994 10238
rect 6453 10235 6519 10238
rect 6821 10235 6887 10238
rect 9857 10298 9923 10301
rect 13077 10298 13143 10301
rect 9857 10296 13143 10298
rect 9857 10240 9862 10296
rect 9918 10240 13082 10296
rect 13138 10240 13143 10296
rect 9857 10238 13143 10240
rect 9857 10235 9923 10238
rect 13077 10235 13143 10238
rect 15561 10298 15627 10301
rect 15694 10298 15700 10300
rect 15561 10296 15700 10298
rect 15561 10240 15566 10296
rect 15622 10240 15700 10296
rect 15561 10238 15700 10240
rect 15561 10235 15627 10238
rect 15694 10236 15700 10238
rect 15764 10236 15770 10300
rect 0 10162 480 10192
rect 3969 10162 4035 10165
rect 0 10160 4035 10162
rect 0 10104 3974 10160
rect 4030 10104 4035 10160
rect 0 10102 4035 10104
rect 0 10072 480 10102
rect 3969 10099 4035 10102
rect 5533 10162 5599 10165
rect 5809 10162 5875 10165
rect 12198 10162 12204 10164
rect 5533 10160 12204 10162
rect 5533 10104 5538 10160
rect 5594 10104 5814 10160
rect 5870 10104 12204 10160
rect 5533 10102 12204 10104
rect 5533 10099 5599 10102
rect 5809 10099 5875 10102
rect 12198 10100 12204 10102
rect 12268 10100 12274 10164
rect 12341 10162 12407 10165
rect 15561 10162 15627 10165
rect 12341 10160 15627 10162
rect 12341 10104 12346 10160
rect 12402 10104 15566 10160
rect 15622 10104 15627 10160
rect 12341 10102 15627 10104
rect 12341 10099 12407 10102
rect 15561 10099 15627 10102
rect 2313 10026 2379 10029
rect 2681 10026 2747 10029
rect 7925 10026 7991 10029
rect 2313 10024 2747 10026
rect 2313 9968 2318 10024
rect 2374 9968 2686 10024
rect 2742 9968 2747 10024
rect 2313 9966 2747 9968
rect 2313 9963 2379 9966
rect 2681 9963 2747 9966
rect 4248 10024 7991 10026
rect 4248 9968 7930 10024
rect 7986 9968 7991 10024
rect 4248 9966 7991 9968
rect 1761 9890 1827 9893
rect 3877 9890 3943 9893
rect 1761 9888 3943 9890
rect 1761 9832 1766 9888
rect 1822 9832 3882 9888
rect 3938 9832 3943 9888
rect 1761 9830 3943 9832
rect 1761 9827 1827 9830
rect 3877 9827 3943 9830
rect 0 9754 480 9784
rect 4248 9754 4308 9966
rect 7925 9963 7991 9966
rect 8293 10026 8359 10029
rect 10961 10026 11027 10029
rect 8293 10024 11027 10026
rect 8293 9968 8298 10024
rect 8354 9968 10966 10024
rect 11022 9968 11027 10024
rect 8293 9966 11027 9968
rect 8293 9963 8359 9966
rect 10961 9963 11027 9966
rect 11145 10026 11211 10029
rect 11513 10026 11579 10029
rect 11145 10024 11579 10026
rect 11145 9968 11150 10024
rect 11206 9968 11518 10024
rect 11574 9968 11579 10024
rect 11145 9966 11579 9968
rect 11145 9963 11211 9966
rect 11513 9963 11579 9966
rect 11697 10026 11763 10029
rect 12382 10026 12388 10028
rect 11697 10024 12388 10026
rect 11697 9968 11702 10024
rect 11758 9968 12388 10024
rect 11697 9966 12388 9968
rect 11697 9963 11763 9966
rect 12382 9964 12388 9966
rect 12452 9964 12458 10028
rect 13721 10026 13787 10029
rect 16113 10026 16179 10029
rect 13721 10024 16179 10026
rect 13721 9968 13726 10024
rect 13782 9968 16118 10024
rect 16174 9968 16179 10024
rect 13721 9966 16179 9968
rect 13721 9963 13787 9966
rect 16113 9963 16179 9966
rect 6126 9828 6132 9892
rect 6196 9890 6202 9892
rect 7097 9890 7163 9893
rect 6196 9888 7163 9890
rect 6196 9832 7102 9888
rect 7158 9832 7163 9888
rect 6196 9830 7163 9832
rect 6196 9828 6202 9830
rect 7097 9827 7163 9830
rect 7465 9890 7531 9893
rect 9857 9890 9923 9893
rect 7465 9888 9923 9890
rect 7465 9832 7470 9888
rect 7526 9832 9862 9888
rect 9918 9832 9923 9888
rect 7465 9830 9923 9832
rect 7465 9827 7531 9830
rect 9857 9827 9923 9830
rect 10501 9890 10567 9893
rect 13537 9890 13603 9893
rect 16757 9890 16823 9893
rect 10501 9888 10610 9890
rect 10501 9832 10506 9888
rect 10562 9832 10610 9888
rect 10501 9827 10610 9832
rect 13537 9888 16823 9890
rect 13537 9832 13542 9888
rect 13598 9832 16762 9888
rect 16818 9832 16823 9888
rect 13537 9830 16823 9832
rect 13537 9827 13603 9830
rect 16757 9827 16823 9830
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 0 9694 4308 9754
rect 0 9664 480 9694
rect 5942 9692 5948 9756
rect 6012 9754 6018 9756
rect 7414 9754 7420 9756
rect 6012 9694 7420 9754
rect 6012 9692 6018 9694
rect 7414 9692 7420 9694
rect 7484 9692 7490 9756
rect 8017 9754 8083 9757
rect 8937 9754 9003 9757
rect 8017 9752 9003 9754
rect 8017 9696 8022 9752
rect 8078 9696 8942 9752
rect 8998 9696 9003 9752
rect 8017 9694 9003 9696
rect 10550 9754 10610 9827
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 10685 9754 10751 9757
rect 10550 9752 10751 9754
rect 10550 9696 10690 9752
rect 10746 9696 10751 9752
rect 10550 9694 10751 9696
rect 8017 9691 8083 9694
rect 8937 9691 9003 9694
rect 10685 9691 10751 9694
rect 12341 9754 12407 9757
rect 17585 9754 17651 9757
rect 12341 9752 17651 9754
rect 12341 9696 12346 9752
rect 12402 9696 17590 9752
rect 17646 9696 17651 9752
rect 12341 9694 17651 9696
rect 12341 9691 12407 9694
rect 17585 9691 17651 9694
rect 15745 9618 15811 9621
rect 2316 9616 15811 9618
rect 2316 9560 15750 9616
rect 15806 9560 15811 9616
rect 2316 9558 15811 9560
rect 2316 9485 2376 9558
rect 15745 9555 15811 9558
rect 1853 9482 1919 9485
rect 2078 9482 2084 9484
rect 1853 9480 2084 9482
rect 1853 9424 1858 9480
rect 1914 9424 2084 9480
rect 1853 9422 2084 9424
rect 1853 9419 1919 9422
rect 2078 9420 2084 9422
rect 2148 9420 2154 9484
rect 2313 9480 2379 9485
rect 2313 9424 2318 9480
rect 2374 9424 2379 9480
rect 2313 9419 2379 9424
rect 3182 9420 3188 9484
rect 3252 9420 3258 9484
rect 4521 9482 4587 9485
rect 4521 9480 8356 9482
rect 4521 9424 4526 9480
rect 4582 9424 8356 9480
rect 4521 9422 8356 9424
rect 3190 9346 3250 9420
rect 4521 9419 4587 9422
rect 4429 9346 4495 9349
rect 3190 9344 4495 9346
rect 3190 9288 4434 9344
rect 4490 9288 4495 9344
rect 3190 9286 4495 9288
rect 4429 9283 4495 9286
rect 6126 9284 6132 9348
rect 6196 9346 6202 9348
rect 6729 9346 6795 9349
rect 6196 9344 6795 9346
rect 6196 9288 6734 9344
rect 6790 9288 6795 9344
rect 6196 9286 6795 9288
rect 8296 9346 8356 9422
rect 9070 9420 9076 9484
rect 9140 9482 9146 9484
rect 9489 9482 9555 9485
rect 9140 9480 9555 9482
rect 9140 9424 9494 9480
rect 9550 9424 9555 9480
rect 9140 9422 9555 9424
rect 9140 9420 9146 9422
rect 9489 9419 9555 9422
rect 10317 9482 10383 9485
rect 14733 9482 14799 9485
rect 10317 9480 14799 9482
rect 10317 9424 10322 9480
rect 10378 9424 14738 9480
rect 14794 9424 14799 9480
rect 10317 9422 14799 9424
rect 10317 9419 10383 9422
rect 14733 9419 14799 9422
rect 12617 9346 12683 9349
rect 8296 9344 12683 9346
rect 8296 9288 12622 9344
rect 12678 9288 12683 9344
rect 8296 9286 12683 9288
rect 6196 9284 6202 9286
rect 6729 9283 6795 9286
rect 12617 9283 12683 9286
rect 7874 9280 8194 9281
rect 0 9210 480 9240
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 2313 9210 2379 9213
rect 0 9208 2379 9210
rect 0 9152 2318 9208
rect 2374 9152 2379 9208
rect 0 9150 2379 9152
rect 0 9120 480 9150
rect 2313 9147 2379 9150
rect 2446 9148 2452 9212
rect 2516 9210 2522 9212
rect 2589 9210 2655 9213
rect 3693 9210 3759 9213
rect 2516 9208 3759 9210
rect 2516 9152 2594 9208
rect 2650 9152 3698 9208
rect 3754 9152 3759 9208
rect 2516 9150 3759 9152
rect 2516 9148 2522 9150
rect 2589 9147 2655 9150
rect 3693 9147 3759 9150
rect 4705 9210 4771 9213
rect 7649 9210 7715 9213
rect 4705 9208 7715 9210
rect 4705 9152 4710 9208
rect 4766 9152 7654 9208
rect 7710 9152 7715 9208
rect 4705 9150 7715 9152
rect 4705 9147 4771 9150
rect 7649 9147 7715 9150
rect 8937 9210 9003 9213
rect 9438 9210 9444 9212
rect 8937 9208 9444 9210
rect 8937 9152 8942 9208
rect 8998 9152 9444 9208
rect 8937 9150 9444 9152
rect 8937 9147 9003 9150
rect 9438 9148 9444 9150
rect 9508 9148 9514 9212
rect 9622 9148 9628 9212
rect 9692 9210 9698 9212
rect 9765 9210 9831 9213
rect 9692 9208 9831 9210
rect 9692 9152 9770 9208
rect 9826 9152 9831 9208
rect 9692 9150 9831 9152
rect 9692 9148 9698 9150
rect 9765 9147 9831 9150
rect 14089 9210 14155 9213
rect 14457 9210 14523 9213
rect 14089 9208 14523 9210
rect 14089 9152 14094 9208
rect 14150 9152 14462 9208
rect 14518 9152 14523 9208
rect 14089 9150 14523 9152
rect 14089 9147 14155 9150
rect 14457 9147 14523 9150
rect 1853 9074 1919 9077
rect 18045 9074 18111 9077
rect 1853 9072 18111 9074
rect 1853 9016 1858 9072
rect 1914 9016 18050 9072
rect 18106 9016 18111 9072
rect 1853 9014 18111 9016
rect 1853 9011 1919 9014
rect 18045 9011 18111 9014
rect 4153 8938 4219 8941
rect 19701 8938 19767 8941
rect 4153 8936 19767 8938
rect 4153 8880 4158 8936
rect 4214 8880 19706 8936
rect 19762 8880 19767 8936
rect 4153 8878 19767 8880
rect 4153 8875 4219 8878
rect 19701 8875 19767 8878
rect 0 8802 480 8832
rect 4153 8804 4219 8805
rect 3182 8802 3188 8804
rect 0 8742 3188 8802
rect 0 8712 480 8742
rect 3182 8740 3188 8742
rect 3252 8740 3258 8804
rect 4102 8740 4108 8804
rect 4172 8802 4219 8804
rect 5073 8802 5139 8805
rect 10358 8802 10364 8804
rect 4172 8800 4264 8802
rect 4214 8744 4264 8800
rect 4172 8742 4264 8744
rect 5073 8800 10364 8802
rect 5073 8744 5078 8800
rect 5134 8744 10364 8800
rect 5073 8742 10364 8744
rect 4172 8740 4219 8742
rect 4153 8739 4219 8740
rect 5073 8739 5139 8742
rect 10358 8740 10364 8742
rect 10428 8740 10434 8804
rect 14222 8740 14228 8804
rect 14292 8802 14298 8804
rect 14365 8802 14431 8805
rect 14292 8800 14431 8802
rect 14292 8744 14370 8800
rect 14426 8744 14431 8800
rect 14292 8742 14431 8744
rect 14292 8740 14298 8742
rect 14365 8739 14431 8742
rect 4409 8736 4729 8737
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 2129 8666 2195 8669
rect 5809 8668 5875 8669
rect 4102 8666 4108 8668
rect 2129 8664 4108 8666
rect 2129 8608 2134 8664
rect 2190 8608 4108 8664
rect 2129 8606 4108 8608
rect 2129 8603 2195 8606
rect 4102 8604 4108 8606
rect 4172 8604 4178 8668
rect 5758 8666 5764 8668
rect 5718 8606 5764 8666
rect 5828 8664 5875 8668
rect 6545 8666 6611 8669
rect 5870 8608 5875 8664
rect 5758 8604 5764 8606
rect 5828 8604 5875 8608
rect 5809 8603 5875 8604
rect 5950 8664 6611 8666
rect 5950 8608 6550 8664
rect 6606 8608 6611 8664
rect 5950 8606 6611 8608
rect 2313 8530 2379 8533
rect 3693 8530 3759 8533
rect 5950 8530 6010 8606
rect 6545 8603 6611 8606
rect 7557 8666 7623 8669
rect 8702 8666 8708 8668
rect 7557 8664 8708 8666
rect 7557 8608 7562 8664
rect 7618 8608 8708 8664
rect 7557 8606 8708 8608
rect 7557 8603 7623 8606
rect 8702 8604 8708 8606
rect 8772 8604 8778 8668
rect 9857 8666 9923 8669
rect 11053 8668 11119 8669
rect 10910 8666 10916 8668
rect 9857 8664 10916 8666
rect 9857 8608 9862 8664
rect 9918 8608 10916 8664
rect 9857 8606 10916 8608
rect 9857 8603 9923 8606
rect 10910 8604 10916 8606
rect 10980 8604 10986 8668
rect 11053 8664 11100 8668
rect 11164 8666 11170 8668
rect 12525 8666 12591 8669
rect 16941 8666 17007 8669
rect 11053 8608 11058 8664
rect 11053 8604 11100 8608
rect 11164 8606 11210 8666
rect 12525 8664 17007 8666
rect 12525 8608 12530 8664
rect 12586 8608 16946 8664
rect 17002 8608 17007 8664
rect 12525 8606 17007 8608
rect 11164 8604 11170 8606
rect 11053 8603 11119 8604
rect 12525 8603 12591 8606
rect 16941 8603 17007 8606
rect 7414 8530 7420 8532
rect 2313 8528 2882 8530
rect 2313 8472 2318 8528
rect 2374 8472 2882 8528
rect 2313 8470 2882 8472
rect 2313 8467 2379 8470
rect 2589 8396 2655 8397
rect 2589 8392 2636 8396
rect 2700 8394 2706 8396
rect 2822 8394 2882 8470
rect 3693 8528 6010 8530
rect 3693 8472 3698 8528
rect 3754 8472 6010 8528
rect 3693 8470 6010 8472
rect 6456 8470 7420 8530
rect 3693 8467 3759 8470
rect 6456 8394 6516 8470
rect 7414 8468 7420 8470
rect 7484 8530 7490 8532
rect 13537 8530 13603 8533
rect 7484 8528 13603 8530
rect 7484 8472 13542 8528
rect 13598 8472 13603 8528
rect 7484 8470 13603 8472
rect 7484 8468 7490 8470
rect 13537 8467 13603 8470
rect 14273 8530 14339 8533
rect 16021 8530 16087 8533
rect 14273 8528 16087 8530
rect 14273 8472 14278 8528
rect 14334 8472 16026 8528
rect 16082 8472 16087 8528
rect 14273 8470 16087 8472
rect 14273 8467 14339 8470
rect 16021 8467 16087 8470
rect 2589 8336 2594 8392
rect 2589 8332 2636 8336
rect 2700 8334 2746 8394
rect 2822 8334 6516 8394
rect 7744 8334 8356 8394
rect 2700 8332 2706 8334
rect 2589 8331 2655 8332
rect 0 8258 480 8288
rect 5758 8258 5764 8260
rect 0 8198 5764 8258
rect 0 8168 480 8198
rect 5758 8196 5764 8198
rect 5828 8196 5834 8260
rect 7744 8122 7804 8334
rect 8296 8258 8356 8334
rect 10542 8332 10548 8396
rect 10612 8394 10618 8396
rect 17125 8394 17191 8397
rect 10612 8392 17191 8394
rect 10612 8336 17130 8392
rect 17186 8336 17191 8392
rect 10612 8334 17191 8336
rect 10612 8332 10618 8334
rect 17125 8331 17191 8334
rect 12014 8258 12020 8260
rect 8296 8198 12020 8258
rect 12014 8196 12020 8198
rect 12084 8196 12090 8260
rect 7874 8192 8194 8193
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 3742 8062 7804 8122
rect 8296 8062 14658 8122
rect 0 7850 480 7880
rect 1853 7850 1919 7853
rect 0 7848 1919 7850
rect 0 7792 1858 7848
rect 1914 7792 1919 7848
rect 0 7790 1919 7792
rect 0 7760 480 7790
rect 1853 7787 1919 7790
rect 2037 7850 2103 7853
rect 3742 7850 3802 8062
rect 3969 7986 4035 7989
rect 8296 7986 8356 8062
rect 3969 7984 8356 7986
rect 3969 7928 3974 7984
rect 4030 7928 8356 7984
rect 3969 7926 8356 7928
rect 3969 7923 4035 7926
rect 8886 7924 8892 7988
rect 8956 7986 8962 7988
rect 11421 7986 11487 7989
rect 8956 7984 11487 7986
rect 8956 7928 11426 7984
rect 11482 7928 11487 7984
rect 8956 7926 11487 7928
rect 8956 7924 8962 7926
rect 11421 7923 11487 7926
rect 12985 7986 13051 7989
rect 13118 7986 13124 7988
rect 12985 7984 13124 7986
rect 12985 7928 12990 7984
rect 13046 7928 13124 7984
rect 12985 7926 13124 7928
rect 12985 7923 13051 7926
rect 13118 7924 13124 7926
rect 13188 7924 13194 7988
rect 14598 7986 14658 8062
rect 15837 7986 15903 7989
rect 14598 7984 15903 7986
rect 14598 7928 15842 7984
rect 15898 7928 15903 7984
rect 14598 7926 15903 7928
rect 15837 7923 15903 7926
rect 2037 7848 3802 7850
rect 2037 7792 2042 7848
rect 2098 7792 3802 7848
rect 4429 7848 4495 7853
rect 4429 7816 4434 7848
rect 2037 7790 3802 7792
rect 4294 7792 4434 7816
rect 4490 7792 4495 7848
rect 2037 7787 2103 7790
rect 4294 7787 4495 7792
rect 4613 7850 4679 7853
rect 4838 7850 4844 7852
rect 4613 7848 4844 7850
rect 4613 7792 4618 7848
rect 4674 7792 4844 7848
rect 4613 7790 4844 7792
rect 4613 7787 4679 7790
rect 4838 7788 4844 7790
rect 4908 7788 4914 7852
rect 5809 7850 5875 7853
rect 6177 7850 6243 7853
rect 5809 7848 6243 7850
rect 5809 7792 5814 7848
rect 5870 7792 6182 7848
rect 6238 7792 6243 7848
rect 5809 7790 6243 7792
rect 5809 7787 5875 7790
rect 6177 7787 6243 7790
rect 6637 7850 6703 7853
rect 7741 7850 7807 7853
rect 6637 7848 7807 7850
rect 6637 7792 6642 7848
rect 6698 7792 7746 7848
rect 7802 7792 7807 7848
rect 6637 7790 7807 7792
rect 6637 7787 6703 7790
rect 7741 7787 7807 7790
rect 8017 7850 8083 7853
rect 8334 7850 8340 7852
rect 8017 7848 8340 7850
rect 8017 7792 8022 7848
rect 8078 7792 8340 7848
rect 8017 7790 8340 7792
rect 8017 7787 8083 7790
rect 8334 7788 8340 7790
rect 8404 7788 8410 7852
rect 8661 7850 8727 7853
rect 18137 7850 18203 7853
rect 8661 7848 18203 7850
rect 8661 7792 8666 7848
rect 8722 7792 18142 7848
rect 18198 7792 18203 7848
rect 8661 7790 18203 7792
rect 8661 7787 8727 7790
rect 18137 7787 18203 7790
rect 4294 7756 4492 7787
rect 4294 7748 4354 7756
rect 3182 7652 3188 7716
rect 3252 7714 3258 7716
rect 4248 7714 4354 7748
rect 3252 7688 4354 7714
rect 3252 7654 4308 7688
rect 4846 7654 11208 7714
rect 3252 7652 3258 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 2865 7578 2931 7581
rect 3325 7578 3391 7581
rect 2865 7576 3391 7578
rect 2865 7520 2870 7576
rect 2926 7520 3330 7576
rect 3386 7520 3391 7576
rect 2865 7518 3391 7520
rect 2865 7515 2931 7518
rect 3325 7515 3391 7518
rect 1761 7442 1827 7445
rect 4846 7442 4906 7654
rect 4981 7578 5047 7581
rect 9029 7578 9095 7581
rect 4981 7576 9095 7578
rect 4981 7520 4986 7576
rect 5042 7520 9034 7576
rect 9090 7520 9095 7576
rect 4981 7518 9095 7520
rect 4981 7515 5047 7518
rect 9029 7515 9095 7518
rect 9765 7578 9831 7581
rect 10593 7578 10659 7581
rect 9765 7576 10659 7578
rect 9765 7520 9770 7576
rect 9826 7520 10598 7576
rect 10654 7520 10659 7576
rect 9765 7518 10659 7520
rect 9765 7515 9831 7518
rect 10593 7515 10659 7518
rect 10726 7516 10732 7580
rect 10796 7578 10802 7580
rect 10961 7578 11027 7581
rect 10796 7576 11027 7578
rect 10796 7520 10966 7576
rect 11022 7520 11027 7576
rect 10796 7518 11027 7520
rect 10796 7516 10802 7518
rect 10961 7515 11027 7518
rect 1761 7440 4906 7442
rect 1761 7384 1766 7440
rect 1822 7384 4906 7440
rect 1761 7382 4906 7384
rect 5073 7442 5139 7445
rect 5206 7442 5212 7444
rect 5073 7440 5212 7442
rect 5073 7384 5078 7440
rect 5134 7384 5212 7440
rect 5073 7382 5212 7384
rect 1761 7379 1827 7382
rect 5073 7379 5139 7382
rect 5206 7380 5212 7382
rect 5276 7380 5282 7444
rect 6085 7442 6151 7445
rect 10961 7444 11027 7445
rect 6085 7440 9874 7442
rect 6085 7384 6090 7440
rect 6146 7384 9874 7440
rect 6085 7382 9874 7384
rect 6085 7379 6151 7382
rect 0 7306 480 7336
rect 5257 7306 5323 7309
rect 9814 7306 9874 7382
rect 10910 7380 10916 7444
rect 10980 7442 11027 7444
rect 11148 7442 11208 7654
rect 12934 7652 12940 7716
rect 13004 7714 13010 7716
rect 13629 7714 13695 7717
rect 13004 7712 13695 7714
rect 13004 7656 13634 7712
rect 13690 7656 13695 7712
rect 13004 7654 13695 7656
rect 13004 7652 13010 7654
rect 13629 7651 13695 7654
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 7583 18590 7584
rect 14457 7578 14523 7581
rect 16665 7578 16731 7581
rect 14457 7576 16731 7578
rect 14457 7520 14462 7576
rect 14518 7520 16670 7576
rect 16726 7520 16731 7576
rect 14457 7518 16731 7520
rect 14457 7515 14523 7518
rect 16665 7515 16731 7518
rect 11830 7442 11836 7444
rect 10980 7440 11072 7442
rect 11022 7384 11072 7440
rect 10980 7382 11072 7384
rect 11148 7382 11836 7442
rect 10980 7380 11027 7382
rect 11830 7380 11836 7382
rect 11900 7442 11906 7444
rect 19333 7442 19399 7445
rect 11900 7440 19399 7442
rect 11900 7384 19338 7440
rect 19394 7384 19399 7440
rect 11900 7382 19399 7384
rect 11900 7380 11906 7382
rect 10961 7379 11027 7380
rect 19333 7379 19399 7382
rect 19793 7306 19859 7309
rect 0 7246 5136 7306
rect 0 7216 480 7246
rect 2129 7170 2195 7173
rect 5076 7170 5136 7246
rect 5257 7304 8356 7306
rect 5257 7248 5262 7304
rect 5318 7248 8356 7304
rect 5257 7246 8356 7248
rect 9814 7304 19859 7306
rect 9814 7248 19798 7304
rect 19854 7248 19859 7304
rect 9814 7246 19859 7248
rect 5257 7243 5323 7246
rect 6453 7170 6519 7173
rect 2129 7168 4906 7170
rect 2129 7112 2134 7168
rect 2190 7112 4906 7168
rect 2129 7110 4906 7112
rect 5076 7168 6519 7170
rect 5076 7112 6458 7168
rect 6514 7112 6519 7168
rect 5076 7110 6519 7112
rect 2129 7107 2195 7110
rect 3366 6972 3372 7036
rect 3436 7034 3442 7036
rect 3601 7034 3667 7037
rect 3436 7032 3667 7034
rect 3436 6976 3606 7032
rect 3662 6976 3667 7032
rect 3436 6974 3667 6976
rect 4846 7034 4906 7110
rect 6453 7107 6519 7110
rect 7281 7170 7347 7173
rect 7741 7170 7807 7173
rect 7281 7168 7807 7170
rect 7281 7112 7286 7168
rect 7342 7112 7746 7168
rect 7802 7112 7807 7168
rect 7281 7110 7807 7112
rect 7281 7107 7347 7110
rect 7741 7107 7807 7110
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 5533 7034 5599 7037
rect 4846 7032 5599 7034
rect 4846 6976 5538 7032
rect 5594 6976 5599 7032
rect 4846 6974 5599 6976
rect 3436 6972 3442 6974
rect 3601 6971 3667 6974
rect 5533 6971 5599 6974
rect 5758 6972 5764 7036
rect 5828 7034 5834 7036
rect 6361 7034 6427 7037
rect 5828 7032 6427 7034
rect 5828 6976 6366 7032
rect 6422 6976 6427 7032
rect 5828 6974 6427 6976
rect 8296 7034 8356 7246
rect 19793 7243 19859 7246
rect 9489 7170 9555 7173
rect 12893 7170 12959 7173
rect 9489 7168 12959 7170
rect 9489 7112 9494 7168
rect 9550 7112 12898 7168
rect 12954 7112 12959 7168
rect 9489 7110 12959 7112
rect 9489 7107 9555 7110
rect 12893 7107 12959 7110
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 7039 15125 7040
rect 9857 7034 9923 7037
rect 10910 7034 10916 7036
rect 8296 6974 9690 7034
rect 5828 6972 5834 6974
rect 6361 6971 6427 6974
rect 0 6898 480 6928
rect 3693 6898 3759 6901
rect 0 6896 3759 6898
rect 0 6840 3698 6896
rect 3754 6840 3759 6896
rect 0 6838 3759 6840
rect 0 6808 480 6838
rect 3693 6835 3759 6838
rect 4102 6836 4108 6900
rect 4172 6898 4178 6900
rect 5206 6898 5212 6900
rect 4172 6838 5212 6898
rect 4172 6836 4178 6838
rect 5206 6836 5212 6838
rect 5276 6898 5282 6900
rect 9121 6898 9187 6901
rect 9305 6900 9371 6901
rect 5276 6896 9187 6898
rect 5276 6840 9126 6896
rect 9182 6840 9187 6896
rect 5276 6838 9187 6840
rect 5276 6836 5282 6838
rect 9121 6835 9187 6838
rect 9254 6836 9260 6900
rect 9324 6898 9371 6900
rect 9630 6898 9690 6974
rect 9857 7032 10916 7034
rect 9857 6976 9862 7032
rect 9918 6976 10916 7032
rect 9857 6974 10916 6976
rect 9857 6971 9923 6974
rect 10910 6972 10916 6974
rect 10980 7034 10986 7036
rect 11697 7034 11763 7037
rect 10980 7032 11763 7034
rect 10980 6976 11702 7032
rect 11758 6976 11763 7032
rect 10980 6974 11763 6976
rect 10980 6972 10986 6974
rect 11697 6971 11763 6974
rect 12382 6972 12388 7036
rect 12452 7034 12458 7036
rect 14549 7034 14615 7037
rect 12452 7032 14615 7034
rect 12452 6976 14554 7032
rect 14610 6976 14615 7032
rect 12452 6974 14615 6976
rect 12452 6972 12458 6974
rect 14549 6971 14615 6974
rect 19609 6898 19675 6901
rect 9324 6896 9416 6898
rect 9366 6840 9416 6896
rect 9324 6838 9416 6840
rect 9630 6896 19675 6898
rect 9630 6840 19614 6896
rect 19670 6840 19675 6896
rect 9630 6838 19675 6840
rect 9324 6836 9371 6838
rect 9305 6835 9371 6836
rect 19609 6835 19675 6838
rect 2957 6762 3023 6765
rect 14549 6762 14615 6765
rect 2957 6760 14615 6762
rect 2957 6704 2962 6760
rect 3018 6704 14554 6760
rect 14610 6704 14615 6760
rect 2957 6702 14615 6704
rect 2957 6699 3023 6702
rect 14549 6699 14615 6702
rect 4102 6564 4108 6628
rect 4172 6626 4178 6628
rect 4245 6626 4311 6629
rect 4172 6624 4311 6626
rect 4172 6568 4250 6624
rect 4306 6568 4311 6624
rect 4172 6566 4311 6568
rect 4172 6564 4178 6566
rect 4245 6563 4311 6566
rect 4981 6626 5047 6629
rect 10726 6626 10732 6628
rect 4981 6624 10732 6626
rect 4981 6568 4986 6624
rect 5042 6568 10732 6624
rect 4981 6566 10732 6568
rect 4981 6563 5047 6566
rect 10726 6564 10732 6566
rect 10796 6564 10802 6628
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 1853 6490 1919 6493
rect 4061 6490 4127 6493
rect 1853 6488 4127 6490
rect 1853 6432 1858 6488
rect 1914 6432 4066 6488
rect 4122 6432 4127 6488
rect 1853 6430 4127 6432
rect 1853 6427 1919 6430
rect 4061 6427 4127 6430
rect 5206 6428 5212 6492
rect 5276 6490 5282 6492
rect 5349 6490 5415 6493
rect 6269 6492 6335 6493
rect 6269 6490 6316 6492
rect 5276 6488 5415 6490
rect 5276 6432 5354 6488
rect 5410 6432 5415 6488
rect 5276 6430 5415 6432
rect 6224 6488 6316 6490
rect 6224 6432 6274 6488
rect 6224 6430 6316 6432
rect 5276 6428 5282 6430
rect 5349 6427 5415 6430
rect 6269 6428 6316 6430
rect 6380 6428 6386 6492
rect 6453 6490 6519 6493
rect 6678 6490 6684 6492
rect 6453 6488 6684 6490
rect 6453 6432 6458 6488
rect 6514 6432 6684 6488
rect 6453 6430 6684 6432
rect 6269 6427 6335 6428
rect 6453 6427 6519 6430
rect 6678 6428 6684 6430
rect 6748 6428 6754 6492
rect 6821 6490 6887 6493
rect 7046 6490 7052 6492
rect 6821 6488 7052 6490
rect 6821 6432 6826 6488
rect 6882 6432 7052 6488
rect 6821 6430 7052 6432
rect 6821 6427 6887 6430
rect 7046 6428 7052 6430
rect 7116 6490 7122 6492
rect 10593 6490 10659 6493
rect 7116 6488 10659 6490
rect 7116 6432 10598 6488
rect 10654 6432 10659 6488
rect 7116 6430 10659 6432
rect 7116 6428 7122 6430
rect 10593 6427 10659 6430
rect 12157 6490 12223 6493
rect 15745 6490 15811 6493
rect 12157 6488 15811 6490
rect 12157 6432 12162 6488
rect 12218 6432 15750 6488
rect 15806 6432 15811 6488
rect 12157 6430 15811 6432
rect 12157 6427 12223 6430
rect 15745 6427 15811 6430
rect 0 6354 480 6384
rect 3969 6354 4035 6357
rect 0 6352 4035 6354
rect 0 6296 3974 6352
rect 4030 6296 4035 6352
rect 0 6294 4035 6296
rect 0 6264 480 6294
rect 3969 6291 4035 6294
rect 5206 6292 5212 6356
rect 5276 6354 5282 6356
rect 5717 6354 5783 6357
rect 5276 6352 5783 6354
rect 5276 6296 5722 6352
rect 5778 6296 5783 6352
rect 5276 6294 5783 6296
rect 5276 6292 5282 6294
rect 5717 6291 5783 6294
rect 7373 6354 7439 6357
rect 18505 6354 18571 6357
rect 7373 6352 18571 6354
rect 7373 6296 7378 6352
rect 7434 6296 18510 6352
rect 18566 6296 18571 6352
rect 7373 6294 18571 6296
rect 7373 6291 7439 6294
rect 18505 6291 18571 6294
rect 4429 6218 4495 6221
rect 18045 6218 18111 6221
rect 2868 6158 4354 6218
rect 2868 6082 2928 6158
rect 3233 6082 3299 6085
rect 1166 6022 2928 6082
rect 3006 6080 3299 6082
rect 3006 6024 3238 6080
rect 3294 6024 3299 6080
rect 3006 6022 3299 6024
rect 4294 6082 4354 6158
rect 4429 6216 11024 6218
rect 4429 6160 4434 6216
rect 4490 6160 11024 6216
rect 4429 6158 11024 6160
rect 4429 6155 4495 6158
rect 6637 6082 6703 6085
rect 7046 6082 7052 6084
rect 4294 6022 6562 6082
rect 0 5946 480 5976
rect 1166 5946 1226 6022
rect 0 5886 1226 5946
rect 0 5856 480 5886
rect 3006 5810 3066 6022
rect 3233 6019 3299 6022
rect 3969 5946 4035 5949
rect 6361 5946 6427 5949
rect 3969 5944 6427 5946
rect 3969 5888 3974 5944
rect 4030 5888 6366 5944
rect 6422 5888 6427 5944
rect 3969 5886 6427 5888
rect 6502 5946 6562 6022
rect 6637 6080 7052 6082
rect 6637 6024 6642 6080
rect 6698 6024 7052 6080
rect 6637 6022 7052 6024
rect 6637 6019 6703 6022
rect 7046 6020 7052 6022
rect 7116 6082 7122 6084
rect 7741 6082 7807 6085
rect 7116 6080 7807 6082
rect 7116 6024 7746 6080
rect 7802 6024 7807 6080
rect 7116 6022 7807 6024
rect 7116 6020 7122 6022
rect 7741 6019 7807 6022
rect 8385 6082 8451 6085
rect 9438 6082 9444 6084
rect 8385 6080 9444 6082
rect 8385 6024 8390 6080
rect 8446 6024 9444 6080
rect 8385 6022 9444 6024
rect 8385 6019 8451 6022
rect 9438 6020 9444 6022
rect 9508 6020 9514 6084
rect 10041 6082 10107 6085
rect 10501 6082 10567 6085
rect 10041 6080 10567 6082
rect 10041 6024 10046 6080
rect 10102 6024 10506 6080
rect 10562 6024 10567 6080
rect 10041 6022 10567 6024
rect 10041 6019 10107 6022
rect 10501 6019 10567 6022
rect 10685 6084 10751 6085
rect 10685 6080 10732 6084
rect 10796 6082 10802 6084
rect 10964 6082 11024 6158
rect 11286 6216 18111 6218
rect 11286 6160 18050 6216
rect 18106 6160 18111 6216
rect 11286 6158 18111 6160
rect 11286 6082 11346 6158
rect 18045 6155 18111 6158
rect 10685 6024 10690 6080
rect 10685 6020 10732 6024
rect 10796 6022 10842 6082
rect 10964 6022 11346 6082
rect 11421 6082 11487 6085
rect 11830 6082 11836 6084
rect 11421 6080 11836 6082
rect 11421 6024 11426 6080
rect 11482 6024 11836 6080
rect 11421 6022 11836 6024
rect 10796 6020 10802 6022
rect 10685 6019 10751 6020
rect 11421 6019 11487 6022
rect 11830 6020 11836 6022
rect 11900 6020 11906 6084
rect 12198 6020 12204 6084
rect 12268 6082 12274 6084
rect 12341 6082 12407 6085
rect 12268 6080 12407 6082
rect 12268 6024 12346 6080
rect 12402 6024 12407 6080
rect 12268 6022 12407 6024
rect 12268 6020 12274 6022
rect 12341 6019 12407 6022
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 7281 5946 7347 5949
rect 6502 5944 7347 5946
rect 6502 5888 7286 5944
rect 7342 5888 7347 5944
rect 6502 5886 7347 5888
rect 3969 5883 4035 5886
rect 6361 5883 6427 5886
rect 7281 5883 7347 5886
rect 8293 5946 8359 5949
rect 8293 5944 13876 5946
rect 8293 5888 8298 5944
rect 8354 5888 13876 5944
rect 8293 5886 13876 5888
rect 8293 5883 8359 5886
rect 13629 5810 13695 5813
rect 3006 5808 13695 5810
rect 3006 5752 13634 5808
rect 13690 5752 13695 5808
rect 3006 5750 13695 5752
rect 13816 5810 13876 5886
rect 17401 5810 17467 5813
rect 13816 5808 17467 5810
rect 13816 5752 17406 5808
rect 17462 5752 17467 5808
rect 13816 5750 17467 5752
rect 13629 5747 13695 5750
rect 17401 5747 17467 5750
rect 1393 5674 1459 5677
rect 5809 5674 5875 5677
rect 6729 5674 6795 5677
rect 16573 5674 16639 5677
rect 20069 5674 20135 5677
rect 1393 5672 5875 5674
rect 1393 5616 1398 5672
rect 1454 5616 5814 5672
rect 5870 5616 5875 5672
rect 1393 5614 5875 5616
rect 1393 5611 1459 5614
rect 5809 5611 5875 5614
rect 5950 5672 6795 5674
rect 5950 5616 6734 5672
rect 6790 5616 6795 5672
rect 5950 5614 6795 5616
rect 3325 5538 3391 5541
rect 3918 5538 3924 5540
rect 3325 5536 3924 5538
rect 3325 5480 3330 5536
rect 3386 5480 3924 5536
rect 3325 5478 3924 5480
rect 3325 5475 3391 5478
rect 3918 5476 3924 5478
rect 3988 5476 3994 5540
rect 5950 5538 6010 5614
rect 6729 5611 6795 5614
rect 7790 5672 20135 5674
rect 7790 5616 16578 5672
rect 16634 5616 20074 5672
rect 20130 5616 20135 5672
rect 7790 5614 20135 5616
rect 5214 5478 6010 5538
rect 4409 5472 4729 5473
rect 0 5402 480 5432
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 3601 5402 3667 5405
rect 0 5400 3667 5402
rect 0 5344 3606 5400
rect 3662 5344 3667 5400
rect 0 5342 3667 5344
rect 0 5312 480 5342
rect 3601 5339 3667 5342
rect 5214 5269 5274 5478
rect 6310 5476 6316 5540
rect 6380 5538 6386 5540
rect 7790 5538 7850 5614
rect 16573 5611 16639 5614
rect 20069 5611 20135 5614
rect 6380 5478 7850 5538
rect 8753 5538 8819 5541
rect 9949 5538 10015 5541
rect 10501 5538 10567 5541
rect 10961 5538 11027 5541
rect 8753 5536 11027 5538
rect 8753 5480 8758 5536
rect 8814 5480 9954 5536
rect 10010 5480 10506 5536
rect 10562 5480 10966 5536
rect 11022 5480 11027 5536
rect 8753 5478 11027 5480
rect 6380 5476 6386 5478
rect 8753 5475 8819 5478
rect 9949 5475 10015 5478
rect 10501 5475 10567 5478
rect 10961 5475 11027 5478
rect 12801 5538 12867 5541
rect 15377 5538 15443 5541
rect 12801 5536 15443 5538
rect 12801 5480 12806 5536
rect 12862 5480 15382 5536
rect 15438 5480 15443 5536
rect 12801 5478 15443 5480
rect 12801 5475 12867 5478
rect 15377 5475 15443 5478
rect 15510 5476 15516 5540
rect 15580 5538 15586 5540
rect 15745 5538 15811 5541
rect 15580 5536 15811 5538
rect 15580 5480 15750 5536
rect 15806 5480 15811 5536
rect 15580 5478 15811 5480
rect 15580 5476 15586 5478
rect 15745 5475 15811 5478
rect 15929 5536 15995 5541
rect 15929 5480 15934 5536
rect 15990 5480 15995 5536
rect 15929 5475 15995 5480
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 5349 5402 5415 5405
rect 9121 5402 9187 5405
rect 5349 5400 9187 5402
rect 5349 5344 5354 5400
rect 5410 5344 9126 5400
rect 9182 5344 9187 5400
rect 5349 5342 9187 5344
rect 5349 5339 5415 5342
rect 9121 5339 9187 5342
rect 9397 5402 9463 5405
rect 11053 5402 11119 5405
rect 9397 5400 11119 5402
rect 9397 5344 9402 5400
rect 9458 5344 11058 5400
rect 11114 5344 11119 5400
rect 9397 5342 11119 5344
rect 9397 5339 9463 5342
rect 11053 5339 11119 5342
rect 12198 5340 12204 5404
rect 12268 5402 12274 5404
rect 15561 5402 15627 5405
rect 12268 5400 15627 5402
rect 12268 5344 15566 5400
rect 15622 5344 15627 5400
rect 12268 5342 15627 5344
rect 12268 5340 12274 5342
rect 15561 5339 15627 5342
rect 15694 5340 15700 5404
rect 15764 5402 15770 5404
rect 15932 5402 15992 5475
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 15764 5342 15992 5402
rect 15764 5340 15770 5342
rect 4102 5204 4108 5268
rect 4172 5266 4178 5268
rect 4245 5266 4311 5269
rect 4172 5264 4311 5266
rect 4172 5208 4250 5264
rect 4306 5208 4311 5264
rect 4172 5206 4311 5208
rect 5214 5264 5323 5269
rect 5214 5208 5262 5264
rect 5318 5208 5323 5264
rect 5214 5206 5323 5208
rect 4172 5204 4178 5206
rect 4245 5203 4311 5206
rect 5257 5203 5323 5206
rect 5942 5204 5948 5268
rect 6012 5266 6018 5268
rect 6361 5266 6427 5269
rect 6012 5264 6427 5266
rect 6012 5208 6366 5264
rect 6422 5208 6427 5264
rect 6012 5206 6427 5208
rect 6012 5204 6018 5206
rect 6361 5203 6427 5206
rect 6862 5204 6868 5268
rect 6932 5266 6938 5268
rect 7925 5266 7991 5269
rect 6932 5264 7991 5266
rect 6932 5208 7930 5264
rect 7986 5208 7991 5264
rect 6932 5206 7991 5208
rect 6932 5204 6938 5206
rect 7925 5203 7991 5206
rect 8201 5266 8267 5269
rect 8334 5266 8340 5268
rect 8201 5264 8340 5266
rect 8201 5208 8206 5264
rect 8262 5208 8340 5264
rect 8201 5206 8340 5208
rect 8201 5203 8267 5206
rect 8334 5204 8340 5206
rect 8404 5204 8410 5268
rect 8661 5266 8727 5269
rect 12566 5266 12572 5268
rect 8661 5264 12572 5266
rect 8661 5208 8666 5264
rect 8722 5208 12572 5264
rect 8661 5206 12572 5208
rect 8661 5203 8727 5206
rect 12566 5204 12572 5206
rect 12636 5204 12642 5268
rect 2497 5130 2563 5133
rect 19609 5130 19675 5133
rect 2497 5128 19675 5130
rect 2497 5072 2502 5128
rect 2558 5072 19614 5128
rect 19670 5072 19675 5128
rect 2497 5070 19675 5072
rect 2497 5067 2563 5070
rect 19609 5067 19675 5070
rect 0 4994 480 5024
rect 6126 4994 6132 4996
rect 0 4934 6132 4994
rect 0 4904 480 4934
rect 6126 4932 6132 4934
rect 6196 4932 6202 4996
rect 6453 4994 6519 4997
rect 7557 4994 7623 4997
rect 6453 4992 7623 4994
rect 6453 4936 6458 4992
rect 6514 4936 7562 4992
rect 7618 4936 7623 4992
rect 6453 4934 7623 4936
rect 6453 4931 6519 4934
rect 7557 4931 7623 4934
rect 8385 4994 8451 4997
rect 13537 4994 13603 4997
rect 8385 4992 13603 4994
rect 8385 4936 8390 4992
rect 8446 4936 13542 4992
rect 13598 4936 13603 4992
rect 8385 4934 13603 4936
rect 8385 4931 8451 4934
rect 13537 4931 13603 4934
rect 7874 4928 8194 4929
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 3325 4858 3391 4861
rect 3550 4858 3556 4860
rect 3325 4856 3556 4858
rect 3325 4800 3330 4856
rect 3386 4800 3556 4856
rect 3325 4798 3556 4800
rect 3325 4795 3391 4798
rect 3550 4796 3556 4798
rect 3620 4796 3626 4860
rect 5349 4858 5415 4861
rect 6494 4858 6500 4860
rect 5349 4856 6500 4858
rect 5349 4800 5354 4856
rect 5410 4800 6500 4856
rect 5349 4798 6500 4800
rect 5349 4795 5415 4798
rect 6494 4796 6500 4798
rect 6564 4796 6570 4860
rect 9489 4858 9555 4861
rect 12433 4858 12499 4861
rect 9489 4856 12499 4858
rect 9489 4800 9494 4856
rect 9550 4800 12438 4856
rect 12494 4800 12499 4856
rect 9489 4798 12499 4800
rect 9489 4795 9555 4798
rect 12433 4795 12499 4798
rect 1669 4722 1735 4725
rect 3785 4722 3851 4725
rect 5390 4722 5396 4724
rect 1669 4720 5396 4722
rect 1669 4664 1674 4720
rect 1730 4664 3790 4720
rect 3846 4664 5396 4720
rect 1669 4662 5396 4664
rect 1669 4659 1735 4662
rect 3785 4659 3851 4662
rect 5390 4660 5396 4662
rect 5460 4660 5466 4724
rect 5625 4722 5691 4725
rect 12198 4722 12204 4724
rect 5625 4720 12204 4722
rect 5625 4664 5630 4720
rect 5686 4664 12204 4720
rect 5625 4662 12204 4664
rect 5625 4659 5691 4662
rect 12198 4660 12204 4662
rect 12268 4660 12274 4724
rect 15561 4722 15627 4725
rect 12574 4720 15627 4722
rect 12574 4664 15566 4720
rect 15622 4664 15627 4720
rect 12574 4662 15627 4664
rect 2129 4586 2195 4589
rect 12574 4586 12634 4662
rect 15561 4659 15627 4662
rect 15837 4722 15903 4725
rect 19057 4722 19123 4725
rect 15837 4720 19123 4722
rect 15837 4664 15842 4720
rect 15898 4664 19062 4720
rect 19118 4664 19123 4720
rect 15837 4662 19123 4664
rect 15837 4659 15903 4662
rect 19057 4659 19123 4662
rect 2129 4584 12634 4586
rect 2129 4528 2134 4584
rect 2190 4528 12634 4584
rect 2129 4526 12634 4528
rect 12801 4586 12867 4589
rect 18873 4586 18939 4589
rect 12801 4584 18939 4586
rect 12801 4528 12806 4584
rect 12862 4528 18878 4584
rect 18934 4528 18939 4584
rect 12801 4526 18939 4528
rect 2129 4523 2195 4526
rect 12801 4523 12867 4526
rect 18873 4523 18939 4526
rect 0 4450 480 4480
rect 2814 4450 2820 4452
rect 0 4390 2820 4450
rect 0 4360 480 4390
rect 2814 4388 2820 4390
rect 2884 4388 2890 4452
rect 5073 4450 5139 4453
rect 5625 4450 5691 4453
rect 5809 4452 5875 4453
rect 6177 4452 6243 4453
rect 5073 4448 5691 4450
rect 5073 4392 5078 4448
rect 5134 4392 5630 4448
rect 5686 4392 5691 4448
rect 5073 4390 5691 4392
rect 5073 4387 5139 4390
rect 5625 4387 5691 4390
rect 5758 4388 5764 4452
rect 5828 4450 5875 4452
rect 5828 4448 5920 4450
rect 5870 4392 5920 4448
rect 5828 4390 5920 4392
rect 5828 4388 5875 4390
rect 6126 4388 6132 4452
rect 6196 4450 6243 4452
rect 6453 4450 6519 4453
rect 6637 4450 6703 4453
rect 11053 4450 11119 4453
rect 12341 4450 12407 4453
rect 6196 4448 6288 4450
rect 6238 4392 6288 4448
rect 6196 4390 6288 4392
rect 6453 4448 11119 4450
rect 6453 4392 6458 4448
rect 6514 4392 6642 4448
rect 6698 4392 11058 4448
rect 11114 4392 11119 4448
rect 6453 4390 11119 4392
rect 6196 4388 6243 4390
rect 5809 4387 5875 4388
rect 6177 4387 6243 4388
rect 6453 4387 6519 4390
rect 6637 4387 6703 4390
rect 11053 4387 11119 4390
rect 12022 4448 12407 4450
rect 12022 4392 12346 4448
rect 12402 4392 12407 4448
rect 12022 4390 12407 4392
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 4797 4314 4863 4317
rect 5993 4314 6059 4317
rect 4797 4312 6059 4314
rect 4797 4256 4802 4312
rect 4858 4256 5998 4312
rect 6054 4256 6059 4312
rect 4797 4254 6059 4256
rect 4797 4251 4863 4254
rect 5993 4251 6059 4254
rect 6361 4314 6427 4317
rect 6729 4314 6795 4317
rect 6361 4312 6795 4314
rect 6361 4256 6366 4312
rect 6422 4256 6734 4312
rect 6790 4256 6795 4312
rect 6361 4254 6795 4256
rect 6361 4251 6427 4254
rect 6729 4251 6795 4254
rect 7741 4314 7807 4317
rect 8886 4314 8892 4316
rect 7741 4312 8892 4314
rect 7741 4256 7746 4312
rect 7802 4256 8892 4312
rect 7741 4254 8892 4256
rect 7741 4251 7807 4254
rect 8886 4252 8892 4254
rect 8956 4252 8962 4316
rect 9121 4314 9187 4317
rect 10593 4314 10659 4317
rect 9121 4312 10659 4314
rect 9121 4256 9126 4312
rect 9182 4256 10598 4312
rect 10654 4256 10659 4312
rect 9121 4254 10659 4256
rect 9121 4251 9187 4254
rect 10593 4251 10659 4254
rect 10777 4314 10843 4317
rect 11145 4314 11211 4317
rect 10777 4312 11211 4314
rect 10777 4256 10782 4312
rect 10838 4256 11150 4312
rect 11206 4256 11211 4312
rect 10777 4254 11211 4256
rect 10777 4251 10843 4254
rect 11145 4251 11211 4254
rect 2865 4178 2931 4181
rect 12022 4178 12082 4390
rect 12341 4387 12407 4390
rect 12617 4450 12683 4453
rect 16757 4450 16823 4453
rect 12617 4448 16823 4450
rect 12617 4392 12622 4448
rect 12678 4392 16762 4448
rect 16818 4392 16823 4448
rect 12617 4390 16823 4392
rect 12617 4387 12683 4390
rect 16757 4387 16823 4390
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 4319 18590 4320
rect 12157 4314 12223 4317
rect 14222 4314 14228 4316
rect 12157 4312 14228 4314
rect 12157 4256 12162 4312
rect 12218 4256 14228 4312
rect 12157 4254 14228 4256
rect 12157 4251 12223 4254
rect 14222 4252 14228 4254
rect 14292 4252 14298 4316
rect 14365 4312 14431 4317
rect 14365 4256 14370 4312
rect 14426 4256 14431 4312
rect 14365 4251 14431 4256
rect 14368 4178 14428 4251
rect 2865 4176 12082 4178
rect 2865 4120 2870 4176
rect 2926 4120 12082 4176
rect 2865 4118 12082 4120
rect 12528 4118 14428 4178
rect 2865 4115 2931 4118
rect 0 4042 480 4072
rect 4521 4042 4587 4045
rect 5574 4042 5580 4044
rect 0 3982 4354 4042
rect 0 3952 480 3982
rect 4294 3906 4354 3982
rect 4521 4040 5580 4042
rect 4521 3984 4526 4040
rect 4582 3984 5580 4040
rect 4521 3982 5580 3984
rect 4521 3979 4587 3982
rect 5574 3980 5580 3982
rect 5644 3980 5650 4044
rect 6637 4042 6703 4045
rect 8017 4042 8083 4045
rect 6637 4040 8083 4042
rect 6637 3984 6642 4040
rect 6698 3984 8022 4040
rect 8078 3984 8083 4040
rect 6637 3982 8083 3984
rect 6637 3979 6703 3982
rect 8017 3979 8083 3982
rect 8201 4042 8267 4045
rect 9397 4042 9463 4045
rect 8201 4040 9463 4042
rect 8201 3984 8206 4040
rect 8262 3984 9402 4040
rect 9458 3984 9463 4040
rect 8201 3982 9463 3984
rect 8201 3979 8267 3982
rect 9397 3979 9463 3982
rect 9673 4042 9739 4045
rect 12528 4042 12588 4118
rect 9673 4040 12588 4042
rect 9673 3984 9678 4040
rect 9734 3984 12588 4040
rect 9673 3982 12588 3984
rect 13905 4042 13971 4045
rect 19057 4042 19123 4045
rect 13905 4040 19123 4042
rect 13905 3984 13910 4040
rect 13966 3984 19062 4040
rect 19118 3984 19123 4040
rect 13905 3982 19123 3984
rect 9673 3979 9739 3982
rect 13905 3979 13971 3982
rect 19057 3979 19123 3982
rect 6862 3906 6868 3908
rect 4294 3846 6868 3906
rect 6862 3844 6868 3846
rect 6932 3844 6938 3908
rect 7281 3906 7347 3909
rect 7414 3906 7420 3908
rect 7281 3904 7420 3906
rect 7281 3848 7286 3904
rect 7342 3848 7420 3904
rect 7281 3846 7420 3848
rect 7281 3843 7347 3846
rect 7414 3844 7420 3846
rect 7484 3844 7490 3908
rect 8293 3904 8359 3909
rect 8293 3848 8298 3904
rect 8354 3848 8359 3904
rect 8293 3843 8359 3848
rect 8518 3844 8524 3908
rect 8588 3906 8594 3908
rect 12801 3906 12867 3909
rect 8588 3904 12867 3906
rect 8588 3848 12806 3904
rect 12862 3848 12867 3904
rect 8588 3846 12867 3848
rect 8588 3844 8594 3846
rect 12801 3843 12867 3846
rect 17677 3906 17743 3909
rect 22520 3906 23000 3936
rect 17677 3904 23000 3906
rect 17677 3848 17682 3904
rect 17738 3848 23000 3904
rect 17677 3846 23000 3848
rect 17677 3843 17743 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 4705 3770 4771 3773
rect 7598 3770 7604 3772
rect 4705 3768 7604 3770
rect 4705 3712 4710 3768
rect 4766 3712 7604 3768
rect 4705 3710 7604 3712
rect 4705 3707 4771 3710
rect 7598 3708 7604 3710
rect 7668 3708 7674 3772
rect 8296 3770 8356 3843
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 22520 3816 23000 3846
rect 14805 3775 15125 3776
rect 9397 3770 9463 3773
rect 8296 3768 9463 3770
rect 8296 3712 9402 3768
rect 9458 3712 9463 3768
rect 8296 3710 9463 3712
rect 9397 3707 9463 3710
rect 10358 3708 10364 3772
rect 10428 3770 10434 3772
rect 10869 3770 10935 3773
rect 10428 3768 10935 3770
rect 10428 3712 10874 3768
rect 10930 3712 10935 3768
rect 10428 3710 10935 3712
rect 10428 3708 10434 3710
rect 10869 3707 10935 3710
rect 11513 3770 11579 3773
rect 11830 3770 11836 3772
rect 11513 3768 11836 3770
rect 11513 3712 11518 3768
rect 11574 3712 11836 3768
rect 11513 3710 11836 3712
rect 11513 3707 11579 3710
rect 11830 3708 11836 3710
rect 11900 3708 11906 3772
rect 12249 3770 12315 3773
rect 12382 3770 12388 3772
rect 12249 3768 12388 3770
rect 12249 3712 12254 3768
rect 12310 3712 12388 3768
rect 12249 3710 12388 3712
rect 12249 3707 12315 3710
rect 12382 3708 12388 3710
rect 12452 3708 12458 3772
rect 12525 3770 12591 3773
rect 13118 3770 13124 3772
rect 12525 3768 13124 3770
rect 12525 3712 12530 3768
rect 12586 3712 13124 3768
rect 12525 3710 13124 3712
rect 12525 3707 12591 3710
rect 13118 3708 13124 3710
rect 13188 3708 13194 3772
rect 4429 3634 4495 3637
rect 5993 3634 6059 3637
rect 8017 3634 8083 3637
rect 4429 3632 5872 3634
rect 4429 3576 4434 3632
rect 4490 3576 5872 3632
rect 4429 3574 5872 3576
rect 4429 3571 4495 3574
rect 0 3498 480 3528
rect 5812 3501 5872 3574
rect 5993 3632 8083 3634
rect 5993 3576 5998 3632
rect 6054 3576 8022 3632
rect 8078 3576 8083 3632
rect 5993 3574 8083 3576
rect 5993 3571 6059 3574
rect 8017 3571 8083 3574
rect 8385 3634 8451 3637
rect 10501 3634 10567 3637
rect 8385 3632 10567 3634
rect 8385 3576 8390 3632
rect 8446 3576 10506 3632
rect 10562 3576 10567 3632
rect 8385 3574 10567 3576
rect 8385 3571 8451 3574
rect 10501 3571 10567 3574
rect 11094 3572 11100 3636
rect 11164 3634 11170 3636
rect 11329 3634 11395 3637
rect 11164 3632 11395 3634
rect 11164 3576 11334 3632
rect 11390 3576 11395 3632
rect 11164 3574 11395 3576
rect 11164 3572 11170 3574
rect 11329 3571 11395 3574
rect 11973 3634 12039 3637
rect 15694 3634 15700 3636
rect 11973 3632 15700 3634
rect 11973 3576 11978 3632
rect 12034 3576 15700 3632
rect 11973 3574 15700 3576
rect 11973 3571 12039 3574
rect 15694 3572 15700 3574
rect 15764 3572 15770 3636
rect 2313 3498 2379 3501
rect 2446 3498 2452 3500
rect 0 3496 2452 3498
rect 0 3440 2318 3496
rect 2374 3440 2452 3496
rect 0 3438 2452 3440
rect 0 3408 480 3438
rect 2313 3435 2379 3438
rect 2446 3436 2452 3438
rect 2516 3436 2522 3500
rect 2773 3498 2839 3501
rect 3182 3498 3188 3500
rect 2773 3496 3188 3498
rect 2773 3440 2778 3496
rect 2834 3440 3188 3496
rect 2773 3438 3188 3440
rect 2773 3435 2839 3438
rect 3182 3436 3188 3438
rect 3252 3436 3258 3500
rect 3325 3498 3391 3501
rect 5022 3498 5028 3500
rect 3325 3496 5028 3498
rect 3325 3440 3330 3496
rect 3386 3440 5028 3496
rect 3325 3438 5028 3440
rect 3325 3435 3391 3438
rect 5022 3436 5028 3438
rect 5092 3436 5098 3500
rect 5809 3498 5875 3501
rect 7649 3498 7715 3501
rect 5809 3496 7715 3498
rect 5809 3440 5814 3496
rect 5870 3440 7654 3496
rect 7710 3440 7715 3496
rect 5809 3438 7715 3440
rect 5809 3435 5875 3438
rect 7649 3435 7715 3438
rect 8293 3498 8359 3501
rect 19425 3498 19491 3501
rect 8293 3496 19491 3498
rect 8293 3440 8298 3496
rect 8354 3440 19430 3496
rect 19486 3440 19491 3496
rect 8293 3438 19491 3440
rect 8293 3435 8359 3438
rect 19425 3435 19491 3438
rect 6085 3362 6151 3365
rect 6678 3362 6684 3364
rect 6085 3360 6684 3362
rect 6085 3304 6090 3360
rect 6146 3304 6684 3360
rect 6085 3302 6684 3304
rect 6085 3299 6151 3302
rect 6678 3300 6684 3302
rect 6748 3300 6754 3364
rect 7373 3362 7439 3365
rect 8334 3362 8340 3364
rect 7373 3360 8340 3362
rect 7373 3304 7378 3360
rect 7434 3304 8340 3360
rect 7373 3302 8340 3304
rect 7373 3299 7439 3302
rect 8334 3300 8340 3302
rect 8404 3362 8410 3364
rect 9765 3362 9831 3365
rect 8404 3360 9831 3362
rect 8404 3304 9770 3360
rect 9826 3304 9831 3360
rect 8404 3302 9831 3304
rect 8404 3300 8410 3302
rect 9765 3299 9831 3302
rect 10041 3362 10107 3365
rect 11145 3362 11211 3365
rect 10041 3360 11211 3362
rect 10041 3304 10046 3360
rect 10102 3304 11150 3360
rect 11206 3304 11211 3360
rect 10041 3302 11211 3304
rect 10041 3299 10107 3302
rect 11145 3299 11211 3302
rect 12157 3362 12223 3365
rect 18045 3362 18111 3365
rect 12157 3360 18111 3362
rect 12157 3304 12162 3360
rect 12218 3304 18050 3360
rect 18106 3304 18111 3360
rect 12157 3302 18111 3304
rect 12157 3299 12223 3302
rect 18045 3299 18111 3302
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 5533 3226 5599 3229
rect 9489 3226 9555 3229
rect 10501 3228 10567 3229
rect 5533 3224 9555 3226
rect 5533 3168 5538 3224
rect 5594 3168 9494 3224
rect 9550 3168 9555 3224
rect 5533 3166 9555 3168
rect 5533 3163 5599 3166
rect 9489 3163 9555 3166
rect 9814 3166 10426 3226
rect 0 3090 480 3120
rect 1577 3090 1643 3093
rect 0 3088 1643 3090
rect 0 3032 1582 3088
rect 1638 3032 1643 3088
rect 0 3030 1643 3032
rect 0 3000 480 3030
rect 1577 3027 1643 3030
rect 2497 3090 2563 3093
rect 9814 3090 9874 3166
rect 2497 3088 9874 3090
rect 2497 3032 2502 3088
rect 2558 3032 9874 3088
rect 2497 3030 9874 3032
rect 10366 3090 10426 3166
rect 10501 3224 10548 3228
rect 10612 3226 10618 3228
rect 12341 3226 12407 3229
rect 12750 3226 12756 3228
rect 10501 3168 10506 3224
rect 10501 3164 10548 3168
rect 10612 3166 10658 3226
rect 11838 3166 12266 3226
rect 10612 3164 10618 3166
rect 10501 3163 10567 3164
rect 11838 3090 11898 3166
rect 10366 3030 11898 3090
rect 12206 3090 12266 3166
rect 12341 3224 12756 3226
rect 12341 3168 12346 3224
rect 12402 3168 12756 3224
rect 12341 3166 12756 3168
rect 12341 3163 12407 3166
rect 12750 3164 12756 3166
rect 12820 3164 12826 3228
rect 18689 3090 18755 3093
rect 12206 3088 18755 3090
rect 12206 3032 18694 3088
rect 18750 3032 18755 3088
rect 12206 3030 18755 3032
rect 2497 3027 2563 3030
rect 18689 3027 18755 3030
rect 2221 2954 2287 2957
rect 18137 2954 18203 2957
rect 2221 2952 18203 2954
rect 2221 2896 2226 2952
rect 2282 2896 18142 2952
rect 18198 2896 18203 2952
rect 2221 2894 18203 2896
rect 2221 2891 2287 2894
rect 18137 2891 18203 2894
rect 1526 2756 1532 2820
rect 1596 2818 1602 2820
rect 5533 2818 5599 2821
rect 6269 2820 6335 2821
rect 6269 2818 6316 2820
rect 1596 2816 5599 2818
rect 1596 2760 5538 2816
rect 5594 2760 5599 2816
rect 1596 2758 5599 2760
rect 6224 2816 6316 2818
rect 6224 2760 6274 2816
rect 6224 2758 6316 2760
rect 1596 2756 1602 2758
rect 5533 2755 5599 2758
rect 6269 2756 6316 2758
rect 6380 2756 6386 2820
rect 6678 2756 6684 2820
rect 6748 2818 6754 2820
rect 7465 2818 7531 2821
rect 6748 2816 7531 2818
rect 6748 2760 7470 2816
rect 7526 2760 7531 2816
rect 6748 2758 7531 2760
rect 6748 2756 6754 2758
rect 6269 2755 6335 2756
rect 7465 2755 7531 2758
rect 9581 2820 9647 2821
rect 9857 2820 9923 2821
rect 9581 2816 9628 2820
rect 9692 2818 9698 2820
rect 9581 2760 9586 2816
rect 9581 2756 9628 2760
rect 9692 2758 9738 2818
rect 9692 2756 9698 2758
rect 9806 2756 9812 2820
rect 9876 2818 9923 2820
rect 9876 2816 9968 2818
rect 9918 2760 9968 2816
rect 9876 2758 9968 2760
rect 9876 2756 9923 2758
rect 10174 2756 10180 2820
rect 10244 2818 10250 2820
rect 10409 2818 10475 2821
rect 10244 2816 10475 2818
rect 10244 2760 10414 2816
rect 10470 2760 10475 2816
rect 10244 2758 10475 2760
rect 10244 2756 10250 2758
rect 9581 2755 9647 2756
rect 9857 2755 9923 2756
rect 10409 2755 10475 2758
rect 10593 2818 10659 2821
rect 10726 2818 10732 2820
rect 10593 2816 10732 2818
rect 10593 2760 10598 2816
rect 10654 2760 10732 2816
rect 10593 2758 10732 2760
rect 10593 2755 10659 2758
rect 10726 2756 10732 2758
rect 10796 2756 10802 2820
rect 11053 2818 11119 2821
rect 12065 2818 12131 2821
rect 11053 2816 12131 2818
rect 11053 2760 11058 2816
rect 11114 2760 12070 2816
rect 12126 2760 12131 2816
rect 11053 2758 12131 2760
rect 11053 2755 11119 2758
rect 12065 2755 12131 2758
rect 15510 2756 15516 2820
rect 15580 2818 15586 2820
rect 21725 2818 21791 2821
rect 15580 2816 21791 2818
rect 15580 2760 21730 2816
rect 21786 2760 21791 2816
rect 15580 2758 21791 2760
rect 15580 2756 15586 2758
rect 21725 2755 21791 2758
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 4429 2682 4495 2685
rect 5942 2682 5948 2684
rect 4429 2680 5948 2682
rect 4429 2624 4434 2680
rect 4490 2624 5948 2680
rect 4429 2622 5948 2624
rect 4429 2619 4495 2622
rect 5942 2620 5948 2622
rect 6012 2620 6018 2684
rect 8886 2620 8892 2684
rect 8956 2682 8962 2684
rect 9029 2682 9095 2685
rect 8956 2680 9095 2682
rect 8956 2624 9034 2680
rect 9090 2624 9095 2680
rect 8956 2622 9095 2624
rect 8956 2620 8962 2622
rect 9029 2619 9095 2622
rect 9213 2682 9279 2685
rect 11053 2682 11119 2685
rect 9213 2680 11119 2682
rect 9213 2624 9218 2680
rect 9274 2624 11058 2680
rect 11114 2624 11119 2680
rect 9213 2622 11119 2624
rect 9213 2619 9279 2622
rect 11053 2619 11119 2622
rect 11513 2682 11579 2685
rect 14273 2682 14339 2685
rect 11513 2680 14339 2682
rect 11513 2624 11518 2680
rect 11574 2624 14278 2680
rect 14334 2624 14339 2680
rect 11513 2622 14339 2624
rect 11513 2619 11579 2622
rect 14273 2619 14339 2622
rect 0 2546 480 2576
rect 1025 2546 1091 2549
rect 0 2544 1091 2546
rect 0 2488 1030 2544
rect 1086 2488 1091 2544
rect 0 2486 1091 2488
rect 0 2456 480 2486
rect 1025 2483 1091 2486
rect 7046 2484 7052 2548
rect 7116 2546 7122 2548
rect 7649 2546 7715 2549
rect 7116 2544 7715 2546
rect 7116 2488 7654 2544
rect 7710 2488 7715 2544
rect 7116 2486 7715 2488
rect 7116 2484 7122 2486
rect 7649 2483 7715 2486
rect 8109 2546 8175 2549
rect 8702 2546 8708 2548
rect 8109 2544 8708 2546
rect 8109 2488 8114 2544
rect 8170 2488 8708 2544
rect 8109 2486 8708 2488
rect 8109 2483 8175 2486
rect 8702 2484 8708 2486
rect 8772 2484 8778 2548
rect 9438 2484 9444 2548
rect 9508 2546 9514 2548
rect 10777 2546 10843 2549
rect 9508 2544 10843 2546
rect 9508 2488 10782 2544
rect 10838 2488 10843 2544
rect 9508 2486 10843 2488
rect 9508 2484 9514 2486
rect 10777 2483 10843 2486
rect 10910 2484 10916 2548
rect 10980 2546 10986 2548
rect 11881 2546 11947 2549
rect 10980 2544 11947 2546
rect 10980 2488 11886 2544
rect 11942 2488 11947 2544
rect 10980 2486 11947 2488
rect 10980 2484 10986 2486
rect 11881 2483 11947 2486
rect 2129 2410 2195 2413
rect 5993 2410 6059 2413
rect 2129 2408 6059 2410
rect 2129 2352 2134 2408
rect 2190 2352 5998 2408
rect 6054 2352 6059 2408
rect 2129 2350 6059 2352
rect 2129 2347 2195 2350
rect 5993 2347 6059 2350
rect 6361 2410 6427 2413
rect 12249 2410 12315 2413
rect 6361 2408 12315 2410
rect 6361 2352 6366 2408
rect 6422 2352 12254 2408
rect 12310 2352 12315 2408
rect 6361 2350 12315 2352
rect 6361 2347 6427 2350
rect 12249 2347 12315 2350
rect 5257 2274 5323 2277
rect 9397 2274 9463 2277
rect 10041 2276 10107 2277
rect 5257 2272 9463 2274
rect 5257 2216 5262 2272
rect 5318 2216 9402 2272
rect 9458 2216 9463 2272
rect 5257 2214 9463 2216
rect 5257 2211 5323 2214
rect 9397 2211 9463 2214
rect 9990 2212 9996 2276
rect 10060 2274 10107 2276
rect 10060 2272 10152 2274
rect 10102 2216 10152 2272
rect 10060 2214 10152 2216
rect 10060 2212 10107 2214
rect 10041 2211 10107 2212
rect 4409 2208 4729 2209
rect 0 2138 480 2168
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 4245 2138 4311 2141
rect 10685 2138 10751 2141
rect 0 2136 4311 2138
rect 0 2080 4250 2136
rect 4306 2080 4311 2136
rect 0 2078 4311 2080
rect 0 2048 480 2078
rect 4245 2075 4311 2078
rect 4800 2136 10751 2138
rect 4800 2080 10690 2136
rect 10746 2080 10751 2136
rect 4800 2078 10751 2080
rect 3601 2002 3667 2005
rect 4800 2002 4860 2078
rect 10685 2075 10751 2078
rect 3601 2000 4860 2002
rect 3601 1944 3606 2000
rect 3662 1944 4860 2000
rect 3601 1942 4860 1944
rect 6177 2002 6243 2005
rect 8661 2002 8727 2005
rect 6177 2000 8727 2002
rect 6177 1944 6182 2000
rect 6238 1944 8666 2000
rect 8722 1944 8727 2000
rect 6177 1942 8727 1944
rect 3601 1939 3667 1942
rect 6177 1939 6243 1942
rect 8661 1939 8727 1942
rect 8886 1940 8892 2004
rect 8956 2002 8962 2004
rect 9029 2002 9095 2005
rect 8956 2000 9095 2002
rect 8956 1944 9034 2000
rect 9090 1944 9095 2000
rect 8956 1942 9095 1944
rect 8956 1940 8962 1942
rect 9029 1939 9095 1942
rect 9213 2002 9279 2005
rect 14181 2002 14247 2005
rect 9213 2000 14247 2002
rect 9213 1944 9218 2000
rect 9274 1944 14186 2000
rect 14242 1944 14247 2000
rect 9213 1942 14247 1944
rect 9213 1939 9279 1942
rect 14181 1939 14247 1942
rect 3366 1804 3372 1868
rect 3436 1866 3442 1868
rect 15469 1866 15535 1869
rect 3436 1864 15535 1866
rect 3436 1808 15474 1864
rect 15530 1808 15535 1864
rect 3436 1806 15535 1808
rect 3436 1804 3442 1806
rect 15469 1803 15535 1806
rect 2262 1668 2268 1732
rect 2332 1730 2338 1732
rect 5809 1730 5875 1733
rect 2332 1728 5875 1730
rect 2332 1672 5814 1728
rect 5870 1672 5875 1728
rect 2332 1670 5875 1672
rect 2332 1668 2338 1670
rect 5809 1667 5875 1670
rect 6729 1730 6795 1733
rect 8293 1730 8359 1733
rect 17769 1730 17835 1733
rect 6729 1728 7804 1730
rect 6729 1672 6734 1728
rect 6790 1672 7804 1728
rect 6729 1670 7804 1672
rect 6729 1667 6795 1670
rect 0 1594 480 1624
rect 5206 1594 5212 1596
rect 0 1534 5212 1594
rect 0 1504 480 1534
rect 5206 1532 5212 1534
rect 5276 1532 5282 1596
rect 7465 1594 7531 1597
rect 7054 1592 7531 1594
rect 7054 1536 7470 1592
rect 7526 1536 7531 1592
rect 7054 1534 7531 1536
rect 2497 1458 2563 1461
rect 7054 1458 7114 1534
rect 7465 1531 7531 1534
rect 2497 1456 7114 1458
rect 2497 1400 2502 1456
rect 2558 1400 7114 1456
rect 2497 1398 7114 1400
rect 7189 1458 7255 1461
rect 7598 1458 7604 1460
rect 7189 1456 7604 1458
rect 7189 1400 7194 1456
rect 7250 1400 7604 1456
rect 7189 1398 7604 1400
rect 2497 1395 2563 1398
rect 7189 1395 7255 1398
rect 7598 1396 7604 1398
rect 7668 1396 7674 1460
rect 7744 1458 7804 1670
rect 8293 1728 17835 1730
rect 8293 1672 8298 1728
rect 8354 1672 17774 1728
rect 17830 1672 17835 1728
rect 8293 1670 17835 1672
rect 8293 1667 8359 1670
rect 17769 1667 17835 1670
rect 8017 1594 8083 1597
rect 8477 1594 8543 1597
rect 8017 1592 8543 1594
rect 8017 1536 8022 1592
rect 8078 1536 8482 1592
rect 8538 1536 8543 1592
rect 8017 1534 8543 1536
rect 8017 1531 8083 1534
rect 8477 1531 8543 1534
rect 8661 1594 8727 1597
rect 12934 1594 12940 1596
rect 8661 1592 12940 1594
rect 8661 1536 8666 1592
rect 8722 1536 12940 1592
rect 8661 1534 12940 1536
rect 8661 1531 8727 1534
rect 12934 1532 12940 1534
rect 13004 1532 13010 1596
rect 9070 1458 9076 1460
rect 7744 1398 9076 1458
rect 9070 1396 9076 1398
rect 9140 1458 9146 1460
rect 12341 1458 12407 1461
rect 9140 1456 12407 1458
rect 9140 1400 12346 1456
rect 12402 1400 12407 1456
rect 9140 1398 12407 1400
rect 9140 1396 9146 1398
rect 12341 1395 12407 1398
rect 0 1186 480 1216
rect 3049 1186 3115 1189
rect 0 1184 3115 1186
rect 0 1128 3054 1184
rect 3110 1128 3115 1184
rect 0 1126 3115 1128
rect 0 1096 480 1126
rect 3049 1123 3115 1126
rect 0 642 480 672
rect 2405 642 2471 645
rect 0 640 2471 642
rect 0 584 2410 640
rect 2466 584 2471 640
rect 0 582 2471 584
rect 0 552 480 582
rect 2405 579 2471 582
rect 0 234 480 264
rect 3734 234 3740 236
rect 0 174 3740 234
rect 0 144 480 174
rect 3734 172 3740 174
rect 3804 172 3810 236
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 9812 19756 9876 19820
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 8524 19408 8588 19412
rect 8524 19352 8538 19408
rect 8538 19352 8588 19408
rect 8524 19348 8588 19352
rect 5028 19212 5092 19276
rect 5580 19212 5644 19276
rect 12020 19076 12084 19140
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 12204 18864 12268 18868
rect 12204 18808 12254 18864
rect 12254 18808 12268 18864
rect 12204 18804 12268 18808
rect 13492 18804 13556 18868
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7052 18396 7116 18460
rect 6500 18260 6564 18324
rect 4108 18124 4172 18188
rect 5580 18124 5644 18188
rect 1532 18048 1596 18052
rect 1532 17992 1546 18048
rect 1546 17992 1596 18048
rect 1532 17988 1596 17992
rect 5028 17988 5092 18052
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 12388 17640 12452 17644
rect 12388 17584 12402 17640
rect 12402 17584 12452 17640
rect 12388 17580 12452 17584
rect 14044 17640 14108 17644
rect 14044 17584 14058 17640
rect 14058 17584 14108 17640
rect 14044 17580 14108 17584
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 10180 17308 10244 17372
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 8340 16764 8404 16828
rect 19196 16900 19260 16964
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 8892 16492 8956 16556
rect 12572 16492 12636 16556
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7604 16008 7668 16012
rect 7604 15952 7654 16008
rect 7654 15952 7668 16008
rect 7604 15948 7668 15952
rect 13860 15872 13924 15876
rect 13860 15816 13910 15872
rect 13910 15816 13924 15872
rect 13860 15812 13924 15816
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 9996 15600 10060 15604
rect 9996 15544 10046 15600
rect 10046 15544 10060 15600
rect 9996 15540 10060 15544
rect 15700 15540 15764 15604
rect 5764 15404 5828 15468
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 6132 15132 6196 15196
rect 13860 15132 13924 15196
rect 19196 14996 19260 15060
rect 2636 14724 2700 14788
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 2084 14316 2148 14380
rect 3188 14240 3252 14244
rect 3188 14184 3202 14240
rect 3202 14184 3252 14240
rect 3188 14180 3252 14184
rect 3740 14180 3804 14244
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 4844 13908 4908 13972
rect 4108 13636 4172 13700
rect 5396 13636 5460 13700
rect 9628 13636 9692 13700
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 6316 13364 6380 13428
rect 12020 13364 12084 13428
rect 12204 13364 12268 13428
rect 13492 13560 13556 13564
rect 13492 13504 13542 13560
rect 13542 13504 13556 13560
rect 13492 13500 13556 13504
rect 3556 13092 3620 13156
rect 4844 13228 4908 13292
rect 10364 13092 10428 13156
rect 14044 13092 14108 13156
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 14228 12820 14292 12884
rect 8892 12744 8956 12748
rect 8892 12688 8906 12744
rect 8906 12688 8956 12744
rect 8892 12684 8956 12688
rect 11836 12548 11900 12612
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4844 12412 4908 12476
rect 8340 12472 8404 12476
rect 8340 12416 8354 12472
rect 8354 12416 8404 12472
rect 8340 12412 8404 12416
rect 12020 12472 12084 12476
rect 12020 12416 12034 12472
rect 12034 12416 12084 12472
rect 12020 12412 12084 12416
rect 19196 12472 19260 12476
rect 19196 12416 19246 12472
rect 19246 12416 19260 12472
rect 19196 12412 19260 12416
rect 2820 12336 2884 12340
rect 2820 12280 2834 12336
rect 2834 12280 2884 12336
rect 2820 12276 2884 12280
rect 4108 12276 4172 12340
rect 6868 12276 6932 12340
rect 12756 12276 12820 12340
rect 14228 12200 14292 12204
rect 14228 12144 14242 12200
rect 14242 12144 14292 12200
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 14228 12140 14292 12144
rect 5212 12004 5276 12068
rect 7052 12064 7116 12068
rect 7052 12008 7066 12064
rect 7066 12008 7116 12064
rect 7052 12004 7116 12008
rect 7236 12004 7300 12068
rect 8340 11732 8404 11796
rect 7420 11596 7484 11660
rect 2820 11460 2884 11524
rect 13860 12004 13924 12068
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 13492 11868 13556 11932
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 9444 11324 9508 11388
rect 5028 11188 5092 11252
rect 6684 11188 6748 11252
rect 5028 11052 5092 11116
rect 12572 10916 12636 10980
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 12572 10780 12636 10844
rect 7052 10372 7116 10436
rect 8708 10372 8772 10436
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 2268 10236 2332 10300
rect 3924 10236 3988 10300
rect 15700 10236 15764 10300
rect 12204 10100 12268 10164
rect 12388 9964 12452 10028
rect 6132 9828 6196 9892
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 5948 9692 6012 9756
rect 7420 9692 7484 9756
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 2084 9420 2148 9484
rect 3188 9420 3252 9484
rect 6132 9284 6196 9348
rect 9076 9420 9140 9484
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 2452 9148 2516 9212
rect 9444 9148 9508 9212
rect 9628 9148 9692 9212
rect 3188 8740 3252 8804
rect 4108 8800 4172 8804
rect 4108 8744 4158 8800
rect 4158 8744 4172 8800
rect 4108 8740 4172 8744
rect 10364 8740 10428 8804
rect 14228 8740 14292 8804
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 4108 8604 4172 8668
rect 5764 8664 5828 8668
rect 5764 8608 5814 8664
rect 5814 8608 5828 8664
rect 5764 8604 5828 8608
rect 8708 8604 8772 8668
rect 10916 8604 10980 8668
rect 11100 8664 11164 8668
rect 11100 8608 11114 8664
rect 11114 8608 11164 8664
rect 11100 8604 11164 8608
rect 2636 8392 2700 8396
rect 7420 8468 7484 8532
rect 2636 8336 2650 8392
rect 2650 8336 2700 8392
rect 2636 8332 2700 8336
rect 5764 8196 5828 8260
rect 10548 8332 10612 8396
rect 12020 8196 12084 8260
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 8892 7924 8956 7988
rect 13124 7924 13188 7988
rect 4844 7788 4908 7852
rect 8340 7788 8404 7852
rect 3188 7652 3252 7716
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 10732 7516 10796 7580
rect 5212 7380 5276 7444
rect 10916 7440 10980 7444
rect 12940 7652 13004 7716
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 10916 7384 10966 7440
rect 10966 7384 10980 7440
rect 10916 7380 10980 7384
rect 11836 7380 11900 7444
rect 3372 6972 3436 7036
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 5764 6972 5828 7036
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4108 6836 4172 6900
rect 5212 6836 5276 6900
rect 9260 6896 9324 6900
rect 10916 6972 10980 7036
rect 12388 6972 12452 7036
rect 9260 6840 9310 6896
rect 9310 6840 9324 6896
rect 9260 6836 9324 6840
rect 4108 6564 4172 6628
rect 10732 6564 10796 6628
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 5212 6428 5276 6492
rect 6316 6488 6380 6492
rect 6316 6432 6330 6488
rect 6330 6432 6380 6488
rect 6316 6428 6380 6432
rect 6684 6428 6748 6492
rect 7052 6428 7116 6492
rect 5212 6292 5276 6356
rect 7052 6020 7116 6084
rect 9444 6020 9508 6084
rect 10732 6080 10796 6084
rect 10732 6024 10746 6080
rect 10746 6024 10796 6080
rect 10732 6020 10796 6024
rect 11836 6020 11900 6084
rect 12204 6020 12268 6084
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 3924 5476 3988 5540
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 6316 5476 6380 5540
rect 15516 5476 15580 5540
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 12204 5340 12268 5404
rect 15700 5340 15764 5404
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 4108 5204 4172 5268
rect 5948 5204 6012 5268
rect 6868 5204 6932 5268
rect 8340 5204 8404 5268
rect 12572 5204 12636 5268
rect 6132 4932 6196 4996
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 3556 4796 3620 4860
rect 6500 4796 6564 4860
rect 5396 4660 5460 4724
rect 12204 4660 12268 4724
rect 2820 4388 2884 4452
rect 5764 4448 5828 4452
rect 5764 4392 5814 4448
rect 5814 4392 5828 4448
rect 5764 4388 5828 4392
rect 6132 4448 6196 4452
rect 6132 4392 6182 4448
rect 6182 4392 6196 4448
rect 6132 4388 6196 4392
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 8892 4252 8956 4316
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 14228 4252 14292 4316
rect 5580 3980 5644 4044
rect 6868 3844 6932 3908
rect 7420 3844 7484 3908
rect 8524 3844 8588 3908
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 7604 3708 7668 3772
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 10364 3708 10428 3772
rect 11836 3708 11900 3772
rect 12388 3708 12452 3772
rect 13124 3708 13188 3772
rect 11100 3572 11164 3636
rect 15700 3572 15764 3636
rect 2452 3436 2516 3500
rect 3188 3436 3252 3500
rect 5028 3436 5092 3500
rect 6684 3300 6748 3364
rect 8340 3300 8404 3364
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 10548 3224 10612 3228
rect 10548 3168 10562 3224
rect 10562 3168 10612 3224
rect 10548 3164 10612 3168
rect 12756 3164 12820 3228
rect 1532 2756 1596 2820
rect 6316 2816 6380 2820
rect 6316 2760 6330 2816
rect 6330 2760 6380 2816
rect 6316 2756 6380 2760
rect 6684 2756 6748 2820
rect 9628 2816 9692 2820
rect 9628 2760 9642 2816
rect 9642 2760 9692 2816
rect 9628 2756 9692 2760
rect 9812 2816 9876 2820
rect 9812 2760 9862 2816
rect 9862 2760 9876 2816
rect 9812 2756 9876 2760
rect 10180 2756 10244 2820
rect 10732 2756 10796 2820
rect 15516 2756 15580 2820
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 5948 2620 6012 2684
rect 8892 2620 8956 2684
rect 7052 2484 7116 2548
rect 8708 2484 8772 2548
rect 9444 2484 9508 2548
rect 10916 2484 10980 2548
rect 9996 2272 10060 2276
rect 9996 2216 10046 2272
rect 10046 2216 10060 2272
rect 9996 2212 10060 2216
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
rect 8892 1940 8956 2004
rect 3372 1804 3436 1868
rect 2268 1668 2332 1732
rect 5212 1532 5276 1596
rect 7604 1396 7668 1460
rect 12940 1532 13004 1596
rect 9076 1396 9140 1460
rect 3740 172 3804 236
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 5027 19276 5093 19277
rect 5027 19212 5028 19276
rect 5092 19212 5093 19276
rect 5027 19211 5093 19212
rect 5579 19276 5645 19277
rect 5579 19212 5580 19276
rect 5644 19212 5645 19276
rect 5579 19211 5645 19212
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4107 18188 4173 18189
rect 4107 18124 4108 18188
rect 4172 18124 4173 18188
rect 4107 18123 4173 18124
rect 1531 18052 1597 18053
rect 1531 17988 1532 18052
rect 1596 17988 1597 18052
rect 1531 17987 1597 17988
rect 1534 2821 1594 17987
rect 2635 14788 2701 14789
rect 2635 14724 2636 14788
rect 2700 14724 2701 14788
rect 2635 14723 2701 14724
rect 2083 14380 2149 14381
rect 2083 14316 2084 14380
rect 2148 14316 2149 14380
rect 2083 14315 2149 14316
rect 2086 9485 2146 14315
rect 2267 10300 2333 10301
rect 2267 10236 2268 10300
rect 2332 10236 2333 10300
rect 2267 10235 2333 10236
rect 2083 9484 2149 9485
rect 2083 9420 2084 9484
rect 2148 9420 2149 9484
rect 2083 9419 2149 9420
rect 1531 2820 1597 2821
rect 1531 2756 1532 2820
rect 1596 2756 1597 2820
rect 1531 2755 1597 2756
rect 2270 1733 2330 10235
rect 2451 9212 2517 9213
rect 2451 9148 2452 9212
rect 2516 9148 2517 9212
rect 2451 9147 2517 9148
rect 2454 3501 2514 9147
rect 2638 8397 2698 14723
rect 3187 14244 3253 14245
rect 3187 14180 3188 14244
rect 3252 14180 3253 14244
rect 3187 14179 3253 14180
rect 3739 14244 3805 14245
rect 3739 14180 3740 14244
rect 3804 14180 3805 14244
rect 3739 14179 3805 14180
rect 2819 12340 2885 12341
rect 2819 12276 2820 12340
rect 2884 12276 2885 12340
rect 2819 12275 2885 12276
rect 2822 11525 2882 12275
rect 2819 11524 2885 11525
rect 2819 11460 2820 11524
rect 2884 11460 2885 11524
rect 2819 11459 2885 11460
rect 2635 8396 2701 8397
rect 2635 8332 2636 8396
rect 2700 8332 2701 8396
rect 2635 8331 2701 8332
rect 2822 4453 2882 11459
rect 3190 9485 3250 14179
rect 3555 13156 3621 13157
rect 3555 13092 3556 13156
rect 3620 13092 3621 13156
rect 3555 13091 3621 13092
rect 3187 9484 3253 9485
rect 3187 9420 3188 9484
rect 3252 9420 3253 9484
rect 3187 9419 3253 9420
rect 3190 8805 3250 9062
rect 3187 8804 3253 8805
rect 3187 8740 3188 8804
rect 3252 8740 3253 8804
rect 3187 8739 3253 8740
rect 3187 7716 3253 7717
rect 3187 7652 3188 7716
rect 3252 7652 3253 7716
rect 3187 7651 3253 7652
rect 2819 4452 2885 4453
rect 2819 4388 2820 4452
rect 2884 4388 2885 4452
rect 2819 4387 2885 4388
rect 3190 3501 3250 7651
rect 3371 7036 3437 7037
rect 3371 6972 3372 7036
rect 3436 6972 3437 7036
rect 3371 6971 3437 6972
rect 2451 3500 2517 3501
rect 2451 3436 2452 3500
rect 2516 3436 2517 3500
rect 2451 3435 2517 3436
rect 3187 3500 3253 3501
rect 3187 3436 3188 3500
rect 3252 3436 3253 3500
rect 3187 3435 3253 3436
rect 3374 1869 3434 6971
rect 3558 4861 3618 13091
rect 3555 4860 3621 4861
rect 3555 4796 3556 4860
rect 3620 4796 3621 4860
rect 3555 4795 3621 4796
rect 3371 1868 3437 1869
rect 3371 1804 3372 1868
rect 3436 1804 3437 1868
rect 3371 1803 3437 1804
rect 2267 1732 2333 1733
rect 2267 1668 2268 1732
rect 2332 1668 2333 1732
rect 2267 1667 2333 1668
rect 3742 237 3802 14179
rect 4110 13701 4170 18123
rect 4409 17440 4729 18464
rect 5030 18053 5090 19211
rect 5582 18189 5642 19211
rect 7874 19072 8195 20096
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 9811 19820 9877 19821
rect 9811 19756 9812 19820
rect 9876 19756 9877 19820
rect 9811 19755 9877 19756
rect 8523 19412 8589 19413
rect 8523 19348 8524 19412
rect 8588 19348 8589 19412
rect 8523 19347 8589 19348
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7051 18460 7117 18461
rect 7051 18396 7052 18460
rect 7116 18396 7117 18460
rect 7051 18395 7117 18396
rect 6499 18324 6565 18325
rect 6499 18260 6500 18324
rect 6564 18260 6565 18324
rect 6499 18259 6565 18260
rect 5579 18188 5645 18189
rect 5579 18124 5580 18188
rect 5644 18124 5645 18188
rect 5579 18123 5645 18124
rect 5027 18052 5093 18053
rect 5027 17988 5028 18052
rect 5092 17988 5093 18052
rect 5027 17987 5093 17988
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4107 13700 4173 13701
rect 4107 13636 4108 13700
rect 4172 13636 4173 13700
rect 4107 13635 4173 13636
rect 4409 13088 4729 14112
rect 4843 13972 4909 13973
rect 4843 13908 4844 13972
rect 4908 13908 4909 13972
rect 4843 13907 4909 13908
rect 4846 13293 4906 13907
rect 4843 13292 4909 13293
rect 4843 13228 4844 13292
rect 4908 13228 4909 13292
rect 4843 13227 4909 13228
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4107 12340 4173 12341
rect 4107 12276 4108 12340
rect 4172 12276 4173 12340
rect 4107 12275 4173 12276
rect 3923 10300 3989 10301
rect 3923 10236 3924 10300
rect 3988 10236 3989 10300
rect 3923 10235 3989 10236
rect 3926 5541 3986 10235
rect 4110 8805 4170 12275
rect 4409 12000 4729 13024
rect 4843 12476 4909 12477
rect 4843 12412 4844 12476
rect 4908 12412 4909 12476
rect 4843 12411 4909 12412
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4107 8804 4173 8805
rect 4107 8740 4108 8804
rect 4172 8740 4173 8804
rect 4107 8739 4173 8740
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4107 8668 4173 8669
rect 4107 8604 4108 8668
rect 4172 8604 4173 8668
rect 4107 8603 4173 8604
rect 4110 6901 4170 8603
rect 4409 7648 4729 8672
rect 4846 7853 4906 12411
rect 5030 11253 5090 17987
rect 5395 13700 5461 13701
rect 5395 13636 5396 13700
rect 5460 13636 5461 13700
rect 5395 13635 5461 13636
rect 5211 12068 5277 12069
rect 5211 12004 5212 12068
rect 5276 12004 5277 12068
rect 5211 12003 5277 12004
rect 5027 11252 5093 11253
rect 5027 11188 5028 11252
rect 5092 11188 5093 11252
rect 5027 11187 5093 11188
rect 5027 11116 5093 11117
rect 5027 11052 5028 11116
rect 5092 11052 5093 11116
rect 5027 11051 5093 11052
rect 4843 7852 4909 7853
rect 4843 7788 4844 7852
rect 4908 7788 4909 7852
rect 4843 7787 4909 7788
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4107 6900 4173 6901
rect 4107 6836 4108 6900
rect 4172 6836 4173 6900
rect 4107 6835 4173 6836
rect 4107 6628 4173 6629
rect 4107 6564 4108 6628
rect 4172 6564 4173 6628
rect 4107 6563 4173 6564
rect 3923 5540 3989 5541
rect 3923 5476 3924 5540
rect 3988 5476 3989 5540
rect 3923 5475 3989 5476
rect 4110 5269 4170 6563
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4107 5268 4173 5269
rect 4107 5204 4108 5268
rect 4172 5204 4173 5268
rect 4107 5203 4173 5204
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 5030 3501 5090 11051
rect 5214 7445 5274 12003
rect 5211 7444 5277 7445
rect 5211 7380 5212 7444
rect 5276 7380 5277 7444
rect 5211 7379 5277 7380
rect 5211 6900 5277 6901
rect 5211 6836 5212 6900
rect 5276 6836 5277 6900
rect 5211 6835 5277 6836
rect 5214 6493 5274 6835
rect 5211 6492 5277 6493
rect 5211 6428 5212 6492
rect 5276 6428 5277 6492
rect 5211 6427 5277 6428
rect 5211 6356 5277 6357
rect 5211 6292 5212 6356
rect 5276 6292 5277 6356
rect 5211 6291 5277 6292
rect 5027 3500 5093 3501
rect 5027 3436 5028 3500
rect 5092 3436 5093 3500
rect 5027 3435 5093 3436
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 5214 1597 5274 6291
rect 5398 4725 5458 13635
rect 5395 4724 5461 4725
rect 5395 4660 5396 4724
rect 5460 4660 5461 4724
rect 5395 4659 5461 4660
rect 5582 4045 5642 18123
rect 5763 15468 5829 15469
rect 5763 15404 5764 15468
rect 5828 15404 5829 15468
rect 5763 15403 5829 15404
rect 5766 8669 5826 15403
rect 6131 15196 6197 15197
rect 6131 15132 6132 15196
rect 6196 15132 6197 15196
rect 6131 15131 6197 15132
rect 6134 9893 6194 15131
rect 6315 13428 6381 13429
rect 6315 13364 6316 13428
rect 6380 13364 6381 13428
rect 6315 13363 6381 13364
rect 6131 9892 6197 9893
rect 6131 9828 6132 9892
rect 6196 9828 6197 9892
rect 6131 9827 6197 9828
rect 5947 9756 6013 9757
rect 5947 9692 5948 9756
rect 6012 9692 6013 9756
rect 5947 9691 6013 9692
rect 5763 8668 5829 8669
rect 5763 8604 5764 8668
rect 5828 8604 5829 8668
rect 5763 8603 5829 8604
rect 5763 8260 5829 8261
rect 5763 8196 5764 8260
rect 5828 8196 5829 8260
rect 5763 8195 5829 8196
rect 5766 7037 5826 8195
rect 5763 7036 5829 7037
rect 5763 6972 5764 7036
rect 5828 6972 5829 7036
rect 5763 6971 5829 6972
rect 5766 4453 5826 6971
rect 5950 5269 6010 9691
rect 6131 9348 6197 9349
rect 6131 9284 6132 9348
rect 6196 9284 6197 9348
rect 6131 9283 6197 9284
rect 5947 5268 6013 5269
rect 5947 5204 5948 5268
rect 6012 5204 6013 5268
rect 5947 5203 6013 5204
rect 5763 4452 5829 4453
rect 5763 4388 5764 4452
rect 5828 4388 5829 4452
rect 5763 4387 5829 4388
rect 5579 4044 5645 4045
rect 5579 3980 5580 4044
rect 5644 3980 5645 4044
rect 5579 3979 5645 3980
rect 5950 2685 6010 5203
rect 6134 4997 6194 9283
rect 6318 6493 6378 13363
rect 6315 6492 6381 6493
rect 6315 6428 6316 6492
rect 6380 6428 6381 6492
rect 6315 6427 6381 6428
rect 6315 5540 6381 5541
rect 6315 5476 6316 5540
rect 6380 5476 6381 5540
rect 6315 5475 6381 5476
rect 6131 4996 6197 4997
rect 6131 4932 6132 4996
rect 6196 4932 6197 4996
rect 6131 4931 6197 4932
rect 6134 4453 6194 4931
rect 6131 4452 6197 4453
rect 6131 4388 6132 4452
rect 6196 4388 6197 4452
rect 6131 4387 6197 4388
rect 6318 2821 6378 5475
rect 6502 4861 6562 18259
rect 6867 12340 6933 12341
rect 6867 12276 6868 12340
rect 6932 12276 6933 12340
rect 6867 12275 6933 12276
rect 6683 11252 6749 11253
rect 6683 11188 6684 11252
rect 6748 11188 6749 11252
rect 6683 11187 6749 11188
rect 6686 6493 6746 11187
rect 6683 6492 6749 6493
rect 6683 6428 6684 6492
rect 6748 6428 6749 6492
rect 6683 6427 6749 6428
rect 6870 5269 6930 12275
rect 7054 12069 7114 18395
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7603 16012 7669 16013
rect 7603 15948 7604 16012
rect 7668 15948 7669 16012
rect 7603 15947 7669 15948
rect 7051 12068 7117 12069
rect 7051 12004 7052 12068
rect 7116 12004 7117 12068
rect 7051 12003 7117 12004
rect 7235 12068 7301 12069
rect 7235 12004 7236 12068
rect 7300 12004 7301 12068
rect 7235 12003 7301 12004
rect 7051 10436 7117 10437
rect 7051 10372 7052 10436
rect 7116 10372 7117 10436
rect 7051 10371 7117 10372
rect 7054 6493 7114 10371
rect 7051 6492 7117 6493
rect 7051 6428 7052 6492
rect 7116 6428 7117 6492
rect 7051 6427 7117 6428
rect 7051 6084 7117 6085
rect 7051 6020 7052 6084
rect 7116 6020 7117 6084
rect 7051 6019 7117 6020
rect 6867 5268 6933 5269
rect 6867 5204 6868 5268
rect 6932 5204 6933 5268
rect 6867 5203 6933 5204
rect 6499 4860 6565 4861
rect 6499 4796 6500 4860
rect 6564 4796 6565 4860
rect 6499 4795 6565 4796
rect 6870 3909 6930 5203
rect 6867 3908 6933 3909
rect 6867 3844 6868 3908
rect 6932 3844 6933 3908
rect 6867 3843 6933 3844
rect 6683 3364 6749 3365
rect 6683 3300 6684 3364
rect 6748 3300 6749 3364
rect 6683 3299 6749 3300
rect 6686 2821 6746 3299
rect 6315 2820 6381 2821
rect 6315 2756 6316 2820
rect 6380 2756 6381 2820
rect 6315 2755 6381 2756
rect 6683 2820 6749 2821
rect 6683 2756 6684 2820
rect 6748 2756 6749 2820
rect 6683 2755 6749 2756
rect 5947 2684 6013 2685
rect 5947 2620 5948 2684
rect 6012 2620 6013 2684
rect 5947 2619 6013 2620
rect 7054 2549 7114 6019
rect 7238 3226 7298 12003
rect 7419 11660 7485 11661
rect 7419 11596 7420 11660
rect 7484 11596 7485 11660
rect 7419 11595 7485 11596
rect 7422 9757 7482 11595
rect 7419 9756 7485 9757
rect 7419 9692 7420 9756
rect 7484 9692 7485 9756
rect 7419 9691 7485 9692
rect 7419 8532 7485 8533
rect 7419 8468 7420 8532
rect 7484 8468 7485 8532
rect 7419 8467 7485 8468
rect 7422 3909 7482 8467
rect 7419 3908 7485 3909
rect 7419 3844 7420 3908
rect 7484 3844 7485 3908
rect 7419 3843 7485 3844
rect 7606 3773 7666 15947
rect 7874 15808 8195 16832
rect 8339 16828 8405 16829
rect 8339 16764 8340 16828
rect 8404 16764 8405 16828
rect 8339 16763 8405 16764
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 8342 12477 8402 16763
rect 8339 12476 8405 12477
rect 8339 12412 8340 12476
rect 8404 12412 8405 12476
rect 8339 12411 8405 12412
rect 8339 11796 8405 11797
rect 8339 11732 8340 11796
rect 8404 11732 8405 11796
rect 8339 11731 8405 11732
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 8342 7853 8402 11731
rect 8339 7852 8405 7853
rect 8339 7788 8340 7852
rect 8404 7788 8405 7852
rect 8339 7787 8405 7788
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 8339 5268 8405 5269
rect 8339 5204 8340 5268
rect 8404 5204 8405 5268
rect 8339 5203 8405 5204
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7603 3772 7669 3773
rect 7603 3708 7604 3772
rect 7668 3708 7669 3772
rect 7603 3707 7669 3708
rect 7238 3166 7666 3226
rect 7051 2548 7117 2549
rect 7051 2484 7052 2548
rect 7116 2484 7117 2548
rect 7051 2483 7117 2484
rect 5211 1596 5277 1597
rect 5211 1532 5212 1596
rect 5276 1532 5277 1596
rect 5211 1531 5277 1532
rect 7606 1461 7666 3166
rect 7874 2752 8195 3776
rect 8342 3365 8402 5203
rect 8526 3909 8586 19347
rect 8891 16556 8957 16557
rect 8891 16492 8892 16556
rect 8956 16492 8957 16556
rect 8891 16491 8957 16492
rect 8894 12749 8954 16491
rect 9627 13700 9693 13701
rect 9627 13636 9628 13700
rect 9692 13636 9693 13700
rect 9627 13635 9693 13636
rect 8891 12748 8957 12749
rect 8891 12684 8892 12748
rect 8956 12684 8957 12748
rect 8891 12683 8957 12684
rect 9443 11388 9509 11389
rect 9443 11324 9444 11388
rect 9508 11324 9509 11388
rect 9443 11323 9509 11324
rect 8707 10436 8773 10437
rect 8707 10372 8708 10436
rect 8772 10372 8773 10436
rect 8707 10371 8773 10372
rect 8710 8669 8770 10371
rect 9075 9484 9141 9485
rect 9075 9420 9076 9484
rect 9140 9420 9141 9484
rect 9075 9419 9141 9420
rect 9078 9298 9138 9419
rect 9446 9346 9506 11323
rect 9308 9286 9506 9346
rect 9308 8802 9368 9286
rect 9630 9213 9690 13635
rect 9443 9212 9509 9213
rect 9443 9148 9444 9212
rect 9508 9148 9509 9212
rect 9443 9147 9509 9148
rect 9627 9212 9693 9213
rect 9627 9148 9628 9212
rect 9692 9148 9693 9212
rect 9627 9147 9693 9148
rect 9078 8742 9368 8802
rect 8707 8668 8773 8669
rect 8707 8604 8708 8668
rect 8772 8604 8773 8668
rect 8707 8603 8773 8604
rect 8523 3908 8589 3909
rect 8523 3844 8524 3908
rect 8588 3844 8589 3908
rect 8523 3843 8589 3844
rect 8339 3364 8405 3365
rect 8339 3300 8340 3364
rect 8404 3300 8405 3364
rect 8339 3299 8405 3300
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 8710 2549 8770 8603
rect 8891 7988 8957 7989
rect 8891 7924 8892 7988
rect 8956 7924 8957 7988
rect 8891 7923 8957 7924
rect 8894 4317 8954 7923
rect 8891 4316 8957 4317
rect 8891 4252 8892 4316
rect 8956 4252 8957 4316
rect 8891 4251 8957 4252
rect 8891 2684 8957 2685
rect 8891 2620 8892 2684
rect 8956 2620 8957 2684
rect 8891 2619 8957 2620
rect 8707 2548 8773 2549
rect 8707 2484 8708 2548
rect 8772 2484 8773 2548
rect 8707 2483 8773 2484
rect 8894 2005 8954 2619
rect 8891 2004 8957 2005
rect 8891 1940 8892 2004
rect 8956 1940 8957 2004
rect 8891 1939 8957 1940
rect 9078 1461 9138 8742
rect 9259 6900 9325 6901
rect 9259 6836 9260 6900
rect 9324 6836 9325 6900
rect 9259 6835 9325 6836
rect 9262 5266 9322 6835
rect 9446 6085 9506 9147
rect 9443 6084 9509 6085
rect 9443 6020 9444 6084
rect 9508 6020 9509 6084
rect 9443 6019 9509 6020
rect 9262 5206 9506 5266
rect 9446 2549 9506 5206
rect 9630 2821 9690 9147
rect 9814 2821 9874 19755
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 12019 19140 12085 19141
rect 12019 19076 12020 19140
rect 12084 19076 12085 19140
rect 12019 19075 12085 19076
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 10179 17372 10245 17373
rect 10179 17308 10180 17372
rect 10244 17308 10245 17372
rect 10179 17307 10245 17308
rect 9995 15604 10061 15605
rect 9995 15540 9996 15604
rect 10060 15540 10061 15604
rect 9995 15539 10061 15540
rect 9627 2820 9693 2821
rect 9627 2756 9628 2820
rect 9692 2756 9693 2820
rect 9627 2755 9693 2756
rect 9811 2820 9877 2821
rect 9811 2756 9812 2820
rect 9876 2756 9877 2820
rect 9811 2755 9877 2756
rect 9443 2548 9509 2549
rect 9443 2484 9444 2548
rect 9508 2484 9509 2548
rect 9443 2483 9509 2484
rect 9998 2277 10058 15539
rect 10182 2821 10242 17307
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 10363 13156 10429 13157
rect 10363 13092 10364 13156
rect 10428 13092 10429 13156
rect 10363 13091 10429 13092
rect 10366 8805 10426 13091
rect 11340 13088 11660 14112
rect 12022 13429 12082 19075
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 12203 18868 12269 18869
rect 12203 18804 12204 18868
rect 12268 18804 12269 18868
rect 12203 18803 12269 18804
rect 13491 18868 13557 18869
rect 13491 18804 13492 18868
rect 13556 18804 13557 18868
rect 13491 18803 13557 18804
rect 12206 13429 12266 18803
rect 12387 17644 12453 17645
rect 12387 17580 12388 17644
rect 12452 17580 12453 17644
rect 12387 17579 12453 17580
rect 12019 13428 12085 13429
rect 12019 13364 12020 13428
rect 12084 13364 12085 13428
rect 12019 13363 12085 13364
rect 12203 13428 12269 13429
rect 12203 13364 12204 13428
rect 12268 13364 12269 13428
rect 12203 13363 12269 13364
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11835 12612 11901 12613
rect 11835 12548 11836 12612
rect 11900 12548 11901 12612
rect 11835 12547 11901 12548
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 10363 8804 10429 8805
rect 10363 8740 10364 8804
rect 10428 8740 10429 8804
rect 10363 8739 10429 8740
rect 10366 3773 10426 8739
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 10915 8668 10981 8669
rect 10915 8604 10916 8668
rect 10980 8604 10981 8668
rect 10915 8603 10981 8604
rect 11099 8668 11165 8669
rect 11099 8604 11100 8668
rect 11164 8604 11165 8668
rect 11099 8603 11165 8604
rect 10547 8396 10613 8397
rect 10547 8332 10548 8396
rect 10612 8332 10613 8396
rect 10547 8331 10613 8332
rect 10363 3772 10429 3773
rect 10363 3708 10364 3772
rect 10428 3708 10429 3772
rect 10363 3707 10429 3708
rect 10550 3229 10610 8331
rect 10731 7580 10797 7581
rect 10731 7516 10732 7580
rect 10796 7516 10797 7580
rect 10731 7515 10797 7516
rect 10734 6629 10794 7515
rect 10918 7445 10978 8603
rect 10915 7444 10981 7445
rect 10915 7380 10916 7444
rect 10980 7380 10981 7444
rect 10915 7379 10981 7380
rect 10915 7036 10981 7037
rect 10915 6972 10916 7036
rect 10980 6972 10981 7036
rect 10915 6971 10981 6972
rect 10731 6628 10797 6629
rect 10731 6564 10732 6628
rect 10796 6564 10797 6628
rect 10731 6563 10797 6564
rect 10731 6084 10797 6085
rect 10731 6020 10732 6084
rect 10796 6020 10797 6084
rect 10731 6019 10797 6020
rect 10547 3228 10613 3229
rect 10547 3164 10548 3228
rect 10612 3164 10613 3228
rect 10547 3163 10613 3164
rect 10734 2821 10794 6019
rect 10179 2820 10245 2821
rect 10179 2756 10180 2820
rect 10244 2756 10245 2820
rect 10179 2755 10245 2756
rect 10731 2820 10797 2821
rect 10731 2756 10732 2820
rect 10796 2756 10797 2820
rect 10731 2755 10797 2756
rect 10918 2549 10978 6971
rect 11102 3637 11162 8603
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11838 7445 11898 12547
rect 12019 12476 12085 12477
rect 12019 12412 12020 12476
rect 12084 12412 12085 12476
rect 12019 12411 12085 12412
rect 12022 8261 12082 12411
rect 12203 10164 12269 10165
rect 12203 10100 12204 10164
rect 12268 10100 12269 10164
rect 12203 10099 12269 10100
rect 12019 8260 12085 8261
rect 12019 8196 12020 8260
rect 12084 8196 12085 8260
rect 12019 8195 12085 8196
rect 11835 7444 11901 7445
rect 11835 7380 11836 7444
rect 11900 7380 11901 7444
rect 11835 7379 11901 7380
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 12206 6085 12266 10099
rect 12390 10029 12450 17579
rect 12571 16556 12637 16557
rect 12571 16492 12572 16556
rect 12636 16492 12637 16556
rect 12571 16491 12637 16492
rect 12574 10981 12634 16491
rect 13494 13565 13554 18803
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14043 17644 14109 17645
rect 14043 17580 14044 17644
rect 14108 17580 14109 17644
rect 14043 17579 14109 17580
rect 13859 15876 13925 15877
rect 13859 15812 13860 15876
rect 13924 15812 13925 15876
rect 13859 15811 13925 15812
rect 13862 15197 13922 15811
rect 13859 15196 13925 15197
rect 13859 15132 13860 15196
rect 13924 15132 13925 15196
rect 13859 15131 13925 15132
rect 13491 13564 13557 13565
rect 13491 13500 13492 13564
rect 13556 13500 13557 13564
rect 13491 13499 13557 13500
rect 12755 12340 12821 12341
rect 12755 12276 12756 12340
rect 12820 12276 12821 12340
rect 12755 12275 12821 12276
rect 12571 10980 12637 10981
rect 12571 10916 12572 10980
rect 12636 10916 12637 10980
rect 12571 10915 12637 10916
rect 12571 10844 12637 10845
rect 12571 10780 12572 10844
rect 12636 10780 12637 10844
rect 12571 10779 12637 10780
rect 12387 10028 12453 10029
rect 12387 9964 12388 10028
rect 12452 9964 12453 10028
rect 12387 9963 12453 9964
rect 12387 7036 12453 7037
rect 12387 6972 12388 7036
rect 12452 6972 12453 7036
rect 12387 6971 12453 6972
rect 11835 6084 11901 6085
rect 11835 6020 11836 6084
rect 11900 6020 11901 6084
rect 11835 6019 11901 6020
rect 12203 6084 12269 6085
rect 12203 6020 12204 6084
rect 12268 6020 12269 6084
rect 12203 6019 12269 6020
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11099 3636 11165 3637
rect 11099 3572 11100 3636
rect 11164 3572 11165 3636
rect 11099 3571 11165 3572
rect 11340 3296 11660 4320
rect 11838 3773 11898 6019
rect 12203 5404 12269 5405
rect 12203 5340 12204 5404
rect 12268 5340 12269 5404
rect 12203 5339 12269 5340
rect 12206 4725 12266 5339
rect 12203 4724 12269 4725
rect 12203 4660 12204 4724
rect 12268 4660 12269 4724
rect 12203 4659 12269 4660
rect 12390 3773 12450 6971
rect 12574 5269 12634 10779
rect 12571 5268 12637 5269
rect 12571 5204 12572 5268
rect 12636 5204 12637 5268
rect 12571 5203 12637 5204
rect 11835 3772 11901 3773
rect 11835 3708 11836 3772
rect 11900 3708 11901 3772
rect 11835 3707 11901 3708
rect 12387 3772 12453 3773
rect 12387 3708 12388 3772
rect 12452 3708 12453 3772
rect 12387 3707 12453 3708
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 10915 2548 10981 2549
rect 10915 2484 10916 2548
rect 10980 2484 10981 2548
rect 10915 2483 10981 2484
rect 9995 2276 10061 2277
rect 9995 2212 9996 2276
rect 10060 2212 10061 2276
rect 9995 2211 10061 2212
rect 11340 2208 11660 3232
rect 12758 3229 12818 12275
rect 13494 11933 13554 13499
rect 13862 12069 13922 15131
rect 14046 13157 14106 17579
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 18270 20704 18590 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 19616 18590 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 18528 18590 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 17440 18590 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 16352 18590 17376
rect 19195 16964 19261 16965
rect 19195 16900 19196 16964
rect 19260 16900 19261 16964
rect 19195 16899 19261 16900
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 15699 15604 15765 15605
rect 15699 15540 15700 15604
rect 15764 15540 15765 15604
rect 15699 15539 15765 15540
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14043 13156 14109 13157
rect 14043 13092 14044 13156
rect 14108 13092 14109 13156
rect 14043 13091 14109 13092
rect 14227 12884 14293 12885
rect 14227 12820 14228 12884
rect 14292 12820 14293 12884
rect 14227 12819 14293 12820
rect 14230 12205 14290 12819
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14227 12204 14293 12205
rect 14227 12140 14228 12204
rect 14292 12140 14293 12204
rect 14227 12139 14293 12140
rect 13859 12068 13925 12069
rect 13859 12004 13860 12068
rect 13924 12004 13925 12068
rect 13859 12003 13925 12004
rect 13491 11932 13557 11933
rect 13491 11868 13492 11932
rect 13556 11868 13557 11932
rect 13491 11867 13557 11868
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 15702 10301 15762 15539
rect 18270 15264 18590 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 14176 18590 15200
rect 19198 15061 19258 16899
rect 19195 15060 19261 15061
rect 19195 14996 19196 15060
rect 19260 14996 19261 15060
rect 19195 14995 19261 14996
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 13088 18590 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 12000 18590 13024
rect 19198 12477 19258 14995
rect 19195 12476 19261 12477
rect 19195 12412 19196 12476
rect 19260 12412 19261 12476
rect 19195 12411 19261 12412
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 10912 18590 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 15699 10300 15765 10301
rect 15699 10236 15700 10300
rect 15764 10236 15765 10300
rect 15699 10235 15765 10236
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14227 8804 14293 8805
rect 14227 8740 14228 8804
rect 14292 8740 14293 8804
rect 14227 8739 14293 8740
rect 13123 7988 13189 7989
rect 13123 7924 13124 7988
rect 13188 7924 13189 7988
rect 13123 7923 13189 7924
rect 12939 7716 13005 7717
rect 12939 7652 12940 7716
rect 13004 7652 13005 7716
rect 12939 7651 13005 7652
rect 12755 3228 12821 3229
rect 12755 3164 12756 3228
rect 12820 3164 12821 3228
rect 12755 3163 12821 3164
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 12942 1597 13002 7651
rect 13126 3773 13186 7923
rect 14230 4317 14290 8739
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 18270 9824 18590 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 8736 18590 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 7648 18590 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 6560 18590 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 15515 5540 15581 5541
rect 15515 5476 15516 5540
rect 15580 5476 15581 5540
rect 15515 5475 15581 5476
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14227 4316 14293 4317
rect 14227 4252 14228 4316
rect 14292 4252 14293 4316
rect 14227 4251 14293 4252
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 13123 3772 13189 3773
rect 13123 3708 13124 3772
rect 13188 3708 13189 3772
rect 13123 3707 13189 3708
rect 14805 2752 15125 3776
rect 15518 2821 15578 5475
rect 18270 5472 18590 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 15699 5404 15765 5405
rect 15699 5340 15700 5404
rect 15764 5340 15765 5404
rect 15699 5339 15765 5340
rect 15702 3637 15762 5339
rect 18270 4384 18590 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 15699 3636 15765 3637
rect 15699 3572 15700 3636
rect 15764 3572 15765 3636
rect 15699 3571 15765 3572
rect 18270 3296 18590 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 15515 2820 15581 2821
rect 15515 2756 15516 2820
rect 15580 2756 15581 2820
rect 15515 2755 15581 2756
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 2208 18590 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2128 18590 2144
rect 12939 1596 13005 1597
rect 12939 1532 12940 1596
rect 13004 1532 13005 1596
rect 12939 1531 13005 1532
rect 7603 1460 7669 1461
rect 7603 1396 7604 1460
rect 7668 1396 7669 1460
rect 7603 1395 7669 1396
rect 9075 1460 9141 1461
rect 9075 1396 9076 1460
rect 9140 1396 9141 1460
rect 9075 1395 9141 1396
rect 3739 236 3805 237
rect 3739 172 3740 236
rect 3804 172 3805 236
rect 3739 171 3805 172
<< via4 >>
rect 3102 9062 3338 9298
rect 8990 9062 9226 9298
<< metal5 >>
rect 3060 9298 9268 9340
rect 3060 9062 3102 9298
rect 3338 9062 8990 9298
rect 9226 9062 9268 9298
rect 3060 9020 9268 9062
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2852 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2852 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4508 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_35 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6348 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5520 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6164 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1604681595
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8280 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 7084 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8372 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10488 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10580 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9752 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1604681595
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_100
timestamp 1604681595
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_3_
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11316 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121
timestamp 1604681595
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1604681595
transform 1 0 13984 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_0_134 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13432 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_132
timestamp 1604681595
transform 1 0 13248 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 15548 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_146
timestamp 1604681595
transform 1 0 14536 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1604681595
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_165
timestamp 1604681595
transform 1 0 16284 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_149
timestamp 1604681595
transform 1 0 14812 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_161
timestamp 1604681595
transform 1 0 15916 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_173
timestamp 1604681595
transform 1 0 17020 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 17020 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 16652 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1604681595
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_177
timestamp 1604681595
transform 1 0 17388 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_187 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1604681595
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 19964 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 18860 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 19136 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20240 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1604681595
transform 1 0 19228 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_188
timestamp 1604681595
transform 1 0 18400 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_200
timestamp 1604681595
transform 1 0 19504 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_209
timestamp 1604681595
transform 1 0 20332 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222
timestamp 1604681595
transform 1 0 21528 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_214
timestamp 1604681595
transform 1 0 20792 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_222
timestamp 1604681595
transform 1 0 21528 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 2852 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_28
timestamp 1604681595
transform 1 0 3680 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 5796 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_2_48
timestamp 1604681595
transform 1 0 5520 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 7636 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_67
timestamp 1604681595
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_80
timestamp 1604681595
transform 1 0 8464 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_4_
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10488 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1604681595
transform 1 0 9108 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_86
timestamp 1604681595
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 12144 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12512 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 11316 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1604681595
transform 1 0 14076 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_130
timestamp 1604681595
transform 1 0 13064 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_138
timestamp 1604681595
transform 1 0 13800 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_145
timestamp 1604681595
transform 1 0 14444 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_158
timestamp 1604681595
transform 1 0 15640 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_166
timestamp 1604681595
transform 1 0 16376 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 16468 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 17572 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_171
timestamp 1604681595
transform 1 0 16836 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 19596 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_188 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 18400 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_200
timestamp 1604681595
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_205
timestamp 1604681595
transform 1 0 19964 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1604681595
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2852 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4324 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1604681595
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7728 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_3_71
timestamp 1604681595
transform 1 0 7636 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9936 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9200 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_94
timestamp 1604681595
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1604681595
transform 1 0 12512 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11592 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_3_
timestamp 1604681595
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1604681595
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 14444 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_3_128
timestamp 1604681595
transform 1 0 12880 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_140
timestamp 1604681595
transform 1 0 13984 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_144
timestamp 1604681595
transform 1 0 14352 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_161
timestamp 1604681595
transform 1 0 15916 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 16652 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_173
timestamp 1604681595
transform 1 0 17020 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 19596 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_193
timestamp 1604681595
transform 1 0 18860 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_210
timestamp 1604681595
transform 1 0 20424 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_222
timestamp 1604681595
transform 1 0 21528 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_3_
timestamp 1604681595
transform 1 0 2852 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_28
timestamp 1604681595
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5520 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6348 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 7176 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8648 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_72
timestamp 1604681595
transform 1 0 7728 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9936 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1604681595
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_5_
timestamp 1604681595
transform 1 0 11592 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_4_111
timestamp 1604681595
transform 1 0 11316 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_123
timestamp 1604681595
transform 1 0 12420 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13156 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_140
timestamp 1604681595
transform 1 0 13984 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15824 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1604681595
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17388 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_4_169
timestamp 1604681595
transform 1 0 16652 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 19688 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_193
timestamp 1604681595
transform 1 0 18860 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_201
timestamp 1604681595
transform 1 0 19596 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_206
timestamp 1604681595
transform 1 0 20056 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2852 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4324 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_60
timestamp 1604681595
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7728 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8648 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_71
timestamp 1604681595
transform 1 0 7636 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_81
timestamp 1604681595
transform 1 0 8556 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9844 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_91
timestamp 1604681595
transform 1 0 9476 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_104
timestamp 1604681595
transform 1 0 10672 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_116
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_139
timestamp 1604681595
transform 1 0 13892 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 14628 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_5_163
timestamp 1604681595
transform 1 0 16100 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_175
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19596 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_193
timestamp 1604681595
transform 1 0 18860 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_210
timestamp 1604681595
transform 1 0 20424 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1604681595
transform 1 0 21528 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2024 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2852 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_9
timestamp 1604681595
transform 1 0 1932 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4232 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4508 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 3496 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_28
timestamp 1604681595
transform 1 0 3680 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_35
timestamp 1604681595
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604681595
transform 1 0 6348 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5704 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6532 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6900 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7452 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8556 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_3_
timestamp 1604681595
transform 1 0 8372 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_78
timestamp 1604681595
transform 1 0 8280 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 9200 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10212 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1604681595
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_92
timestamp 1604681595
transform 1 0 9568 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_98
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11868 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_109
timestamp 1604681595
transform 1 0 11132 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_108
timestamp 1604681595
transform 1 0 11040 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 13432 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_6_126
timestamp 1604681595
transform 1 0 12696 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_143
timestamp 1604681595
transform 1 0 14260 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_139
timestamp 1604681595
transform 1 0 13892 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15824 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16192 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14628 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1604681595
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_156
timestamp 1604681595
transform 1 0 15456 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18308 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_176
timestamp 1604681595
transform 1 0 17296 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_184
timestamp 1604681595
transform 1 0 18032 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_173
timestamp 1604681595
transform 1 0 17020 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19596 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_6_203
timestamp 1604681595
transform 1 0 19780 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_193
timestamp 1604681595
transform 1 0 18860 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_211
timestamp 1604681595
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_210
timestamp 1604681595
transform 1 0 20424 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_222
timestamp 1604681595
transform 1 0 21528 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2852 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4876 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_28
timestamp 1604681595
transform 1 0 3680 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 6532 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5704 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_8_62
timestamp 1604681595
transform 1 0 6808 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7268 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_66
timestamp 1604681595
transform 1 0 7176 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_76
timestamp 1604681595
transform 1 0 8096 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10028 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_88
timestamp 1604681595
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 11592 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_106
timestamp 1604681595
transform 1 0 10856 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1604681595
transform 1 0 12420 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_135
timestamp 1604681595
transform 1 0 13524 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_145
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16192 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_162
timestamp 1604681595
transform 1 0 16008 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_180
timestamp 1604681595
transform 1 0 17664 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 18400 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_8_204
timestamp 1604681595
transform 1 0 19872 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1604681595
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1604681595
transform 1 0 2208 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4048 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4876 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1604681595
transform 1 0 3864 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_21
timestamp 1604681595
transform 1 0 3036 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_29
timestamp 1604681595
transform 1 0 3772 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5704 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_78
timestamp 1604681595
transform 1 0 8280 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 10120 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_9_89
timestamp 1604681595
transform 1 0 9292 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_97
timestamp 1604681595
transform 1 0 10028 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_139
timestamp 1604681595
transform 1 0 13892 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 14996 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_160
timestamp 1604681595
transform 1 0 15824 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16560 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18308 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_174
timestamp 1604681595
transform 1 0 17112 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1604681595
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1604681595
transform 1 0 19596 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1604681595
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_193
timestamp 1604681595
transform 1 0 18860 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_210
timestamp 1604681595
transform 1 0 20424 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_222
timestamp 1604681595
transform 1 0 21528 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1604681595
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_23
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_41
timestamp 1604681595
transform 1 0 4876 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 6440 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4968 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_62
timestamp 1604681595
transform 1 0 6808 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7176 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8740 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_75
timestamp 1604681595
transform 1 0 8004 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_86
timestamp 1604681595
transform 1 0 9016 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_6_
timestamp 1604681595
transform 1 0 12052 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_109
timestamp 1604681595
transform 1 0 11132 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_117
timestamp 1604681595
transform 1 0 11868 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_128
timestamp 1604681595
transform 1 0 12880 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_145
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_163
timestamp 1604681595
transform 1 0 16100 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 17480 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_10_175
timestamp 1604681595
transform 1 0 17204 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 19688 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_194
timestamp 1604681595
transform 1 0 18952 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_206
timestamp 1604681595
transform 1 0 20056 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1472 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2944 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 3680 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_26
timestamp 1604681595
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5704 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 5428 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_44
timestamp 1604681595
transform 1 0 5152 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7544 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_79
timestamp 1604681595
transform 1 0 8372 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 9200 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1604681595
transform 1 0 10212 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_87
timestamp 1604681595
transform 1 0 9108 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_91
timestamp 1604681595
transform 1 0 9476 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_102
timestamp 1604681595
transform 1 0 10488 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_110
timestamp 1604681595
transform 1 0 11224 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_114
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 12880 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 14076 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_127
timestamp 1604681595
transform 1 0 12788 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_131
timestamp 1604681595
transform 1 0 13156 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_139
timestamp 1604681595
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_157
timestamp 1604681595
transform 1 0 15548 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_165
timestamp 1604681595
transform 1 0 16284 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_175
timestamp 1604681595
transform 1 0 17204 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_200
timestamp 1604681595
transform 1 0 19504 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_211
timestamp 1604681595
transform 1 0 20516 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_12
timestamp 1604681595
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4876 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_26
timestamp 1604681595
transform 1 0 3496 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1604681595
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5428 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_56
timestamp 1604681595
transform 1 0 6256 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6992 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_73
timestamp 1604681595
transform 1 0 7820 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 9844 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_84
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_104
timestamp 1604681595
transform 1 0 10672 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12328 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 11684 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_112
timestamp 1604681595
transform 1 0 11408 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_118
timestamp 1604681595
transform 1 0 11960 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 14168 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 13892 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_131
timestamp 1604681595
transform 1 0 13156 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_145
timestamp 1604681595
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_163
timestamp 1604681595
transform 1 0 16100 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1604681595
transform 1 0 17388 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_175
timestamp 1604681595
transform 1 0 17204 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_180
timestamp 1604681595
transform 1 0 17664 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 18400 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1604681595
transform 1 0 19228 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_209
timestamp 1604681595
transform 1 0 20332 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1604681595
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1472 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1604681595
transform 1 0 2116 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_20
timestamp 1604681595
transform 1 0 2944 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1604681595
transform 1 0 2944 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3680 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_37
timestamp 1604681595
transform 1 0 4508 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_28
timestamp 1604681595
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_38
timestamp 1604681595
transform 1 0 4600 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5336 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5244 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_62
timestamp 1604681595
transform 1 0 6808 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1604681595
transform 1 0 7912 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7544 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_66
timestamp 1604681595
transform 1 0 7176 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_83
timestamp 1604681595
transform 1 0 8740 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_79
timestamp 1604681595
transform 1 0 8372 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10212 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 9844 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 9476 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_94
timestamp 1604681595
transform 1 0 9752 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_104
timestamp 1604681595
transform 1 0 10672 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1604681595
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12420 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12512 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_116
timestamp 1604681595
transform 1 0 11776 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_115
timestamp 1604681595
transform 1 0 11684 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 14076 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_133
timestamp 1604681595
transform 1 0 13340 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_144
timestamp 1604681595
transform 1 0 14352 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_139
timestamp 1604681595
transform 1 0 13892 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 14720 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_164
timestamp 1604681595
transform 1 0 16192 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1604681595
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_163
timestamp 1604681595
transform 1 0 16100 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 16928 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1604681595
transform 1 0 16836 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_175
timestamp 1604681595
transform 1 0 17204 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_180
timestamp 1604681595
transform 1 0 17664 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18400 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_200
timestamp 1604681595
transform 1 0 19504 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1604681595
transform 1 0 19228 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_211
timestamp 1604681595
transform 1 0 20516 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1604681595
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1604681595
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2024 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 1604681595
transform 1 0 1932 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4232 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_26
timestamp 1604681595
transform 1 0 3496 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_43
timestamp 1604681595
transform 1 0 5060 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_55
timestamp 1604681595
transform 1 0 6164 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_78
timestamp 1604681595
transform 1 0 8280 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9568 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_89
timestamp 1604681595
transform 1 0 9292 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_108
timestamp 1604681595
transform 1 0 11040 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_116
timestamp 1604681595
transform 1 0 11776 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 14444 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_15_132
timestamp 1604681595
transform 1 0 13248 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_144
timestamp 1604681595
transform 1 0 14352 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_161
timestamp 1604681595
transform 1 0 15916 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16652 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_175
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 19596 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1604681595
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1604681595
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_195
timestamp 1604681595
transform 1 0 19044 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1604681595
transform 1 0 20424 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_212
timestamp 1604681595
transform 1 0 20608 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_220
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_6
timestamp 1604681595
transform 1 0 1656 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4508 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_36
timestamp 1604681595
transform 1 0 4416 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1604681595
transform 1 0 5980 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_65
timestamp 1604681595
transform 1 0 7084 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10396 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_16_84
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12236 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_130
timestamp 1604681595
transform 1 0 13064 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_145
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_160
timestamp 1604681595
transform 1 0 15824 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 16744 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_168
timestamp 1604681595
transform 1 0 16560 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_186
timestamp 1604681595
transform 1 0 18216 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 18952 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_203
timestamp 1604681595
transform 1 0 19780 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_211
timestamp 1604681595
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2392 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_6
timestamp 1604681595
transform 1 0 1656 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4600 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_30
timestamp 1604681595
transform 1 0 3864 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_47
timestamp 1604681595
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6992 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8556 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_73
timestamp 1604681595
transform 1 0 7820 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_90
timestamp 1604681595
transform 1 0 9384 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11132 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1604681595
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 13984 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_132
timestamp 1604681595
transform 1 0 13248 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_143
timestamp 1604681595
transform 1 0 14260 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 14904 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_149
timestamp 1604681595
transform 1 0 14812 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_159
timestamp 1604681595
transform 1 0 15732 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16468 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_173
timestamp 1604681595
transform 1 0 17020 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1604681595
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 19596 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_193
timestamp 1604681595
transform 1 0 18860 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_210
timestamp 1604681595
transform 1 0 20424 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_222
timestamp 1604681595
transform 1 0 21528 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2116 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1604681595
transform 1 0 2944 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4140 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_28
timestamp 1604681595
transform 1 0 3680 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 6348 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_49
timestamp 1604681595
transform 1 0 5612 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7912 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_66
timestamp 1604681595
transform 1 0 7176 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_83
timestamp 1604681595
transform 1 0 8740 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1604681595
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_102
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_119
timestamp 1604681595
transform 1 0 12052 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12972 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_127
timestamp 1604681595
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_145
timestamp 1604681595
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_163
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 17020 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_171
timestamp 1604681595
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_189
timestamp 1604681595
transform 1 0 18492 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_206
timestamp 1604681595
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_9
timestamp 1604681595
transform 1 0 1932 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_10
timestamp 1604681595
transform 1 0 2024 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2024 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 1656 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2760 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_20_16
timestamp 1604681595
transform 1 0 2576 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4324 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_27
timestamp 1604681595
transform 1 0 3588 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_28
timestamp 1604681595
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_41
timestamp 1604681595
transform 1 0 4876 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6348 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 5796 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_44
timestamp 1604681595
transform 1 0 5152 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_56
timestamp 1604681595
transform 1 0 6256 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_49
timestamp 1604681595
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_54
timestamp 1604681595
transform 1 0 6072 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 8556 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8372 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_19_71
timestamp 1604681595
transform 1 0 7636 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_73
timestamp 1604681595
transform 1 0 7820 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_88
timestamp 1604681595
transform 1 0 9200 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_96
timestamp 1604681595
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11868 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_109
timestamp 1604681595
transform 1 0 11132 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_19_139
timestamp 1604681595
transform 1 0 13892 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_126
timestamp 1604681595
transform 1 0 12696 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_134
timestamp 1604681595
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 14628 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_163
timestamp 1604681595
transform 1 0 16100 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_160
timestamp 1604681595
transform 1 0 15824 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 16836 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 16744 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_175
timestamp 1604681595
transform 1 0 17204 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_168
timestamp 1604681595
transform 1 0 16560 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_186
timestamp 1604681595
transform 1 0 18216 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19596 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18952 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_19_193
timestamp 1604681595
transform 1 0 18860 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_203
timestamp 1604681595
transform 1 0 19780 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_210
timestamp 1604681595
transform 1 0 20424 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_222
timestamp 1604681595
transform 1 0 21528 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_211
timestamp 1604681595
transform 1 0 20516 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1472 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_20
timestamp 1604681595
transform 1 0 2944 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3680 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_37
timestamp 1604681595
transform 1 0 4508 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 5244 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_49
timestamp 1604681595
transform 1 0 5612 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7452 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_68
timestamp 1604681595
transform 1 0 7360 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_85
timestamp 1604681595
transform 1 0 8924 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_102
timestamp 1604681595
transform 1 0 10488 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 11224 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13064 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_129
timestamp 1604681595
transform 1 0 12972 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_139
timestamp 1604681595
transform 1 0 13892 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 14628 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_21_163
timestamp 1604681595
transform 1 0 16100 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 16836 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_175
timestamp 1604681595
transform 1 0 17204 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19412 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_21_190
timestamp 1604681595
transform 1 0 18584 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_198
timestamp 1604681595
transform 1 0 19320 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_215
timestamp 1604681595
transform 1 0 20884 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1748 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4416 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6440 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_22_45
timestamp 1604681595
transform 1 0 5244 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_57
timestamp 1604681595
transform 1 0 6348 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_67
timestamp 1604681595
transform 1 0 7268 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1604681595
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_84
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_104
timestamp 1604681595
transform 1 0 10672 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11868 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 11224 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_113
timestamp 1604681595
transform 1 0 11500 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 14076 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_133
timestamp 1604681595
transform 1 0 13340 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_160
timestamp 1604681595
transform 1 0 15824 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18216 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16652 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_168
timestamp 1604681595
transform 1 0 16560 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_178
timestamp 1604681595
transform 1 0 17480 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 19780 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_195
timestamp 1604681595
transform 1 0 19044 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_206
timestamp 1604681595
transform 1 0 20056 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1604681595
transform 1 0 2208 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_11
timestamp 1604681595
transform 1 0 2116 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 3772 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_23_21
timestamp 1604681595
transform 1 0 3036 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_45
timestamp 1604681595
transform 1 0 5244 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8556 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_23_71
timestamp 1604681595
transform 1 0 7636 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_79
timestamp 1604681595
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_97
timestamp 1604681595
transform 1 0 10028 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_114
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12696 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 14904 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 14628 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_159
timestamp 1604681595
transform 1 0 15732 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16652 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_167
timestamp 1604681595
transform 1 0 16468 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_175
timestamp 1604681595
transform 1 0 17204 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_5_
timestamp 1604681595
transform 1 0 19596 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_193
timestamp 1604681595
transform 1 0 18860 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_210
timestamp 1604681595
transform 1 0 20424 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_222
timestamp 1604681595
transform 1 0 21528 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_6
timestamp 1604681595
transform 1 0 1656 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4232 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_23
timestamp 1604681595
transform 1 0 3220 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 5796 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_43
timestamp 1604681595
transform 1 0 5060 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_67
timestamp 1604681595
transform 1 0 7268 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_84
timestamp 1604681595
transform 1 0 8832 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_102
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11224 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_119
timestamp 1604681595
transform 1 0 12052 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_131
timestamp 1604681595
transform 1 0 13156 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_135
timestamp 1604681595
transform 1 0 13524 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_145
timestamp 1604681595
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_160
timestamp 1604681595
transform 1 0 15824 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16560 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_184
timestamp 1604681595
transform 1 0 18032 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_6_
timestamp 1604681595
transform 1 0 18768 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_201
timestamp 1604681595
transform 1 0 19596 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1604681595
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2116 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_17
timestamp 1604681595
transform 1 0 2668 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 3404 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_31
timestamp 1604681595
transform 1 0 3956 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_48
timestamp 1604681595
transform 1 0 5520 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_60
timestamp 1604681595
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8556 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 6992 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_73
timestamp 1604681595
transform 1 0 7820 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_97
timestamp 1604681595
transform 1 0 10028 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12788 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_25_143
timestamp 1604681595
transform 1 0 14260 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 14996 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_160
timestamp 1604681595
transform 1 0 15824 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16560 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_174
timestamp 1604681595
transform 1 0 17112 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1604681595
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_4_
timestamp 1604681595
transform 1 0 19596 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_193
timestamp 1604681595
transform 1 0 18860 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_210
timestamp 1604681595
transform 1 0 20424 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_222
timestamp 1604681595
transform 1 0 21528 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2208 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2024 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_9
timestamp 1604681595
transform 1 0 1932 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_16
timestamp 1604681595
transform 1 0 2576 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_11
timestamp 1604681595
transform 1 0 2116 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4416 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_28
timestamp 1604681595
transform 1 0 3680 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1604681595
transform 1 0 4876 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_28
timestamp 1604681595
transform 1 0 3680 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1604681595
transform 1 0 6348 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_53
timestamp 1604681595
transform 1 0 5980 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_60
timestamp 1604681595
transform 1 0 6624 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_45
timestamp 1604681595
transform 1 0 5244 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1604681595
transform 1 0 6348 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7636 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_70
timestamp 1604681595
transform 1 0 7544 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_80
timestamp 1604681595
transform 1 0 8464 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604681595
transform 1 0 9200 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10120 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10212 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_84
timestamp 1604681595
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_97
timestamp 1604681595
transform 1 0 10028 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_91
timestamp 1604681595
transform 1 0 9476 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12236 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_107
timestamp 1604681595
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_119
timestamp 1604681595
transform 1 0 12052 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_108
timestamp 1604681595
transform 1 0 11040 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1604681595
transform 1 0 13800 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13708 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1604681595
transform 1 0 13616 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_130
timestamp 1604681595
transform 1 0 13064 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1604681595
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_126
timestamp 1604681595
transform 1 0 12696 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_134
timestamp 1604681595
transform 1 0 13432 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 15272 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15824 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_146
timestamp 1604681595
transform 1 0 14536 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18032 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_176
timestamp 1604681595
transform 1 0 17296 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_170
timestamp 1604681595
transform 1 0 16744 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1604681595
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 19596 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 19596 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_26_193
timestamp 1604681595
transform 1 0 18860 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_205
timestamp 1604681595
transform 1 0 19964 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_193
timestamp 1604681595
transform 1 0 18860 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1604681595
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_210
timestamp 1604681595
transform 1 0 20424 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_222
timestamp 1604681595
transform 1 0 21528 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2024 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_9
timestamp 1604681595
transform 1 0 1932 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_16
timestamp 1604681595
transform 1 0 2576 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_28
timestamp 1604681595
transform 1 0 3680 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1604681595
transform 1 0 6256 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_48
timestamp 1604681595
transform 1 0 5520 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_59
timestamp 1604681595
transform 1 0 6532 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_28_67
timestamp 1604681595
transform 1 0 7268 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604681595
transform 1 0 10580 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_101
timestamp 1604681595
transform 1 0 10396 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11592 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_106
timestamp 1604681595
transform 1 0 10856 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1604681595
transform 1 0 12420 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604681595
transform 1 0 14076 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_135
timestamp 1604681595
transform 1 0 13524 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_145
timestamp 1604681595
transform 1 0 14444 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_163
timestamp 1604681595
transform 1 0 16100 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16836 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1604681595
transform 1 0 18216 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_180
timestamp 1604681595
transform 1 0 17664 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18400 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1604681595
transform 1 0 19228 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_199
timestamp 1604681595
transform 1 0 19412 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_211
timestamp 1604681595
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2944 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_11
timestamp 1604681595
transform 1 0 2116 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_19
timestamp 1604681595
transform 1 0 2852 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4508 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_29_29
timestamp 1604681595
transform 1 0 3772 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_53
timestamp 1604681595
transform 1 0 5980 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8188 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_29_65
timestamp 1604681595
transform 1 0 7084 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1604681595
transform 1 0 10396 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_93
timestamp 1604681595
transform 1 0 9660 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_104
timestamp 1604681595
transform 1 0 10672 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_116
timestamp 1604681595
transform 1 0 11776 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_132
timestamp 1604681595
transform 1 0 13248 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15548 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_29_149
timestamp 1604681595
transform 1 0 14812 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_173
timestamp 1604681595
transform 1 0 17020 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1604681595
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1604681595
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_195
timestamp 1604681595
transform 1 0 19044 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_207
timestamp 1604681595
transform 1 0 20148 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 20516 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_215
timestamp 1604681595
transform 1 0 20884 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604681595
transform 1 0 2852 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_11
timestamp 1604681595
transform 1 0 2116 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_23
timestamp 1604681595
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_41
timestamp 1604681595
transform 1 0 4876 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5612 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_58
timestamp 1604681595
transform 1 0 6440 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7176 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_82
timestamp 1604681595
transform 1 0 8648 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_102
timestamp 1604681595
transform 1 0 10488 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1604681595
transform 1 0 11224 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_113
timestamp 1604681595
transform 1 0 11500 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_125
timestamp 1604681595
transform 1 0 12604 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604681595
transform 1 0 14076 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_133
timestamp 1604681595
transform 1 0 13340 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_145
timestamp 1604681595
transform 1 0 14444 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_163
timestamp 1604681595
transform 1 0 16100 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1604681595
transform 1 0 16836 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_180
timestamp 1604681595
transform 1 0 17664 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 18400 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 19688 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_191
timestamp 1604681595
transform 1 0 18676 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_199
timestamp 1604681595
transform 1 0 19412 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_206
timestamp 1604681595
transform 1 0 20056 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604681595
transform 1 0 1472 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2576 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_8
timestamp 1604681595
transform 1 0 1840 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4140 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_25
timestamp 1604681595
transform 1 0 3404 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_49
timestamp 1604681595
transform 1 0 5612 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7084 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1604681595
transform 1 0 8556 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_93
timestamp 1604681595
transform 1 0 9660 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_97
timestamp 1604681595
transform 1 0 10028 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_114
timestamp 1604681595
transform 1 0 11592 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 13708 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_129
timestamp 1604681595
transform 1 0 12972 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_141
timestamp 1604681595
transform 1 0 14076 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16100 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14812 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_155
timestamp 1604681595
transform 1 0 15364 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1604681595
transform 1 0 16652 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1604681595
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_187
timestamp 1604681595
transform 1 0 18308 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604681595
transform 1 0 19504 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_199
timestamp 1604681595
transform 1 0 19412 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_204
timestamp 1604681595
transform 1 0 19872 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 20608 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_215
timestamp 1604681595
transform 1 0 20884 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604681595
transform 1 0 2852 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_11
timestamp 1604681595
transform 1 0 2116 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_23
timestamp 1604681595
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1604681595
transform 1 0 4876 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6348 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_32_53
timestamp 1604681595
transform 1 0 5980 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 8556 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_73
timestamp 1604681595
transform 1 0 7820 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10580 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_84
timestamp 1604681595
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_101
timestamp 1604681595
transform 1 0 10396 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12144 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_112
timestamp 1604681595
transform 1 0 11408 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1604681595
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_145
timestamp 1604681595
transform 1 0 14444 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1604681595
transform 1 0 15548 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_161
timestamp 1604681595
transform 1 0 15916 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604681595
transform 1 0 17480 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_173
timestamp 1604681595
transform 1 0 17020 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_177
timestamp 1604681595
transform 1 0 17388 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_182
timestamp 1604681595
transform 1 0 17848 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 19688 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 18584 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_194
timestamp 1604681595
transform 1 0 18952 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_206
timestamp 1604681595
transform 1 0 20056 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1748 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604681595
transform 1 0 4048 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 3956 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_23
timestamp 1604681595
transform 1 0 3220 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_36
timestamp 1604681595
transform 1 0 4416 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5244 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_44
timestamp 1604681595
transform 1 0 5152 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_54
timestamp 1604681595
transform 1 0 6072 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 8464 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6900 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_33_72
timestamp 1604681595
transform 1 0 7728 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9752 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9660 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_84
timestamp 1604681595
transform 1 0 8832 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_92
timestamp 1604681595
transform 1 0 9568 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_103
timestamp 1604681595
transform 1 0 10580 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 11316 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12604 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12512 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_115
timestamp 1604681595
transform 1 0 11684 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 14168 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_134
timestamp 1604681595
transform 1 0 13432 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1604681595
transform 1 0 15548 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 15364 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_146
timestamp 1604681595
transform 1 0 14536 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_154
timestamp 1604681595
transform 1 0 15272 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_156
timestamp 1604681595
transform 1 0 15456 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_161
timestamp 1604681595
transform 1 0 15916 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16652 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 18216 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_175
timestamp 1604681595
transform 1 0 17204 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_183
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_187
timestamp 1604681595
transform 1 0 18308 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 19964 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 18584 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_194
timestamp 1604681595
transform 1 0 18952 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_202
timestamp 1604681595
transform 1 0 19688 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_209
timestamp 1604681595
transform 1 0 20332 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1604681595
transform 1 0 21160 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1604681595
transform 1 0 21528 0 1 20128
box -38 -48 130 592
<< labels >>
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 0 nsew default input
rlabel metal2 s 662 0 718 480 6 bottom_left_grid_pin_43_
port 1 nsew default input
rlabel metal2 s 1122 0 1178 480 6 bottom_left_grid_pin_44_
port 2 nsew default input
rlabel metal2 s 1582 0 1638 480 6 bottom_left_grid_pin_45_
port 3 nsew default input
rlabel metal2 s 2042 0 2098 480 6 bottom_left_grid_pin_46_
port 4 nsew default input
rlabel metal2 s 2502 0 2558 480 6 bottom_left_grid_pin_47_
port 5 nsew default input
rlabel metal2 s 2962 0 3018 480 6 bottom_left_grid_pin_48_
port 6 nsew default input
rlabel metal2 s 3422 0 3478 480 6 bottom_left_grid_pin_49_
port 7 nsew default input
rlabel metal2 s 22650 0 22706 480 6 bottom_right_grid_pin_1_
port 8 nsew default input
rlabel metal3 s 22520 11432 23000 11552 6 ccff_head
port 9 nsew default input
rlabel metal3 s 22520 19048 23000 19168 6 ccff_tail
port 10 nsew default tristate
rlabel metal3 s 0 3952 480 4072 6 chanx_left_in[0]
port 11 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[10]
port 12 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_left_in[11]
port 13 nsew default input
rlabel metal3 s 0 9664 480 9784 6 chanx_left_in[12]
port 14 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[13]
port 15 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_left_in[14]
port 16 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chanx_left_in[15]
port 17 nsew default input
rlabel metal3 s 0 11568 480 11688 6 chanx_left_in[16]
port 18 nsew default input
rlabel metal3 s 0 12112 480 12232 6 chanx_left_in[17]
port 19 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[18]
port 20 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_in[19]
port 21 nsew default input
rlabel metal3 s 0 4360 480 4480 6 chanx_left_in[1]
port 22 nsew default input
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[2]
port 23 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[3]
port 24 nsew default input
rlabel metal3 s 0 5856 480 5976 6 chanx_left_in[4]
port 25 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_left_in[5]
port 26 nsew default input
rlabel metal3 s 0 6808 480 6928 6 chanx_left_in[6]
port 27 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[7]
port 28 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[8]
port 29 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[9]
port 30 nsew default input
rlabel metal3 s 0 13472 480 13592 6 chanx_left_out[0]
port 31 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[10]
port 32 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[11]
port 33 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[12]
port 34 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[13]
port 35 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[14]
port 36 nsew default tristate
rlabel metal3 s 0 20680 480 20800 6 chanx_left_out[15]
port 37 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[16]
port 38 nsew default tristate
rlabel metal3 s 0 21632 480 21752 6 chanx_left_out[17]
port 39 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[18]
port 40 nsew default tristate
rlabel metal3 s 0 22584 480 22704 6 chanx_left_out[19]
port 41 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chanx_left_out[1]
port 42 nsew default tristate
rlabel metal3 s 0 14424 480 14544 6 chanx_left_out[2]
port 43 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[3]
port 44 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chanx_left_out[4]
port 45 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[5]
port 46 nsew default tristate
rlabel metal3 s 0 16328 480 16448 6 chanx_left_out[6]
port 47 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chanx_left_out[7]
port 48 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[8]
port 49 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[9]
port 50 nsew default tristate
rlabel metal2 s 3882 0 3938 480 6 chany_bottom_in[0]
port 51 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[10]
port 52 nsew default input
rlabel metal2 s 9034 0 9090 480 6 chany_bottom_in[11]
port 53 nsew default input
rlabel metal2 s 9586 0 9642 480 6 chany_bottom_in[12]
port 54 nsew default input
rlabel metal2 s 10046 0 10102 480 6 chany_bottom_in[13]
port 55 nsew default input
rlabel metal2 s 10506 0 10562 480 6 chany_bottom_in[14]
port 56 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[15]
port 57 nsew default input
rlabel metal2 s 11426 0 11482 480 6 chany_bottom_in[16]
port 58 nsew default input
rlabel metal2 s 11886 0 11942 480 6 chany_bottom_in[17]
port 59 nsew default input
rlabel metal2 s 12346 0 12402 480 6 chany_bottom_in[18]
port 60 nsew default input
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_in[19]
port 61 nsew default input
rlabel metal2 s 4342 0 4398 480 6 chany_bottom_in[1]
port 62 nsew default input
rlabel metal2 s 4894 0 4950 480 6 chany_bottom_in[2]
port 63 nsew default input
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_in[3]
port 64 nsew default input
rlabel metal2 s 5814 0 5870 480 6 chany_bottom_in[4]
port 65 nsew default input
rlabel metal2 s 6274 0 6330 480 6 chany_bottom_in[5]
port 66 nsew default input
rlabel metal2 s 6734 0 6790 480 6 chany_bottom_in[6]
port 67 nsew default input
rlabel metal2 s 7194 0 7250 480 6 chany_bottom_in[7]
port 68 nsew default input
rlabel metal2 s 7654 0 7710 480 6 chany_bottom_in[8]
port 69 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chany_bottom_in[9]
port 70 nsew default input
rlabel metal2 s 13266 0 13322 480 6 chany_bottom_out[0]
port 71 nsew default tristate
rlabel metal2 s 17958 0 18014 480 6 chany_bottom_out[10]
port 72 nsew default tristate
rlabel metal2 s 18418 0 18474 480 6 chany_bottom_out[11]
port 73 nsew default tristate
rlabel metal2 s 18970 0 19026 480 6 chany_bottom_out[12]
port 74 nsew default tristate
rlabel metal2 s 19430 0 19486 480 6 chany_bottom_out[13]
port 75 nsew default tristate
rlabel metal2 s 19890 0 19946 480 6 chany_bottom_out[14]
port 76 nsew default tristate
rlabel metal2 s 20350 0 20406 480 6 chany_bottom_out[15]
port 77 nsew default tristate
rlabel metal2 s 20810 0 20866 480 6 chany_bottom_out[16]
port 78 nsew default tristate
rlabel metal2 s 21270 0 21326 480 6 chany_bottom_out[17]
port 79 nsew default tristate
rlabel metal2 s 21730 0 21786 480 6 chany_bottom_out[18]
port 80 nsew default tristate
rlabel metal2 s 22190 0 22246 480 6 chany_bottom_out[19]
port 81 nsew default tristate
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_out[1]
port 82 nsew default tristate
rlabel metal2 s 14278 0 14334 480 6 chany_bottom_out[2]
port 83 nsew default tristate
rlabel metal2 s 14738 0 14794 480 6 chany_bottom_out[3]
port 84 nsew default tristate
rlabel metal2 s 15198 0 15254 480 6 chany_bottom_out[4]
port 85 nsew default tristate
rlabel metal2 s 15658 0 15714 480 6 chany_bottom_out[5]
port 86 nsew default tristate
rlabel metal2 s 16118 0 16174 480 6 chany_bottom_out[6]
port 87 nsew default tristate
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_out[7]
port 88 nsew default tristate
rlabel metal2 s 17038 0 17094 480 6 chany_bottom_out[8]
port 89 nsew default tristate
rlabel metal2 s 17498 0 17554 480 6 chany_bottom_out[9]
port 90 nsew default tristate
rlabel metal2 s 3882 22520 3938 23000 6 chany_top_in[0]
port 91 nsew default input
rlabel metal2 s 8574 22520 8630 23000 6 chany_top_in[10]
port 92 nsew default input
rlabel metal2 s 9034 22520 9090 23000 6 chany_top_in[11]
port 93 nsew default input
rlabel metal2 s 9586 22520 9642 23000 6 chany_top_in[12]
port 94 nsew default input
rlabel metal2 s 10046 22520 10102 23000 6 chany_top_in[13]
port 95 nsew default input
rlabel metal2 s 10506 22520 10562 23000 6 chany_top_in[14]
port 96 nsew default input
rlabel metal2 s 10966 22520 11022 23000 6 chany_top_in[15]
port 97 nsew default input
rlabel metal2 s 11426 22520 11482 23000 6 chany_top_in[16]
port 98 nsew default input
rlabel metal2 s 11886 22520 11942 23000 6 chany_top_in[17]
port 99 nsew default input
rlabel metal2 s 12346 22520 12402 23000 6 chany_top_in[18]
port 100 nsew default input
rlabel metal2 s 12806 22520 12862 23000 6 chany_top_in[19]
port 101 nsew default input
rlabel metal2 s 4342 22520 4398 23000 6 chany_top_in[1]
port 102 nsew default input
rlabel metal2 s 4894 22520 4950 23000 6 chany_top_in[2]
port 103 nsew default input
rlabel metal2 s 5354 22520 5410 23000 6 chany_top_in[3]
port 104 nsew default input
rlabel metal2 s 5814 22520 5870 23000 6 chany_top_in[4]
port 105 nsew default input
rlabel metal2 s 6274 22520 6330 23000 6 chany_top_in[5]
port 106 nsew default input
rlabel metal2 s 6734 22520 6790 23000 6 chany_top_in[6]
port 107 nsew default input
rlabel metal2 s 7194 22520 7250 23000 6 chany_top_in[7]
port 108 nsew default input
rlabel metal2 s 7654 22520 7710 23000 6 chany_top_in[8]
port 109 nsew default input
rlabel metal2 s 8114 22520 8170 23000 6 chany_top_in[9]
port 110 nsew default input
rlabel metal2 s 13266 22520 13322 23000 6 chany_top_out[0]
port 111 nsew default tristate
rlabel metal2 s 17958 22520 18014 23000 6 chany_top_out[10]
port 112 nsew default tristate
rlabel metal2 s 18418 22520 18474 23000 6 chany_top_out[11]
port 113 nsew default tristate
rlabel metal2 s 18970 22520 19026 23000 6 chany_top_out[12]
port 114 nsew default tristate
rlabel metal2 s 19430 22520 19486 23000 6 chany_top_out[13]
port 115 nsew default tristate
rlabel metal2 s 19890 22520 19946 23000 6 chany_top_out[14]
port 116 nsew default tristate
rlabel metal2 s 20350 22520 20406 23000 6 chany_top_out[15]
port 117 nsew default tristate
rlabel metal2 s 20810 22520 20866 23000 6 chany_top_out[16]
port 118 nsew default tristate
rlabel metal2 s 21270 22520 21326 23000 6 chany_top_out[17]
port 119 nsew default tristate
rlabel metal2 s 21730 22520 21786 23000 6 chany_top_out[18]
port 120 nsew default tristate
rlabel metal2 s 22190 22520 22246 23000 6 chany_top_out[19]
port 121 nsew default tristate
rlabel metal2 s 13726 22520 13782 23000 6 chany_top_out[1]
port 122 nsew default tristate
rlabel metal2 s 14278 22520 14334 23000 6 chany_top_out[2]
port 123 nsew default tristate
rlabel metal2 s 14738 22520 14794 23000 6 chany_top_out[3]
port 124 nsew default tristate
rlabel metal2 s 15198 22520 15254 23000 6 chany_top_out[4]
port 125 nsew default tristate
rlabel metal2 s 15658 22520 15714 23000 6 chany_top_out[5]
port 126 nsew default tristate
rlabel metal2 s 16118 22520 16174 23000 6 chany_top_out[6]
port 127 nsew default tristate
rlabel metal2 s 16578 22520 16634 23000 6 chany_top_out[7]
port 128 nsew default tristate
rlabel metal2 s 17038 22520 17094 23000 6 chany_top_out[8]
port 129 nsew default tristate
rlabel metal2 s 17498 22520 17554 23000 6 chany_top_out[9]
port 130 nsew default tristate
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_34_
port 131 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_35_
port 132 nsew default input
rlabel metal3 s 0 1096 480 1216 6 left_bottom_grid_pin_36_
port 133 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_37_
port 134 nsew default input
rlabel metal3 s 0 2048 480 2168 6 left_bottom_grid_pin_38_
port 135 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_39_
port 136 nsew default input
rlabel metal3 s 0 3000 480 3120 6 left_bottom_grid_pin_40_
port 137 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_41_
port 138 nsew default input
rlabel metal3 s 22520 3816 23000 3936 6 prog_clk
port 139 nsew default input
rlabel metal2 s 202 22520 258 23000 6 top_left_grid_pin_42_
port 140 nsew default input
rlabel metal2 s 662 22520 718 23000 6 top_left_grid_pin_43_
port 141 nsew default input
rlabel metal2 s 1122 22520 1178 23000 6 top_left_grid_pin_44_
port 142 nsew default input
rlabel metal2 s 1582 22520 1638 23000 6 top_left_grid_pin_45_
port 143 nsew default input
rlabel metal2 s 2042 22520 2098 23000 6 top_left_grid_pin_46_
port 144 nsew default input
rlabel metal2 s 2502 22520 2558 23000 6 top_left_grid_pin_47_
port 145 nsew default input
rlabel metal2 s 2962 22520 3018 23000 6 top_left_grid_pin_48_
port 146 nsew default input
rlabel metal2 s 3422 22520 3478 23000 6 top_left_grid_pin_49_
port 147 nsew default input
rlabel metal2 s 22650 22520 22706 23000 6 top_right_grid_pin_1_
port 148 nsew default input
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 149 nsew default input
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 150 nsew default input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
