* NGSPICE file created from sb_0__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxbp_1 abstract view
.subckt sky130_fd_sc_hd__dfxbp_1 D Q Q_N CLK VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A X VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VNB VPB VPWR
.ends

.subckt sb_0__1_ bottom_left_grid_pin_1_ ccff_head ccff_tail chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9]
+ chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] prog_clk right_bottom_grid_pin_34_ right_bottom_grid_pin_35_ right_bottom_grid_pin_36_
+ right_bottom_grid_pin_37_ right_bottom_grid_pin_38_ right_bottom_grid_pin_39_ right_bottom_grid_pin_40_
+ right_bottom_grid_pin_41_ top_left_grid_pin_1_ VPWR VGND
XFILLER_22_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_18.mux_l1_in_0__S mux_right_track_18.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l1_in_1_ chanx_right_in[11] chanx_right_in[4] mux_bottom_track_3.mux_l1_in_0_/S
+ mux_bottom_track_3.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l3_in_0__A0 mux_right_track_2.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_1.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__124__A _124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_12.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_36.mux_l2_in_0__A1 mux_right_track_36.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A1 chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_36.sky130_fd_sc_hd__buf_4_0_ mux_right_track_36.mux_l2_in_0_/X _067_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_track_0.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_062_ _062_/HI _062_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_6.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l3_in_0__S mux_bottom_track_1.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__119__A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0_prog_clk clkbuf_3_5_0_prog_clk/A clkbuf_3_4_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_20.mux_l2_in_0_/S
+ mux_right_track_22.mux_l1_in_0_/S mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_2.mux_l1_in_2__A1 right_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_114_ chany_bottom_in[10] chany_top_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_045_ _045_/HI _045_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l3_in_0__S mux_bottom_track_25.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_17.mux_l1_in_0_ chany_top_in[17] chany_top_in[8] mux_bottom_track_17.mux_l1_in_1_/S
+ mux_bottom_track_17.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l1_in_1__S mux_right_track_0.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l2_in_1__A1 mux_right_track_2.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_22.sky130_fd_sc_hd__buf_4_0__A mux_right_track_22.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_28.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_3.mux_l3_in_0_/X _104_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
Xmem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_28.mux_l1_in_0_/S
+ mux_right_track_28.mux_l2_in_0_/S mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A0 chanx_right_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l2_in_1__S mux_top_track_0.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l1_in_0_ chany_top_in[13] chany_top_in[4] mux_bottom_track_3.mux_l1_in_0_/S
+ mux_bottom_track_3.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_36_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_2.mux_l3_in_0__A1 mux_right_track_2.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_0__A0 mux_bottom_track_3.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_10.mux_l2_in_0__A0 right_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 top_left_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_061_ _061_/HI _061_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_14_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_5.mux_l2_in_0_/S
+ mux_bottom_track_5.mux_l3_in_0_/S mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_113_ _113_/A chany_top_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_044_ _044_/HI _044_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_24.mux_l1_in_0__S mux_top_track_24.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l3_in_0__S mux_right_track_8.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_26.mux_l2_in_0_/S
+ mux_right_track_28.mux_l1_in_0_/S mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_3.mux_l1_in_1__A1 chanx_right_in[4] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_31_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_6.mux_l1_in_1__A0 right_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_22.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_20.mux_l2_in_0__S mux_right_track_20.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_0__A1 mux_bottom_track_3.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_10.mux_l2_in_0__A1 mux_right_track_10.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_3__A0 _043_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_28.sky130_fd_sc_hd__buf_4_0__A mux_right_track_28.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0__A0 mux_right_track_6.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0__S mux_right_track_14.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_10.mux_l3_in_0_ mux_right_track_10.mux_l2_in_1_/X mux_right_track_10.mux_l2_in_0_/X
+ mux_right_track_10.mux_l3_in_0_/S mux_right_track_10.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_060_ _060_/HI _060_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0__S mux_top_track_16.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_5.mux_l1_in_0_/S
+ mux_bottom_track_5.mux_l2_in_0_/S mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_112_ chany_bottom_in[12] chany_top_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_043_ _043_/HI _043_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_right_track_10.mux_l2_in_1_ _061_/HI chany_bottom_in[9] mux_right_track_10.mux_l2_in_0_/S
+ mux_right_track_10.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__D mux_top_track_2.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_3.mux_l2_in_1__S mux_bottom_track_3.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2__S mux_bottom_track_9.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_12.mux_l3_in_0__S mux_right_track_12.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_1_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_3_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_6.mux_l1_in_1__A1 right_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1__A0 chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_3.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A mux_top_track_0.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_3__A1 chany_bottom_in[5] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_14.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_6.mux_l1_in_0__S mux_right_track_6.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_6.mux_l2_in_0__A1 mux_right_track_6.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l2_in_0__A0 mux_top_track_2.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_8.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0__A0 chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_track_14.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_14.mux_l2_in_1_/S
+ mux_right_track_14.mux_l3_in_0_/S mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_3.mux_l3_in_0_/S
+ mux_bottom_track_5.mux_l1_in_0_/S mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_111_ chany_bottom_in[13] chany_top_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_042_ _042_/HI _042_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A0 bottom_left_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_10.mux_l2_in_0_ right_bottom_grid_pin_35_ mux_right_track_10.mux_l1_in_0_/X
+ mux_right_track_10.mux_l2_in_0_/S mux_right_track_10.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_8.mux_l3_in_0_ mux_right_track_8.mux_l2_in_1_/X mux_right_track_8.mux_l2_in_0_/X
+ mux_right_track_8.mux_l3_in_0_/S mux_right_track_8.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_37_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_0_/S mux_top_track_0.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA__072__A _072_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_3_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_3_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A0 _058_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__067__A _067_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_12.mux_l2_in_1__A0 _062_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_5.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_6.mux_l1_in_3__S mux_right_track_6.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l2_in_1_ _045_/HI chany_bottom_in[8] mux_right_track_8.mux_l2_in_1_/S
+ mux_right_track_8.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_4.mux_l3_in_0__S mux_right_track_4.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1_ _046_/HI mux_top_track_0.mux_l1_in_2_/X mux_top_track_0.mux_l2_in_1_/S
+ mux_top_track_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l1_in_1__A1 chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l3_in_0__A0 mux_bottom_track_5.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_12.mux_l3_in_0__A0 mux_right_track_12.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_22.mux_l1_in_0__A0 right_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__080__A _080_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l1_in_2_ chany_bottom_in[12] chany_bottom_in[2] mux_top_track_0.mux_l1_in_2_/S
+ mux_top_track_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2__D mux_top_track_32.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l2_in_0__A1 mux_top_track_2.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l3_in_0_/X _117_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_23_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__075__A _075_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0__A1 chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_14.mux_l1_in_0_/S
+ mux_right_track_14.mux_l2_in_1_/S mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_22.mux_l1_in_1__S mux_right_track_22.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_10.mux_l1_in_0__S mux_right_track_10.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_110_ chany_bottom_in[14] chany_top_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_041_ _041_/HI _041_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_track_5.mux_l1_in_2__A1 chanx_right_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_24.mux_l2_in_1__S mux_top_track_24.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_0.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_17.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_16.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_1__A1 mux_bottom_track_5.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_12.mux_l2_in_1__A1 chany_bottom_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_33_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l3_in_0_/X _125_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA__083__A _083_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_2.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_10.mux_l1_in_0_ chany_top_in[11] chany_top_in[9] mux_right_track_10.mux_l1_in_0_/S
+ mux_right_track_10.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.mux_l2_in_0_ right_bottom_grid_pin_34_ mux_right_track_8.mux_l1_in_0_/X
+ mux_right_track_8.mux_l2_in_1_/S mux_right_track_8.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_8.mux_l2_in_1__A0 _045_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_24.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l2_in_0_ mux_top_track_0.mux_l1_in_1_/X mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_1_/S mux_top_track_0.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_22.mux_l2_in_0_ mux_right_track_22.mux_l1_in_1_/X mux_right_track_22.mux_l1_in_0_/X
+ mux_right_track_22.mux_l2_in_0_/S mux_right_track_22.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_30.mux_l1_in_0__A0 chany_bottom_in[7] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__078__A _078_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_2__S mux_bottom_track_5.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l3_in_0__A1 mux_bottom_track_5.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_12.mux_l3_in_0__A1 mux_right_track_12.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_22.mux_l1_in_0__A1 chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.mux_l3_in_0__A0 mux_right_track_8.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__S mux_bottom_track_9.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_0.mux_l1_in_1_ chanx_right_in[15] chanx_right_in[8] mux_top_track_0.mux_l1_in_2_/S
+ mux_top_track_0.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_22.mux_l1_in_1_ _035_/HI chany_bottom_in[17] mux_right_track_22.mux_l1_in_0_/S
+ mux_right_track_22.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_3.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A0 chany_top_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_14.mux_l2_in_1__S mux_right_track_14.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_1__S mux_bottom_track_17.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__091__A chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_12.mux_l3_in_0_/S
+ mux_right_track_14.mux_l1_in_0_/S mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_14.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0__S mux_right_track_2.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__086__A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_040_ _040_/HI _040_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_3_3_0_prog_clk_A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0__S mux_top_track_2.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_10.sky130_fd_sc_hd__buf_4_0_ mux_right_track_10.mux_l3_in_0_/X _080_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l1_in_2__A0 chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_8.mux_l1_in_1__S mux_top_track_8.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_14.sky130_fd_sc_hd__buf_4_0__A mux_right_track_14.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_16.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_8.mux_l2_in_1__A1 chany_bottom_in[8] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l2_in_1__A0 _051_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_30.mux_l1_in_0__A1 right_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1__A0 chanx_right_in[9] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1__A0 _064_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__094__A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_33.mux_l2_in_0_/X
+ _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A0 chany_top_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l1_in_3__S mux_right_track_2.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l3_in_0__S mux_right_track_0.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ mux_bottom_track_25.mux_l3_in_0_/S mux_bottom_track_25.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_35_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_8.mux_l1_in_0_ chany_top_in[8] chany_top_in[7] mux_right_track_8.mux_l1_in_0_/S
+ mux_right_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_8.mux_l3_in_0__A1 mux_right_track_8.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__089__A _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_4.mux_l3_in_0__A0 mux_top_track_4.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_0.mux_l1_in_0_ chanx_right_in[1] top_left_grid_pin_1_ mux_top_track_0.mux_l1_in_2_/S
+ mux_top_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_6.mux_l2_in_1__S mux_right_track_6.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_22.mux_l1_in_0_ right_bottom_grid_pin_41_ chany_top_in[17] mux_right_track_22.mux_l1_in_0_/S
+ mux_right_track_22.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_1_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A1 chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A0 mux_bottom_track_9.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_34.mux_l2_in_0_ _041_/HI mux_right_track_34.mux_l1_in_0_/X mux_right_track_34.mux_l2_in_0_/S
+ mux_right_track_34.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_16.mux_l2_in_0__A0 mux_right_track_16.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_8.sky130_fd_sc_hd__buf_4_0_ mux_right_track_8.mux_l3_in_0_/X _081_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_25.mux_l2_in_1_ _055_/HI chanx_right_in[14] mux_bottom_track_25.mux_l2_in_1_/S
+ mux_bottom_track_25.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_0_/S mux_bottom_track_9.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_099_ chany_top_in[5] chany_bottom_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_37_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_4.mux_l1_in_2__A1 chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A mux_right_track_0.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__097__A _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l2_in_1_ _059_/HI mux_bottom_track_9.mux_l1_in_2_/X mux_bottom_track_9.mux_l2_in_1_/S
+ mux_bottom_track_9.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_34.mux_l2_in_0__S mux_right_track_34.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_0.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_32.sky130_fd_sc_hd__buf_4_0_ mux_right_track_32.mux_l2_in_0_/X _069_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_40_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_ mux_top_track_0.mux_l2_in_1_/S mux_top_track_0.mux_l3_in_0_/S
+ mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_0_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A0 chanx_right_in[6] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_28.mux_l1_in_0__S mux_right_track_28.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_track_4.mux_l2_in_1__A1 mux_top_track_4.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_16.mux_l1_in_1__A0 chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_9.mux_l1_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0_prog_clk clkbuf_3_3_0_prog_clk/A clkbuf_3_2_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_right_track_16.mux_l1_in_1__A1 chany_bottom_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l1_in_2_ bottom_left_grid_pin_1_ chanx_right_in[16] mux_bottom_track_9.mux_l1_in_2_/S
+ mux_bottom_track_9.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A1 chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l2_in_0_/S mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_29_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l2_in_0__A0 chany_bottom_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_26.sky130_fd_sc_hd__buf_4_0_ mux_right_track_26.mux_l2_in_0_/X _072_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_24.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_4.mux_l3_in_0__A1 mux_top_track_4.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_16.mux_l2_in_0__A0 mux_top_track_16.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0__A1 mux_bottom_track_9.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2__S mux_bottom_track_1.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0__A1 mux_right_track_16.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_0__S mux_bottom_track_5.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l2_in_0_ mux_bottom_track_25.mux_l1_in_1_/X mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_1_/S mux_bottom_track_25.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_10.mux_l2_in_1__S mux_right_track_10.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_34.mux_l1_in_0_ chany_bottom_in[1] right_bottom_grid_pin_39_ mux_right_track_34.mux_l1_in_0_/S
+ mux_right_track_34.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_098_ chany_top_in[6] chany_bottom_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l1_in_1_ chanx_right_in[7] chanx_right_in[0] mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_9.mux_l2_in_0_ mux_bottom_track_9.mux_l1_in_1_/X mux_bottom_track_9.mux_l1_in_0_/X
+ mux_bottom_track_9.mux_l2_in_1_/S mux_bottom_track_9.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_2_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_0.mux_l1_in_2_/S mux_top_track_0.mux_l2_in_1_/S
+ mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_0_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A1 chany_top_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_32.mux_l2_in_0__A0 _040_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_1__S mux_top_track_4.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A0 right_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1__A1 chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_24.mux_l2_in_0__A0 chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_9.mux_l1_in_1_ chanx_right_in[9] chanx_right_in[2] mux_bottom_track_9.mux_l1_in_2_/S
+ mux_bottom_track_9.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_6.sky130_fd_sc_hd__buf_4_0__A mux_right_track_6.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_30.mux_l2_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/S mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.mux_l2_in_0__A1 mux_right_track_24.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1__A0 chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0__A1 mux_top_track_16.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_18.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.mux_l3_in_0_ mux_top_track_16.mux_l2_in_1_/X mux_top_track_16.mux_l2_in_0_/X
+ mux_top_track_16.mux_l3_in_0_/S mux_top_track_16.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_8.mux_l2_in_0__A0 mux_top_track_8.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A mux_right_track_32.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l2_in_1__S mux_right_track_2.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_0.mux_l2_in_1_/S mux_right_track_0.mux_l3_in_0_/S
+ mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_6_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_097_ _097_/A chany_bottom_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_16.mux_l2_in_1_ _047_/HI chany_bottom_in[17] mux_top_track_16.mux_l2_in_1_/S
+ mux_top_track_16.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_25.mux_l1_in_0_ chany_top_in[18] chany_top_in[9] mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_3_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_32.mux_l2_in_0__A0 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_ ccff_head mux_top_track_0.mux_l1_in_2_/S
+ mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_0_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_33_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_32.mux_l2_in_0__A1 mux_right_track_32.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_34.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_0__A1 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_30.mux_l2_in_0__S mux_right_track_30.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_24.mux_l2_in_0__A1 mux_top_track_24.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_33.mux_l1_in_0__S mux_bottom_track_33.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_9.mux_l1_in_0_ chany_top_in[16] chany_top_in[6] mux_bottom_track_9.mux_l1_in_2_/S
+ mux_bottom_track_9.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_21_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1__A1 chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_32.mux_l3_in_0__S mux_top_track_32.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l1_in_0__S mux_right_track_24.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l3_in_0_/X _101_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_28.mux_l1_in_0__A0 chany_bottom_in[11] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_8.mux_l2_in_0__A1 mux_top_track_8.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__100__A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_096_ chany_top_in[8] chany_bottom_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0__S mux_bottom_track_1.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_0.mux_l1_in_0_/S mux_right_track_0.mux_l2_in_1_/S
+ mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_6_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_37_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_1_/S mux_top_track_16.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_4.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_079_ _079_/A chanx_right_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_32.mux_l2_in_0__A1 mux_top_track_32.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__S mux_bottom_track_25.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_4.mux_l1_in_3_ _043_/HI chany_bottom_in[5] mux_right_track_4.mux_l1_in_1_/S
+ mux_right_track_4.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_16.mux_l1_in_1_ chany_bottom_in[8] chanx_right_in[19] mux_top_track_16.mux_l1_in_1_/S
+ mux_top_track_16.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_16.mux_l2_in_0__S mux_right_track_16.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_6.mux_l2_in_0_/S mux_right_track_6.mux_l3_in_0_/S
+ mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_7_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_28.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_36.mux_l1_in_0__A0 chany_bottom_in[0] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1__S mux_top_track_0.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__103__A _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_28.mux_l1_in_0__A1 right_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_1_0_prog_clk clkbuf_3_1_0_prog_clk/A clkbuf_3_1_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
Xmux_right_track_4.mux_l3_in_0_ mux_right_track_4.mux_l2_in_1_/X mux_right_track_4.mux_l2_in_0_/X
+ mux_right_track_4.mux_l3_in_0_/S mux_right_track_4.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_25.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l1_in_1__A0 right_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_1_ mux_right_track_4.mux_l1_in_3_/X mux_right_track_4.mux_l1_in_2_/X
+ mux_right_track_4.mux_l2_in_1_/S mux_right_track_4.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_095_ chany_top_in[9] chany_bottom_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_32.mux_l3_in_0_/S mux_right_track_0.mux_l1_in_0_/S
+ mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_6_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA__111__A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_17.mux_l3_in_0__S mux_bottom_track_17.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__D mux_top_track_8.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_2__S mux_right_track_4.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__106__A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_078_ _078_/A chanx_right_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l2_in_0__A0 mux_right_track_2.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l1_in_2_ right_bottom_grid_pin_40_ right_bottom_grid_pin_38_
+ mux_right_track_4.mux_l1_in_1_/S mux_right_track_4.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0__S mux_right_track_8.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_16.mux_l1_in_0_ chanx_right_in[12] chanx_right_in[5] mux_top_track_16.mux_l1_in_1_/S
+ mux_top_track_16.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_24.mux_l2_in_0_/S
+ mux_right_track_24.mux_l3_in_0_/S mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_6.mux_l1_in_1_/S mux_right_track_6.mux_l2_in_0_/S
+ mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_5_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_top_track_8.mux_l3_in_0__S mux_top_track_8.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_36.mux_l1_in_0__A1 right_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__114__A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_20.mux_l1_in_0__S mux_right_track_20.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_20.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__109__A _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_25.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_16.mux_l2_in_0_ mux_right_track_16.mux_l1_in_1_/X mux_right_track_16.mux_l1_in_0_/X
+ mux_right_track_16.mux_l2_in_0_/S mux_right_track_16.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1__A1 right_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l2_in_0_ mux_right_track_4.mux_l1_in_1_/X mux_right_track_4.mux_l1_in_0_/X
+ mux_right_track_4.mux_l2_in_1_/S mux_right_track_4.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_094_ chany_top_in[10] chany_bottom_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0__S mux_top_track_16.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__122__A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_077_ _077_/A chanx_right_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_33_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_16.mux_l1_in_1_ _064_/HI chany_bottom_in[13] mux_right_track_16.mux_l1_in_0_/S
+ mux_right_track_16.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l2_in_0__A1 mux_right_track_2.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_4.mux_l1_in_1_ right_bottom_grid_pin_36_ right_bottom_grid_pin_34_
+ mux_right_track_4.mux_l1_in_1_/S mux_right_track_4.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A0 chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_24.mux_l1_in_0_/S
+ mux_right_track_24.mux_l2_in_0_/S mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__D mux_top_track_0.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_1__S mux_bottom_track_3.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__117__A _117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0__A0 chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_4.mux_l3_in_0_/S mux_right_track_6.mux_l1_in_1_/S
+ mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_5_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A0 bottom_left_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l2_in_1__S mux_right_track_24.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_12.mux_l2_in_0__S mux_right_track_12.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_18.mux_l1_in_1__S mux_right_track_18.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_1.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_1__A0 _053_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__125__A _125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_12.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_1.mux_l2_in_1_/S
+ mux_bottom_track_1.mux_l3_in_0_/S mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_093_ _093_/A chany_bottom_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_6.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_17.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l3_in_0__A0 mux_bottom_track_1.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_0_prog_clk prog_clk clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_076_ _076_/A chanx_right_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_16.mux_l1_in_0_ right_bottom_grid_pin_38_ chany_top_in[13] mux_right_track_16.mux_l1_in_0_/S
+ mux_right_track_16.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_4.mux_l1_in_0_ chany_top_in[5] chany_top_in[1] mux_right_track_4.mux_l1_in_1_/S
+ mux_right_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_4_0_prog_clk_A clkbuf_3_5_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_4.sky130_fd_sc_hd__buf_4_0_ mux_right_track_4.mux_l3_in_0_/X _083_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_28.mux_l2_in_0_ _038_/HI mux_right_track_28.mux_l1_in_0_/X mux_right_track_28.mux_l2_in_0_/S
+ mux_right_track_28.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A1 chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_22.mux_l2_in_0_/S
+ mux_right_track_24.mux_l1_in_0_/S mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_10.mux_l1_in_0__A1 chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_059_ _059_/HI _059_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_right_track_30.mux_l2_in_0_ _039_/HI mux_right_track_30.mux_l1_in_0_/X mux_right_track_30.mux_l2_in_0_/S
+ mux_right_track_30.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_0.mux_l1_in_2__S mux_right_track_0.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0__A0 chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_17.mux_l3_in_0_/X
+ _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_30.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.mux_l2_in_0__S mux_right_track_4.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2__A1 chanx_right_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_7_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_0_/S mux_bottom_track_5.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_41_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l1_in_2__A0 right_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_4.mux_l3_in_0__S mux_top_track_4.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A mux_right_track_24.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_1.mux_l2_in_1__A1 mux_bottom_track_1.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l2_in_1_ _058_/HI mux_bottom_track_5.mux_l1_in_2_/X mux_bottom_track_5.mux_l2_in_0_/S
+ mux_bottom_track_5.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_1__A0 mux_right_track_4.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_prog_clk clkbuf_3_1_0_prog_clk/A clkbuf_3_0_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l2_in_1_/S mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_22.sky130_fd_sc_hd__buf_4_0_ mux_right_track_22.mux_l2_in_0_/X _074_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
X_092_ chany_top_in[12] chany_bottom_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_5_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_track_1.mux_l3_in_0__A1 mux_bottom_track_1.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_5.mux_l1_in_2_ bottom_left_grid_pin_1_ chanx_right_in[17] mux_bottom_track_5.mux_l1_in_0_/S
+ mux_bottom_track_5.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_075_ _075_/A chanx_right_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_4.mux_l3_in_0__A0 mux_right_track_4.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_16.sky130_fd_sc_hd__buf_4_0_ mux_right_track_16.mux_l2_in_0_/X _077_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_058_ _058_/HI _058_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l1_in_0__A1 chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A0 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_28.mux_l1_in_0_ chany_bottom_in[11] right_bottom_grid_pin_36_ mux_right_track_28.mux_l1_in_0_/S
+ mux_right_track_28.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_0.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.mux_l1_in_2__A1 right_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2__A0 chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_30.mux_l1_in_0_ chany_bottom_in[7] right_bottom_grid_pin_37_ mux_right_track_30.mux_l1_in_0_/S
+ mux_right_track_30.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__S mux_bottom_track_9.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_0_/S mux_bottom_track_5.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_10.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_10.mux_l2_in_0_/S
+ mux_right_track_10.mux_l3_in_0_/S mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_9_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_1__A1 mux_right_track_4.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l2_in_1__A0 _046_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_1.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_091_ chany_top_in[13] chany_bottom_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_36.mux_l2_in_0_/S
+ mux_bottom_track_1.mux_l1_in_1_/S mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_1__A0 chanx_right_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l2_in_1__S mux_top_track_16.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_5.mux_l1_in_1_ chanx_right_in[10] chanx_right_in[3] mux_bottom_track_5.mux_l1_in_0_/S
+ mux_bottom_track_5.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_12.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_074_ _074_/A chanx_right_out[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_4.mux_l3_in_0__A1 mux_right_track_4.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__S mux_top_track_2.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_0.mux_l3_in_0__A0 mux_top_track_0.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_6.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A0 mux_bottom_track_5.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_12.mux_l2_in_0__A0 right_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_1.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_057_ _057_/HI _057_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_3_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_109_ _109_/A chany_top_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA__070__A _070_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2__A1 chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0__S mux_right_track_0.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_20.mux_l1_in_1__A0 _034_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l1_in_1__S mux_right_track_6.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_10.mux_l1_in_0_/S
+ mux_right_track_10.mux_l2_in_0_/S mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_top_track_0.mux_l3_in_0__S mux_top_track_0.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_33.mux_l2_in_0_ mux_bottom_track_33.mux_l1_in_1_/X mux_bottom_track_33.mux_l1_in_0_/X
+ ccff_tail mux_bottom_track_33.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_0.mux_l2_in_1__A1 mux_top_track_0.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_090_ chany_top_in[14] chany_bottom_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_1__A1 chanx_right_in[3] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A mux_top_track_2.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l3_in_0_/X _103_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_20.mux_l2_in_0__A0 mux_right_track_20.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l1_in_0_ chany_top_in[14] chany_top_in[5] mux_bottom_track_5.mux_l1_in_0_/S
+ mux_bottom_track_5.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_27_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_33.mux_l1_in_1_ _057_/HI chanx_right_in[13] mux_bottom_track_33.mux_l1_in_1_/S
+ mux_bottom_track_33.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_073_ _073_/A chanx_right_out[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_24.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l3_in_0__A1 mux_top_track_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_5.mux_l2_in_0__A1 mux_bottom_track_5.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_6.mux_l1_in_3__A0 _044_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__073__A _073_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_12.mux_l2_in_0__A1 mux_right_track_12.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_125_ _125_/A chany_top_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_8.mux_l2_in_0__A0 right_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_34.mux_l1_in_0__S mux_right_track_34.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_056_ _056_/HI _056_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2_ mux_top_track_32.mux_l2_in_0_/S mux_top_track_32.mux_l3_in_0_/S
+ mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_3_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA__068__A _068_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_32.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_108_ chany_bottom_in[16] chany_top_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_039_ _039_/HI _039_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_20.mux_l1_in_1__A1 chany_bottom_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__081__A _081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l3_in_0_ mux_top_track_24.mux_l2_in_1_/X mux_top_track_24.mux_l2_in_0_/X
+ mux_top_track_24.mux_l3_in_0_/S mux_top_track_24.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_8.mux_l3_in_0_/S mux_right_track_10.mux_l1_in_0_/S
+ mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_5_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_22.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__076__A _076_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__S mux_bottom_track_5.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_20.mux_l2_in_0__A1 mux_right_track_20.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_1__A0 chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l2_in_1_ _049_/HI chany_bottom_in[18] mux_top_track_24.mux_l2_in_0_/S
+ mux_top_track_24.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_33.mux_l1_in_0_ chanx_right_in[6] chany_top_in[10] mux_bottom_track_33.mux_l1_in_1_/S
+ mux_bottom_track_33.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_2_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_072_ _072_/A chanx_right_out[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_10.sky130_fd_sc_hd__buf_4_0__A mux_right_track_10.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_26.mux_l2_in_0__S mux_right_track_26.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_16.mux_l1_in_0_/S
+ mux_right_track_16.mux_l2_in_0_/S mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_24_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_6.mux_l1_in_3__A1 chany_bottom_in[6] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_124_ _124_/A chany_top_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0__A1 mux_right_track_8.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_055_ _055_/HI _055_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_right_track_12.mux_l3_in_0_ mux_right_track_12.mux_l2_in_1_/X mux_right_track_12.mux_l2_in_0_/X
+ mux_right_track_12.mux_l3_in_0_/S mux_right_track_12.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l2_in_0__A0 mux_top_track_4.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l3_in_0_ mux_right_track_0.mux_l2_in_1_/X mux_right_track_0.mux_l2_in_0_/X
+ mux_right_track_0.mux_l3_in_0_/S mux_right_track_0.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A mux_top_track_8.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_32.mux_l1_in_0_/S mux_top_track_32.mux_l2_in_0_/S
+ mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_3_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_29_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A0 chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A0 right_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__084__A _084_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_4.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_107_ chany_bottom_in[17] chany_top_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_038_ _038_/HI _038_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_7_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__079__A _079_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_12.mux_l2_in_1_ _062_/HI chany_bottom_in[10] mux_right_track_12.mux_l2_in_0_/S
+ mux_right_track_12.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_4_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_0.mux_l2_in_1_ _060_/HI mux_right_track_0.mux_l1_in_2_/X mux_right_track_0.mux_l2_in_1_/S
+ mux_right_track_0.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_3.mux_l3_in_0__S mux_bottom_track_3.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_1__S mux_bottom_track_9.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_right_track_14.mux_l2_in_1__A0 _063_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l1_in_2_ chany_bottom_in[2] right_bottom_grid_pin_40_ mux_right_track_0.mux_l1_in_0_/S
+ mux_right_track_0.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__092__A chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_16.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_2.mux_l1_in_1__S mux_right_track_2.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l2_in_0_ chany_bottom_in[9] mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_0_/S mux_top_track_24.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l1_in_1__A1 chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__087__A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_071_ _071_/A chanx_right_out[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_2_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_2.mux_l2_in_1__S mux_top_track_2.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_14.mux_l3_in_0__A0 mux_right_track_14.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_14.mux_l3_in_0_/S
+ mux_right_track_16.mux_l1_in_0_/S mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_24.mux_l1_in_0__A0 right_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2__S mux_top_track_8.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_123_ _123_/A chany_top_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_054_ _054_/HI _054_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_4.mux_l2_in_0__A1 mux_top_track_4.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0__A0 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_24.mux_l3_in_0_/S mux_top_track_32.mux_l1_in_0_/S
+ mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_3_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_37_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A1 chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0__A1 chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2__D mux_top_track_16.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_106_ chany_bottom_in[18] chany_top_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_037_ _037_/HI _037_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_30.mux_l1_in_0__S mux_right_track_30.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A mux_right_track_16.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_32.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_12.mux_l2_in_0_ right_bottom_grid_pin_36_ mux_right_track_12.mux_l1_in_0_/X
+ mux_right_track_12.mux_l2_in_0_/S mux_right_track_12.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__095__A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_0.mux_l2_in_0_ mux_right_track_0.mux_l1_in_1_/X mux_right_track_0.mux_l1_in_0_/X
+ mux_right_track_0.mux_l2_in_1_/S mux_right_track_0.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_0_/S mux_top_track_2.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l3_in_0_ mux_right_track_24.mux_l2_in_1_/X mux_right_track_24.mux_l2_in_0_/X
+ mux_right_track_24.mux_l3_in_0_/S mux_right_track_24.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_32.mux_l2_in_0__S mux_top_track_32.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_14.mux_l2_in_1__A1 chany_bottom_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_right_track_0.mux_l1_in_1_ right_bottom_grid_pin_38_ right_bottom_grid_pin_36_
+ mux_right_track_0.mux_l1_in_0_/S mux_right_track_0.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_1_ _048_/HI chany_bottom_in[13] mux_top_track_2.mux_l2_in_1_/S
+ mux_top_track_2.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_1_ _036_/HI chany_bottom_in[19] mux_right_track_24.mux_l2_in_0_/S
+ mux_right_track_24.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_32.mux_l1_in_0__A0 chany_bottom_in[3] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_070_ _070_/A chanx_right_out[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_24.mux_l1_in_0__A0 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l3_in_0_/X _113_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_14.mux_l3_in_0__A1 mux_right_track_14.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__S mux_bottom_track_1.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.mux_l1_in_0__A1 chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__098__A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_122_ chany_bottom_in[2] chany_top_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_053_ _053_/HI _053_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_24.mux_l1_in_0_ chanx_right_in[13] chanx_right_in[6] mux_top_track_24.mux_l1_in_0_/S
+ mux_top_track_24.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_16.mux_l1_in_0__A1 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_22.mux_l2_in_0__S mux_right_track_22.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__S mux_bottom_track_25.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A mux_right_track_2.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_105_ _105_/A chany_bottom_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_24.mux_l3_in_0__S mux_top_track_24.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_036_ _036_/HI _036_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_track_16.mux_l1_in_0__S mux_right_track_16.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_ mux_top_track_2.mux_l2_in_1_/S mux_top_track_2.mux_l3_in_0_/S
+ mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_1_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_track_0.sky130_fd_sc_hd__buf_4_0_ mux_right_track_0.mux_l3_in_0_/X _085_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_26.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_1__A0 _054_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_12.mux_l1_in_0_ chany_top_in[15] chany_top_in[10] mux_right_track_12.mux_l1_in_0_/S
+ mux_right_track_12.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_34.mux_l1_in_0_/S
+ mux_right_track_34.mux_l2_in_0_/S mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_right_track_0.mux_l1_in_0_ right_bottom_grid_pin_34_ chany_top_in[2] mux_right_track_0.mux_l1_in_0_/S
+ mux_right_track_0.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_32.mux_l1_in_0__A0 chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_prog_clk_A clkbuf_3_1_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_1_/S mux_top_track_2.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l2_in_0_ chany_bottom_in[18] mux_right_track_24.mux_l1_in_0_/X
+ mux_right_track_24.mux_l2_in_0_/S mux_right_track_24.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l3_in_0_/X _124_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l2_in_1__S mux_bottom_track_5.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_32.mux_l1_in_0__A1 right_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_17.mux_l3_in_0__A0 mux_bottom_track_17.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_18.mux_l1_in_1__A0 _065_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_24.mux_l1_in_0__A1 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_33.mux_l1_in_1_/S
+ ccff_tail mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_14.mux_l3_in_0__S mux_right_track_14.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_0_/S mux_bottom_track_1.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l1_in_1_ chany_bottom_in[4] chanx_right_in[16] mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_32_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_17.mux_l2_in_0__S mux_bottom_track_17.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_121_ _121_/A chany_top_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_23_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_052_ _052_/HI _052_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_18.mux_l2_in_0__A0 mux_right_track_18.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_8.mux_l1_in_0__S mux_right_track_8.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_4.mux_l1_in_2__S mux_top_track_4.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_035_ _035_/HI _035_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
X_104_ _104_/A chany_bottom_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l2_in_1_ _053_/HI mux_bottom_track_1.mux_l1_in_2_/X mux_bottom_track_1.mux_l2_in_1_/S
+ mux_bottom_track_1.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 top_left_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_34_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_5_0_prog_clk_A clkbuf_3_5_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_25.mux_l2_in_1__A0 _055_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_8.mux_l2_in_0__S mux_top_track_8.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_2.mux_l1_in_1_/S mux_top_track_2.mux_l2_in_1_/S
+ mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_1_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_12.sky130_fd_sc_hd__buf_4_0_ mux_right_track_12.mux_l3_in_0_/X _079_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_1__A1 chanx_right_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l1_in_2_ bottom_left_grid_pin_1_ chanx_right_in[19] mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_9_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l3_in_0__A0 mux_bottom_track_25.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A mux_right_track_8.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_32.mux_l2_in_0_/S
+ mux_right_track_34.mux_l1_in_0_/S mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_32.mux_l1_in_0__A1 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2_ mux_top_track_8.mux_l2_in_0_/S mux_top_track_8.mux_l3_in_0_/S
+ mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_6_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_17.mux_l3_in_0__A1 mux_bottom_track_17.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_18.mux_l1_in_1__A1 chany_bottom_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_42_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_25.mux_l3_in_0_/S
+ mux_bottom_track_33.mux_l1_in_1_/S mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_26.mux_l2_in_0__A0 _037_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_6.mux_l3_in_0__S mux_right_track_6.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_2.mux_l1_in_0_ chanx_right_in[9] chanx_right_in[2] mux_top_track_2.mux_l1_in_1_/S
+ mux_top_track_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_24.mux_l1_in_0_ right_bottom_grid_pin_34_ chany_top_in[18] mux_right_track_24.mux_l1_in_0_/S
+ mux_right_track_24.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_34.sky130_fd_sc_hd__buf_4_0__A mux_right_track_34.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2_ mux_top_track_24.mux_l2_in_0_/S mux_top_track_24.mux_l3_in_0_/S
+ mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_3_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_120_ chany_bottom_in[4] chany_top_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_36.mux_l2_in_0_ _042_/HI mux_right_track_36.mux_l1_in_0_/X mux_right_track_36.mux_l2_in_0_/S
+ mux_right_track_36.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_051_ _051_/HI _051_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_18.mux_l2_in_0__A1 mux_right_track_18.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_2.mux_l2_in_0_/S mux_right_track_2.mux_l3_in_0_/S
+ mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_6_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_034_ _034_/HI _034_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_36.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_103_ _103_/A chany_bottom_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_1_/S mux_bottom_track_1.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_25.mux_l2_in_1__A1 chanx_right_in[14] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_33.mux_l1_in_1__S mux_bottom_track_33.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_0.mux_l3_in_0_/S mux_top_track_2.mux_l1_in_1_/S
+ mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_0_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_6_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_12.mux_l1_in_0__S mux_right_track_12.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_1.mux_l1_in_1_ chanx_right_in[12] chanx_right_in[5] mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_25.mux_l3_in_0__A1 mux_bottom_track_25.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_34.sky130_fd_sc_hd__buf_4_0_ mux_right_track_34.mux_l2_in_0_/X _068_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mux_right_track_34.mux_l2_in_0__A0 _041_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0__A0 chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__101__A _101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_8.mux_l1_in_2_/S mux_top_track_8.mux_l2_in_0_/S
+ mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_4_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_35_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_26.mux_l2_in_0__A1 mux_right_track_26.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_10.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2__A0 chany_bottom_in[2] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_1__S mux_bottom_track_1.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_28.sky130_fd_sc_hd__buf_4_0_ mux_right_track_28.mux_l2_in_0_/X _071_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_24.mux_l1_in_0_/S mux_top_track_24.mux_l2_in_0_/S
+ mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_3_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_050_ _050_/HI _050_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A mux_top_track_32.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_25.mux_l2_in_1__S mux_bottom_track_25.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_10.mux_l3_in_0__S mux_right_track_10.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_2.mux_l1_in_1_/S mux_right_track_2.mux_l2_in_0_/S
+ mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_4_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_0.mux_l2_in_1__A0 _060_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l3_in_0_/X _105_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_11_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_102_ chany_top_in[2] chany_bottom_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_033_ _033_/HI _033_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_36.mux_l1_in_0_ chany_bottom_in[0] right_bottom_grid_pin_40_ mux_right_track_36.mux_l1_in_0_/S
+ mux_right_track_36.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_4.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_4.mux_l1_in_0__S mux_right_track_4.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__104__A _104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2__S mux_top_track_0.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A0 mux_right_track_0.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l1_in_0_ chany_top_in[12] chany_top_in[2] mux_bottom_track_1.mux_l1_in_1_/S
+ mux_bottom_track_1.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_4.mux_l2_in_0__S mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_8.mux_l2_in_1_/S mux_right_track_8.mux_l3_in_0_/S
+ mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_5_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_33.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_34.mux_l2_in_0__A1 mux_right_track_34.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_5.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0__A1 chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_4.mux_l3_in_0_/S mux_top_track_8.mux_l1_in_2_/S
+ mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_4_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_0.mux_l1_in_2__A1 right_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__112__A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_16.mux_l3_in_0_/S mux_top_track_24.mux_l1_in_0_/S
+ mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_3_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__107__A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_3__S mux_right_track_4.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_20.mux_l1_in_1_/S
+ mux_right_track_20.mux_l2_in_0_/S mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_2.mux_l3_in_0__S mux_right_track_2.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_0.mux_l3_in_0_/S mux_right_track_2.mux_l1_in_1_/S
+ mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_6_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l2_in_1__A1 mux_right_track_0.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l2_in_1__S mux_right_track_8.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_101_ _101_/A chany_bottom_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A0 chanx_right_in[12] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__120__A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l3_in_0__A1 mux_right_track_0.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A0 mux_bottom_track_1.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_8.mux_l1_in_0_/S mux_right_track_8.mux_l2_in_1_/S
+ mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_5_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__D ccff_head VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__115__A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_20.mux_l1_in_1__S mux_right_track_20.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_36.mux_l2_in_0__S mux_right_track_36.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_25.mux_l2_in_1_/S
+ mux_bottom_track_25.mux_l3_in_0_/S mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_25.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_16.mux_l1_in_1__S mux_top_track_16.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_36.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__123__A _123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_18.mux_l2_in_0_/S
+ mux_right_track_20.mux_l1_in_1_/S mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_37_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_10.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_100_ chany_top_in[4] chany_bottom_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_11_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__118__A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_4.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_9.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1__A1 chanx_right_in[5] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_4.mux_l1_in_1__A0 right_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_20.sky130_fd_sc_hd__buf_4_0__A mux_right_track_20.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_12.mux_l2_in_1__S mux_right_track_12.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_26.mux_l1_in_0_/S
+ mux_right_track_26.mux_l2_in_0_/S mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_6.mux_l3_in_0_/S mux_right_track_8.mux_l1_in_0_/S
+ mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_5_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_0_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0__A1 mux_bottom_track_1.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_32.mux_l3_in_0_ mux_top_track_32.mux_l2_in_1_/X mux_top_track_32.mux_l2_in_0_/X
+ mux_top_track_32.mux_l3_in_0_/S mux_top_track_32.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_2.mux_l1_in_3__A0 _033_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_6.mux_l1_in_3_ _044_/HI chany_bottom_in[6] mux_right_track_6.mux_l1_in_1_/S
+ mux_right_track_6.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_4.mux_l2_in_0__A0 mux_right_track_4.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0__S mux_right_track_0.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_0.mux_l2_in_0__S mux_top_track_0.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_25.mux_l1_in_0_/S
+ mux_bottom_track_25.mux_l2_in_1_/S mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_35_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_32.mux_l2_in_1_ _050_/HI chany_bottom_in[10] mux_top_track_32.mux_l2_in_0_/S
+ mux_top_track_32.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_6.mux_l3_in_0_ mux_right_track_6.mux_l2_in_1_/X mux_right_track_6.mux_l2_in_0_/X
+ mux_right_track_6.mux_l3_in_0_/S mux_right_track_6.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_3.mux_l2_in_1_/S
+ mux_bottom_track_3.mux_l3_in_0_/S mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_6.mux_l2_in_1_ mux_right_track_6.mux_l1_in_3_/X mux_right_track_6.mux_l1_in_2_/X
+ mux_right_track_6.mux_l2_in_0_/S mux_right_track_6.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_4.mux_l1_in_1__A1 right_bottom_grid_pin_34_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1__A0 chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_4.mux_l2_in_1__S mux_right_track_4.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_24.mux_l3_in_0_/S
+ mux_right_track_26.mux_l1_in_0_/S mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_4_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_3__A1 chany_bottom_in[4] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_8_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_6.mux_l1_in_2_ right_bottom_grid_pin_41_ right_bottom_grid_pin_39_
+ mux_right_track_6.mux_l1_in_1_/S mux_right_track_6.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_4.mux_l2_in_0__A1 mux_right_track_4.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0__A0 mux_top_track_0.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A0 chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0__A0 chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_17.mux_l3_in_0_/S
+ mux_bottom_track_25.mux_l1_in_0_/S mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_35_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_32.mux_l2_in_0_ chanx_right_in[14] mux_top_track_32.mux_l1_in_0_/X
+ mux_top_track_32.mux_l2_in_0_/S mux_top_track_32.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_26.sky130_fd_sc_hd__buf_4_0__A mux_right_track_26.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_20.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2_ mux_top_track_16.mux_l2_in_1_/S mux_top_track_16.mux_l3_in_0_/S
+ mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_3_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_32.mux_l2_in_0__S mux_right_track_32.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_26.mux_l1_in_0__S mux_right_track_26.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_3.mux_l1_in_0_/S
+ mux_bottom_track_3.mux_l2_in_1_/S mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_3_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_9_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_0_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A0 _056_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_10.mux_l2_in_1__A0 _061_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_18.mux_l2_in_0_ mux_right_track_18.mux_l1_in_1_/X mux_right_track_18.mux_l1_in_0_/X
+ mux_right_track_18.mux_l2_in_0_/S mux_right_track_18.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
X_089_ _089_/A chany_bottom_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_6.mux_l2_in_0_ mux_right_track_6.mux_l1_in_1_/X mux_right_track_6.mux_l1_in_0_/X
+ mux_right_track_6.mux_l2_in_0_/S mux_right_track_6.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_33_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_0_/S mux_top_track_8.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_20.mux_l2_in_0_ mux_right_track_20.mux_l1_in_1_/X mux_right_track_20.mux_l1_in_0_/X
+ mux_right_track_20.mux_l2_in_0_/S mux_right_track_20.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_0.mux_l1_in_1__A1 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_0_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l3_in_0__A0 mux_bottom_track_3.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_10.mux_l3_in_0__A0 mux_right_track_10.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_2.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_9.mux_l2_in_1_/S
+ mux_bottom_track_9.mux_l3_in_0_/S mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_20.mux_l1_in_0__A0 right_bottom_grid_pin_40_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_18.mux_l1_in_1_ _065_/HI chany_bottom_in[14] mux_right_track_18.mux_l1_in_1_/S
+ mux_right_track_18.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_3.mux_l2_in_0__S mux_bottom_track_3.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_6.mux_l1_in_1_ right_bottom_grid_pin_37_ right_bottom_grid_pin_35_
+ mux_right_track_6.mux_l1_in_1_/S mux_right_track_6.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_8.mux_l2_in_1_ _052_/HI mux_top_track_8.mux_l1_in_2_/X mux_top_track_8.mux_l2_in_0_/S
+ mux_top_track_8.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_20.mux_l1_in_1_ _034_/HI chany_bottom_in[16] mux_right_track_20.mux_l1_in_1_/S
+ mux_right_track_20.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_0.mux_l2_in_0__A1 mux_top_track_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_1__S mux_bottom_track_9.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_7_0_prog_clk clkbuf_3_7_0_prog_clk/A clkbuf_3_7_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A1 chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0__A1 chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l3_in_0__S mux_right_track_24.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A0 chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_3.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_8.mux_l1_in_2_ chany_bottom_in[16] chany_bottom_in[6] mux_top_track_8.mux_l1_in_2_/S
+ mux_top_track_8.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_16.mux_l1_in_1_/S mux_top_track_16.mux_l2_in_1_/S
+ mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_3_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_18.mux_l2_in_0__S mux_right_track_18.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A mux_top_track_24.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_1_0_prog_clk_A clkbuf_3_1_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_12.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_12.mux_l2_in_0_/S
+ mux_right_track_12.mux_l3_in_0_/S mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_23_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_6.mux_l1_in_2__A0 right_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l1_in_1__S mux_top_track_2.mux_l1_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_32.mux_l1_in_0_ chanx_right_in[7] chanx_right_in[0] mux_top_track_32.mux_l1_in_0_/S
+ mux_top_track_32.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_1.mux_l3_in_0_/S
+ mux_bottom_track_3.mux_l1_in_0_/S mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_1_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_8.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_3.mux_l2_in_1__A1 chanx_right_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_10.mux_l2_in_1__A1 chany_bottom_in[9] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_34_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_6.mux_l2_in_1__A0 mux_right_track_6.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_088_ chany_top_in[16] chany_bottom_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_3.mux_l3_in_0__A1 mux_bottom_track_3.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_10.mux_l3_in_0__A1 mux_right_track_10.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_3.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_20.mux_l1_in_0__A1 chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_9.mux_l1_in_2_/S
+ mux_bottom_track_9.mux_l2_in_1_/S mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__071__A _071_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_18.mux_l1_in_0_ right_bottom_grid_pin_39_ chany_top_in[14] mux_right_track_18.mux_l1_in_1_/S
+ mux_right_track_18.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_right_track_6.mux_l3_in_0__A0 mux_right_track_6.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_6.mux_l1_in_0_ chany_top_in[6] chany_top_in[3] mux_right_track_6.mux_l1_in_1_/S
+ mux_right_track_6.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_32.mux_l1_in_0__S mux_top_track_32.mux_l1_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_prog_clk_A clkbuf_3_7_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_8.mux_l2_in_0_ mux_top_track_8.mux_l1_in_1_/X mux_top_track_8.mux_l1_in_0_/X
+ mux_top_track_8.mux_l2_in_0_/S mux_top_track_8.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l3_in_0_/X
+ _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_30.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l2_in_1__S mux_right_track_0.mux_l2_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_20.mux_l1_in_0_ right_bottom_grid_pin_40_ chany_top_in[16] mux_right_track_20.mux_l1_in_1_/S
+ mux_right_track_20.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__066__A right_bottom_grid_pin_41_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_right_track_6.sky130_fd_sc_hd__buf_4_0_ mux_right_track_6.mux_l3_in_0_/X _082_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_30_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_track_32.mux_l2_in_0_ _040_/HI mux_right_track_32.mux_l1_in_0_/X mux_right_track_32.mux_l2_in_0_/S
+ mux_right_track_32.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_6.mux_l1_in_2__S mux_right_track_6.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0__A1 chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_1_ chanx_right_in[18] chanx_right_in[11] mux_top_track_8.mux_l1_in_2_/S
+ mux_top_track_8.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_8.mux_l3_in_0_/S mux_top_track_16.mux_l1_in_1_/S
+ mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_3_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l3_in_0_/X _121_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_17_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_12.mux_l1_in_0_/S
+ mux_right_track_12.mux_l2_in_0_/S mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_6.mux_l1_in_2__A1 right_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_32.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A mux_top_track_4.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_30.sky130_fd_sc_hd__buf_4_0_ mux_right_track_30.mux_l2_in_0_/X _070_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA__074__A _074_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_087_ chany_top_in[17] chany_bottom_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_6.mux_l2_in_1__A1 mux_right_track_6.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l2_in_1__A0 _048_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_22.mux_l1_in_0__S mux_right_track_22.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__069__A _069_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_24.mux_l2_in_0__S mux_top_track_24.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_0.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_24.sky130_fd_sc_hd__buf_4_0_ mux_right_track_24.mux_l3_in_0_/X _073_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_5.mux_l3_in_0_/S
+ mux_bottom_track_9.mux_l1_in_2_/S mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_9_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_6.mux_l3_in_0__A1 mux_right_track_6.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l3_in_0__A0 mux_top_track_2.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2_ mux_bottom_track_17.mux_l2_in_1_/S
+ mux_bottom_track_17.mux_l3_in_0_/S mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2_/Q_N
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_38_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_14.mux_l2_in_0__A0 right_bottom_grid_pin_37_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_18.sky130_fd_sc_hd__buf_4_0_ mux_right_track_18.mux_l2_in_0_/X _076_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__082__A _082_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_24.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 top_left_grid_pin_1_ VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__077__A _077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_9.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmux_top_track_8.mux_l1_in_0_ chanx_right_in[4] top_left_grid_pin_1_ mux_top_track_8.mux_l1_in_2_/S
+ mux_top_track_8.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_1_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_5.mux_l1_in_1__S mux_bottom_track_5.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_10.mux_l3_in_0_/S
+ mux_right_track_12.mux_l1_in_0_/S mem_right_track_12.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_5_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_right_track_32.mux_l1_in_0_ chany_bottom_in[3] right_bottom_grid_pin_38_ mux_right_track_32.mux_l1_in_0_/S
+ mux_right_track_32.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_14.mux_l2_in_0__S mux_right_track_14.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0__S mux_bottom_track_17.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_22.mux_l1_in_1__A0 _035_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_0_0_prog_clk_A clkbuf_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__090__A chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2__D mux_top_track_24.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l3_in_0__S mux_top_track_16.mux_l3_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_086_ chany_top_in[18] chany_bottom_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l2_in_1__A1 chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_12.sky130_fd_sc_hd__buf_4_0__A mux_right_track_12.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__085__A _085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_18.mux_l1_in_1_/S
+ mux_right_track_18.mux_l2_in_0_/S mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_3_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__D mux_top_track_4.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_069_ _069_/A chanx_right_out[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_22.mux_l2_in_0__A0 mux_right_track_22.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_8.mux_l1_in_0__S mux_top_track_8.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_2.mux_l3_in_0__A1 mux_top_track_2.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1_ mux_bottom_track_17.mux_l1_in_1_/S
+ mux_bottom_track_17.mux_l2_in_1_/S mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_14.mux_l2_in_0__A1 mux_right_track_14.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__D mux_top_track_8.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__D mux_bottom_track_5.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__093__A _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l1_in_2__S mux_right_track_2.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_6_0_prog_clk clkbuf_3_7_0_prog_clk/A clkbuf_3_6_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_23_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__088__A chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_6.mux_l2_in_0__S mux_right_track_6.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_22.mux_l1_in_1__A1 chany_bottom_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_30.mux_l2_in_0__A0 _039_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A0 chanx_right_in[8] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_085_ _085_/A chanx_right_out[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_18_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_16.mux_l2_in_0_/S
+ mux_right_track_18.mux_l1_in_1_/S mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_7_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_068_ _068_/A chanx_right_out[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_22.mux_l2_in_0__A1 mux_right_track_22.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxbp_1_1__D mux_right_track_34.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0__A0 mux_bottom_track_17.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__096__A chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_32.mux_l2_in_1__S mux_top_track_32.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0_ mux_bottom_track_9.mux_l3_in_0_/S
+ mux_bottom_track_17.mux_l1_in_1_/S mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_38_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_30.mux_l1_in_0_/S
+ mux_right_track_30.mux_l2_in_0_/S mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_18.sky130_fd_sc_hd__buf_4_0__A mux_right_track_18.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_18.mux_l1_in_0__A0 right_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_33.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_2__A0 bottom_left_grid_pin_1_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_25.mux_l1_in_1__A0 chanx_right_in[7] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_2_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_1__S mux_bottom_track_1.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__099__A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_30.mux_l2_in_0__A1 mux_right_track_30.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_1__A1 chanx_right_in[1] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_084_ _084_/A chanx_right_out[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_3_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l1_in_3_ _033_/HI chany_bottom_in[4] mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_3_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_9.mux_l2_in_1__A0 _059_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__D mux_right_track_2.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l1_in_1__S mux_bottom_track_25.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A0 mux_bottom_track_25.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_10.mux_l2_in_0__S mux_right_track_10.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_067_ _067_/A chanx_right_out[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_16.mux_l1_in_1__S mux_right_track_16.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0__A1 mux_bottom_track_17.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l3_in_0__A0 mux_bottom_track_9.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_119_ chany_bottom_in[5] chany_top_out[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_right_track_26.mux_l1_in_0__A0 chany_bottom_in[15] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A mux_right_track_4.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_28.mux_l2_in_0_/S
+ mux_right_track_30.mux_l1_in_0_/S mem_right_track_30.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_0_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
Xmux_right_track_14.mux_l3_in_0_ mux_right_track_14.mux_l2_in_1_/X mux_right_track_14.mux_l2_in_0_/X
+ mux_right_track_14.mux_l3_in_0_/S mux_right_track_14.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_2.mux_l3_in_0_ mux_right_track_2.mux_l2_in_1_/X mux_right_track_2.mux_l2_in_0_/X
+ mux_right_track_2.mux_l3_in_0_/S mux_right_track_2.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_29_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_4.mux_l1_in_0__S mux_top_track_4.mux_l1_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A mux_top_track_16.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_ mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l3_in_0_/S
+ mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_1_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_right_track_18.mux_l1_in_0__A1 chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_33.mux_l1_in_1__A0 _057_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_14.mux_l2_in_1_ _063_/HI chany_bottom_in[12] mux_right_track_14.mux_l2_in_1_/S
+ mux_right_track_14.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l2_in_1_ mux_right_track_2.mux_l1_in_3_/X mux_right_track_2.mux_l1_in_2_/X
+ mux_right_track_2.mux_l2_in_0_/S mux_right_track_2.mux_l2_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2__A1 chanx_right_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_39_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_30.sky130_fd_sc_hd__buf_4_0__A mux_right_track_30.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_bottom_track_9.mux_l3_in_0__S mux_bottom_track_9.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_36.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_36.mux_l1_in_0_/S
+ mux_right_track_36.mux_l2_in_0_/S mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_bottom_track_25.mux_l1_in_1__A1 chanx_right_in[0] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_33.mux_l2_in_0__A0 mux_bottom_track_33.mux_l1_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_24.mux_l2_in_1__A0 _036_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_17.mux_l2_in_1__S mux_bottom_track_17.mux_l2_in_1_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_16.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_16.mux_l2_in_1__A0 _047_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_083_ _083_/A chanx_right_out[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
Xmux_right_track_2.mux_l1_in_2_ right_bottom_grid_pin_41_ right_bottom_grid_pin_39_
+ mux_right_track_2.mux_l1_in_1_/S mux_right_track_2.mux_l1_in_2_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_2.mux_l2_in_0__S mux_right_track_2.mux_l2_in_0_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_1__A1 mux_bottom_track_9.mux_l1_in_2_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.mux_l2_in_0__A1 mux_bottom_track_25.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_24.mux_l3_in_0__A0 mux_right_track_24.mux_l2_in_1_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_34.mux_l1_in_0__A0 chany_bottom_in[1] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l3_in_0__S mux_top_track_2.mux_l3_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
X_066_ right_bottom_grid_pin_41_ chanx_right_out[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_4_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_3_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_7_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_16.mux_l3_in_0__A0 mux_top_track_16.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_8.mux_l2_in_1__S mux_top_track_8.mux_l2_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_9.mux_l3_in_0__A1 mux_bottom_track_9.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_118_ chany_bottom_in[6] chany_top_out[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
X_049_ _049_/HI _049_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_right_track_26.mux_l1_in_0__A1 right_bottom_grid_pin_35_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_ mux_top_track_4.mux_l1_in_0_/S mux_top_track_4.mux_l2_in_1_/S
+ mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_1_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_26_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_33.mux_l1_in_1__A1 chanx_right_in[13] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_36.mux_l1_in_0__S mux_right_track_36.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1__A0 right_bottom_grid_pin_38_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_14.mux_l2_in_0_ right_bottom_grid_pin_37_ mux_right_track_14.mux_l1_in_0_/X
+ mux_right_track_14.mux_l2_in_1_/S mux_right_track_14.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.mux_l2_in_0_ mux_right_track_2.mux_l1_in_1_/X mux_right_track_2.mux_l1_in_0_/X
+ mux_right_track_2.mux_l2_in_0_/S mux_right_track_2.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_39_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_0_/S mux_top_track_4.mux_l3_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_24.mux_l2_in_1__A0 _049_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_6_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_right_track_36.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_34.mux_l2_in_0_/S
+ mux_right_track_36.mux_l1_in_0_/S mem_right_track_36.sky130_fd_sc_hd__dfxbp_1_0_/Q_N
+ clkbuf_3_2_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l2_in_1__A1 chany_bottom_in[19] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_33.mux_l2_in_0__A1 mux_bottom_track_33.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2__A0 chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0__A0 mux_right_track_0.mux_l1_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l2_in_1__A1 chany_bottom_in[17] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_082_ _082_/A chanx_right_out[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_10_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_5_0_prog_clk clkbuf_3_5_0_prog_clk/A clkbuf_3_5_0_prog_clk/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_33_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l1_in_1_ right_bottom_grid_pin_37_ right_bottom_grid_pin_35_
+ mux_right_track_2.mux_l1_in_1_/S mux_right_track_2.mux_l1_in_1_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_24.mux_l3_in_0__A0 mux_top_track_24.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l2_in_1_ _051_/HI mux_top_track_4.mux_l1_in_2_/X mux_top_track_4.mux_l2_in_1_/S
+ mux_top_track_4.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_32.sky130_fd_sc_hd__buf_4_0_ mux_top_track_32.mux_l3_in_0_/X _109_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_right_track_24.mux_l3_in_0__A1 mux_right_track_24.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_8.mux_l2_in_1__A0 _052_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_36.sky130_fd_sc_hd__buf_4_0__A mux_right_track_36.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_34.mux_l1_in_0__A1 right_bottom_grid_pin_39_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_065_ _065_/HI _065_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_8.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_track_16.mux_l3_in_0__A1 mux_top_track_16.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_2.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_5_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l1_in_2_ chany_bottom_in[14] chany_bottom_in[5] mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_2_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_117_ _117_/A chany_top_out[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_ mux_right_track_4.mux_l2_in_1_/S mux_right_track_4.mux_l3_in_0_/S
+ mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_/Q_N clkbuf_3_4_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_7_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_048_ _048_/HI _048_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_38_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_8.mux_l3_in_0__A0 mux_top_track_8.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_28.mux_l2_in_0__S mux_right_track_28.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_ mux_top_track_2.mux_l3_in_0_/S mux_top_track_4.mux_l1_in_0_/S
+ mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_1_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XANTENNA_mux_top_track_32.mux_l2_in_1__A0 _050_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_26.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1__A1 right_bottom_grid_pin_36_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0__S mux_top_track_0.mux_l1_in_2_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA__102__A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_24.mux_l2_in_1__A1 chany_bottom_in[18] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxbp_1_0__CLK clkbuf_3_4_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_32.mux_l3_in_0__A0 mux_top_track_32.mux_l2_in_1_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_8.mux_l1_in_2__A1 chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_17.mux_l3_in_0_ mux_bottom_track_17.mux_l2_in_1_/X mux_bottom_track_17.mux_l2_in_0_/X
+ mux_bottom_track_17.mux_l3_in_0_/S mux_bottom_track_17.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
Xmux_right_track_2.sky130_fd_sc_hd__buf_4_0_ mux_right_track_2.mux_l3_in_0_/X _084_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_27_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_right_track_0.mux_l2_in_0__A1 mux_right_track_0.mux_l1_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_right_track_14.mux_l1_in_0_ chany_top_in[19] chany_top_in[12] mux_right_track_14.mux_l1_in_0_/S
+ mux_right_track_14.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_081_ _081_/A chanx_right_out[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_5.mux_l3_in_0__S mux_bottom_track_5.mux_l3_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_2.mux_l1_in_0_ chany_top_in[4] chany_top_in[0] mux_right_track_2.mux_l1_in_1_/S
+ mux_right_track_2.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_2_0_prog_clk_A clkbuf_3_3_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A0 chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_24.mux_l3_in_0__A1 mux_top_track_24.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_1_/S mux_top_track_4.mux_l2_in_0_/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__mux2_1
Xmux_right_track_26.mux_l2_in_0_ _037_/HI mux_right_track_26.mux_l1_in_0_/X mux_right_track_26.mux_l2_in_0_/S
+ mux_right_track_26.mux_l2_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_7_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_track_8.mux_l2_in_1__A1 mux_top_track_8.mux_l1_in_2_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l3_in_0_/X _123_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK clkbuf_3_1_0_prog_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_064_ _064_/HI _064_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_2_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_17.mux_l2_in_1_ _054_/HI chanx_right_in[15] mux_bottom_track_17.mux_l2_in_1_/S
+ mux_bottom_track_17.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA__110__A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_28.mux_l2_in_0__A0 _038_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_0_/S mux_bottom_track_3.mux_l3_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l1_in_1_ chanx_right_in[17] chanx_right_in[10] mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xmem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_4.mux_l1_in_1_/S mux_right_track_4.mux_l2_in_1_/S
+ mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_/Q_N clkbuf_3_5_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
X_116_ chany_bottom_in[8] chany_top_out[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XANTENNA_mux_right_track_4.mux_l1_in_1__S mux_right_track_4.mux_l1_in_1_/S VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__105__A _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK clkbuf_3_1_0_prog_clk/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_047_ _047_/HI _047_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_8.mux_l3_in_0__A1 mux_top_track_8.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l2_in_1__S mux_top_track_4.mux_l2_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_mux_top_track_32.mux_l2_in_1__A1 chany_bottom_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_34_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_3.mux_l2_in_1_ _056_/HI chanx_right_in[18] mux_bottom_track_3.mux_l2_in_1_/S
+ mux_bottom_track_3.mux_l2_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__D mux_bottom_track_9.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_7_0_prog_clk_A clkbuf_3_7_0_prog_clk/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_20.sky130_fd_sc_hd__buf_4_0_ mux_right_track_20.mux_l2_in_0_/X _075_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_32.mux_l3_in_0__A1 mux_top_track_32.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__113__A _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_right_track_32.mux_l1_in_0__S mux_right_track_32.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxbp_1_0__D mux_right_track_18.mux_l2_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_track_14.sky130_fd_sc_hd__buf_4_0_ mux_right_track_14.mux_l3_in_0_/X _078_/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_4
XFILLER_27_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_080_ _080_/A chanx_right_out[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__108__A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A1 chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__D mux_bottom_track_17.mux_l3_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_36.mux_l2_in_0__A0 _042_/HI VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_4.mux_l1_in_0__A0 chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_063_ _063_/HI _063_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_1_/S mux_bottom_track_17.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1_ mux_right_track_22.mux_l1_in_0_/S
+ mux_right_track_22.mux_l2_in_0_/S mem_right_track_22.sky130_fd_sc_hd__dfxbp_1_1_/Q_N
+ clkbuf_3_6_0_prog_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_20_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_right_track_28.mux_l2_in_0__A1 mux_right_track_28.mux_l1_in_0_/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_right_track_2.mux_l1_in_2__A0 right_bottom_grid_pin_41_ VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l1_in_0_ chanx_right_in[3] top_left_grid_pin_1_ mux_top_track_4.mux_l1_in_0_/S
+ mux_top_track_4.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
XFILLER_34_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_ mux_right_track_2.mux_l3_in_0_/S mux_right_track_4.mux_l1_in_1_/S
+ mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_/Q_N clkbuf_3_7_0_prog_clk/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__dfxbp_1
XFILLER_11_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_track_26.mux_l1_in_0_ chany_bottom_in[15] right_bottom_grid_pin_35_ mux_right_track_26.mux_l1_in_0_/S
+ mux_right_track_26.mux_l1_in_0_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
X_115_ chany_bottom_in[9] chany_top_out[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__buf_2
XFILLER_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_046_ _046_/HI _046_/LO VGND VGND VPWR VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__121__A _121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_17.mux_l1_in_1_ chanx_right_in[8] chanx_right_in[1] mux_bottom_track_17.mux_l1_in_1_/S
+ mux_bottom_track_17.mux_l1_in_1_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__mux2_1
Xclkbuf_2_2_0_prog_clk clkbuf_0_prog_clk/X clkbuf_3_5_0_prog_clk/A VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__S mux_bottom_track_3.mux_l1_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__116__A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__D mux_top_track_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_1_/S mux_bottom_track_3.mux_l2_in_0_/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__mux2_1
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_2.mux_l2_in_1__A0 mux_right_track_2.mux_l1_in_3_/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_33.mux_l2_in_0__S ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A mux_bottom_track_25.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_right_track_24.mux_l2_in_0__S mux_right_track_24.mux_l2_in_0_/S VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

