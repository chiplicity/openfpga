version https://git-lfs.github.com/spec/v1
oid sha256:c084d554143877b453c074f833fe0e7b5540900d5d866b0b259c9bfbb9c3fe44
size 217124165
