magic
tech sky130A
magscale 1 2
timestamp 1605003539
<< locali >>
rect 17509 25143 17543 25313
rect 5273 23579 5307 23817
rect 21741 22423 21775 22525
rect 23673 16983 23707 17153
rect 2881 14807 2915 15113
rect 6469 13855 6503 13957
rect 11989 11679 12023 11849
rect 27077 9707 27111 27421
<< viali >>
rect 27077 27421 27111 27455
rect 4261 25449 4295 25483
rect 5365 25449 5399 25483
rect 10517 25449 10551 25483
rect 15945 25449 15979 25483
rect 17325 25449 17359 25483
rect 18153 25449 18187 25483
rect 18797 25449 18831 25483
rect 24777 25449 24811 25483
rect 8677 25381 8711 25415
rect 13645 25381 13679 25415
rect 14933 25381 14967 25415
rect 1409 25313 1443 25347
rect 2513 25313 2547 25347
rect 4077 25313 4111 25347
rect 5181 25313 5215 25347
rect 7481 25313 7515 25347
rect 7573 25313 7607 25347
rect 10333 25313 10367 25347
rect 11437 25313 11471 25347
rect 13001 25313 13035 25347
rect 14289 25313 14323 25347
rect 17141 25313 17175 25347
rect 17509 25313 17543 25347
rect 17785 25313 17819 25347
rect 18705 25313 18739 25347
rect 19993 25313 20027 25347
rect 21925 25313 21959 25347
rect 24593 25313 24627 25347
rect 7757 25245 7791 25279
rect 13093 25245 13127 25279
rect 13277 25245 13311 25279
rect 15301 25245 15335 25279
rect 16037 25245 16071 25279
rect 16221 25245 16255 25279
rect 1593 25177 1627 25211
rect 6745 25177 6779 25211
rect 14105 25177 14139 25211
rect 14473 25177 14507 25211
rect 18889 25245 18923 25279
rect 22201 25245 22235 25279
rect 20177 25177 20211 25211
rect 2697 25109 2731 25143
rect 4721 25109 4755 25143
rect 7113 25109 7147 25143
rect 8585 25109 8619 25143
rect 11621 25109 11655 25143
rect 12633 25109 12667 25143
rect 15577 25109 15611 25143
rect 16589 25109 16623 25143
rect 17049 25109 17083 25143
rect 17509 25109 17543 25143
rect 18337 25109 18371 25143
rect 19349 25109 19383 25143
rect 19901 25109 19935 25143
rect 21465 25109 21499 25143
rect 21741 25109 21775 25143
rect 3801 24905 3835 24939
rect 4905 24905 4939 24939
rect 10517 24905 10551 24939
rect 19809 24837 19843 24871
rect 20821 24837 20855 24871
rect 25145 24837 25179 24871
rect 4261 24769 4295 24803
rect 6653 24769 6687 24803
rect 7389 24769 7423 24803
rect 7573 24769 7607 24803
rect 8953 24769 8987 24803
rect 9137 24769 9171 24803
rect 11253 24769 11287 24803
rect 12265 24769 12299 24803
rect 14289 24769 14323 24803
rect 15761 24769 15795 24803
rect 17785 24769 17819 24803
rect 18797 24769 18831 24803
rect 20361 24769 20395 24803
rect 21925 24769 21959 24803
rect 24409 24769 24443 24803
rect 1409 24701 1443 24735
rect 2513 24701 2547 24735
rect 3433 24701 3467 24735
rect 3617 24701 3651 24735
rect 4721 24701 4755 24735
rect 5917 24701 5951 24735
rect 7297 24701 7331 24735
rect 11069 24701 11103 24735
rect 12541 24701 12575 24735
rect 13185 24701 13219 24735
rect 14013 24701 14047 24735
rect 18705 24701 18739 24735
rect 19349 24701 19383 24735
rect 24593 24701 24627 24735
rect 8401 24633 8435 24667
rect 8861 24633 8895 24667
rect 10057 24633 10091 24667
rect 13461 24633 13495 24667
rect 14105 24633 14139 24667
rect 15577 24633 15611 24667
rect 18613 24633 18647 24667
rect 19717 24633 19751 24667
rect 21189 24633 21223 24667
rect 21741 24633 21775 24667
rect 1593 24565 1627 24599
rect 2053 24565 2087 24599
rect 2421 24565 2455 24599
rect 2697 24565 2731 24599
rect 3157 24565 3191 24599
rect 4537 24565 4571 24599
rect 5273 24565 5307 24599
rect 6193 24565 6227 24599
rect 6929 24565 6963 24599
rect 7941 24565 7975 24599
rect 8493 24565 8527 24599
rect 9597 24565 9631 24599
rect 10977 24565 11011 24599
rect 11897 24565 11931 24599
rect 12725 24565 12759 24599
rect 13645 24565 13679 24599
rect 14749 24565 14783 24599
rect 15117 24565 15151 24599
rect 15209 24565 15243 24599
rect 15669 24565 15703 24599
rect 16221 24565 16255 24599
rect 16589 24565 16623 24599
rect 17049 24565 17083 24599
rect 17509 24565 17543 24599
rect 18245 24565 18279 24599
rect 20177 24565 20211 24599
rect 20269 24565 20303 24599
rect 21373 24565 21407 24599
rect 21833 24565 21867 24599
rect 22477 24565 22511 24599
rect 24777 24565 24811 24599
rect 2053 24361 2087 24395
rect 4261 24361 4295 24395
rect 8677 24361 8711 24395
rect 10149 24361 10183 24395
rect 12909 24361 12943 24395
rect 13277 24361 13311 24395
rect 14657 24361 14691 24395
rect 15485 24361 15519 24395
rect 16221 24361 16255 24395
rect 19441 24361 19475 24395
rect 20913 24361 20947 24395
rect 24777 24361 24811 24395
rect 10057 24293 10091 24327
rect 11713 24293 11747 24327
rect 12173 24293 12207 24327
rect 15853 24293 15887 24327
rect 18429 24293 18463 24327
rect 22937 24293 22971 24327
rect 1409 24225 1443 24259
rect 2513 24225 2547 24259
rect 4077 24225 4111 24259
rect 6081 24225 6115 24259
rect 8493 24225 8527 24259
rect 12265 24225 12299 24259
rect 13737 24225 13771 24259
rect 13829 24225 13863 24259
rect 15301 24225 15335 24259
rect 16497 24225 16531 24259
rect 16764 24225 16798 24259
rect 19349 24225 19383 24259
rect 19993 24225 20027 24259
rect 21281 24225 21315 24259
rect 22385 24225 22419 24259
rect 22845 24225 22879 24259
rect 24593 24225 24627 24259
rect 5825 24157 5859 24191
rect 10241 24157 10275 24191
rect 11069 24157 11103 24191
rect 12357 24157 12391 24191
rect 13921 24157 13955 24191
rect 19533 24157 19567 24191
rect 21373 24157 21407 24191
rect 21465 24157 21499 24191
rect 23029 24157 23063 24191
rect 18981 24089 19015 24123
rect 1593 24021 1627 24055
rect 2697 24021 2731 24055
rect 4721 24021 4755 24055
rect 7205 24021 7239 24055
rect 7849 24021 7883 24055
rect 9689 24021 9723 24055
rect 10793 24021 10827 24055
rect 11805 24021 11839 24055
rect 13369 24021 13403 24055
rect 15025 24021 15059 24055
rect 17877 24021 17911 24055
rect 18797 24021 18831 24055
rect 20545 24021 20579 24055
rect 22017 24021 22051 24055
rect 22477 24021 22511 24055
rect 23765 24021 23799 24055
rect 2605 23817 2639 23851
rect 5273 23817 5307 23851
rect 8401 23817 8435 23851
rect 9689 23817 9723 23851
rect 10057 23817 10091 23851
rect 11897 23817 11931 23851
rect 12265 23817 12299 23851
rect 14749 23817 14783 23851
rect 15393 23817 15427 23851
rect 16497 23817 16531 23851
rect 16773 23817 16807 23851
rect 19441 23817 19475 23851
rect 19993 23817 20027 23851
rect 20453 23817 20487 23851
rect 23489 23817 23523 23851
rect 4169 23749 4203 23783
rect 1869 23681 1903 23715
rect 3801 23681 3835 23715
rect 4997 23681 5031 23715
rect 1593 23613 1627 23647
rect 2881 23613 2915 23647
rect 4905 23613 4939 23647
rect 10425 23749 10459 23783
rect 14473 23749 14507 23783
rect 17417 23749 17451 23783
rect 20545 23749 20579 23783
rect 6285 23681 6319 23715
rect 7297 23681 7331 23715
rect 7481 23681 7515 23715
rect 7941 23681 7975 23715
rect 8861 23681 8895 23715
rect 8953 23681 8987 23715
rect 11069 23681 11103 23715
rect 16037 23681 16071 23715
rect 21097 23681 21131 23715
rect 24225 23681 24259 23715
rect 5549 23613 5583 23647
rect 8769 23613 8803 23647
rect 10885 23613 10919 23647
rect 12449 23613 12483 23647
rect 15853 23613 15887 23647
rect 18061 23613 18095 23647
rect 22293 23613 22327 23647
rect 24133 23613 24167 23647
rect 25237 23613 25271 23647
rect 25789 23613 25823 23647
rect 5273 23545 5307 23579
rect 6653 23545 6687 23579
rect 12716 23545 12750 23579
rect 15761 23545 15795 23579
rect 17877 23545 17911 23579
rect 18328 23545 18362 23579
rect 21005 23545 21039 23579
rect 22569 23545 22603 23579
rect 24685 23545 24719 23579
rect 3065 23477 3099 23511
rect 4445 23477 4479 23511
rect 4813 23477 4847 23511
rect 5825 23477 5859 23511
rect 6837 23477 6871 23511
rect 7205 23477 7239 23511
rect 8309 23477 8343 23511
rect 10793 23477 10827 23511
rect 11437 23477 11471 23511
rect 13829 23477 13863 23511
rect 15209 23477 15243 23511
rect 16957 23477 16991 23511
rect 20913 23477 20947 23511
rect 21557 23477 21591 23511
rect 22201 23477 22235 23511
rect 23029 23477 23063 23511
rect 23673 23477 23707 23511
rect 24041 23477 24075 23511
rect 25421 23477 25455 23511
rect 2881 23273 2915 23307
rect 6469 23273 6503 23307
rect 8033 23273 8067 23307
rect 8585 23273 8619 23307
rect 12357 23273 12391 23307
rect 13461 23273 13495 23307
rect 13921 23273 13955 23307
rect 16681 23273 16715 23307
rect 17233 23273 17267 23307
rect 19073 23273 19107 23307
rect 20637 23273 20671 23307
rect 23213 23273 23247 23307
rect 23857 23273 23891 23307
rect 24225 23273 24259 23307
rect 2053 23205 2087 23239
rect 17877 23205 17911 23239
rect 22100 23205 22134 23239
rect 24685 23205 24719 23239
rect 1777 23137 1811 23171
rect 4997 23137 5031 23171
rect 5089 23137 5123 23171
rect 5356 23137 5390 23171
rect 7941 23137 7975 23171
rect 9689 23137 9723 23171
rect 11244 23137 11278 23171
rect 13829 23137 13863 23171
rect 15301 23137 15335 23171
rect 15568 23137 15602 23171
rect 17969 23137 18003 23171
rect 19625 23137 19659 23171
rect 24777 23137 24811 23171
rect 4077 23069 4111 23103
rect 8125 23069 8159 23103
rect 9045 23069 9079 23103
rect 9965 23069 9999 23103
rect 10977 23069 11011 23103
rect 14013 23069 14047 23103
rect 18245 23069 18279 23103
rect 19717 23069 19751 23103
rect 19901 23069 19935 23103
rect 21465 23069 21499 23103
rect 21833 23069 21867 23103
rect 24869 23069 24903 23103
rect 7113 23001 7147 23035
rect 7389 23001 7423 23035
rect 14473 23001 14507 23035
rect 19257 23001 19291 23035
rect 25329 23001 25363 23035
rect 1685 22933 1719 22967
rect 3709 22933 3743 22967
rect 4629 22933 4663 22967
rect 7573 22933 7607 22967
rect 9413 22933 9447 22967
rect 10425 22933 10459 22967
rect 10793 22933 10827 22967
rect 12909 22933 12943 22967
rect 13277 22933 13311 22967
rect 15025 22933 15059 22967
rect 21097 22933 21131 22967
rect 24317 22933 24351 22967
rect 4721 22729 4755 22763
rect 9689 22729 9723 22763
rect 14381 22729 14415 22763
rect 14749 22729 14783 22763
rect 16405 22729 16439 22763
rect 17509 22729 17543 22763
rect 19165 22729 19199 22763
rect 20729 22729 20763 22763
rect 22017 22729 22051 22763
rect 23029 22729 23063 22763
rect 25605 22729 25639 22763
rect 25973 22729 26007 22763
rect 2513 22661 2547 22695
rect 5181 22661 5215 22695
rect 9597 22661 9631 22695
rect 11437 22661 11471 22695
rect 1685 22593 1719 22627
rect 4169 22593 4203 22627
rect 5089 22593 5123 22627
rect 5825 22593 5859 22627
rect 10333 22593 10367 22627
rect 12265 22593 12299 22627
rect 15393 22593 15427 22627
rect 15485 22593 15519 22627
rect 16865 22593 16899 22627
rect 22661 22593 22695 22627
rect 1409 22525 1443 22559
rect 2145 22525 2179 22559
rect 3525 22525 3559 22559
rect 3985 22525 4019 22559
rect 6929 22525 6963 22559
rect 10149 22525 10183 22559
rect 11253 22525 11287 22559
rect 12449 22525 12483 22559
rect 12716 22525 12750 22559
rect 16681 22525 16715 22559
rect 17877 22525 17911 22559
rect 18061 22525 18095 22559
rect 19349 22525 19383 22559
rect 21741 22525 21775 22559
rect 21833 22525 21867 22559
rect 23673 22525 23707 22559
rect 23940 22525 23974 22559
rect 5549 22457 5583 22491
rect 6653 22457 6687 22491
rect 7174 22457 7208 22491
rect 18337 22457 18371 22491
rect 19594 22457 19628 22491
rect 22477 22457 22511 22491
rect 3157 22389 3191 22423
rect 3617 22389 3651 22423
rect 4077 22389 4111 22423
rect 5641 22389 5675 22423
rect 6193 22389 6227 22423
rect 8309 22389 8343 22423
rect 9137 22389 9171 22423
rect 10057 22389 10091 22423
rect 10793 22389 10827 22423
rect 11161 22389 11195 22423
rect 11897 22389 11931 22423
rect 13829 22389 13863 22423
rect 14933 22389 14967 22423
rect 15301 22389 15335 22423
rect 16037 22389 16071 22423
rect 18797 22389 18831 22423
rect 21465 22389 21499 22423
rect 21741 22389 21775 22423
rect 22385 22389 22419 22423
rect 23489 22389 23523 22423
rect 25053 22389 25087 22423
rect 26341 22389 26375 22423
rect 2789 22185 2823 22219
rect 3709 22185 3743 22219
rect 5457 22185 5491 22219
rect 6009 22185 6043 22219
rect 6561 22185 6595 22219
rect 6929 22185 6963 22219
rect 7021 22185 7055 22219
rect 7941 22185 7975 22219
rect 10057 22185 10091 22219
rect 12357 22185 12391 22219
rect 13553 22185 13587 22219
rect 17141 22185 17175 22219
rect 19441 22185 19475 22219
rect 19809 22185 19843 22219
rect 20545 22185 20579 22219
rect 22293 22185 22327 22219
rect 22937 22185 22971 22219
rect 1409 22117 1443 22151
rect 2881 22117 2915 22151
rect 7665 22117 7699 22151
rect 12725 22117 12759 22151
rect 18613 22117 18647 22151
rect 21158 22117 21192 22151
rect 24010 22117 24044 22151
rect 1961 22049 1995 22083
rect 4077 22049 4111 22083
rect 4344 22049 4378 22083
rect 8125 22049 8159 22083
rect 9505 22049 9539 22083
rect 11253 22049 11287 22083
rect 12265 22049 12299 22083
rect 13921 22049 13955 22083
rect 14197 22049 14231 22083
rect 15025 22049 15059 22083
rect 16028 22049 16062 22083
rect 18705 22049 18739 22083
rect 3065 21981 3099 22015
rect 7113 21981 7147 22015
rect 10149 21981 10183 22015
rect 10241 21981 10275 22015
rect 12817 21981 12851 22015
rect 13001 21981 13035 22015
rect 15761 21981 15795 22015
rect 18797 21981 18831 22015
rect 20913 21981 20947 22015
rect 23305 21981 23339 22015
rect 23673 21981 23707 22015
rect 23765 21981 23799 22015
rect 2329 21913 2363 21947
rect 8309 21913 8343 21947
rect 9689 21913 9723 21947
rect 11069 21913 11103 21947
rect 11437 21913 11471 21947
rect 18245 21913 18279 21947
rect 2421 21845 2455 21879
rect 6469 21845 6503 21879
rect 8769 21845 8803 21879
rect 9137 21845 9171 21879
rect 10793 21845 10827 21879
rect 11897 21845 11931 21879
rect 15485 21845 15519 21879
rect 17693 21845 17727 21879
rect 18153 21845 18187 21879
rect 25145 21845 25179 21879
rect 1869 21641 1903 21675
rect 2237 21641 2271 21675
rect 5089 21641 5123 21675
rect 6285 21641 6319 21675
rect 7113 21641 7147 21675
rect 9689 21641 9723 21675
rect 10517 21641 10551 21675
rect 11805 21641 11839 21675
rect 12449 21641 12483 21675
rect 13461 21641 13495 21675
rect 17049 21641 17083 21675
rect 17785 21641 17819 21675
rect 20453 21641 20487 21675
rect 22017 21641 22051 21675
rect 24777 21641 24811 21675
rect 25145 21641 25179 21675
rect 6561 21573 6595 21607
rect 13829 21573 13863 21607
rect 17509 21573 17543 21607
rect 2329 21505 2363 21539
rect 5641 21505 5675 21539
rect 7573 21505 7607 21539
rect 10977 21505 11011 21539
rect 11161 21505 11195 21539
rect 13001 21505 13035 21539
rect 14381 21505 14415 21539
rect 18613 21505 18647 21539
rect 19533 21505 19567 21539
rect 21005 21505 21039 21539
rect 21465 21505 21499 21539
rect 21925 21505 21959 21539
rect 22661 21505 22695 21539
rect 24317 21505 24351 21539
rect 25421 21505 25455 21539
rect 2596 21437 2630 21471
rect 7840 21437 7874 21471
rect 12265 21437 12299 21471
rect 12909 21437 12943 21471
rect 16865 21437 16899 21471
rect 18521 21437 18555 21471
rect 19809 21437 19843 21471
rect 22477 21437 22511 21471
rect 24041 21437 24075 21471
rect 25237 21437 25271 21471
rect 25973 21437 26007 21471
rect 4997 21369 5031 21403
rect 5549 21369 5583 21403
rect 7481 21369 7515 21403
rect 14289 21369 14323 21403
rect 14648 21369 14682 21403
rect 18429 21369 18463 21403
rect 20821 21369 20855 21403
rect 23121 21369 23155 21403
rect 24133 21369 24167 21403
rect 3709 21301 3743 21335
rect 4261 21301 4295 21335
rect 5457 21301 5491 21335
rect 8953 21301 8987 21335
rect 10057 21301 10091 21335
rect 10885 21301 10919 21335
rect 12817 21301 12851 21335
rect 15761 21301 15795 21335
rect 16405 21301 16439 21335
rect 16773 21301 16807 21335
rect 18061 21301 18095 21335
rect 19073 21301 19107 21335
rect 20361 21301 20395 21335
rect 20913 21301 20947 21335
rect 22385 21301 22419 21335
rect 23489 21301 23523 21335
rect 23673 21301 23707 21335
rect 26341 21301 26375 21335
rect 2053 21097 2087 21131
rect 2513 21097 2547 21131
rect 4077 21097 4111 21131
rect 4537 21097 4571 21131
rect 5181 21097 5215 21131
rect 5457 21097 5491 21131
rect 6469 21097 6503 21131
rect 7665 21097 7699 21131
rect 8493 21097 8527 21131
rect 9045 21097 9079 21131
rect 9413 21097 9447 21131
rect 14565 21097 14599 21131
rect 14841 21097 14875 21131
rect 16681 21097 16715 21131
rect 19165 21097 19199 21131
rect 20453 21097 20487 21131
rect 22201 21097 22235 21131
rect 22661 21097 22695 21131
rect 23673 21097 23707 21131
rect 3157 21029 3191 21063
rect 4445 21029 4479 21063
rect 8401 21029 8435 21063
rect 13093 21029 13127 21063
rect 15568 21029 15602 21063
rect 19717 21029 19751 21063
rect 24032 21029 24066 21063
rect 2421 20961 2455 20995
rect 10497 20961 10531 20995
rect 17233 20961 17267 20995
rect 17601 20961 17635 20995
rect 17785 20961 17819 20995
rect 18052 20961 18086 20995
rect 20913 20961 20947 20995
rect 22569 20961 22603 20995
rect 23765 20961 23799 20995
rect 2605 20893 2639 20927
rect 4629 20893 4663 20927
rect 6561 20893 6595 20927
rect 6653 20893 6687 20927
rect 7297 20893 7331 20927
rect 8585 20893 8619 20927
rect 10241 20893 10275 20927
rect 12449 20893 12483 20927
rect 13185 20893 13219 20927
rect 13369 20893 13403 20927
rect 15301 20893 15335 20927
rect 21097 20893 21131 20927
rect 22109 20893 22143 20927
rect 22845 20893 22879 20927
rect 1869 20757 1903 20791
rect 3525 20757 3559 20791
rect 3893 20757 3927 20791
rect 5825 20757 5859 20791
rect 6101 20757 6135 20791
rect 8033 20757 8067 20791
rect 9965 20757 9999 20791
rect 11621 20757 11655 20791
rect 12725 20757 12759 20791
rect 13829 20757 13863 20791
rect 14197 20757 14231 20791
rect 20085 20757 20119 20791
rect 21741 20757 21775 20791
rect 23305 20757 23339 20791
rect 25145 20757 25179 20791
rect 2145 20553 2179 20587
rect 3617 20553 3651 20587
rect 4169 20553 4203 20587
rect 5825 20553 5859 20587
rect 6193 20553 6227 20587
rect 7757 20553 7791 20587
rect 10609 20553 10643 20587
rect 12265 20553 12299 20587
rect 15117 20553 15151 20587
rect 15761 20553 15795 20587
rect 16037 20553 16071 20587
rect 17877 20553 17911 20587
rect 20545 20553 20579 20587
rect 21189 20553 21223 20587
rect 22753 20553 22787 20587
rect 23673 20553 23707 20587
rect 24685 20553 24719 20587
rect 25421 20553 25455 20587
rect 26249 20553 26283 20587
rect 6285 20485 6319 20519
rect 10149 20485 10183 20519
rect 18245 20485 18279 20519
rect 25145 20485 25179 20519
rect 5273 20417 5307 20451
rect 7849 20417 7883 20451
rect 11069 20417 11103 20451
rect 11253 20417 11287 20451
rect 11621 20417 11655 20451
rect 12725 20417 12759 20451
rect 16773 20417 16807 20451
rect 22201 20417 22235 20451
rect 24317 20417 24351 20451
rect 2237 20349 2271 20383
rect 2504 20349 2538 20383
rect 5089 20349 5123 20383
rect 6469 20349 6503 20383
rect 6837 20349 6871 20383
rect 12449 20349 12483 20383
rect 13277 20349 13311 20383
rect 13737 20349 13771 20383
rect 16681 20349 16715 20383
rect 18061 20349 18095 20383
rect 19165 20349 19199 20383
rect 21557 20349 21591 20383
rect 23489 20349 23523 20383
rect 24133 20349 24167 20383
rect 25237 20349 25271 20383
rect 25789 20349 25823 20383
rect 1777 20281 1811 20315
rect 7389 20281 7423 20315
rect 8094 20281 8128 20315
rect 14004 20281 14038 20315
rect 16589 20281 16623 20315
rect 17233 20281 17267 20315
rect 19073 20281 19107 20315
rect 19432 20281 19466 20315
rect 22017 20281 22051 20315
rect 22109 20281 22143 20315
rect 24041 20281 24075 20315
rect 4537 20213 4571 20247
rect 4721 20213 4755 20247
rect 5181 20213 5215 20247
rect 9229 20213 9263 20247
rect 10425 20213 10459 20247
rect 10977 20213 11011 20247
rect 13553 20213 13587 20247
rect 16221 20213 16255 20247
rect 18613 20213 18647 20247
rect 21649 20213 21683 20247
rect 23029 20213 23063 20247
rect 2237 20009 2271 20043
rect 2973 20009 3007 20043
rect 4353 20009 4387 20043
rect 8125 20009 8159 20043
rect 10149 20009 10183 20043
rect 12725 20009 12759 20043
rect 13737 20009 13771 20043
rect 14473 20009 14507 20043
rect 15301 20009 15335 20043
rect 15761 20009 15795 20043
rect 16681 20009 16715 20043
rect 17601 20009 17635 20043
rect 19717 20009 19751 20043
rect 20269 20009 20303 20043
rect 20913 20009 20947 20043
rect 24317 20009 24351 20043
rect 4874 19941 4908 19975
rect 7481 19941 7515 19975
rect 12449 19941 12483 19975
rect 13185 19941 13219 19975
rect 16313 19941 16347 19975
rect 20729 19941 20763 19975
rect 22170 19941 22204 19975
rect 2329 19873 2363 19907
rect 3341 19873 3375 19907
rect 4629 19873 4663 19907
rect 9505 19873 9539 19907
rect 10497 19873 10531 19907
rect 13093 19873 13127 19907
rect 15117 19873 15151 19907
rect 15669 19873 15703 19907
rect 16865 19873 16899 19907
rect 18604 19873 18638 19907
rect 24777 19873 24811 19907
rect 2421 19805 2455 19839
rect 3893 19805 3927 19839
rect 7573 19805 7607 19839
rect 7665 19805 7699 19839
rect 8677 19805 8711 19839
rect 10241 19805 10275 19839
rect 13369 19805 13403 19839
rect 15945 19805 15979 19839
rect 17141 19805 17175 19839
rect 18337 19805 18371 19839
rect 21925 19805 21959 19839
rect 24869 19805 24903 19839
rect 24961 19805 24995 19839
rect 7021 19737 7055 19771
rect 23305 19737 23339 19771
rect 24409 19737 24443 19771
rect 1777 19669 1811 19703
rect 1869 19669 1903 19703
rect 6009 19669 6043 19703
rect 6561 19669 6595 19703
rect 7113 19669 7147 19703
rect 9045 19669 9079 19703
rect 9321 19669 9355 19703
rect 11621 19669 11655 19703
rect 14105 19669 14139 19703
rect 14933 19669 14967 19703
rect 18153 19669 18187 19703
rect 21649 19669 21683 19703
rect 23949 19669 23983 19703
rect 25421 19669 25455 19703
rect 1869 19465 1903 19499
rect 4169 19465 4203 19499
rect 5641 19465 5675 19499
rect 9689 19465 9723 19499
rect 11897 19465 11931 19499
rect 15577 19465 15611 19499
rect 17417 19465 17451 19499
rect 3341 19397 3375 19431
rect 19165 19397 19199 19431
rect 2513 19329 2547 19363
rect 7389 19329 7423 19363
rect 9137 19329 9171 19363
rect 10057 19329 10091 19363
rect 10701 19329 10735 19363
rect 13461 19329 13495 19363
rect 15025 19329 15059 19363
rect 16497 19329 16531 19363
rect 16589 19329 16623 19363
rect 18705 19329 18739 19363
rect 24225 19329 24259 19363
rect 2329 19261 2363 19295
rect 2881 19261 2915 19295
rect 4261 19261 4295 19295
rect 6193 19261 6227 19295
rect 7205 19261 7239 19295
rect 12173 19261 12207 19295
rect 14289 19261 14323 19295
rect 14933 19261 14967 19295
rect 17141 19261 17175 19295
rect 19625 19261 19659 19295
rect 20361 19261 20395 19295
rect 21097 19261 21131 19295
rect 23489 19261 23523 19295
rect 25237 19261 25271 19295
rect 2237 19193 2271 19227
rect 3617 19193 3651 19227
rect 4528 19193 4562 19227
rect 7297 19193 7331 19227
rect 8493 19193 8527 19227
rect 10517 19193 10551 19227
rect 11253 19193 11287 19227
rect 12725 19193 12759 19227
rect 13277 19193 13311 19227
rect 17785 19193 17819 19227
rect 18521 19193 18555 19227
rect 19901 19193 19935 19227
rect 21005 19193 21039 19227
rect 21342 19193 21376 19227
rect 23121 19193 23155 19227
rect 24133 19193 24167 19227
rect 25789 19193 25823 19227
rect 1777 19125 1811 19159
rect 6561 19125 6595 19159
rect 6837 19125 6871 19159
rect 7849 19125 7883 19159
rect 8585 19125 8619 19159
rect 8953 19125 8987 19159
rect 9045 19125 9079 19159
rect 10149 19125 10183 19159
rect 10609 19125 10643 19159
rect 12909 19125 12943 19159
rect 13369 19125 13403 19159
rect 13921 19125 13955 19159
rect 14473 19125 14507 19159
rect 14841 19125 14875 19159
rect 15853 19125 15887 19159
rect 16037 19125 16071 19159
rect 16405 19125 16439 19159
rect 18061 19125 18095 19159
rect 18429 19125 18463 19159
rect 19533 19125 19567 19159
rect 22477 19125 22511 19159
rect 23673 19125 23707 19159
rect 24041 19125 24075 19159
rect 24685 19125 24719 19159
rect 25145 19125 25179 19159
rect 25421 19125 25455 19159
rect 26157 19125 26191 19159
rect 2053 18921 2087 18955
rect 2513 18921 2547 18955
rect 4353 18921 4387 18955
rect 6101 18921 6135 18955
rect 7481 18921 7515 18955
rect 8493 18921 8527 18955
rect 13277 18921 13311 18955
rect 15301 18921 15335 18955
rect 16313 18921 16347 18955
rect 16957 18921 16991 18955
rect 18153 18921 18187 18955
rect 18981 18921 19015 18955
rect 20085 18921 20119 18955
rect 21281 18921 21315 18955
rect 22017 18921 22051 18955
rect 22753 18921 22787 18955
rect 25053 18921 25087 18955
rect 1961 18853 1995 18887
rect 3525 18853 3559 18887
rect 3893 18853 3927 18887
rect 6653 18853 6687 18887
rect 7205 18853 7239 18887
rect 8401 18853 8435 18887
rect 10578 18853 10612 18887
rect 13185 18853 13219 18887
rect 15761 18853 15795 18887
rect 16773 18853 16807 18887
rect 23489 18853 23523 18887
rect 2421 18785 2455 18819
rect 4721 18785 4755 18819
rect 4988 18785 5022 18819
rect 7849 18785 7883 18819
rect 10333 18785 10367 18819
rect 15669 18785 15703 18819
rect 17325 18785 17359 18819
rect 17417 18785 17451 18819
rect 18889 18785 18923 18819
rect 19901 18785 19935 18819
rect 20269 18785 20303 18819
rect 21373 18785 21407 18819
rect 22569 18785 22603 18819
rect 23673 18785 23707 18819
rect 23940 18785 23974 18819
rect 2605 18717 2639 18751
rect 8677 18717 8711 18751
rect 13369 18717 13403 18751
rect 14197 18717 14231 18751
rect 15945 18717 15979 18751
rect 17509 18717 17543 18751
rect 19073 18717 19107 18751
rect 21465 18717 21499 18751
rect 12817 18649 12851 18683
rect 15025 18649 15059 18683
rect 3065 18581 3099 18615
rect 8033 18581 8067 18615
rect 9321 18581 9355 18615
rect 10241 18581 10275 18615
rect 11713 18581 11747 18615
rect 12541 18581 12575 18615
rect 14565 18581 14599 18615
rect 18521 18581 18555 18615
rect 19533 18581 19567 18615
rect 20729 18581 20763 18615
rect 20913 18581 20947 18615
rect 22293 18581 22327 18615
rect 23121 18581 23155 18615
rect 25605 18581 25639 18615
rect 2053 18377 2087 18411
rect 4721 18377 4755 18411
rect 6561 18377 6595 18411
rect 7757 18377 7791 18411
rect 9689 18377 9723 18411
rect 10241 18377 10275 18411
rect 12265 18377 12299 18411
rect 13829 18377 13863 18411
rect 16313 18377 16347 18411
rect 17049 18377 17083 18411
rect 19073 18377 19107 18411
rect 19717 18377 19751 18411
rect 21005 18377 21039 18411
rect 21281 18377 21315 18411
rect 22569 18377 22603 18411
rect 23121 18377 23155 18411
rect 25053 18377 25087 18411
rect 8125 18309 8159 18343
rect 21465 18309 21499 18343
rect 2145 18241 2179 18275
rect 4261 18241 4295 18275
rect 5365 18241 5399 18275
rect 11345 18241 11379 18275
rect 18521 18241 18555 18275
rect 18613 18241 18647 18275
rect 20361 18241 20395 18275
rect 20545 18241 20579 18275
rect 21925 18241 21959 18275
rect 22109 18241 22143 18275
rect 23673 18241 23707 18275
rect 4629 18173 4663 18207
rect 6837 18173 6871 18207
rect 8309 18173 8343 18207
rect 10701 18173 10735 18207
rect 11161 18173 11195 18207
rect 12449 18173 12483 18207
rect 14933 18173 14967 18207
rect 17785 18173 17819 18207
rect 18429 18173 18463 18207
rect 20269 18173 20303 18207
rect 2390 18105 2424 18139
rect 5089 18105 5123 18139
rect 6101 18105 6135 18139
rect 7113 18105 7147 18139
rect 8576 18105 8610 18139
rect 11253 18105 11287 18139
rect 11805 18105 11839 18139
rect 12716 18105 12750 18139
rect 14381 18105 14415 18139
rect 14841 18105 14875 18139
rect 15200 18105 15234 18139
rect 21833 18105 21867 18139
rect 23489 18105 23523 18139
rect 23940 18105 23974 18139
rect 1685 18037 1719 18071
rect 3525 18037 3559 18071
rect 5181 18037 5215 18071
rect 5733 18037 5767 18071
rect 10793 18037 10827 18071
rect 17509 18037 17543 18071
rect 18061 18037 18095 18071
rect 19901 18037 19935 18071
rect 2145 17833 2179 17867
rect 2789 17833 2823 17867
rect 6101 17833 6135 17867
rect 6377 17833 6411 17867
rect 6745 17833 6779 17867
rect 7573 17833 7607 17867
rect 8493 17833 8527 17867
rect 10517 17833 10551 17867
rect 12909 17833 12943 17867
rect 14473 17833 14507 17867
rect 15025 17833 15059 17867
rect 15301 17833 15335 17867
rect 16589 17833 16623 17867
rect 16957 17833 16991 17867
rect 19349 17833 19383 17867
rect 22845 17833 22879 17867
rect 24869 17833 24903 17867
rect 11244 17765 11278 17799
rect 13921 17765 13955 17799
rect 17316 17765 17350 17799
rect 18981 17765 19015 17799
rect 19809 17765 19843 17799
rect 25237 17765 25271 17799
rect 1685 17697 1719 17731
rect 2237 17697 2271 17731
rect 3525 17697 3559 17731
rect 4077 17697 4111 17731
rect 4333 17697 4367 17731
rect 6561 17697 6595 17731
rect 7205 17697 7239 17731
rect 8401 17697 8435 17731
rect 9689 17697 9723 17731
rect 10885 17697 10919 17731
rect 13829 17697 13863 17731
rect 15669 17697 15703 17731
rect 15761 17697 15795 17731
rect 19533 17697 19567 17731
rect 21169 17697 21203 17731
rect 23765 17697 23799 17731
rect 24961 17697 24995 17731
rect 2329 17629 2363 17663
rect 8677 17629 8711 17663
rect 9965 17629 9999 17663
rect 10977 17629 11011 17663
rect 14105 17629 14139 17663
rect 15945 17629 15979 17663
rect 17049 17629 17083 17663
rect 20913 17629 20947 17663
rect 23857 17629 23891 17663
rect 23949 17629 23983 17663
rect 8033 17561 8067 17595
rect 9413 17561 9447 17595
rect 12357 17561 12391 17595
rect 13461 17561 13495 17595
rect 23397 17561 23431 17595
rect 1777 17493 1811 17527
rect 3157 17493 3191 17527
rect 5457 17493 5491 17527
rect 7941 17493 7975 17527
rect 9137 17493 9171 17527
rect 13277 17493 13311 17527
rect 18429 17493 18463 17527
rect 20361 17493 20395 17527
rect 20729 17493 20763 17527
rect 22293 17493 22327 17527
rect 23305 17493 23339 17527
rect 24501 17493 24535 17527
rect 1869 17289 1903 17323
rect 4169 17289 4203 17323
rect 5089 17289 5123 17323
rect 7757 17289 7791 17323
rect 8125 17289 8159 17323
rect 10701 17289 10735 17323
rect 13921 17289 13955 17323
rect 15393 17289 15427 17323
rect 16313 17289 16347 17323
rect 19441 17289 19475 17323
rect 20085 17289 20119 17323
rect 22753 17289 22787 17323
rect 23489 17289 23523 17323
rect 25145 17289 25179 17323
rect 25697 17289 25731 17323
rect 26157 17289 26191 17323
rect 9597 17221 9631 17255
rect 15945 17221 15979 17255
rect 5641 17153 5675 17187
rect 6101 17153 6135 17187
rect 10241 17153 10275 17187
rect 11345 17153 11379 17187
rect 12265 17153 12299 17187
rect 13093 17153 13127 17187
rect 20637 17153 20671 17187
rect 23673 17153 23707 17187
rect 23765 17153 23799 17187
rect 1961 17085 1995 17119
rect 4997 17085 5031 17119
rect 5549 17085 5583 17119
rect 6837 17085 6871 17119
rect 8217 17085 8251 17119
rect 8484 17085 8518 17119
rect 10609 17085 10643 17119
rect 11161 17085 11195 17119
rect 11897 17085 11931 17119
rect 12817 17085 12851 17119
rect 14013 17085 14047 17119
rect 14280 17085 14314 17119
rect 16497 17085 16531 17119
rect 18061 17085 18095 17119
rect 20904 17085 20938 17119
rect 2228 17017 2262 17051
rect 7113 17017 7147 17051
rect 16773 17017 16807 17051
rect 18306 17017 18340 17051
rect 23121 17017 23155 17051
rect 24010 17017 24044 17051
rect 3341 16949 3375 16983
rect 4629 16949 4663 16983
rect 5457 16949 5491 16983
rect 6653 16949 6687 16983
rect 11069 16949 11103 16983
rect 12449 16949 12483 16983
rect 12909 16949 12943 16983
rect 13553 16949 13587 16983
rect 17325 16949 17359 16983
rect 17785 16949 17819 16983
rect 20545 16949 20579 16983
rect 22017 16949 22051 16983
rect 23673 16949 23707 16983
rect 1685 16745 1719 16779
rect 3525 16745 3559 16779
rect 4077 16745 4111 16779
rect 7021 16745 7055 16779
rect 7573 16745 7607 16779
rect 8677 16745 8711 16779
rect 9873 16745 9907 16779
rect 10425 16745 10459 16779
rect 13645 16745 13679 16779
rect 14013 16745 14047 16779
rect 14105 16745 14139 16779
rect 15301 16745 15335 16779
rect 16497 16745 16531 16779
rect 17325 16745 17359 16779
rect 17877 16745 17911 16779
rect 18981 16745 19015 16779
rect 20729 16745 20763 16779
rect 24041 16745 24075 16779
rect 24225 16745 24259 16779
rect 3801 16677 3835 16711
rect 9505 16677 9539 16711
rect 10701 16677 10735 16711
rect 15025 16677 15059 16711
rect 19349 16677 19383 16711
rect 21465 16677 21499 16711
rect 22008 16677 22042 16711
rect 24593 16677 24627 16711
rect 2053 16609 2087 16643
rect 2145 16609 2179 16643
rect 3157 16609 3191 16643
rect 5356 16609 5390 16643
rect 7941 16609 7975 16643
rect 9689 16609 9723 16643
rect 11161 16609 11195 16643
rect 11428 16609 11462 16643
rect 14749 16609 14783 16643
rect 15669 16609 15703 16643
rect 17785 16609 17819 16643
rect 18521 16609 18555 16643
rect 2237 16541 2271 16575
rect 2789 16541 2823 16575
rect 5089 16541 5123 16575
rect 7481 16541 7515 16575
rect 8033 16541 8067 16575
rect 8125 16541 8159 16575
rect 14289 16541 14323 16575
rect 15761 16541 15795 16575
rect 15853 16541 15887 16575
rect 17969 16541 18003 16575
rect 19441 16541 19475 16575
rect 19533 16541 19567 16575
rect 21741 16541 21775 16575
rect 24685 16541 24719 16575
rect 24777 16541 24811 16575
rect 6469 16473 6503 16507
rect 17417 16473 17451 16507
rect 4629 16405 4663 16439
rect 4905 16405 4939 16439
rect 9045 16405 9079 16439
rect 12541 16405 12575 16439
rect 13185 16405 13219 16439
rect 13461 16405 13495 16439
rect 16865 16405 16899 16439
rect 18797 16405 18831 16439
rect 20085 16405 20119 16439
rect 21097 16405 21131 16439
rect 23121 16405 23155 16439
rect 23673 16405 23707 16439
rect 25237 16405 25271 16439
rect 2513 16201 2547 16235
rect 2697 16201 2731 16235
rect 4813 16201 4847 16235
rect 4997 16201 5031 16235
rect 7665 16201 7699 16235
rect 9965 16201 9999 16235
rect 14381 16201 14415 16235
rect 14933 16201 14967 16235
rect 15945 16201 15979 16235
rect 19901 16201 19935 16235
rect 21281 16201 21315 16235
rect 23121 16201 23155 16235
rect 23489 16201 23523 16235
rect 25053 16201 25087 16235
rect 2237 16133 2271 16167
rect 7021 16133 7055 16167
rect 10701 16133 10735 16167
rect 14749 16133 14783 16167
rect 21741 16133 21775 16167
rect 3157 16065 3191 16099
rect 3341 16065 3375 16099
rect 5457 16065 5491 16099
rect 5549 16065 5583 16099
rect 6101 16065 6135 16099
rect 11253 16065 11287 16099
rect 11437 16065 11471 16099
rect 15577 16065 15611 16099
rect 16957 16065 16991 16099
rect 18613 16065 18647 16099
rect 20545 16065 20579 16099
rect 22477 16065 22511 16099
rect 22661 16065 22695 16099
rect 1409 15997 1443 16031
rect 4169 15997 4203 16031
rect 6653 15997 6687 16031
rect 6837 15997 6871 16031
rect 8033 15997 8067 16031
rect 8300 15997 8334 16031
rect 11161 15997 11195 16031
rect 12449 15997 12483 16031
rect 12716 15997 12750 16031
rect 16681 15997 16715 16031
rect 18429 15997 18463 16031
rect 20361 15997 20395 16031
rect 21925 15997 21959 16031
rect 23673 15997 23707 16031
rect 23929 15997 23963 16031
rect 1685 15929 1719 15963
rect 3065 15929 3099 15963
rect 5365 15929 5399 15963
rect 12265 15929 12299 15963
rect 15301 15929 15335 15963
rect 16313 15929 16347 15963
rect 18521 15929 18555 15963
rect 20269 15929 20303 15963
rect 21557 15929 21591 15963
rect 22385 15929 22419 15963
rect 3801 15861 3835 15895
rect 4445 15861 4479 15895
rect 9413 15861 9447 15895
rect 10793 15861 10827 15895
rect 11897 15861 11931 15895
rect 13829 15861 13863 15895
rect 15393 15861 15427 15895
rect 17417 15861 17451 15895
rect 17785 15861 17819 15895
rect 18061 15861 18095 15895
rect 19165 15861 19199 15895
rect 19441 15861 19475 15895
rect 22017 15861 22051 15895
rect 25605 15861 25639 15895
rect 1777 15657 1811 15691
rect 2789 15657 2823 15691
rect 6837 15657 6871 15691
rect 7941 15657 7975 15691
rect 8309 15657 8343 15691
rect 10057 15657 10091 15691
rect 13461 15657 13495 15691
rect 14105 15657 14139 15691
rect 17141 15657 17175 15691
rect 17693 15657 17727 15691
rect 20913 15657 20947 15691
rect 22661 15657 22695 15691
rect 23489 15657 23523 15691
rect 24041 15657 24075 15691
rect 24961 15657 24995 15691
rect 4997 15589 5031 15623
rect 6193 15589 6227 15623
rect 6469 15589 6503 15623
rect 7481 15589 7515 15623
rect 10425 15589 10459 15623
rect 10762 15589 10796 15623
rect 12817 15589 12851 15623
rect 18512 15589 18546 15623
rect 23029 15589 23063 15623
rect 24593 15589 24627 15623
rect 1685 15521 1719 15555
rect 2145 15521 2179 15555
rect 4077 15521 4111 15555
rect 5457 15521 5491 15555
rect 6653 15521 6687 15555
rect 8401 15521 8435 15555
rect 9045 15521 9079 15555
rect 9505 15521 9539 15555
rect 10517 15521 10551 15555
rect 13369 15521 13403 15555
rect 15025 15521 15059 15555
rect 16028 15521 16062 15555
rect 20729 15521 20763 15555
rect 21281 15521 21315 15555
rect 22477 15521 22511 15555
rect 23949 15521 23983 15555
rect 25145 15521 25179 15555
rect 2237 15453 2271 15487
rect 2421 15453 2455 15487
rect 5549 15453 5583 15487
rect 5641 15453 5675 15487
rect 8585 15453 8619 15487
rect 13553 15453 13587 15487
rect 15761 15453 15795 15487
rect 18245 15453 18279 15487
rect 21373 15453 21407 15487
rect 21557 15453 21591 15487
rect 24225 15453 24259 15487
rect 4629 15385 4663 15419
rect 7849 15385 7883 15419
rect 20177 15385 20211 15419
rect 23581 15385 23615 15419
rect 25329 15385 25363 15419
rect 3249 15317 3283 15351
rect 3525 15317 3559 15351
rect 5089 15317 5123 15351
rect 11897 15317 11931 15351
rect 12541 15317 12575 15351
rect 13001 15317 13035 15351
rect 14565 15317 14599 15351
rect 15485 15317 15519 15351
rect 18061 15317 18095 15351
rect 19625 15317 19659 15351
rect 22017 15317 22051 15351
rect 1593 15113 1627 15147
rect 2881 15113 2915 15147
rect 3065 15113 3099 15147
rect 7665 15113 7699 15147
rect 9229 15113 9263 15147
rect 12449 15113 12483 15147
rect 13553 15113 13587 15147
rect 13921 15113 13955 15147
rect 16221 15113 16255 15147
rect 16773 15113 16807 15147
rect 17509 15113 17543 15147
rect 19073 15113 19107 15147
rect 21741 15113 21775 15147
rect 22201 15113 22235 15147
rect 23029 15113 23063 15147
rect 23673 15113 23707 15147
rect 24685 15113 24719 15147
rect 25421 15113 25455 15147
rect 2053 14977 2087 15011
rect 2237 14977 2271 15011
rect 1961 14841 1995 14875
rect 4537 15045 4571 15079
rect 10057 15045 10091 15079
rect 14197 15045 14231 15079
rect 18061 15045 18095 15079
rect 25053 15045 25087 15079
rect 6561 14977 6595 15011
rect 11069 14977 11103 15011
rect 11253 14977 11287 15011
rect 13093 14977 13127 15011
rect 18613 14977 18647 15011
rect 24133 14977 24167 15011
rect 24225 14977 24259 15011
rect 3157 14909 3191 14943
rect 3413 14909 3447 14943
rect 5181 14909 5215 14943
rect 5641 14909 5675 14943
rect 7849 14909 7883 14943
rect 8116 14909 8150 14943
rect 10517 14909 10551 14943
rect 10977 14909 11011 14943
rect 14841 14909 14875 14943
rect 17877 14909 17911 14943
rect 18429 14909 18463 14943
rect 19809 14909 19843 14943
rect 22293 14909 22327 14943
rect 24041 14909 24075 14943
rect 25237 14909 25271 14943
rect 25789 14909 25823 14943
rect 12817 14841 12851 14875
rect 15086 14841 15120 14875
rect 18521 14841 18555 14875
rect 20054 14841 20088 14875
rect 23489 14841 23523 14875
rect 2605 14773 2639 14807
rect 2881 14773 2915 14807
rect 5549 14773 5583 14807
rect 5825 14773 5859 14807
rect 6193 14773 6227 14807
rect 6837 14773 6871 14807
rect 7297 14773 7331 14807
rect 10609 14773 10643 14807
rect 11621 14773 11655 14807
rect 12265 14773 12299 14807
rect 12909 14773 12943 14807
rect 14657 14773 14691 14807
rect 17693 14773 17727 14807
rect 19625 14773 19659 14807
rect 21189 14773 21223 14807
rect 22477 14773 22511 14807
rect 2881 14569 2915 14603
rect 4537 14569 4571 14603
rect 5181 14569 5215 14603
rect 7665 14569 7699 14603
rect 8677 14569 8711 14603
rect 9413 14569 9447 14603
rect 11069 14569 11103 14603
rect 12173 14569 12207 14603
rect 15761 14569 15795 14603
rect 16773 14569 16807 14603
rect 20269 14569 20303 14603
rect 20913 14569 20947 14603
rect 21925 14569 21959 14603
rect 22293 14569 22327 14603
rect 22477 14569 22511 14603
rect 23765 14569 23799 14603
rect 25513 14569 25547 14603
rect 1768 14501 1802 14535
rect 8033 14501 8067 14535
rect 9045 14501 9079 14535
rect 9934 14501 9968 14535
rect 12633 14501 12667 14535
rect 20729 14501 20763 14535
rect 22937 14501 22971 14535
rect 25145 14501 25179 14535
rect 4445 14433 4479 14467
rect 5457 14433 5491 14467
rect 5908 14433 5942 14467
rect 8125 14433 8159 14467
rect 12541 14433 12575 14467
rect 13553 14433 13587 14467
rect 13921 14433 13955 14467
rect 14657 14433 14691 14467
rect 15669 14433 15703 14467
rect 17141 14433 17175 14467
rect 18153 14433 18187 14467
rect 18604 14433 18638 14467
rect 21281 14433 21315 14467
rect 22845 14433 22879 14467
rect 24041 14433 24075 14467
rect 24777 14433 24811 14467
rect 25329 14433 25363 14467
rect 1501 14365 1535 14399
rect 4721 14365 4755 14399
rect 5641 14365 5675 14399
rect 9689 14365 9723 14399
rect 11713 14365 11747 14399
rect 12725 14365 12759 14399
rect 14197 14365 14231 14399
rect 16497 14365 16531 14399
rect 17233 14365 17267 14399
rect 17417 14365 17451 14399
rect 18337 14365 18371 14399
rect 21373 14365 21407 14399
rect 21465 14365 21499 14399
rect 23121 14365 23155 14399
rect 24225 14365 24259 14399
rect 8309 14297 8343 14331
rect 12081 14297 12115 14331
rect 19717 14297 19751 14331
rect 3525 14229 3559 14263
rect 3893 14229 3927 14263
rect 4077 14229 4111 14263
rect 7021 14229 7055 14263
rect 13185 14229 13219 14263
rect 15025 14229 15059 14263
rect 1869 14025 1903 14059
rect 6837 14025 6871 14059
rect 7849 14025 7883 14059
rect 10149 14025 10183 14059
rect 10701 14025 10735 14059
rect 11805 14025 11839 14059
rect 12449 14025 12483 14059
rect 14013 14025 14047 14059
rect 15577 14025 15611 14059
rect 17417 14025 17451 14059
rect 20085 14025 20119 14059
rect 21005 14025 21039 14059
rect 23029 14025 23063 14059
rect 23489 14025 23523 14059
rect 25605 14025 25639 14059
rect 4353 13957 4387 13991
rect 6469 13957 6503 13991
rect 6561 13957 6595 13991
rect 13553 13957 13587 13991
rect 16405 13957 16439 13991
rect 19441 13957 19475 13991
rect 22017 13957 22051 13991
rect 25053 13957 25087 13991
rect 4813 13889 4847 13923
rect 5733 13889 5767 13923
rect 6285 13889 6319 13923
rect 7297 13889 7331 13923
rect 7481 13889 7515 13923
rect 8677 13889 8711 13923
rect 13093 13889 13127 13923
rect 14565 13889 14599 13923
rect 15025 13889 15059 13923
rect 15945 13889 15979 13923
rect 17049 13889 17083 13923
rect 18061 13889 18095 13923
rect 21557 13889 21591 13923
rect 2237 13821 2271 13855
rect 2421 13821 2455 13855
rect 2677 13821 2711 13855
rect 5089 13821 5123 13855
rect 6469 13821 6503 13855
rect 7205 13821 7239 13855
rect 8217 13821 8251 13855
rect 8769 13821 8803 13855
rect 9025 13821 9059 13855
rect 12173 13821 12207 13855
rect 12909 13821 12943 13855
rect 14473 13821 14507 13855
rect 16865 13821 16899 13855
rect 20545 13821 20579 13855
rect 22385 13821 22419 13855
rect 22569 13821 22603 13855
rect 23673 13821 23707 13855
rect 23929 13821 23963 13855
rect 5641 13753 5675 13787
rect 11345 13753 11379 13787
rect 16221 13753 16255 13787
rect 16773 13753 16807 13787
rect 17877 13753 17911 13787
rect 18328 13753 18362 13787
rect 21465 13753 21499 13787
rect 3801 13685 3835 13719
rect 4905 13685 4939 13719
rect 5181 13685 5215 13719
rect 5549 13685 5583 13719
rect 11069 13685 11103 13719
rect 12817 13685 12851 13719
rect 13829 13685 13863 13719
rect 14381 13685 14415 13719
rect 20821 13685 20855 13719
rect 21373 13685 21407 13719
rect 1961 13481 1995 13515
rect 2881 13481 2915 13515
rect 3525 13481 3559 13515
rect 3893 13481 3927 13515
rect 4813 13481 4847 13515
rect 6929 13481 6963 13515
rect 8033 13481 8067 13515
rect 8401 13481 8435 13515
rect 8493 13481 8527 13515
rect 9137 13481 9171 13515
rect 9413 13481 9447 13515
rect 18061 13481 18095 13515
rect 19533 13481 19567 13515
rect 20177 13481 20211 13515
rect 20729 13481 20763 13515
rect 21557 13481 21591 13515
rect 22293 13481 22327 13515
rect 22753 13481 22787 13515
rect 4353 13413 4387 13447
rect 5273 13413 5307 13447
rect 9965 13413 9999 13447
rect 12541 13413 12575 13447
rect 21925 13413 21959 13447
rect 2789 13345 2823 13379
rect 4077 13345 4111 13379
rect 5816 13345 5850 13379
rect 10241 13345 10275 13379
rect 10497 13345 10531 13379
rect 12725 13345 12759 13379
rect 15568 13345 15602 13379
rect 17601 13345 17635 13379
rect 18429 13345 18463 13379
rect 21005 13345 21039 13379
rect 22109 13345 22143 13379
rect 24133 13345 24167 13379
rect 24869 13345 24903 13379
rect 1409 13277 1443 13311
rect 2973 13277 3007 13311
rect 5549 13277 5583 13311
rect 8585 13277 8619 13311
rect 15301 13277 15335 13311
rect 17969 13277 18003 13311
rect 18521 13277 18555 13311
rect 18613 13277 18647 13311
rect 19073 13277 19107 13311
rect 19625 13277 19659 13311
rect 24317 13277 24351 13311
rect 25421 13277 25455 13311
rect 21189 13209 21223 13243
rect 2237 13141 2271 13175
rect 2421 13141 2455 13175
rect 7481 13141 7515 13175
rect 11621 13141 11655 13175
rect 14013 13141 14047 13175
rect 14749 13141 14783 13175
rect 16681 13141 16715 13175
rect 23673 13141 23707 13175
rect 3157 12937 3191 12971
rect 3341 12937 3375 12971
rect 4997 12937 5031 12971
rect 5181 12937 5215 12971
rect 6193 12937 6227 12971
rect 6561 12937 6595 12971
rect 8769 12937 8803 12971
rect 9321 12937 9355 12971
rect 10609 12937 10643 12971
rect 13553 12937 13587 12971
rect 15761 12937 15795 12971
rect 16313 12937 16347 12971
rect 18245 12937 18279 12971
rect 19809 12937 19843 12971
rect 21005 12937 21039 12971
rect 21557 12937 21591 12971
rect 22109 12937 22143 12971
rect 22661 12937 22695 12971
rect 1685 12869 1719 12903
rect 10333 12869 10367 12903
rect 17509 12869 17543 12903
rect 19349 12869 19383 12903
rect 2237 12801 2271 12835
rect 2421 12801 2455 12835
rect 3893 12801 3927 12835
rect 5641 12801 5675 12835
rect 5825 12801 5859 12835
rect 9781 12801 9815 12835
rect 11253 12801 11287 12835
rect 11345 12801 11379 12835
rect 12909 12801 12943 12835
rect 13001 12801 13035 12835
rect 14105 12801 14139 12835
rect 14381 12801 14415 12835
rect 17877 12801 17911 12835
rect 18705 12801 18739 12835
rect 18889 12801 18923 12835
rect 19717 12801 19751 12835
rect 20361 12801 20395 12835
rect 23029 12801 23063 12835
rect 23489 12801 23523 12835
rect 3801 12733 3835 12767
rect 5549 12733 5583 12767
rect 6837 12733 6871 12767
rect 7093 12733 7127 12767
rect 9229 12733 9263 12767
rect 9505 12733 9539 12767
rect 11805 12733 11839 12767
rect 12817 12733 12851 12767
rect 18613 12733 18647 12767
rect 20177 12733 20211 12767
rect 21373 12733 21407 12767
rect 22477 12733 22511 12767
rect 23857 12733 23891 12767
rect 24124 12733 24158 12767
rect 4721 12665 4755 12699
rect 14626 12665 14660 12699
rect 16865 12665 16899 12699
rect 1777 12597 1811 12631
rect 2145 12597 2179 12631
rect 2789 12597 2823 12631
rect 3709 12597 3743 12631
rect 8217 12597 8251 12631
rect 10793 12597 10827 12631
rect 11161 12597 11195 12631
rect 12173 12597 12207 12631
rect 12449 12597 12483 12631
rect 13921 12597 13955 12631
rect 14013 12597 14047 12631
rect 16681 12597 16715 12631
rect 20269 12597 20303 12631
rect 25237 12597 25271 12631
rect 2053 12393 2087 12427
rect 3525 12393 3559 12427
rect 4629 12393 4663 12427
rect 5089 12393 5123 12427
rect 6101 12393 6135 12427
rect 6561 12393 6595 12427
rect 6837 12393 6871 12427
rect 7573 12393 7607 12427
rect 8217 12393 8251 12427
rect 8585 12393 8619 12427
rect 9965 12393 9999 12427
rect 12449 12393 12483 12427
rect 13461 12393 13495 12427
rect 15301 12393 15335 12427
rect 17325 12393 17359 12427
rect 18337 12393 18371 12427
rect 18705 12393 18739 12427
rect 19809 12393 19843 12427
rect 20177 12393 20211 12427
rect 21649 12393 21683 12427
rect 22753 12393 22787 12427
rect 3157 12325 3191 12359
rect 4353 12325 4387 12359
rect 10793 12325 10827 12359
rect 17969 12325 18003 12359
rect 19073 12325 19107 12359
rect 23940 12325 23974 12359
rect 2421 12257 2455 12291
rect 5457 12257 5491 12291
rect 7481 12257 7515 12291
rect 9505 12257 9539 12291
rect 11069 12257 11103 12291
rect 11336 12257 11370 12291
rect 13921 12257 13955 12291
rect 15669 12257 15703 12291
rect 17233 12257 17267 12291
rect 21465 12257 21499 12291
rect 22569 12257 22603 12291
rect 2513 12189 2547 12223
rect 2697 12189 2731 12223
rect 5549 12189 5583 12223
rect 5733 12189 5767 12223
rect 7757 12189 7791 12223
rect 10057 12189 10091 12223
rect 14013 12189 14047 12223
rect 14197 12189 14231 12223
rect 15761 12189 15795 12223
rect 15853 12189 15887 12223
rect 17417 12189 17451 12223
rect 19165 12189 19199 12223
rect 19257 12189 19291 12223
rect 23673 12189 23707 12223
rect 1961 12121 1995 12155
rect 3801 12121 3835 12155
rect 13553 12121 13587 12155
rect 16865 12121 16899 12155
rect 7113 12053 7147 12087
rect 13001 12053 13035 12087
rect 14565 12053 14599 12087
rect 15025 12053 15059 12087
rect 16405 12053 16439 12087
rect 16773 12053 16807 12087
rect 23581 12053 23615 12087
rect 25053 12053 25087 12087
rect 2421 11849 2455 11883
rect 3985 11849 4019 11883
rect 7205 11849 7239 11883
rect 7481 11849 7515 11883
rect 7849 11849 7883 11883
rect 10793 11849 10827 11883
rect 11805 11849 11839 11883
rect 11989 11849 12023 11883
rect 12449 11849 12483 11883
rect 14013 11849 14047 11883
rect 15945 11849 15979 11883
rect 17417 11849 17451 11883
rect 17693 11849 17727 11883
rect 18797 11849 18831 11883
rect 19441 11849 19475 11883
rect 21925 11849 21959 11883
rect 22385 11849 22419 11883
rect 22661 11849 22695 11883
rect 23949 11849 23983 11883
rect 24961 11849 24995 11883
rect 25697 11849 25731 11883
rect 1777 11713 1811 11747
rect 2145 11713 2179 11747
rect 2881 11713 2915 11747
rect 3065 11713 3099 11747
rect 3893 11713 3927 11747
rect 4445 11713 4479 11747
rect 4537 11713 4571 11747
rect 5549 11713 5583 11747
rect 8585 11713 8619 11747
rect 11253 11713 11287 11747
rect 11437 11713 11471 11747
rect 18337 11781 18371 11815
rect 13001 11713 13035 11747
rect 14381 11713 14415 11747
rect 15577 11713 15611 11747
rect 16497 11713 16531 11747
rect 19625 11713 19659 11747
rect 21465 11713 21499 11747
rect 23029 11713 23063 11747
rect 24501 11713 24535 11747
rect 10609 11645 10643 11679
rect 11989 11645 12023 11679
rect 12909 11645 12943 11679
rect 13645 11645 13679 11679
rect 14841 11645 14875 11679
rect 16405 11645 16439 11679
rect 22477 11645 22511 11679
rect 23489 11645 23523 11679
rect 24317 11645 24351 11679
rect 25513 11645 25547 11679
rect 26065 11645 26099 11679
rect 2789 11577 2823 11611
rect 10333 11577 10367 11611
rect 11161 11577 11195 11611
rect 12817 11577 12851 11611
rect 15301 11577 15335 11611
rect 24409 11577 24443 11611
rect 3525 11509 3559 11543
rect 4353 11509 4387 11543
rect 5089 11509 5123 11543
rect 12173 11509 12207 11543
rect 14933 11509 14967 11543
rect 15393 11509 15427 11543
rect 17049 11509 17083 11543
rect 19165 11509 19199 11543
rect 1869 11305 1903 11339
rect 2053 11305 2087 11339
rect 3801 11305 3835 11339
rect 4077 11305 4111 11339
rect 4445 11305 4479 11339
rect 5549 11305 5583 11339
rect 10885 11305 10919 11339
rect 12081 11305 12115 11339
rect 12449 11305 12483 11339
rect 13093 11305 13127 11339
rect 14105 11305 14139 11339
rect 15025 11305 15059 11339
rect 15301 11305 15335 11339
rect 16405 11305 16439 11339
rect 22385 11305 22419 11339
rect 22937 11305 22971 11339
rect 23673 11305 23707 11339
rect 24777 11305 24811 11339
rect 3433 11237 3467 11271
rect 13553 11237 13587 11271
rect 24133 11237 24167 11271
rect 2421 11169 2455 11203
rect 3065 11169 3099 11203
rect 12541 11169 12575 11203
rect 14013 11169 14047 11203
rect 15669 11169 15703 11203
rect 15761 11169 15795 11203
rect 23489 11169 23523 11203
rect 24593 11169 24627 11203
rect 2513 11101 2547 11135
rect 2605 11101 2639 11135
rect 4537 11101 4571 11135
rect 4721 11101 4755 11135
rect 12725 11101 12759 11135
rect 14197 11101 14231 11135
rect 15945 11101 15979 11135
rect 16865 11101 16899 11135
rect 5089 11033 5123 11067
rect 11253 11033 11287 11067
rect 13645 11033 13679 11067
rect 24409 11033 24443 11067
rect 2421 10761 2455 10795
rect 4169 10761 4203 10795
rect 4537 10761 4571 10795
rect 4813 10761 4847 10795
rect 12173 10761 12207 10795
rect 14013 10761 14047 10795
rect 14289 10761 14323 10795
rect 14565 10761 14599 10795
rect 23949 10761 23983 10795
rect 24501 10761 24535 10795
rect 3065 10625 3099 10659
rect 11805 10625 11839 10659
rect 13185 10625 13219 10659
rect 15117 10625 15151 10659
rect 16313 10625 16347 10659
rect 12909 10557 12943 10591
rect 14933 10557 14967 10591
rect 24593 10557 24627 10591
rect 25145 10557 25179 10591
rect 1777 10489 1811 10523
rect 2881 10489 2915 10523
rect 15025 10489 15059 10523
rect 16681 10489 16715 10523
rect 2053 10421 2087 10455
rect 2789 10421 2823 10455
rect 3433 10421 3467 10455
rect 12541 10421 12575 10455
rect 13001 10421 13035 10455
rect 13553 10421 13587 10455
rect 15577 10421 15611 10455
rect 16037 10421 16071 10455
rect 24777 10421 24811 10455
rect 1593 10217 1627 10251
rect 2053 10217 2087 10251
rect 3065 10217 3099 10251
rect 12265 10217 12299 10251
rect 12633 10217 12667 10251
rect 12725 10217 12759 10251
rect 13277 10217 13311 10251
rect 14657 10217 14691 10251
rect 15025 10217 15059 10251
rect 15301 10217 15335 10251
rect 15669 10217 15703 10251
rect 24777 10217 24811 10251
rect 12173 10149 12207 10183
rect 1409 10081 1443 10115
rect 2513 10081 2547 10115
rect 15761 10081 15795 10115
rect 24593 10081 24627 10115
rect 12909 10013 12943 10047
rect 14105 10013 14139 10047
rect 15853 10013 15887 10047
rect 2697 9945 2731 9979
rect 13737 9877 13771 9911
rect 2605 9673 2639 9707
rect 12633 9673 12667 9707
rect 13001 9673 13035 9707
rect 15761 9673 15795 9707
rect 16037 9673 16071 9707
rect 24685 9673 24719 9707
rect 27077 9673 27111 9707
rect 14105 9605 14139 9639
rect 15393 9605 15427 9639
rect 12265 9537 12299 9571
rect 14657 9537 14691 9571
rect 1409 9469 1443 9503
rect 1961 9469 1995 9503
rect 14565 9401 14599 9435
rect 1593 9333 1627 9367
rect 14013 9333 14047 9367
rect 14473 9333 14507 9367
rect 1685 9129 1719 9163
rect 14197 8789 14231 8823
rect 23857 8585 23891 8619
rect 23673 8381 23707 8415
rect 24225 8381 24259 8415
rect 24225 5865 24259 5899
rect 24041 5729 24075 5763
rect 24041 5321 24075 5355
rect 24133 4777 24167 4811
rect 24593 4709 24627 4743
rect 24501 4641 24535 4675
rect 24777 4573 24811 4607
rect 24133 4165 24167 4199
rect 24869 4097 24903 4131
rect 24593 3893 24627 3927
rect 11989 2601 12023 2635
rect 12449 2601 12483 2635
rect 14013 2601 14047 2635
rect 25329 2601 25363 2635
rect 12878 2533 12912 2567
rect 12633 2465 12667 2499
rect 25145 2465 25179 2499
rect 25697 2465 25731 2499
rect 24225 2261 24259 2295
<< metal1 >>
rect 8662 27412 8668 27464
rect 8720 27452 8726 27464
rect 8754 27452 8760 27464
rect 8720 27424 8760 27452
rect 8720 27412 8726 27424
rect 8754 27412 8760 27424
rect 8812 27412 8818 27464
rect 27062 27452 27068 27464
rect 27023 27424 27068 27452
rect 27062 27412 27068 27424
rect 27120 27412 27126 27464
rect 3510 26256 3516 26308
rect 3568 26296 3574 26308
rect 8386 26296 8392 26308
rect 3568 26268 8392 26296
rect 3568 26256 3574 26268
rect 8386 26256 8392 26268
rect 8444 26256 8450 26308
rect 4246 25984 4252 26036
rect 4304 26024 4310 26036
rect 17770 26024 17776 26036
rect 4304 25996 17776 26024
rect 4304 25984 4310 25996
rect 17770 25984 17776 25996
rect 17828 25984 17834 26036
rect 14366 25916 14372 25968
rect 14424 25956 14430 25968
rect 20346 25956 20352 25968
rect 14424 25928 20352 25956
rect 14424 25916 14430 25928
rect 20346 25916 20352 25928
rect 20404 25916 20410 25968
rect 14550 25848 14556 25900
rect 14608 25888 14614 25900
rect 24026 25888 24032 25900
rect 14608 25860 24032 25888
rect 14608 25848 14614 25860
rect 24026 25848 24032 25860
rect 24084 25848 24090 25900
rect 16850 25820 16856 25832
rect 13372 25792 16856 25820
rect 3602 25644 3608 25696
rect 3660 25684 3666 25696
rect 13372 25684 13400 25792
rect 16850 25780 16856 25792
rect 16908 25780 16914 25832
rect 13446 25712 13452 25764
rect 13504 25752 13510 25764
rect 25038 25752 25044 25764
rect 13504 25724 25044 25752
rect 13504 25712 13510 25724
rect 25038 25712 25044 25724
rect 25096 25712 25102 25764
rect 3660 25656 13400 25684
rect 3660 25644 3666 25656
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 4154 25440 4160 25492
rect 4212 25480 4218 25492
rect 4249 25483 4307 25489
rect 4249 25480 4261 25483
rect 4212 25452 4261 25480
rect 4212 25440 4218 25452
rect 4249 25449 4261 25452
rect 4295 25449 4307 25483
rect 4249 25443 4307 25449
rect 4338 25440 4344 25492
rect 4396 25480 4402 25492
rect 5353 25483 5411 25489
rect 5353 25480 5365 25483
rect 4396 25452 5365 25480
rect 4396 25440 4402 25452
rect 5353 25449 5365 25452
rect 5399 25449 5411 25483
rect 5353 25443 5411 25449
rect 10505 25483 10563 25489
rect 10505 25449 10517 25483
rect 10551 25480 10563 25483
rect 14366 25480 14372 25492
rect 10551 25452 14372 25480
rect 10551 25449 10563 25452
rect 10505 25443 10563 25449
rect 14366 25440 14372 25452
rect 14424 25440 14430 25492
rect 15933 25483 15991 25489
rect 15933 25449 15945 25483
rect 15979 25480 15991 25483
rect 16114 25480 16120 25492
rect 15979 25452 16120 25480
rect 15979 25449 15991 25452
rect 15933 25443 15991 25449
rect 16114 25440 16120 25452
rect 16172 25440 16178 25492
rect 16482 25440 16488 25492
rect 16540 25480 16546 25492
rect 17313 25483 17371 25489
rect 17313 25480 17325 25483
rect 16540 25452 17325 25480
rect 16540 25440 16546 25452
rect 17313 25449 17325 25452
rect 17359 25449 17371 25483
rect 17313 25443 17371 25449
rect 18141 25483 18199 25489
rect 18141 25449 18153 25483
rect 18187 25480 18199 25483
rect 18785 25483 18843 25489
rect 18785 25480 18797 25483
rect 18187 25452 18797 25480
rect 18187 25449 18199 25452
rect 18141 25443 18199 25449
rect 18785 25449 18797 25452
rect 18831 25480 18843 25483
rect 20898 25480 20904 25492
rect 18831 25452 20904 25480
rect 18831 25449 18843 25452
rect 18785 25443 18843 25449
rect 20898 25440 20904 25452
rect 20956 25440 20962 25492
rect 24762 25480 24768 25492
rect 24723 25452 24768 25480
rect 24762 25440 24768 25452
rect 24820 25440 24826 25492
rect 8665 25415 8723 25421
rect 8665 25381 8677 25415
rect 8711 25412 8723 25415
rect 13633 25415 13691 25421
rect 13633 25412 13645 25415
rect 8711 25384 13645 25412
rect 8711 25381 8723 25384
rect 8665 25375 8723 25381
rect 13633 25381 13645 25384
rect 13679 25412 13691 25415
rect 13998 25412 14004 25424
rect 13679 25384 14004 25412
rect 13679 25381 13691 25384
rect 13633 25375 13691 25381
rect 13998 25372 14004 25384
rect 14056 25372 14062 25424
rect 14921 25415 14979 25421
rect 14921 25412 14933 25415
rect 14292 25384 14933 25412
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 2038 25344 2044 25356
rect 1443 25316 2044 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 2038 25304 2044 25316
rect 2096 25304 2102 25356
rect 2501 25347 2559 25353
rect 2501 25313 2513 25347
rect 2547 25344 2559 25347
rect 3418 25344 3424 25356
rect 2547 25316 3424 25344
rect 2547 25313 2559 25316
rect 2501 25307 2559 25313
rect 3418 25304 3424 25316
rect 3476 25304 3482 25356
rect 4065 25347 4123 25353
rect 4065 25313 4077 25347
rect 4111 25344 4123 25347
rect 4522 25344 4528 25356
rect 4111 25316 4528 25344
rect 4111 25313 4123 25316
rect 4065 25307 4123 25313
rect 4522 25304 4528 25316
rect 4580 25304 4586 25356
rect 5166 25344 5172 25356
rect 5127 25316 5172 25344
rect 5166 25304 5172 25316
rect 5224 25304 5230 25356
rect 6178 25304 6184 25356
rect 6236 25344 6242 25356
rect 7469 25347 7527 25353
rect 7469 25344 7481 25347
rect 6236 25316 7481 25344
rect 6236 25304 6242 25316
rect 7469 25313 7481 25316
rect 7515 25313 7527 25347
rect 7469 25307 7527 25313
rect 7561 25347 7619 25353
rect 7561 25313 7573 25347
rect 7607 25344 7619 25347
rect 7926 25344 7932 25356
rect 7607 25316 7932 25344
rect 7607 25313 7619 25316
rect 7561 25307 7619 25313
rect 7926 25304 7932 25316
rect 7984 25304 7990 25356
rect 10318 25344 10324 25356
rect 10279 25316 10324 25344
rect 10318 25304 10324 25316
rect 10376 25304 10382 25356
rect 11425 25347 11483 25353
rect 11425 25313 11437 25347
rect 11471 25344 11483 25347
rect 12066 25344 12072 25356
rect 11471 25316 12072 25344
rect 11471 25313 11483 25316
rect 11425 25307 11483 25313
rect 12066 25304 12072 25316
rect 12124 25304 12130 25356
rect 12986 25344 12992 25356
rect 12947 25316 12992 25344
rect 12986 25304 12992 25316
rect 13044 25304 13050 25356
rect 14292 25353 14320 25384
rect 14921 25381 14933 25384
rect 14967 25412 14979 25415
rect 20254 25412 20260 25424
rect 14967 25384 20260 25412
rect 14967 25381 14979 25384
rect 14921 25375 14979 25381
rect 20254 25372 20260 25384
rect 20312 25372 20318 25424
rect 14277 25347 14335 25353
rect 14277 25313 14289 25347
rect 14323 25313 14335 25347
rect 14277 25307 14335 25313
rect 17129 25347 17187 25353
rect 17129 25313 17141 25347
rect 17175 25344 17187 25347
rect 17497 25347 17555 25353
rect 17497 25344 17509 25347
rect 17175 25316 17509 25344
rect 17175 25313 17187 25316
rect 17129 25307 17187 25313
rect 17497 25313 17509 25316
rect 17543 25313 17555 25347
rect 17497 25307 17555 25313
rect 17773 25347 17831 25353
rect 17773 25313 17785 25347
rect 17819 25344 17831 25347
rect 18693 25347 18751 25353
rect 18693 25344 18705 25347
rect 17819 25316 18705 25344
rect 17819 25313 17831 25316
rect 17773 25307 17831 25313
rect 18693 25313 18705 25316
rect 18739 25344 18751 25347
rect 19794 25344 19800 25356
rect 18739 25316 19800 25344
rect 18739 25313 18751 25316
rect 18693 25307 18751 25313
rect 19794 25304 19800 25316
rect 19852 25304 19858 25356
rect 19981 25347 20039 25353
rect 19981 25313 19993 25347
rect 20027 25344 20039 25347
rect 20070 25344 20076 25356
rect 20027 25316 20076 25344
rect 20027 25313 20039 25316
rect 19981 25307 20039 25313
rect 20070 25304 20076 25316
rect 20128 25304 20134 25356
rect 21913 25347 21971 25353
rect 21913 25313 21925 25347
rect 21959 25344 21971 25347
rect 22462 25344 22468 25356
rect 21959 25316 22468 25344
rect 21959 25313 21971 25316
rect 21913 25307 21971 25313
rect 22462 25304 22468 25316
rect 22520 25304 22526 25356
rect 23842 25304 23848 25356
rect 23900 25344 23906 25356
rect 24581 25347 24639 25353
rect 24581 25344 24593 25347
rect 23900 25316 24593 25344
rect 23900 25304 23906 25316
rect 24581 25313 24593 25316
rect 24627 25344 24639 25347
rect 25130 25344 25136 25356
rect 24627 25316 25136 25344
rect 24627 25313 24639 25316
rect 24581 25307 24639 25313
rect 25130 25304 25136 25316
rect 25188 25304 25194 25356
rect 7742 25276 7748 25288
rect 7703 25248 7748 25276
rect 7742 25236 7748 25248
rect 7800 25236 7806 25288
rect 13081 25279 13139 25285
rect 13081 25245 13093 25279
rect 13127 25245 13139 25279
rect 13262 25276 13268 25288
rect 13223 25248 13268 25276
rect 13081 25239 13139 25245
rect 1581 25211 1639 25217
rect 1581 25177 1593 25211
rect 1627 25208 1639 25211
rect 2958 25208 2964 25220
rect 1627 25180 2964 25208
rect 1627 25177 1639 25180
rect 1581 25171 1639 25177
rect 2958 25168 2964 25180
rect 3016 25168 3022 25220
rect 6733 25211 6791 25217
rect 6733 25177 6745 25211
rect 6779 25208 6791 25211
rect 7374 25208 7380 25220
rect 6779 25180 7380 25208
rect 6779 25177 6791 25180
rect 6733 25171 6791 25177
rect 7374 25168 7380 25180
rect 7432 25168 7438 25220
rect 12250 25168 12256 25220
rect 12308 25208 12314 25220
rect 13096 25208 13124 25239
rect 13262 25236 13268 25248
rect 13320 25236 13326 25288
rect 15289 25279 15347 25285
rect 15289 25245 15301 25279
rect 15335 25276 15347 25279
rect 15838 25276 15844 25288
rect 15335 25248 15844 25276
rect 15335 25245 15347 25248
rect 15289 25239 15347 25245
rect 15838 25236 15844 25248
rect 15896 25236 15902 25288
rect 16022 25276 16028 25288
rect 15983 25248 16028 25276
rect 16022 25236 16028 25248
rect 16080 25236 16086 25288
rect 16209 25279 16267 25285
rect 16209 25245 16221 25279
rect 16255 25276 16267 25279
rect 16390 25276 16396 25288
rect 16255 25248 16396 25276
rect 16255 25245 16267 25248
rect 16209 25239 16267 25245
rect 16390 25236 16396 25248
rect 16448 25236 16454 25288
rect 17678 25236 17684 25288
rect 17736 25276 17742 25288
rect 18877 25279 18935 25285
rect 18877 25276 18889 25279
rect 17736 25248 18889 25276
rect 17736 25236 17742 25248
rect 18877 25245 18889 25248
rect 18923 25245 18935 25279
rect 18877 25239 18935 25245
rect 22189 25279 22247 25285
rect 22189 25245 22201 25279
rect 22235 25276 22247 25279
rect 22278 25276 22284 25288
rect 22235 25248 22284 25276
rect 22235 25245 22247 25248
rect 22189 25239 22247 25245
rect 22278 25236 22284 25248
rect 22336 25236 22342 25288
rect 14093 25211 14151 25217
rect 12308 25180 13952 25208
rect 12308 25168 12314 25180
rect 2685 25143 2743 25149
rect 2685 25109 2697 25143
rect 2731 25140 2743 25143
rect 2866 25140 2872 25152
rect 2731 25112 2872 25140
rect 2731 25109 2743 25112
rect 2685 25103 2743 25109
rect 2866 25100 2872 25112
rect 2924 25100 2930 25152
rect 4706 25140 4712 25152
rect 4667 25112 4712 25140
rect 4706 25100 4712 25112
rect 4764 25100 4770 25152
rect 7098 25140 7104 25152
rect 7059 25112 7104 25140
rect 7098 25100 7104 25112
rect 7156 25100 7162 25152
rect 8573 25143 8631 25149
rect 8573 25109 8585 25143
rect 8619 25140 8631 25143
rect 8938 25140 8944 25152
rect 8619 25112 8944 25140
rect 8619 25109 8631 25112
rect 8573 25103 8631 25109
rect 8938 25100 8944 25112
rect 8996 25100 9002 25152
rect 11606 25140 11612 25152
rect 11567 25112 11612 25140
rect 11606 25100 11612 25112
rect 11664 25100 11670 25152
rect 12621 25143 12679 25149
rect 12621 25109 12633 25143
rect 12667 25140 12679 25143
rect 13814 25140 13820 25152
rect 12667 25112 13820 25140
rect 12667 25109 12679 25112
rect 12621 25103 12679 25109
rect 13814 25100 13820 25112
rect 13872 25100 13878 25152
rect 13924 25140 13952 25180
rect 14093 25177 14105 25211
rect 14139 25208 14151 25211
rect 14366 25208 14372 25220
rect 14139 25180 14372 25208
rect 14139 25177 14151 25180
rect 14093 25171 14151 25177
rect 14366 25168 14372 25180
rect 14424 25168 14430 25220
rect 14461 25211 14519 25217
rect 14461 25177 14473 25211
rect 14507 25208 14519 25211
rect 17586 25208 17592 25220
rect 14507 25180 17592 25208
rect 14507 25177 14519 25180
rect 14461 25171 14519 25177
rect 17586 25168 17592 25180
rect 17644 25168 17650 25220
rect 19426 25208 19432 25220
rect 17880 25180 19432 25208
rect 15470 25140 15476 25152
rect 13924 25112 15476 25140
rect 15470 25100 15476 25112
rect 15528 25100 15534 25152
rect 15565 25143 15623 25149
rect 15565 25109 15577 25143
rect 15611 25140 15623 25143
rect 16206 25140 16212 25152
rect 15611 25112 16212 25140
rect 15611 25109 15623 25112
rect 15565 25103 15623 25109
rect 16206 25100 16212 25112
rect 16264 25100 16270 25152
rect 16574 25140 16580 25152
rect 16535 25112 16580 25140
rect 16574 25100 16580 25112
rect 16632 25100 16638 25152
rect 17037 25143 17095 25149
rect 17037 25109 17049 25143
rect 17083 25140 17095 25143
rect 17497 25143 17555 25149
rect 17497 25140 17509 25143
rect 17083 25112 17509 25140
rect 17083 25109 17095 25112
rect 17037 25103 17095 25109
rect 17497 25109 17509 25112
rect 17543 25140 17555 25143
rect 17880 25140 17908 25180
rect 19426 25168 19432 25180
rect 19484 25168 19490 25220
rect 20165 25211 20223 25217
rect 20165 25177 20177 25211
rect 20211 25208 20223 25211
rect 24762 25208 24768 25220
rect 20211 25180 24768 25208
rect 20211 25177 20223 25180
rect 20165 25171 20223 25177
rect 24762 25168 24768 25180
rect 24820 25168 24826 25220
rect 18322 25140 18328 25152
rect 17543 25112 17908 25140
rect 18283 25112 18328 25140
rect 17543 25109 17555 25112
rect 17497 25103 17555 25109
rect 18322 25100 18328 25112
rect 18380 25100 18386 25152
rect 18690 25100 18696 25152
rect 18748 25140 18754 25152
rect 19337 25143 19395 25149
rect 19337 25140 19349 25143
rect 18748 25112 19349 25140
rect 18748 25100 18754 25112
rect 19337 25109 19349 25112
rect 19383 25109 19395 25143
rect 19337 25103 19395 25109
rect 19889 25143 19947 25149
rect 19889 25109 19901 25143
rect 19935 25140 19947 25143
rect 19978 25140 19984 25152
rect 19935 25112 19984 25140
rect 19935 25109 19947 25112
rect 19889 25103 19947 25109
rect 19978 25100 19984 25112
rect 20036 25100 20042 25152
rect 21453 25143 21511 25149
rect 21453 25109 21465 25143
rect 21499 25140 21511 25143
rect 21542 25140 21548 25152
rect 21499 25112 21548 25140
rect 21499 25109 21511 25112
rect 21453 25103 21511 25109
rect 21542 25100 21548 25112
rect 21600 25100 21606 25152
rect 21726 25140 21732 25152
rect 21687 25112 21732 25140
rect 21726 25100 21732 25112
rect 21784 25100 21790 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 3786 24936 3792 24948
rect 3747 24908 3792 24936
rect 3786 24896 3792 24908
rect 3844 24896 3850 24948
rect 3878 24896 3884 24948
rect 3936 24936 3942 24948
rect 4893 24939 4951 24945
rect 4893 24936 4905 24939
rect 3936 24908 4905 24936
rect 3936 24896 3942 24908
rect 4893 24905 4905 24908
rect 4939 24905 4951 24939
rect 4893 24899 4951 24905
rect 10318 24896 10324 24948
rect 10376 24936 10382 24948
rect 10505 24939 10563 24945
rect 10505 24936 10517 24939
rect 10376 24908 10517 24936
rect 10376 24896 10382 24908
rect 10505 24905 10517 24908
rect 10551 24905 10563 24939
rect 10505 24899 10563 24905
rect 1854 24828 1860 24880
rect 1912 24868 1918 24880
rect 4706 24868 4712 24880
rect 1912 24840 4712 24868
rect 1912 24828 1918 24840
rect 4706 24828 4712 24840
rect 4764 24828 4770 24880
rect 7834 24868 7840 24880
rect 6840 24840 7840 24868
rect 4246 24800 4252 24812
rect 4207 24772 4252 24800
rect 4246 24760 4252 24772
rect 4304 24760 4310 24812
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24732 1455 24735
rect 2501 24735 2559 24741
rect 1443 24704 2452 24732
rect 1443 24701 1455 24704
rect 1397 24695 1455 24701
rect 2424 24608 2452 24704
rect 2501 24701 2513 24735
rect 2547 24732 2559 24735
rect 2590 24732 2596 24744
rect 2547 24704 2596 24732
rect 2547 24701 2559 24704
rect 2501 24695 2559 24701
rect 2590 24692 2596 24704
rect 2648 24732 2654 24744
rect 3421 24735 3479 24741
rect 3421 24732 3433 24735
rect 2648 24704 3433 24732
rect 2648 24692 2654 24704
rect 3421 24701 3433 24704
rect 3467 24701 3479 24735
rect 3421 24695 3479 24701
rect 3605 24735 3663 24741
rect 3605 24701 3617 24735
rect 3651 24732 3663 24735
rect 4154 24732 4160 24744
rect 3651 24704 4160 24732
rect 3651 24701 3663 24704
rect 3605 24695 3663 24701
rect 4154 24692 4160 24704
rect 4212 24732 4218 24744
rect 4264 24732 4292 24760
rect 4724 24741 4752 24828
rect 4798 24760 4804 24812
rect 4856 24800 4862 24812
rect 5350 24800 5356 24812
rect 4856 24772 5356 24800
rect 4856 24760 4862 24772
rect 5350 24760 5356 24772
rect 5408 24760 5414 24812
rect 6641 24803 6699 24809
rect 6641 24769 6653 24803
rect 6687 24800 6699 24803
rect 6840 24800 6868 24840
rect 7374 24800 7380 24812
rect 6687 24772 6868 24800
rect 7335 24772 7380 24800
rect 6687 24769 6699 24772
rect 6641 24763 6699 24769
rect 7374 24760 7380 24772
rect 7432 24760 7438 24812
rect 7576 24809 7604 24840
rect 7834 24828 7840 24840
rect 7892 24828 7898 24880
rect 7561 24803 7619 24809
rect 7561 24769 7573 24803
rect 7607 24769 7619 24803
rect 8938 24800 8944 24812
rect 8899 24772 8944 24800
rect 7561 24763 7619 24769
rect 8938 24760 8944 24772
rect 8996 24760 9002 24812
rect 9125 24803 9183 24809
rect 9125 24769 9137 24803
rect 9171 24800 9183 24803
rect 10520 24800 10548 24899
rect 11606 24896 11612 24948
rect 11664 24936 11670 24948
rect 11664 24908 16160 24936
rect 11664 24896 11670 24908
rect 13170 24828 13176 24880
rect 13228 24868 13234 24880
rect 13630 24868 13636 24880
rect 13228 24840 13636 24868
rect 13228 24828 13234 24840
rect 13630 24828 13636 24840
rect 13688 24828 13694 24880
rect 16132 24868 16160 24908
rect 18322 24896 18328 24948
rect 18380 24936 18386 24948
rect 25406 24936 25412 24948
rect 18380 24908 25412 24936
rect 18380 24896 18386 24908
rect 25406 24896 25412 24908
rect 25464 24896 25470 24948
rect 19518 24868 19524 24880
rect 16132 24840 19524 24868
rect 19518 24828 19524 24840
rect 19576 24828 19582 24880
rect 19794 24868 19800 24880
rect 19755 24840 19800 24868
rect 19794 24828 19800 24840
rect 19852 24828 19858 24880
rect 20070 24828 20076 24880
rect 20128 24868 20134 24880
rect 20809 24871 20867 24877
rect 20809 24868 20821 24871
rect 20128 24840 20821 24868
rect 20128 24828 20134 24840
rect 20809 24837 20821 24840
rect 20855 24837 20867 24871
rect 20809 24831 20867 24837
rect 21726 24828 21732 24880
rect 21784 24868 21790 24880
rect 25130 24868 25136 24880
rect 21784 24840 21956 24868
rect 25091 24840 25136 24868
rect 21784 24828 21790 24840
rect 11241 24803 11299 24809
rect 11241 24800 11253 24803
rect 9171 24772 9628 24800
rect 10520 24772 11253 24800
rect 9171 24769 9183 24772
rect 9125 24763 9183 24769
rect 4212 24704 4292 24732
rect 4709 24735 4767 24741
rect 4212 24692 4218 24704
rect 4709 24701 4721 24735
rect 4755 24701 4767 24735
rect 4709 24695 4767 24701
rect 5905 24735 5963 24741
rect 5905 24701 5917 24735
rect 5951 24732 5963 24735
rect 7098 24732 7104 24744
rect 5951 24704 7104 24732
rect 5951 24701 5963 24704
rect 5905 24695 5963 24701
rect 7098 24692 7104 24704
rect 7156 24732 7162 24744
rect 7285 24735 7343 24741
rect 7285 24732 7297 24735
rect 7156 24704 7297 24732
rect 7156 24692 7162 24704
rect 7285 24701 7297 24704
rect 7331 24701 7343 24735
rect 7285 24695 7343 24701
rect 8389 24667 8447 24673
rect 8389 24633 8401 24667
rect 8435 24664 8447 24667
rect 8846 24664 8852 24676
rect 8435 24636 8852 24664
rect 8435 24633 8447 24636
rect 8389 24627 8447 24633
rect 8846 24624 8852 24636
rect 8904 24624 8910 24676
rect 1578 24596 1584 24608
rect 1539 24568 1584 24596
rect 1578 24556 1584 24568
rect 1636 24556 1642 24608
rect 2038 24596 2044 24608
rect 1999 24568 2044 24596
rect 2038 24556 2044 24568
rect 2096 24556 2102 24608
rect 2406 24596 2412 24608
rect 2367 24568 2412 24596
rect 2406 24556 2412 24568
rect 2464 24556 2470 24608
rect 2682 24596 2688 24608
rect 2643 24568 2688 24596
rect 2682 24556 2688 24568
rect 2740 24556 2746 24608
rect 3145 24599 3203 24605
rect 3145 24565 3157 24599
rect 3191 24596 3203 24599
rect 3418 24596 3424 24608
rect 3191 24568 3424 24596
rect 3191 24565 3203 24568
rect 3145 24559 3203 24565
rect 3418 24556 3424 24568
rect 3476 24556 3482 24608
rect 4522 24596 4528 24608
rect 4483 24568 4528 24596
rect 4522 24556 4528 24568
rect 4580 24556 4586 24608
rect 5166 24556 5172 24608
rect 5224 24596 5230 24608
rect 5261 24599 5319 24605
rect 5261 24596 5273 24599
rect 5224 24568 5273 24596
rect 5224 24556 5230 24568
rect 5261 24565 5273 24568
rect 5307 24565 5319 24599
rect 6178 24596 6184 24608
rect 6139 24568 6184 24596
rect 5261 24559 5319 24565
rect 6178 24556 6184 24568
rect 6236 24556 6242 24608
rect 6917 24599 6975 24605
rect 6917 24565 6929 24599
rect 6963 24596 6975 24599
rect 7006 24596 7012 24608
rect 6963 24568 7012 24596
rect 6963 24565 6975 24568
rect 6917 24559 6975 24565
rect 7006 24556 7012 24568
rect 7064 24556 7070 24608
rect 7926 24596 7932 24608
rect 7887 24568 7932 24596
rect 7926 24556 7932 24568
rect 7984 24556 7990 24608
rect 8478 24596 8484 24608
rect 8439 24568 8484 24596
rect 8478 24556 8484 24568
rect 8536 24556 8542 24608
rect 9600 24605 9628 24772
rect 11241 24769 11253 24772
rect 11287 24769 11299 24803
rect 12250 24800 12256 24812
rect 12211 24772 12256 24800
rect 11241 24763 11299 24769
rect 12250 24760 12256 24772
rect 12308 24760 12314 24812
rect 13446 24800 13452 24812
rect 12544 24772 13452 24800
rect 12544 24741 12572 24772
rect 13446 24760 13452 24772
rect 13504 24760 13510 24812
rect 14277 24803 14335 24809
rect 14277 24769 14289 24803
rect 14323 24800 14335 24803
rect 14366 24800 14372 24812
rect 14323 24772 14372 24800
rect 14323 24769 14335 24772
rect 14277 24763 14335 24769
rect 14366 24760 14372 24772
rect 14424 24760 14430 24812
rect 15749 24803 15807 24809
rect 15749 24769 15761 24803
rect 15795 24769 15807 24803
rect 17770 24800 17776 24812
rect 17731 24772 17776 24800
rect 15749 24763 15807 24769
rect 11057 24735 11115 24741
rect 11057 24732 11069 24735
rect 10980 24704 11069 24732
rect 9858 24624 9864 24676
rect 9916 24664 9922 24676
rect 10045 24667 10103 24673
rect 10045 24664 10057 24667
rect 9916 24636 10057 24664
rect 9916 24624 9922 24636
rect 10045 24633 10057 24636
rect 10091 24633 10103 24667
rect 10045 24627 10103 24633
rect 10980 24608 11008 24704
rect 11057 24701 11069 24704
rect 11103 24701 11115 24735
rect 11057 24695 11115 24701
rect 12529 24735 12587 24741
rect 12529 24701 12541 24735
rect 12575 24701 12587 24735
rect 12529 24695 12587 24701
rect 13173 24735 13231 24741
rect 13173 24701 13185 24735
rect 13219 24732 13231 24735
rect 13262 24732 13268 24744
rect 13219 24704 13268 24732
rect 13219 24701 13231 24704
rect 13173 24695 13231 24701
rect 13262 24692 13268 24704
rect 13320 24732 13326 24744
rect 13630 24732 13636 24744
rect 13320 24704 13636 24732
rect 13320 24692 13326 24704
rect 13630 24692 13636 24704
rect 13688 24692 13694 24744
rect 13998 24732 14004 24744
rect 13959 24704 14004 24732
rect 13998 24692 14004 24704
rect 14056 24692 14062 24744
rect 14734 24692 14740 24744
rect 14792 24732 14798 24744
rect 15764 24732 15792 24763
rect 17770 24760 17776 24772
rect 17828 24760 17834 24812
rect 18782 24800 18788 24812
rect 18743 24772 18788 24800
rect 18782 24760 18788 24772
rect 18840 24760 18846 24812
rect 21928 24809 21956 24840
rect 25130 24828 25136 24840
rect 25188 24828 25194 24880
rect 20349 24803 20407 24809
rect 20349 24769 20361 24803
rect 20395 24800 20407 24803
rect 21913 24803 21971 24809
rect 20395 24772 20429 24800
rect 20395 24769 20407 24772
rect 20349 24763 20407 24769
rect 21913 24769 21925 24803
rect 21959 24769 21971 24803
rect 21913 24763 21971 24769
rect 14792 24704 15792 24732
rect 14792 24692 14798 24704
rect 12618 24624 12624 24676
rect 12676 24664 12682 24676
rect 13449 24667 13507 24673
rect 13449 24664 13461 24667
rect 12676 24636 13461 24664
rect 12676 24624 12682 24636
rect 13449 24633 13461 24636
rect 13495 24664 13507 24667
rect 14090 24664 14096 24676
rect 13495 24636 14096 24664
rect 13495 24633 13507 24636
rect 13449 24627 13507 24633
rect 14090 24624 14096 24636
rect 14148 24624 14154 24676
rect 15565 24667 15623 24673
rect 15565 24664 15577 24667
rect 15120 24636 15577 24664
rect 15120 24608 15148 24636
rect 15565 24633 15577 24636
rect 15611 24633 15623 24667
rect 17788 24664 17816 24760
rect 18414 24692 18420 24744
rect 18472 24732 18478 24744
rect 18693 24735 18751 24741
rect 18693 24732 18705 24735
rect 18472 24704 18705 24732
rect 18472 24692 18478 24704
rect 18693 24701 18705 24704
rect 18739 24701 18751 24735
rect 18693 24695 18751 24701
rect 19337 24735 19395 24741
rect 19337 24701 19349 24735
rect 19383 24732 19395 24735
rect 20364 24732 20392 24763
rect 22646 24760 22652 24812
rect 22704 24800 22710 24812
rect 23198 24800 23204 24812
rect 22704 24772 23204 24800
rect 22704 24760 22710 24772
rect 23198 24760 23204 24772
rect 23256 24760 23262 24812
rect 24026 24760 24032 24812
rect 24084 24800 24090 24812
rect 24397 24803 24455 24809
rect 24397 24800 24409 24803
rect 24084 24772 24409 24800
rect 24084 24760 24090 24772
rect 24397 24769 24409 24772
rect 24443 24769 24455 24803
rect 24397 24763 24455 24769
rect 21450 24732 21456 24744
rect 19383 24704 21456 24732
rect 19383 24701 19395 24704
rect 19337 24695 19395 24701
rect 21450 24692 21456 24704
rect 21508 24692 21514 24744
rect 24412 24732 24440 24763
rect 24581 24735 24639 24741
rect 24581 24732 24593 24735
rect 24412 24704 24593 24732
rect 24581 24701 24593 24704
rect 24627 24701 24639 24735
rect 24581 24695 24639 24701
rect 18322 24664 18328 24676
rect 17788 24636 18328 24664
rect 15565 24627 15623 24633
rect 18322 24624 18328 24636
rect 18380 24664 18386 24676
rect 18601 24667 18659 24673
rect 18601 24664 18613 24667
rect 18380 24636 18613 24664
rect 18380 24624 18386 24636
rect 18601 24633 18613 24636
rect 18647 24633 18659 24667
rect 18601 24627 18659 24633
rect 19705 24667 19763 24673
rect 19705 24633 19717 24667
rect 19751 24664 19763 24667
rect 21174 24664 21180 24676
rect 19751 24636 20300 24664
rect 21135 24636 21180 24664
rect 19751 24633 19763 24636
rect 19705 24627 19763 24633
rect 9585 24599 9643 24605
rect 9585 24565 9597 24599
rect 9631 24596 9643 24599
rect 9950 24596 9956 24608
rect 9631 24568 9956 24596
rect 9631 24565 9643 24568
rect 9585 24559 9643 24565
rect 9950 24556 9956 24568
rect 10008 24556 10014 24608
rect 10962 24596 10968 24608
rect 10923 24568 10968 24596
rect 10962 24556 10968 24568
rect 11020 24556 11026 24608
rect 11885 24599 11943 24605
rect 11885 24565 11897 24599
rect 11931 24596 11943 24599
rect 11974 24596 11980 24608
rect 11931 24568 11980 24596
rect 11931 24565 11943 24568
rect 11885 24559 11943 24565
rect 11974 24556 11980 24568
rect 12032 24556 12038 24608
rect 12710 24596 12716 24608
rect 12671 24568 12716 24596
rect 12710 24556 12716 24568
rect 12768 24556 12774 24608
rect 13633 24599 13691 24605
rect 13633 24565 13645 24599
rect 13679 24596 13691 24599
rect 13998 24596 14004 24608
rect 13679 24568 14004 24596
rect 13679 24565 13691 24568
rect 13633 24559 13691 24565
rect 13998 24556 14004 24568
rect 14056 24556 14062 24608
rect 14734 24596 14740 24608
rect 14695 24568 14740 24596
rect 14734 24556 14740 24568
rect 14792 24556 14798 24608
rect 15102 24596 15108 24608
rect 15063 24568 15108 24596
rect 15102 24556 15108 24568
rect 15160 24556 15166 24608
rect 15197 24599 15255 24605
rect 15197 24565 15209 24599
rect 15243 24596 15255 24599
rect 15470 24596 15476 24608
rect 15243 24568 15476 24596
rect 15243 24565 15255 24568
rect 15197 24559 15255 24565
rect 15470 24556 15476 24568
rect 15528 24556 15534 24608
rect 15657 24599 15715 24605
rect 15657 24565 15669 24599
rect 15703 24596 15715 24599
rect 15838 24596 15844 24608
rect 15703 24568 15844 24596
rect 15703 24565 15715 24568
rect 15657 24559 15715 24565
rect 15838 24556 15844 24568
rect 15896 24556 15902 24608
rect 16114 24556 16120 24608
rect 16172 24596 16178 24608
rect 16209 24599 16267 24605
rect 16209 24596 16221 24599
rect 16172 24568 16221 24596
rect 16172 24556 16178 24568
rect 16209 24565 16221 24568
rect 16255 24565 16267 24599
rect 16209 24559 16267 24565
rect 16390 24556 16396 24608
rect 16448 24596 16454 24608
rect 16577 24599 16635 24605
rect 16577 24596 16589 24599
rect 16448 24568 16589 24596
rect 16448 24556 16454 24568
rect 16577 24565 16589 24568
rect 16623 24565 16635 24599
rect 16577 24559 16635 24565
rect 17037 24599 17095 24605
rect 17037 24565 17049 24599
rect 17083 24596 17095 24599
rect 17310 24596 17316 24608
rect 17083 24568 17316 24596
rect 17083 24565 17095 24568
rect 17037 24559 17095 24565
rect 17310 24556 17316 24568
rect 17368 24556 17374 24608
rect 17497 24599 17555 24605
rect 17497 24565 17509 24599
rect 17543 24596 17555 24599
rect 17678 24596 17684 24608
rect 17543 24568 17684 24596
rect 17543 24565 17555 24568
rect 17497 24559 17555 24565
rect 17678 24556 17684 24568
rect 17736 24556 17742 24608
rect 18230 24596 18236 24608
rect 18191 24568 18236 24596
rect 18230 24556 18236 24568
rect 18288 24556 18294 24608
rect 19334 24556 19340 24608
rect 19392 24596 19398 24608
rect 19978 24596 19984 24608
rect 19392 24568 19984 24596
rect 19392 24556 19398 24568
rect 19978 24556 19984 24568
rect 20036 24596 20042 24608
rect 20272 24605 20300 24636
rect 21174 24624 21180 24636
rect 21232 24664 21238 24676
rect 21542 24664 21548 24676
rect 21232 24636 21548 24664
rect 21232 24624 21238 24636
rect 21542 24624 21548 24636
rect 21600 24664 21606 24676
rect 21729 24667 21787 24673
rect 21729 24664 21741 24667
rect 21600 24636 21741 24664
rect 21600 24624 21606 24636
rect 21729 24633 21741 24636
rect 21775 24633 21787 24667
rect 21729 24627 21787 24633
rect 22646 24624 22652 24676
rect 22704 24664 22710 24676
rect 23106 24664 23112 24676
rect 22704 24636 23112 24664
rect 22704 24624 22710 24636
rect 23106 24624 23112 24636
rect 23164 24624 23170 24676
rect 20165 24599 20223 24605
rect 20165 24596 20177 24599
rect 20036 24568 20177 24596
rect 20036 24556 20042 24568
rect 20165 24565 20177 24568
rect 20211 24565 20223 24599
rect 20165 24559 20223 24565
rect 20257 24599 20315 24605
rect 20257 24565 20269 24599
rect 20303 24596 20315 24599
rect 20714 24596 20720 24608
rect 20303 24568 20720 24596
rect 20303 24565 20315 24568
rect 20257 24559 20315 24565
rect 20714 24556 20720 24568
rect 20772 24556 20778 24608
rect 21358 24596 21364 24608
rect 21319 24568 21364 24596
rect 21358 24556 21364 24568
rect 21416 24556 21422 24608
rect 21634 24556 21640 24608
rect 21692 24596 21698 24608
rect 21818 24596 21824 24608
rect 21692 24568 21824 24596
rect 21692 24556 21698 24568
rect 21818 24556 21824 24568
rect 21876 24556 21882 24608
rect 22462 24596 22468 24608
rect 22375 24568 22468 24596
rect 22462 24556 22468 24568
rect 22520 24596 22526 24608
rect 23382 24596 23388 24608
rect 22520 24568 23388 24596
rect 22520 24556 22526 24568
rect 23382 24556 23388 24568
rect 23440 24556 23446 24608
rect 24670 24556 24676 24608
rect 24728 24596 24734 24608
rect 24765 24599 24823 24605
rect 24765 24596 24777 24599
rect 24728 24568 24777 24596
rect 24728 24556 24734 24568
rect 24765 24565 24777 24568
rect 24811 24565 24823 24599
rect 24765 24559 24823 24565
rect 24854 24556 24860 24608
rect 24912 24596 24918 24608
rect 25130 24596 25136 24608
rect 24912 24568 25136 24596
rect 24912 24556 24918 24568
rect 25130 24556 25136 24568
rect 25188 24556 25194 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 2038 24392 2044 24404
rect 1999 24364 2044 24392
rect 2038 24352 2044 24364
rect 2096 24352 2102 24404
rect 4246 24392 4252 24404
rect 4207 24364 4252 24392
rect 4246 24352 4252 24364
rect 4304 24352 4310 24404
rect 8665 24395 8723 24401
rect 8665 24361 8677 24395
rect 8711 24392 8723 24395
rect 9582 24392 9588 24404
rect 8711 24364 9588 24392
rect 8711 24361 8723 24364
rect 8665 24355 8723 24361
rect 9582 24352 9588 24364
rect 9640 24352 9646 24404
rect 9674 24352 9680 24404
rect 9732 24392 9738 24404
rect 10137 24395 10195 24401
rect 10137 24392 10149 24395
rect 9732 24364 10149 24392
rect 9732 24352 9738 24364
rect 10137 24361 10149 24364
rect 10183 24361 10195 24395
rect 10137 24355 10195 24361
rect 12434 24352 12440 24404
rect 12492 24392 12498 24404
rect 12897 24395 12955 24401
rect 12897 24392 12909 24395
rect 12492 24364 12909 24392
rect 12492 24352 12498 24364
rect 12897 24361 12909 24364
rect 12943 24392 12955 24395
rect 12986 24392 12992 24404
rect 12943 24364 12992 24392
rect 12943 24361 12955 24364
rect 12897 24355 12955 24361
rect 12986 24352 12992 24364
rect 13044 24352 13050 24404
rect 13265 24395 13323 24401
rect 13265 24361 13277 24395
rect 13311 24392 13323 24395
rect 13446 24392 13452 24404
rect 13311 24364 13452 24392
rect 13311 24361 13323 24364
rect 13265 24355 13323 24361
rect 13446 24352 13452 24364
rect 13504 24352 13510 24404
rect 13998 24352 14004 24404
rect 14056 24392 14062 24404
rect 14645 24395 14703 24401
rect 14645 24392 14657 24395
rect 14056 24364 14657 24392
rect 14056 24352 14062 24364
rect 14645 24361 14657 24364
rect 14691 24392 14703 24395
rect 15286 24392 15292 24404
rect 14691 24364 15292 24392
rect 14691 24361 14703 24364
rect 14645 24355 14703 24361
rect 15286 24352 15292 24364
rect 15344 24352 15350 24404
rect 15473 24395 15531 24401
rect 15473 24361 15485 24395
rect 15519 24392 15531 24395
rect 15930 24392 15936 24404
rect 15519 24364 15936 24392
rect 15519 24361 15531 24364
rect 15473 24355 15531 24361
rect 15930 24352 15936 24364
rect 15988 24352 15994 24404
rect 16206 24392 16212 24404
rect 16167 24364 16212 24392
rect 16206 24352 16212 24364
rect 16264 24352 16270 24404
rect 18230 24352 18236 24404
rect 18288 24392 18294 24404
rect 19429 24395 19487 24401
rect 19429 24392 19441 24395
rect 18288 24364 19441 24392
rect 18288 24352 18294 24364
rect 19429 24361 19441 24364
rect 19475 24392 19487 24395
rect 19978 24392 19984 24404
rect 19475 24364 19984 24392
rect 19475 24361 19487 24364
rect 19429 24355 19487 24361
rect 19978 24352 19984 24364
rect 20036 24352 20042 24404
rect 20898 24392 20904 24404
rect 20859 24364 20904 24392
rect 20898 24352 20904 24364
rect 20956 24352 20962 24404
rect 22094 24352 22100 24404
rect 22152 24392 22158 24404
rect 23106 24392 23112 24404
rect 22152 24364 23112 24392
rect 22152 24352 22158 24364
rect 23106 24352 23112 24364
rect 23164 24352 23170 24404
rect 24118 24352 24124 24404
rect 24176 24392 24182 24404
rect 24765 24395 24823 24401
rect 24765 24392 24777 24395
rect 24176 24364 24777 24392
rect 24176 24352 24182 24364
rect 24765 24361 24777 24364
rect 24811 24361 24823 24395
rect 24765 24355 24823 24361
rect 9214 24284 9220 24336
rect 9272 24324 9278 24336
rect 9490 24324 9496 24336
rect 9272 24296 9496 24324
rect 9272 24284 9278 24296
rect 9490 24284 9496 24296
rect 9548 24324 9554 24336
rect 10042 24324 10048 24336
rect 9548 24296 10048 24324
rect 9548 24284 9554 24296
rect 10042 24284 10048 24296
rect 10100 24284 10106 24336
rect 11701 24327 11759 24333
rect 11701 24293 11713 24327
rect 11747 24324 11759 24327
rect 12066 24324 12072 24336
rect 11747 24296 12072 24324
rect 11747 24293 11759 24296
rect 11701 24287 11759 24293
rect 12066 24284 12072 24296
rect 12124 24324 12130 24336
rect 12161 24327 12219 24333
rect 12161 24324 12173 24327
rect 12124 24296 12173 24324
rect 12124 24284 12130 24296
rect 12161 24293 12173 24296
rect 12207 24293 12219 24327
rect 12161 24287 12219 24293
rect 15562 24284 15568 24336
rect 15620 24324 15626 24336
rect 15841 24327 15899 24333
rect 15841 24324 15853 24327
rect 15620 24296 15853 24324
rect 15620 24284 15626 24296
rect 15841 24293 15853 24296
rect 15887 24324 15899 24327
rect 16022 24324 16028 24336
rect 15887 24296 16028 24324
rect 15887 24293 15899 24296
rect 15841 24287 15899 24293
rect 16022 24284 16028 24296
rect 16080 24324 16086 24336
rect 16298 24324 16304 24336
rect 16080 24296 16304 24324
rect 16080 24284 16086 24296
rect 16298 24284 16304 24296
rect 16356 24284 16362 24336
rect 18414 24324 18420 24336
rect 18375 24296 18420 24324
rect 18414 24284 18420 24296
rect 18472 24284 18478 24336
rect 22738 24284 22744 24336
rect 22796 24324 22802 24336
rect 22925 24327 22983 24333
rect 22925 24324 22937 24327
rect 22796 24296 22937 24324
rect 22796 24284 22802 24296
rect 22925 24293 22937 24296
rect 22971 24293 22983 24327
rect 22925 24287 22983 24293
rect 1397 24259 1455 24265
rect 1397 24225 1409 24259
rect 1443 24256 1455 24259
rect 1670 24256 1676 24268
rect 1443 24228 1676 24256
rect 1443 24225 1455 24228
rect 1397 24219 1455 24225
rect 1670 24216 1676 24228
rect 1728 24216 1734 24268
rect 2498 24256 2504 24268
rect 2459 24228 2504 24256
rect 2498 24216 2504 24228
rect 2556 24216 2562 24268
rect 4062 24256 4068 24268
rect 4023 24228 4068 24256
rect 4062 24216 4068 24228
rect 4120 24216 4126 24268
rect 5534 24216 5540 24268
rect 5592 24256 5598 24268
rect 6069 24259 6127 24265
rect 6069 24256 6081 24259
rect 5592 24228 6081 24256
rect 5592 24216 5598 24228
rect 6069 24225 6081 24228
rect 6115 24225 6127 24259
rect 6069 24219 6127 24225
rect 8481 24259 8539 24265
rect 8481 24225 8493 24259
rect 8527 24256 8539 24259
rect 9030 24256 9036 24268
rect 8527 24228 9036 24256
rect 8527 24225 8539 24228
rect 8481 24219 8539 24225
rect 9030 24216 9036 24228
rect 9088 24216 9094 24268
rect 10134 24216 10140 24268
rect 10192 24256 10198 24268
rect 10870 24256 10876 24268
rect 10192 24228 10876 24256
rect 10192 24216 10198 24228
rect 10870 24216 10876 24228
rect 10928 24216 10934 24268
rect 11422 24216 11428 24268
rect 11480 24256 11486 24268
rect 12253 24259 12311 24265
rect 12253 24256 12265 24259
rect 11480 24228 12265 24256
rect 11480 24216 11486 24228
rect 12253 24225 12265 24228
rect 12299 24225 12311 24259
rect 12253 24219 12311 24225
rect 13538 24216 13544 24268
rect 13596 24256 13602 24268
rect 13725 24259 13783 24265
rect 13725 24256 13737 24259
rect 13596 24228 13737 24256
rect 13596 24216 13602 24228
rect 13725 24225 13737 24228
rect 13771 24225 13783 24259
rect 13725 24219 13783 24225
rect 13817 24259 13875 24265
rect 13817 24225 13829 24259
rect 13863 24256 13875 24259
rect 14550 24256 14556 24268
rect 13863 24228 14556 24256
rect 13863 24225 13875 24228
rect 13817 24219 13875 24225
rect 14550 24216 14556 24228
rect 14608 24216 14614 24268
rect 15289 24259 15347 24265
rect 15289 24256 15301 24259
rect 15028 24228 15301 24256
rect 5813 24191 5871 24197
rect 5813 24157 5825 24191
rect 5859 24157 5871 24191
rect 5813 24151 5871 24157
rect 10229 24191 10287 24197
rect 10229 24157 10241 24191
rect 10275 24157 10287 24191
rect 10229 24151 10287 24157
rect 1394 24012 1400 24064
rect 1452 24052 1458 24064
rect 1581 24055 1639 24061
rect 1581 24052 1593 24055
rect 1452 24024 1593 24052
rect 1452 24012 1458 24024
rect 1581 24021 1593 24024
rect 1627 24021 1639 24055
rect 1581 24015 1639 24021
rect 1762 24012 1768 24064
rect 1820 24052 1826 24064
rect 2685 24055 2743 24061
rect 2685 24052 2697 24055
rect 1820 24024 2697 24052
rect 1820 24012 1826 24024
rect 2685 24021 2697 24024
rect 2731 24021 2743 24055
rect 2685 24015 2743 24021
rect 4709 24055 4767 24061
rect 4709 24021 4721 24055
rect 4755 24052 4767 24055
rect 4890 24052 4896 24064
rect 4755 24024 4896 24052
rect 4755 24021 4767 24024
rect 4709 24015 4767 24021
rect 4890 24012 4896 24024
rect 4948 24012 4954 24064
rect 5828 24052 5856 24151
rect 9950 24080 9956 24132
rect 10008 24120 10014 24132
rect 10244 24120 10272 24151
rect 10686 24148 10692 24200
rect 10744 24188 10750 24200
rect 11057 24191 11115 24197
rect 11057 24188 11069 24191
rect 10744 24160 11069 24188
rect 10744 24148 10750 24160
rect 11057 24157 11069 24160
rect 11103 24157 11115 24191
rect 12342 24188 12348 24200
rect 12303 24160 12348 24188
rect 11057 24151 11115 24157
rect 12342 24148 12348 24160
rect 12400 24148 12406 24200
rect 13909 24191 13967 24197
rect 13909 24157 13921 24191
rect 13955 24157 13967 24191
rect 13909 24151 13967 24157
rect 10008 24092 10272 24120
rect 10008 24080 10014 24092
rect 13722 24080 13728 24132
rect 13780 24120 13786 24132
rect 13924 24120 13952 24151
rect 13780 24092 13952 24120
rect 13780 24080 13786 24092
rect 5994 24052 6000 24064
rect 5828 24024 6000 24052
rect 5994 24012 6000 24024
rect 6052 24012 6058 24064
rect 7098 24012 7104 24064
rect 7156 24052 7162 24064
rect 7193 24055 7251 24061
rect 7193 24052 7205 24055
rect 7156 24024 7205 24052
rect 7156 24012 7162 24024
rect 7193 24021 7205 24024
rect 7239 24021 7251 24055
rect 7193 24015 7251 24021
rect 7742 24012 7748 24064
rect 7800 24052 7806 24064
rect 7837 24055 7895 24061
rect 7837 24052 7849 24055
rect 7800 24024 7849 24052
rect 7800 24012 7806 24024
rect 7837 24021 7849 24024
rect 7883 24052 7895 24055
rect 8294 24052 8300 24064
rect 7883 24024 8300 24052
rect 7883 24021 7895 24024
rect 7837 24015 7895 24021
rect 8294 24012 8300 24024
rect 8352 24012 8358 24064
rect 8846 24012 8852 24064
rect 8904 24052 8910 24064
rect 9677 24055 9735 24061
rect 9677 24052 9689 24055
rect 8904 24024 9689 24052
rect 8904 24012 8910 24024
rect 9677 24021 9689 24024
rect 9723 24021 9735 24055
rect 9677 24015 9735 24021
rect 10781 24055 10839 24061
rect 10781 24021 10793 24055
rect 10827 24052 10839 24055
rect 11330 24052 11336 24064
rect 10827 24024 11336 24052
rect 10827 24021 10839 24024
rect 10781 24015 10839 24021
rect 11330 24012 11336 24024
rect 11388 24012 11394 24064
rect 11790 24052 11796 24064
rect 11751 24024 11796 24052
rect 11790 24012 11796 24024
rect 11848 24012 11854 24064
rect 13354 24052 13360 24064
rect 13315 24024 13360 24052
rect 13354 24012 13360 24024
rect 13412 24012 13418 24064
rect 14826 24012 14832 24064
rect 14884 24052 14890 24064
rect 15028 24061 15056 24228
rect 15289 24225 15301 24228
rect 15335 24225 15347 24259
rect 15289 24219 15347 24225
rect 16485 24259 16543 24265
rect 16485 24225 16497 24259
rect 16531 24256 16543 24259
rect 16574 24256 16580 24268
rect 16531 24228 16580 24256
rect 16531 24225 16543 24228
rect 16485 24219 16543 24225
rect 16574 24216 16580 24228
rect 16632 24216 16638 24268
rect 16758 24265 16764 24268
rect 16752 24219 16764 24265
rect 16816 24256 16822 24268
rect 19334 24256 19340 24268
rect 16816 24228 16852 24256
rect 19295 24228 19340 24256
rect 16758 24216 16764 24219
rect 16816 24216 16822 24228
rect 19334 24216 19340 24228
rect 19392 24256 19398 24268
rect 19981 24259 20039 24265
rect 19981 24256 19993 24259
rect 19392 24228 19993 24256
rect 19392 24216 19398 24228
rect 19981 24225 19993 24228
rect 20027 24225 20039 24259
rect 19981 24219 20039 24225
rect 21082 24216 21088 24268
rect 21140 24256 21146 24268
rect 21269 24259 21327 24265
rect 21269 24256 21281 24259
rect 21140 24228 21281 24256
rect 21140 24216 21146 24228
rect 21269 24225 21281 24228
rect 21315 24225 21327 24259
rect 21269 24219 21327 24225
rect 22373 24259 22431 24265
rect 22373 24225 22385 24259
rect 22419 24256 22431 24259
rect 22830 24256 22836 24268
rect 22419 24228 22836 24256
rect 22419 24225 22431 24228
rect 22373 24219 22431 24225
rect 22830 24216 22836 24228
rect 22888 24216 22894 24268
rect 24581 24259 24639 24265
rect 24581 24225 24593 24259
rect 24627 24256 24639 24259
rect 24670 24256 24676 24268
rect 24627 24228 24676 24256
rect 24627 24225 24639 24228
rect 24581 24219 24639 24225
rect 24670 24216 24676 24228
rect 24728 24216 24734 24268
rect 15102 24148 15108 24200
rect 15160 24188 15166 24200
rect 15930 24188 15936 24200
rect 15160 24160 15936 24188
rect 15160 24148 15166 24160
rect 15930 24148 15936 24160
rect 15988 24148 15994 24200
rect 19518 24188 19524 24200
rect 19479 24160 19524 24188
rect 19518 24148 19524 24160
rect 19576 24148 19582 24200
rect 20438 24148 20444 24200
rect 20496 24188 20502 24200
rect 21361 24191 21419 24197
rect 21361 24188 21373 24191
rect 20496 24160 21373 24188
rect 20496 24148 20502 24160
rect 21284 24132 21312 24160
rect 21361 24157 21373 24160
rect 21407 24157 21419 24191
rect 21361 24151 21419 24157
rect 21450 24148 21456 24200
rect 21508 24188 21514 24200
rect 23014 24188 23020 24200
rect 21508 24160 21553 24188
rect 22975 24160 23020 24188
rect 21508 24148 21514 24160
rect 23014 24148 23020 24160
rect 23072 24148 23078 24200
rect 17770 24080 17776 24132
rect 17828 24120 17834 24132
rect 18969 24123 19027 24129
rect 18969 24120 18981 24123
rect 17828 24092 18981 24120
rect 17828 24080 17834 24092
rect 18969 24089 18981 24092
rect 19015 24089 19027 24123
rect 18969 24083 19027 24089
rect 21266 24080 21272 24132
rect 21324 24080 21330 24132
rect 15013 24055 15071 24061
rect 15013 24052 15025 24055
rect 14884 24024 15025 24052
rect 14884 24012 14890 24024
rect 15013 24021 15025 24024
rect 15059 24021 15071 24055
rect 17862 24052 17868 24064
rect 17823 24024 17868 24052
rect 15013 24015 15071 24021
rect 17862 24012 17868 24024
rect 17920 24012 17926 24064
rect 18782 24052 18788 24064
rect 18743 24024 18788 24052
rect 18782 24012 18788 24024
rect 18840 24012 18846 24064
rect 20530 24052 20536 24064
rect 20491 24024 20536 24052
rect 20530 24012 20536 24024
rect 20588 24012 20594 24064
rect 22005 24055 22063 24061
rect 22005 24021 22017 24055
rect 22051 24052 22063 24055
rect 22186 24052 22192 24064
rect 22051 24024 22192 24052
rect 22051 24021 22063 24024
rect 22005 24015 22063 24021
rect 22186 24012 22192 24024
rect 22244 24012 22250 24064
rect 22370 24012 22376 24064
rect 22428 24052 22434 24064
rect 22465 24055 22523 24061
rect 22465 24052 22477 24055
rect 22428 24024 22477 24052
rect 22428 24012 22434 24024
rect 22465 24021 22477 24024
rect 22511 24021 22523 24055
rect 22465 24015 22523 24021
rect 23753 24055 23811 24061
rect 23753 24021 23765 24055
rect 23799 24052 23811 24055
rect 24026 24052 24032 24064
rect 23799 24024 24032 24052
rect 23799 24021 23811 24024
rect 23753 24015 23811 24021
rect 24026 24012 24032 24024
rect 24084 24012 24090 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2498 23808 2504 23860
rect 2556 23848 2562 23860
rect 2593 23851 2651 23857
rect 2593 23848 2605 23851
rect 2556 23820 2605 23848
rect 2556 23808 2562 23820
rect 2593 23817 2605 23820
rect 2639 23848 2651 23851
rect 5261 23851 5319 23857
rect 5261 23848 5273 23851
rect 2639 23820 5273 23848
rect 2639 23817 2651 23820
rect 2593 23811 2651 23817
rect 5261 23817 5273 23820
rect 5307 23817 5319 23851
rect 5261 23811 5319 23817
rect 7374 23808 7380 23860
rect 7432 23848 7438 23860
rect 8389 23851 8447 23857
rect 8389 23848 8401 23851
rect 7432 23820 8401 23848
rect 7432 23808 7438 23820
rect 8389 23817 8401 23820
rect 8435 23817 8447 23851
rect 9674 23848 9680 23860
rect 9635 23820 9680 23848
rect 8389 23811 8447 23817
rect 9674 23808 9680 23820
rect 9732 23808 9738 23860
rect 10042 23848 10048 23860
rect 10003 23820 10048 23848
rect 10042 23808 10048 23820
rect 10100 23808 10106 23860
rect 11885 23851 11943 23857
rect 11885 23817 11897 23851
rect 11931 23848 11943 23851
rect 12253 23851 12311 23857
rect 12253 23848 12265 23851
rect 11931 23820 12265 23848
rect 11931 23817 11943 23820
rect 11885 23811 11943 23817
rect 12253 23817 12265 23820
rect 12299 23848 12311 23851
rect 12342 23848 12348 23860
rect 12299 23820 12348 23848
rect 12299 23817 12311 23820
rect 12253 23811 12311 23817
rect 12342 23808 12348 23820
rect 12400 23808 12406 23860
rect 13538 23808 13544 23860
rect 13596 23848 13602 23860
rect 14737 23851 14795 23857
rect 14737 23848 14749 23851
rect 13596 23820 14749 23848
rect 13596 23808 13602 23820
rect 14737 23817 14749 23820
rect 14783 23817 14795 23851
rect 15378 23848 15384 23860
rect 15339 23820 15384 23848
rect 14737 23811 14795 23817
rect 15378 23808 15384 23820
rect 15436 23808 15442 23860
rect 16485 23851 16543 23857
rect 16485 23817 16497 23851
rect 16531 23848 16543 23851
rect 16758 23848 16764 23860
rect 16531 23820 16764 23848
rect 16531 23817 16543 23820
rect 16485 23811 16543 23817
rect 4062 23740 4068 23792
rect 4120 23780 4126 23792
rect 4157 23783 4215 23789
rect 4157 23780 4169 23783
rect 4120 23752 4169 23780
rect 4120 23740 4126 23752
rect 4157 23749 4169 23752
rect 4203 23780 4215 23783
rect 5074 23780 5080 23792
rect 4203 23752 5080 23780
rect 4203 23749 4215 23752
rect 4157 23743 4215 23749
rect 5074 23740 5080 23752
rect 5132 23780 5138 23792
rect 6638 23780 6644 23792
rect 5132 23752 6644 23780
rect 5132 23740 5138 23752
rect 6638 23740 6644 23752
rect 6696 23740 6702 23792
rect 10413 23783 10471 23789
rect 10413 23749 10425 23783
rect 10459 23780 10471 23783
rect 10870 23780 10876 23792
rect 10459 23752 10876 23780
rect 10459 23749 10471 23752
rect 10413 23743 10471 23749
rect 10870 23740 10876 23752
rect 10928 23740 10934 23792
rect 14366 23740 14372 23792
rect 14424 23780 14430 23792
rect 14461 23783 14519 23789
rect 14461 23780 14473 23783
rect 14424 23752 14473 23780
rect 14424 23740 14430 23752
rect 14461 23749 14473 23752
rect 14507 23780 14519 23783
rect 14550 23780 14556 23792
rect 14507 23752 14556 23780
rect 14507 23749 14519 23752
rect 14461 23743 14519 23749
rect 14550 23740 14556 23752
rect 14608 23740 14614 23792
rect 1854 23712 1860 23724
rect 1815 23684 1860 23712
rect 1854 23672 1860 23684
rect 1912 23672 1918 23724
rect 3786 23712 3792 23724
rect 3699 23684 3792 23712
rect 3786 23672 3792 23684
rect 3844 23712 3850 23724
rect 4985 23715 5043 23721
rect 4985 23712 4997 23715
rect 3844 23684 4997 23712
rect 3844 23672 3850 23684
rect 4985 23681 4997 23684
rect 5031 23681 5043 23715
rect 4985 23675 5043 23681
rect 6273 23715 6331 23721
rect 6273 23681 6285 23715
rect 6319 23712 6331 23715
rect 7282 23712 7288 23724
rect 6319 23684 7288 23712
rect 6319 23681 6331 23684
rect 6273 23675 6331 23681
rect 7282 23672 7288 23684
rect 7340 23672 7346 23724
rect 7466 23712 7472 23724
rect 7427 23684 7472 23712
rect 7466 23672 7472 23684
rect 7524 23672 7530 23724
rect 7929 23715 7987 23721
rect 7929 23681 7941 23715
rect 7975 23712 7987 23715
rect 8846 23712 8852 23724
rect 7975 23684 8852 23712
rect 7975 23681 7987 23684
rect 7929 23675 7987 23681
rect 8846 23672 8852 23684
rect 8904 23672 8910 23724
rect 8941 23715 8999 23721
rect 8941 23681 8953 23715
rect 8987 23681 8999 23715
rect 8941 23675 8999 23681
rect 11057 23715 11115 23721
rect 11057 23681 11069 23715
rect 11103 23712 11115 23715
rect 11330 23712 11336 23724
rect 11103 23684 11336 23712
rect 11103 23681 11115 23684
rect 11057 23675 11115 23681
rect 1581 23647 1639 23653
rect 1581 23613 1593 23647
rect 1627 23644 1639 23647
rect 2038 23644 2044 23656
rect 1627 23616 2044 23644
rect 1627 23613 1639 23616
rect 1581 23607 1639 23613
rect 2038 23604 2044 23616
rect 2096 23604 2102 23656
rect 2866 23644 2872 23656
rect 2827 23616 2872 23644
rect 2866 23604 2872 23616
rect 2924 23604 2930 23656
rect 4890 23644 4896 23656
rect 4851 23616 4896 23644
rect 4890 23604 4896 23616
rect 4948 23604 4954 23656
rect 5166 23604 5172 23656
rect 5224 23644 5230 23656
rect 5537 23647 5595 23653
rect 5537 23644 5549 23647
rect 5224 23616 5549 23644
rect 5224 23604 5230 23616
rect 5537 23613 5549 23616
rect 5583 23644 5595 23647
rect 5994 23644 6000 23656
rect 5583 23616 6000 23644
rect 5583 23613 5595 23616
rect 5537 23607 5595 23613
rect 5994 23604 6000 23616
rect 6052 23644 6058 23656
rect 6730 23644 6736 23656
rect 6052 23616 6736 23644
rect 6052 23604 6058 23616
rect 6730 23604 6736 23616
rect 6788 23604 6794 23656
rect 8478 23604 8484 23656
rect 8536 23644 8542 23656
rect 8757 23647 8815 23653
rect 8757 23644 8769 23647
rect 8536 23616 8769 23644
rect 8536 23604 8542 23616
rect 8757 23613 8769 23616
rect 8803 23613 8815 23647
rect 8757 23607 8815 23613
rect 2406 23536 2412 23588
rect 2464 23576 2470 23588
rect 5261 23579 5319 23585
rect 2464 23548 4844 23576
rect 2464 23536 2470 23548
rect 3050 23508 3056 23520
rect 3011 23480 3056 23508
rect 3050 23468 3056 23480
rect 3108 23468 3114 23520
rect 4430 23508 4436 23520
rect 4391 23480 4436 23508
rect 4430 23468 4436 23480
rect 4488 23468 4494 23520
rect 4816 23517 4844 23548
rect 5261 23545 5273 23579
rect 5307 23576 5319 23579
rect 6641 23579 6699 23585
rect 6641 23576 6653 23579
rect 5307 23548 6653 23576
rect 5307 23545 5319 23548
rect 5261 23539 5319 23545
rect 6641 23545 6653 23548
rect 6687 23576 6699 23579
rect 6687 23548 7236 23576
rect 6687 23545 6699 23548
rect 6641 23539 6699 23545
rect 4801 23511 4859 23517
rect 4801 23477 4813 23511
rect 4847 23508 4859 23511
rect 4890 23508 4896 23520
rect 4847 23480 4896 23508
rect 4847 23477 4859 23480
rect 4801 23471 4859 23477
rect 4890 23468 4896 23480
rect 4948 23468 4954 23520
rect 5534 23468 5540 23520
rect 5592 23508 5598 23520
rect 5813 23511 5871 23517
rect 5813 23508 5825 23511
rect 5592 23480 5825 23508
rect 5592 23468 5598 23480
rect 5813 23477 5825 23480
rect 5859 23477 5871 23511
rect 6822 23508 6828 23520
rect 6783 23480 6828 23508
rect 5813 23471 5871 23477
rect 6822 23468 6828 23480
rect 6880 23468 6886 23520
rect 7208 23517 7236 23548
rect 7282 23536 7288 23588
rect 7340 23576 7346 23588
rect 7926 23576 7932 23588
rect 7340 23548 7932 23576
rect 7340 23536 7346 23548
rect 7926 23536 7932 23548
rect 7984 23536 7990 23588
rect 8956 23576 8984 23675
rect 11330 23672 11336 23684
rect 11388 23672 11394 23724
rect 16025 23715 16083 23721
rect 16025 23681 16037 23715
rect 16071 23712 16083 23715
rect 16500 23712 16528 23811
rect 16758 23808 16764 23820
rect 16816 23808 16822 23860
rect 19429 23851 19487 23857
rect 19429 23817 19441 23851
rect 19475 23848 19487 23851
rect 19518 23848 19524 23860
rect 19475 23820 19524 23848
rect 19475 23817 19487 23820
rect 19429 23811 19487 23817
rect 19518 23808 19524 23820
rect 19576 23808 19582 23860
rect 19978 23848 19984 23860
rect 19939 23820 19984 23848
rect 19978 23808 19984 23820
rect 20036 23808 20042 23860
rect 20438 23848 20444 23860
rect 20399 23820 20444 23848
rect 20438 23808 20444 23820
rect 20496 23808 20502 23860
rect 23477 23851 23535 23857
rect 23477 23817 23489 23851
rect 23523 23848 23535 23851
rect 23934 23848 23940 23860
rect 23523 23820 23940 23848
rect 23523 23817 23535 23820
rect 23477 23811 23535 23817
rect 23934 23808 23940 23820
rect 23992 23808 23998 23860
rect 16574 23740 16580 23792
rect 16632 23780 16638 23792
rect 17218 23780 17224 23792
rect 16632 23752 17224 23780
rect 16632 23740 16638 23752
rect 17218 23740 17224 23752
rect 17276 23780 17282 23792
rect 17405 23783 17463 23789
rect 17405 23780 17417 23783
rect 17276 23752 17417 23780
rect 17276 23740 17282 23752
rect 17405 23749 17417 23752
rect 17451 23749 17463 23783
rect 17405 23743 17463 23749
rect 19334 23740 19340 23792
rect 19392 23780 19398 23792
rect 20533 23783 20591 23789
rect 20533 23780 20545 23783
rect 19392 23752 20545 23780
rect 19392 23740 19398 23752
rect 20533 23749 20545 23752
rect 20579 23749 20591 23783
rect 20533 23743 20591 23749
rect 16071 23684 16528 23712
rect 16071 23681 16083 23684
rect 16025 23675 16083 23681
rect 20714 23672 20720 23724
rect 20772 23712 20778 23724
rect 21085 23715 21143 23721
rect 21085 23712 21097 23715
rect 20772 23684 21097 23712
rect 20772 23672 20778 23684
rect 21085 23681 21097 23684
rect 21131 23712 21143 23715
rect 22002 23712 22008 23724
rect 21131 23684 22008 23712
rect 21131 23681 21143 23684
rect 21085 23675 21143 23681
rect 22002 23672 22008 23684
rect 22060 23672 22066 23724
rect 10778 23604 10784 23656
rect 10836 23644 10842 23656
rect 10873 23647 10931 23653
rect 10873 23644 10885 23647
rect 10836 23616 10885 23644
rect 10836 23604 10842 23616
rect 10873 23613 10885 23616
rect 10919 23613 10931 23647
rect 12434 23644 12440 23656
rect 12395 23616 12440 23644
rect 10873 23607 10931 23613
rect 12434 23604 12440 23616
rect 12492 23604 12498 23656
rect 15841 23647 15899 23653
rect 15841 23613 15853 23647
rect 15887 23644 15899 23647
rect 16206 23644 16212 23656
rect 15887 23616 16212 23644
rect 15887 23613 15899 23616
rect 15841 23607 15899 23613
rect 16206 23604 16212 23616
rect 16264 23604 16270 23656
rect 18049 23647 18107 23653
rect 18049 23613 18061 23647
rect 18095 23644 18107 23647
rect 18690 23644 18696 23656
rect 18095 23616 18696 23644
rect 18095 23613 18107 23616
rect 18049 23607 18107 23613
rect 18690 23604 18696 23616
rect 18748 23604 18754 23656
rect 22186 23604 22192 23656
rect 22244 23644 22250 23656
rect 22281 23647 22339 23653
rect 22281 23644 22293 23647
rect 22244 23616 22293 23644
rect 22244 23604 22250 23616
rect 22281 23613 22293 23616
rect 22327 23613 22339 23647
rect 23952 23644 23980 23808
rect 24210 23712 24216 23724
rect 24171 23684 24216 23712
rect 24210 23672 24216 23684
rect 24268 23672 24274 23724
rect 24121 23647 24179 23653
rect 24121 23644 24133 23647
rect 23952 23616 24133 23644
rect 22281 23607 22339 23613
rect 24121 23613 24133 23616
rect 24167 23613 24179 23647
rect 24121 23607 24179 23613
rect 24762 23604 24768 23656
rect 24820 23644 24826 23656
rect 25225 23647 25283 23653
rect 25225 23644 25237 23647
rect 24820 23616 25237 23644
rect 24820 23604 24826 23616
rect 25225 23613 25237 23616
rect 25271 23644 25283 23647
rect 25777 23647 25835 23653
rect 25777 23644 25789 23647
rect 25271 23616 25789 23644
rect 25271 23613 25283 23616
rect 25225 23607 25283 23613
rect 25777 23613 25789 23616
rect 25823 23613 25835 23647
rect 25777 23607 25835 23613
rect 8312 23548 8984 23576
rect 12704 23579 12762 23585
rect 8312 23520 8340 23548
rect 12704 23545 12716 23579
rect 12750 23545 12762 23579
rect 12704 23539 12762 23545
rect 7193 23511 7251 23517
rect 7193 23477 7205 23511
rect 7239 23508 7251 23511
rect 7374 23508 7380 23520
rect 7239 23480 7380 23508
rect 7239 23477 7251 23480
rect 7193 23471 7251 23477
rect 7374 23468 7380 23480
rect 7432 23468 7438 23520
rect 8294 23508 8300 23520
rect 8255 23480 8300 23508
rect 8294 23468 8300 23480
rect 8352 23468 8358 23520
rect 10686 23468 10692 23520
rect 10744 23508 10750 23520
rect 10781 23511 10839 23517
rect 10781 23508 10793 23511
rect 10744 23480 10793 23508
rect 10744 23468 10750 23480
rect 10781 23477 10793 23480
rect 10827 23477 10839 23511
rect 10781 23471 10839 23477
rect 10962 23468 10968 23520
rect 11020 23508 11026 23520
rect 11422 23508 11428 23520
rect 11020 23480 11428 23508
rect 11020 23468 11026 23480
rect 11422 23468 11428 23480
rect 11480 23468 11486 23520
rect 12342 23468 12348 23520
rect 12400 23508 12406 23520
rect 12728 23508 12756 23539
rect 15286 23536 15292 23588
rect 15344 23576 15350 23588
rect 15749 23579 15807 23585
rect 15749 23576 15761 23579
rect 15344 23548 15761 23576
rect 15344 23536 15350 23548
rect 15749 23545 15761 23548
rect 15795 23545 15807 23579
rect 17862 23576 17868 23588
rect 17775 23548 17868 23576
rect 15749 23539 15807 23545
rect 17862 23536 17868 23548
rect 17920 23576 17926 23588
rect 18316 23579 18374 23585
rect 18316 23576 18328 23579
rect 17920 23548 18328 23576
rect 17920 23536 17926 23548
rect 18316 23545 18328 23548
rect 18362 23576 18374 23579
rect 18782 23576 18788 23588
rect 18362 23548 18788 23576
rect 18362 23545 18374 23548
rect 18316 23539 18374 23545
rect 18782 23536 18788 23548
rect 18840 23536 18846 23588
rect 19150 23536 19156 23588
rect 19208 23576 19214 23588
rect 20530 23576 20536 23588
rect 19208 23548 20536 23576
rect 19208 23536 19214 23548
rect 20530 23536 20536 23548
rect 20588 23576 20594 23588
rect 20993 23579 21051 23585
rect 20993 23576 21005 23579
rect 20588 23548 21005 23576
rect 20588 23536 20594 23548
rect 20993 23545 21005 23548
rect 21039 23545 21051 23579
rect 22554 23576 22560 23588
rect 22515 23548 22560 23576
rect 20993 23539 21051 23545
rect 22554 23536 22560 23548
rect 22612 23536 22618 23588
rect 23934 23536 23940 23588
rect 23992 23576 23998 23588
rect 24670 23576 24676 23588
rect 23992 23548 24676 23576
rect 23992 23536 23998 23548
rect 24670 23536 24676 23548
rect 24728 23536 24734 23588
rect 12986 23508 12992 23520
rect 12400 23480 12992 23508
rect 12400 23468 12406 23480
rect 12986 23468 12992 23480
rect 13044 23468 13050 23520
rect 13817 23511 13875 23517
rect 13817 23477 13829 23511
rect 13863 23508 13875 23511
rect 13998 23508 14004 23520
rect 13863 23480 14004 23508
rect 13863 23477 13875 23480
rect 13817 23471 13875 23477
rect 13998 23468 14004 23480
rect 14056 23468 14062 23520
rect 15197 23511 15255 23517
rect 15197 23477 15209 23511
rect 15243 23508 15255 23511
rect 15378 23508 15384 23520
rect 15243 23480 15384 23508
rect 15243 23477 15255 23480
rect 15197 23471 15255 23477
rect 15378 23468 15384 23480
rect 15436 23468 15442 23520
rect 16942 23508 16948 23520
rect 16903 23480 16948 23508
rect 16942 23468 16948 23480
rect 17000 23468 17006 23520
rect 20806 23468 20812 23520
rect 20864 23508 20870 23520
rect 20901 23511 20959 23517
rect 20901 23508 20913 23511
rect 20864 23480 20913 23508
rect 20864 23468 20870 23480
rect 20901 23477 20913 23480
rect 20947 23477 20959 23511
rect 20901 23471 20959 23477
rect 21082 23468 21088 23520
rect 21140 23508 21146 23520
rect 21545 23511 21603 23517
rect 21545 23508 21557 23511
rect 21140 23480 21557 23508
rect 21140 23468 21146 23480
rect 21545 23477 21557 23480
rect 21591 23477 21603 23511
rect 21545 23471 21603 23477
rect 22189 23511 22247 23517
rect 22189 23477 22201 23511
rect 22235 23508 22247 23511
rect 22738 23508 22744 23520
rect 22235 23480 22744 23508
rect 22235 23477 22247 23480
rect 22189 23471 22247 23477
rect 22738 23468 22744 23480
rect 22796 23468 22802 23520
rect 22922 23468 22928 23520
rect 22980 23508 22986 23520
rect 23017 23511 23075 23517
rect 23017 23508 23029 23511
rect 22980 23480 23029 23508
rect 22980 23468 22986 23480
rect 23017 23477 23029 23480
rect 23063 23477 23075 23511
rect 23658 23508 23664 23520
rect 23619 23480 23664 23508
rect 23017 23471 23075 23477
rect 23658 23468 23664 23480
rect 23716 23468 23722 23520
rect 24026 23508 24032 23520
rect 23987 23480 24032 23508
rect 24026 23468 24032 23480
rect 24084 23468 24090 23520
rect 25406 23508 25412 23520
rect 25367 23480 25412 23508
rect 25406 23468 25412 23480
rect 25464 23468 25470 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 2866 23304 2872 23316
rect 2827 23276 2872 23304
rect 2866 23264 2872 23276
rect 2924 23264 2930 23316
rect 5534 23264 5540 23316
rect 5592 23304 5598 23316
rect 6457 23307 6515 23313
rect 6457 23304 6469 23307
rect 5592 23276 6469 23304
rect 5592 23264 5598 23276
rect 6457 23273 6469 23276
rect 6503 23273 6515 23307
rect 8018 23304 8024 23316
rect 7979 23276 8024 23304
rect 6457 23267 6515 23273
rect 8018 23264 8024 23276
rect 8076 23264 8082 23316
rect 8478 23264 8484 23316
rect 8536 23304 8542 23316
rect 8573 23307 8631 23313
rect 8573 23304 8585 23307
rect 8536 23276 8585 23304
rect 8536 23264 8542 23276
rect 8573 23273 8585 23276
rect 8619 23273 8631 23307
rect 8573 23267 8631 23273
rect 9674 23264 9680 23316
rect 9732 23304 9738 23316
rect 10134 23304 10140 23316
rect 9732 23276 10140 23304
rect 9732 23264 9738 23276
rect 10134 23264 10140 23276
rect 10192 23264 10198 23316
rect 12342 23304 12348 23316
rect 12303 23276 12348 23304
rect 12342 23264 12348 23276
rect 12400 23264 12406 23316
rect 13449 23307 13507 23313
rect 13449 23273 13461 23307
rect 13495 23273 13507 23307
rect 13906 23304 13912 23316
rect 13867 23276 13912 23304
rect 13449 23267 13507 23273
rect 2041 23239 2099 23245
rect 2041 23205 2053 23239
rect 2087 23236 2099 23239
rect 2590 23236 2596 23248
rect 2087 23208 2596 23236
rect 2087 23205 2099 23208
rect 2041 23199 2099 23205
rect 2590 23196 2596 23208
rect 2648 23196 2654 23248
rect 5442 23196 5448 23248
rect 5500 23196 5506 23248
rect 13464 23236 13492 23267
rect 13906 23264 13912 23276
rect 13964 23264 13970 23316
rect 16669 23307 16727 23313
rect 16669 23273 16681 23307
rect 16715 23304 16727 23307
rect 16758 23304 16764 23316
rect 16715 23276 16764 23304
rect 16715 23273 16727 23276
rect 16669 23267 16727 23273
rect 16758 23264 16764 23276
rect 16816 23264 16822 23316
rect 17218 23304 17224 23316
rect 17179 23276 17224 23304
rect 17218 23264 17224 23276
rect 17276 23264 17282 23316
rect 19061 23307 19119 23313
rect 19061 23273 19073 23307
rect 19107 23304 19119 23307
rect 19518 23304 19524 23316
rect 19107 23276 19524 23304
rect 19107 23273 19119 23276
rect 19061 23267 19119 23273
rect 19518 23264 19524 23276
rect 19576 23264 19582 23316
rect 20625 23307 20683 23313
rect 20625 23273 20637 23307
rect 20671 23304 20683 23307
rect 20714 23304 20720 23316
rect 20671 23276 20720 23304
rect 20671 23273 20683 23276
rect 20625 23267 20683 23273
rect 20714 23264 20720 23276
rect 20772 23264 20778 23316
rect 23201 23307 23259 23313
rect 23201 23273 23213 23307
rect 23247 23304 23259 23307
rect 23845 23307 23903 23313
rect 23845 23304 23857 23307
rect 23247 23276 23857 23304
rect 23247 23273 23259 23276
rect 23201 23267 23259 23273
rect 23845 23273 23857 23276
rect 23891 23304 23903 23307
rect 24210 23304 24216 23316
rect 23891 23276 24216 23304
rect 23891 23273 23903 23276
rect 23845 23267 23903 23273
rect 24210 23264 24216 23276
rect 24268 23264 24274 23316
rect 25130 23264 25136 23316
rect 25188 23304 25194 23316
rect 25314 23304 25320 23316
rect 25188 23276 25320 23304
rect 25188 23264 25194 23276
rect 25314 23264 25320 23276
rect 25372 23264 25378 23316
rect 16574 23236 16580 23248
rect 9692 23208 13492 23236
rect 15304 23208 16580 23236
rect 1765 23171 1823 23177
rect 1765 23137 1777 23171
rect 1811 23168 1823 23171
rect 2498 23168 2504 23180
rect 1811 23140 2504 23168
rect 1811 23137 1823 23140
rect 1765 23131 1823 23137
rect 2498 23128 2504 23140
rect 2556 23128 2562 23180
rect 3878 23128 3884 23180
rect 3936 23168 3942 23180
rect 4985 23171 5043 23177
rect 4985 23168 4997 23171
rect 3936 23140 4997 23168
rect 3936 23128 3942 23140
rect 4985 23137 4997 23140
rect 5031 23168 5043 23171
rect 5077 23171 5135 23177
rect 5077 23168 5089 23171
rect 5031 23140 5089 23168
rect 5031 23137 5043 23140
rect 4985 23131 5043 23137
rect 5077 23137 5089 23140
rect 5123 23168 5135 23171
rect 5166 23168 5172 23180
rect 5123 23140 5172 23168
rect 5123 23137 5135 23140
rect 5077 23131 5135 23137
rect 5166 23128 5172 23140
rect 5224 23128 5230 23180
rect 5344 23171 5402 23177
rect 5344 23137 5356 23171
rect 5390 23168 5402 23171
rect 5460 23168 5488 23196
rect 7926 23168 7932 23180
rect 5390 23140 7144 23168
rect 7887 23140 7932 23168
rect 5390 23137 5402 23140
rect 5344 23131 5402 23137
rect 3970 23060 3976 23112
rect 4028 23100 4034 23112
rect 4065 23103 4123 23109
rect 4065 23100 4077 23103
rect 4028 23072 4077 23100
rect 4028 23060 4034 23072
rect 4065 23069 4077 23072
rect 4111 23069 4123 23103
rect 4065 23063 4123 23069
rect 7116 23041 7144 23140
rect 7926 23128 7932 23140
rect 7984 23128 7990 23180
rect 9582 23128 9588 23180
rect 9640 23168 9646 23180
rect 9692 23177 9720 23208
rect 9677 23171 9735 23177
rect 9677 23168 9689 23171
rect 9640 23140 9689 23168
rect 9640 23128 9646 23140
rect 9677 23137 9689 23140
rect 9723 23137 9735 23171
rect 9677 23131 9735 23137
rect 11232 23171 11290 23177
rect 11232 23137 11244 23171
rect 11278 23168 11290 23171
rect 11606 23168 11612 23180
rect 11278 23140 11612 23168
rect 11278 23137 11290 23140
rect 11232 23131 11290 23137
rect 11606 23128 11612 23140
rect 11664 23128 11670 23180
rect 13262 23128 13268 23180
rect 13320 23168 13326 23180
rect 15304 23177 15332 23208
rect 16574 23196 16580 23208
rect 16632 23196 16638 23248
rect 17865 23239 17923 23245
rect 17865 23205 17877 23239
rect 17911 23236 17923 23239
rect 19242 23236 19248 23248
rect 17911 23208 19248 23236
rect 17911 23205 17923 23208
rect 17865 23199 17923 23205
rect 13817 23171 13875 23177
rect 13817 23168 13829 23171
rect 13320 23140 13829 23168
rect 13320 23128 13326 23140
rect 13817 23137 13829 23140
rect 13863 23137 13875 23171
rect 13817 23131 13875 23137
rect 15289 23171 15347 23177
rect 15289 23137 15301 23171
rect 15335 23137 15347 23171
rect 15289 23131 15347 23137
rect 15556 23171 15614 23177
rect 15556 23137 15568 23171
rect 15602 23168 15614 23171
rect 16022 23168 16028 23180
rect 15602 23140 16028 23168
rect 15602 23137 15614 23140
rect 15556 23131 15614 23137
rect 16022 23128 16028 23140
rect 16080 23168 16086 23180
rect 16390 23168 16396 23180
rect 16080 23140 16396 23168
rect 16080 23128 16086 23140
rect 16390 23128 16396 23140
rect 16448 23128 16454 23180
rect 17972 23177 18000 23208
rect 19242 23196 19248 23208
rect 19300 23196 19306 23248
rect 22094 23245 22100 23248
rect 22088 23199 22100 23245
rect 22152 23236 22158 23248
rect 22152 23208 22188 23236
rect 22094 23196 22100 23199
rect 22152 23196 22158 23208
rect 23658 23196 23664 23248
rect 23716 23236 23722 23248
rect 24673 23239 24731 23245
rect 24673 23236 24685 23239
rect 23716 23208 24685 23236
rect 23716 23196 23722 23208
rect 24673 23205 24685 23208
rect 24719 23236 24731 23239
rect 25866 23236 25872 23248
rect 24719 23208 25872 23236
rect 24719 23205 24731 23208
rect 24673 23199 24731 23205
rect 25866 23196 25872 23208
rect 25924 23196 25930 23248
rect 17957 23171 18015 23177
rect 17957 23137 17969 23171
rect 18003 23168 18015 23171
rect 19610 23168 19616 23180
rect 18003 23140 18037 23168
rect 19571 23140 19616 23168
rect 18003 23137 18015 23140
rect 17957 23131 18015 23137
rect 19610 23128 19616 23140
rect 19668 23128 19674 23180
rect 20070 23128 20076 23180
rect 20128 23168 20134 23180
rect 24026 23168 24032 23180
rect 20128 23140 24032 23168
rect 20128 23128 20134 23140
rect 24026 23128 24032 23140
rect 24084 23128 24090 23180
rect 24762 23168 24768 23180
rect 24723 23140 24768 23168
rect 24762 23128 24768 23140
rect 24820 23128 24826 23180
rect 7466 23060 7472 23112
rect 7524 23060 7530 23112
rect 8113 23103 8171 23109
rect 8113 23069 8125 23103
rect 8159 23069 8171 23103
rect 9030 23100 9036 23112
rect 8991 23072 9036 23100
rect 8113 23063 8171 23069
rect 7101 23035 7159 23041
rect 7101 23001 7113 23035
rect 7147 23032 7159 23035
rect 7377 23035 7435 23041
rect 7377 23032 7389 23035
rect 7147 23004 7389 23032
rect 7147 23001 7159 23004
rect 7101 22995 7159 23001
rect 7377 23001 7389 23004
rect 7423 23032 7435 23035
rect 7484 23032 7512 23060
rect 8128 23032 8156 23063
rect 9030 23060 9036 23072
rect 9088 23060 9094 23112
rect 9953 23103 10011 23109
rect 9953 23069 9965 23103
rect 9999 23100 10011 23103
rect 10134 23100 10140 23112
rect 9999 23072 10140 23100
rect 9999 23069 10011 23072
rect 9953 23063 10011 23069
rect 10134 23060 10140 23072
rect 10192 23060 10198 23112
rect 10965 23103 11023 23109
rect 10965 23069 10977 23103
rect 11011 23069 11023 23103
rect 13998 23100 14004 23112
rect 13959 23072 14004 23100
rect 10965 23063 11023 23069
rect 10980 23032 11008 23063
rect 13998 23060 14004 23072
rect 14056 23060 14062 23112
rect 18233 23103 18291 23109
rect 18233 23069 18245 23103
rect 18279 23100 18291 23103
rect 18966 23100 18972 23112
rect 18279 23072 18972 23100
rect 18279 23069 18291 23072
rect 18233 23063 18291 23069
rect 18966 23060 18972 23072
rect 19024 23060 19030 23112
rect 19702 23100 19708 23112
rect 19663 23072 19708 23100
rect 19702 23060 19708 23072
rect 19760 23060 19766 23112
rect 19889 23103 19947 23109
rect 19889 23069 19901 23103
rect 19935 23100 19947 23103
rect 20530 23100 20536 23112
rect 19935 23072 20536 23100
rect 19935 23069 19947 23072
rect 19889 23063 19947 23069
rect 20530 23060 20536 23072
rect 20588 23060 20594 23112
rect 20806 23060 20812 23112
rect 20864 23100 20870 23112
rect 21453 23103 21511 23109
rect 21453 23100 21465 23103
rect 20864 23072 21465 23100
rect 20864 23060 20870 23072
rect 21453 23069 21465 23072
rect 21499 23069 21511 23103
rect 21453 23063 21511 23069
rect 21634 23060 21640 23112
rect 21692 23100 21698 23112
rect 21821 23103 21879 23109
rect 21821 23100 21833 23103
rect 21692 23072 21833 23100
rect 21692 23060 21698 23072
rect 21821 23069 21833 23072
rect 21867 23069 21879 23103
rect 24854 23100 24860 23112
rect 24815 23072 24860 23100
rect 21821 23063 21879 23069
rect 24854 23060 24860 23072
rect 24912 23060 24918 23112
rect 14461 23035 14519 23041
rect 14461 23032 14473 23035
rect 7423 23004 8156 23032
rect 9416 23004 11008 23032
rect 7423 23001 7435 23004
rect 7377 22995 7435 23001
rect 1670 22964 1676 22976
rect 1631 22936 1676 22964
rect 1670 22924 1676 22936
rect 1728 22924 1734 22976
rect 3694 22964 3700 22976
rect 3655 22936 3700 22964
rect 3694 22924 3700 22936
rect 3752 22924 3758 22976
rect 4617 22967 4675 22973
rect 4617 22933 4629 22967
rect 4663 22964 4675 22967
rect 4890 22964 4896 22976
rect 4663 22936 4896 22964
rect 4663 22933 4675 22936
rect 4617 22927 4675 22933
rect 4890 22924 4896 22936
rect 4948 22924 4954 22976
rect 7466 22924 7472 22976
rect 7524 22964 7530 22976
rect 7561 22967 7619 22973
rect 7561 22964 7573 22967
rect 7524 22936 7573 22964
rect 7524 22924 7530 22936
rect 7561 22933 7573 22936
rect 7607 22933 7619 22967
rect 7561 22927 7619 22933
rect 9306 22924 9312 22976
rect 9364 22964 9370 22976
rect 9416 22973 9444 23004
rect 9401 22967 9459 22973
rect 9401 22964 9413 22967
rect 9364 22936 9413 22964
rect 9364 22924 9370 22936
rect 9401 22933 9413 22936
rect 9447 22933 9459 22967
rect 9401 22927 9459 22933
rect 9950 22924 9956 22976
rect 10008 22964 10014 22976
rect 10410 22964 10416 22976
rect 10008 22936 10416 22964
rect 10008 22924 10014 22936
rect 10410 22924 10416 22936
rect 10468 22924 10474 22976
rect 10778 22964 10784 22976
rect 10739 22936 10784 22964
rect 10778 22924 10784 22936
rect 10836 22924 10842 22976
rect 10980 22964 11008 23004
rect 12912 23004 14473 23032
rect 12434 22964 12440 22976
rect 10980 22936 12440 22964
rect 12434 22924 12440 22936
rect 12492 22964 12498 22976
rect 12912 22973 12940 23004
rect 14461 23001 14473 23004
rect 14507 23032 14519 23035
rect 14550 23032 14556 23044
rect 14507 23004 14556 23032
rect 14507 23001 14519 23004
rect 14461 22995 14519 23001
rect 14550 22992 14556 23004
rect 14608 22992 14614 23044
rect 14734 22992 14740 23044
rect 14792 22992 14798 23044
rect 19150 22992 19156 23044
rect 19208 23032 19214 23044
rect 19245 23035 19303 23041
rect 19245 23032 19257 23035
rect 19208 23004 19257 23032
rect 19208 22992 19214 23004
rect 19245 23001 19257 23004
rect 19291 23001 19303 23035
rect 19245 22995 19303 23001
rect 23566 22992 23572 23044
rect 23624 23032 23630 23044
rect 25317 23035 25375 23041
rect 25317 23032 25329 23035
rect 23624 23004 25329 23032
rect 23624 22992 23630 23004
rect 25317 23001 25329 23004
rect 25363 23001 25375 23035
rect 25317 22995 25375 23001
rect 12897 22967 12955 22973
rect 12897 22964 12909 22967
rect 12492 22936 12909 22964
rect 12492 22924 12498 22936
rect 12897 22933 12909 22936
rect 12943 22933 12955 22967
rect 13262 22964 13268 22976
rect 13223 22936 13268 22964
rect 12897 22927 12955 22933
rect 13262 22924 13268 22936
rect 13320 22924 13326 22976
rect 14752 22964 14780 22992
rect 15013 22967 15071 22973
rect 15013 22964 15025 22967
rect 14752 22936 15025 22964
rect 15013 22933 15025 22936
rect 15059 22964 15071 22967
rect 15286 22964 15292 22976
rect 15059 22936 15292 22964
rect 15059 22933 15071 22936
rect 15013 22927 15071 22933
rect 15286 22924 15292 22936
rect 15344 22924 15350 22976
rect 20346 22924 20352 22976
rect 20404 22964 20410 22976
rect 21085 22967 21143 22973
rect 21085 22964 21097 22967
rect 20404 22936 21097 22964
rect 20404 22924 20410 22936
rect 21085 22933 21097 22936
rect 21131 22964 21143 22967
rect 21450 22964 21456 22976
rect 21131 22936 21456 22964
rect 21131 22933 21143 22936
rect 21085 22927 21143 22933
rect 21450 22924 21456 22936
rect 21508 22924 21514 22976
rect 23382 22924 23388 22976
rect 23440 22964 23446 22976
rect 24305 22967 24363 22973
rect 24305 22964 24317 22967
rect 23440 22936 24317 22964
rect 23440 22924 23446 22936
rect 24305 22933 24317 22936
rect 24351 22933 24363 22967
rect 24305 22927 24363 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 4709 22763 4767 22769
rect 4709 22729 4721 22763
rect 4755 22760 4767 22763
rect 5442 22760 5448 22772
rect 4755 22732 5448 22760
rect 4755 22729 4767 22732
rect 4709 22723 4767 22729
rect 5442 22720 5448 22732
rect 5500 22720 5506 22772
rect 9677 22763 9735 22769
rect 9677 22729 9689 22763
rect 9723 22760 9735 22763
rect 10962 22760 10968 22772
rect 9723 22732 10968 22760
rect 9723 22729 9735 22732
rect 9677 22723 9735 22729
rect 10962 22720 10968 22732
rect 11020 22720 11026 22772
rect 13906 22720 13912 22772
rect 13964 22760 13970 22772
rect 14369 22763 14427 22769
rect 14369 22760 14381 22763
rect 13964 22732 14381 22760
rect 13964 22720 13970 22732
rect 14369 22729 14381 22732
rect 14415 22729 14427 22763
rect 14734 22760 14740 22772
rect 14695 22732 14740 22760
rect 14369 22723 14427 22729
rect 14734 22720 14740 22732
rect 14792 22760 14798 22772
rect 16393 22763 16451 22769
rect 14792 22732 15424 22760
rect 14792 22720 14798 22732
rect 2498 22692 2504 22704
rect 2459 22664 2504 22692
rect 2498 22652 2504 22664
rect 2556 22692 2562 22704
rect 5169 22695 5227 22701
rect 5169 22692 5181 22695
rect 2556 22664 5181 22692
rect 2556 22652 2562 22664
rect 5169 22661 5181 22664
rect 5215 22661 5227 22695
rect 5169 22655 5227 22661
rect 9585 22695 9643 22701
rect 9585 22661 9597 22695
rect 9631 22692 9643 22695
rect 9950 22692 9956 22704
rect 9631 22664 9956 22692
rect 9631 22661 9643 22664
rect 9585 22655 9643 22661
rect 9950 22652 9956 22664
rect 10008 22652 10014 22704
rect 11422 22692 11428 22704
rect 11383 22664 11428 22692
rect 11422 22652 11428 22664
rect 11480 22652 11486 22704
rect 1673 22627 1731 22633
rect 1673 22593 1685 22627
rect 1719 22624 1731 22627
rect 2866 22624 2872 22636
rect 1719 22596 2872 22624
rect 1719 22593 1731 22596
rect 1673 22587 1731 22593
rect 2866 22584 2872 22596
rect 2924 22584 2930 22636
rect 4154 22584 4160 22636
rect 4212 22624 4218 22636
rect 15396 22633 15424 22732
rect 16393 22729 16405 22763
rect 16439 22760 16451 22763
rect 16574 22760 16580 22772
rect 16439 22732 16580 22760
rect 16439 22729 16451 22732
rect 16393 22723 16451 22729
rect 16574 22720 16580 22732
rect 16632 22720 16638 22772
rect 17497 22763 17555 22769
rect 17497 22729 17509 22763
rect 17543 22760 17555 22763
rect 17770 22760 17776 22772
rect 17543 22732 17776 22760
rect 17543 22729 17555 22732
rect 17497 22723 17555 22729
rect 5077 22627 5135 22633
rect 4212 22596 4257 22624
rect 4212 22584 4218 22596
rect 5077 22593 5089 22627
rect 5123 22624 5135 22627
rect 5813 22627 5871 22633
rect 5813 22624 5825 22627
rect 5123 22596 5825 22624
rect 5123 22593 5135 22596
rect 5077 22587 5135 22593
rect 5813 22593 5825 22596
rect 5859 22624 5871 22627
rect 10321 22627 10379 22633
rect 5859 22596 6684 22624
rect 5859 22593 5871 22596
rect 5813 22587 5871 22593
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22556 1455 22559
rect 2038 22556 2044 22568
rect 1443 22528 2044 22556
rect 1443 22525 1455 22528
rect 1397 22519 1455 22525
rect 2038 22516 2044 22528
rect 2096 22556 2102 22568
rect 2133 22559 2191 22565
rect 2133 22556 2145 22559
rect 2096 22528 2145 22556
rect 2096 22516 2102 22528
rect 2133 22525 2145 22528
rect 2179 22525 2191 22559
rect 2133 22519 2191 22525
rect 3513 22559 3571 22565
rect 3513 22525 3525 22559
rect 3559 22556 3571 22559
rect 3970 22556 3976 22568
rect 3559 22528 3976 22556
rect 3559 22525 3571 22528
rect 3513 22519 3571 22525
rect 3970 22516 3976 22528
rect 4028 22516 4034 22568
rect 5537 22491 5595 22497
rect 5537 22488 5549 22491
rect 3620 22460 5549 22488
rect 3142 22420 3148 22432
rect 3103 22392 3148 22420
rect 3142 22380 3148 22392
rect 3200 22380 3206 22432
rect 3620 22429 3648 22460
rect 5537 22457 5549 22460
rect 5583 22488 5595 22491
rect 5994 22488 6000 22500
rect 5583 22460 6000 22488
rect 5583 22457 5595 22460
rect 5537 22451 5595 22457
rect 5994 22448 6000 22460
rect 6052 22448 6058 22500
rect 6656 22497 6684 22596
rect 10321 22593 10333 22627
rect 10367 22624 10379 22627
rect 12253 22627 12311 22633
rect 10367 22596 10824 22624
rect 10367 22593 10379 22596
rect 10321 22587 10379 22593
rect 6730 22516 6736 22568
rect 6788 22556 6794 22568
rect 6917 22559 6975 22565
rect 6917 22556 6929 22559
rect 6788 22528 6929 22556
rect 6788 22516 6794 22528
rect 6917 22525 6929 22528
rect 6963 22556 6975 22559
rect 7650 22556 7656 22568
rect 6963 22528 7656 22556
rect 6963 22525 6975 22528
rect 6917 22519 6975 22525
rect 7650 22516 7656 22528
rect 7708 22516 7714 22568
rect 9122 22516 9128 22568
rect 9180 22556 9186 22568
rect 10137 22559 10195 22565
rect 10137 22556 10149 22559
rect 9180 22528 10149 22556
rect 9180 22516 9186 22528
rect 10137 22525 10149 22528
rect 10183 22525 10195 22559
rect 10137 22519 10195 22525
rect 6641 22491 6699 22497
rect 6641 22457 6653 22491
rect 6687 22488 6699 22491
rect 7098 22488 7104 22500
rect 6687 22460 7104 22488
rect 6687 22457 6699 22460
rect 6641 22451 6699 22457
rect 7098 22448 7104 22460
rect 7156 22497 7162 22500
rect 7156 22491 7220 22497
rect 7156 22457 7174 22491
rect 7208 22457 7220 22491
rect 10410 22488 10416 22500
rect 7156 22451 7220 22457
rect 8312 22460 10416 22488
rect 7156 22448 7162 22451
rect 3605 22423 3663 22429
rect 3605 22389 3617 22423
rect 3651 22389 3663 22423
rect 3605 22383 3663 22389
rect 3694 22380 3700 22432
rect 3752 22420 3758 22432
rect 4065 22423 4123 22429
rect 4065 22420 4077 22423
rect 3752 22392 4077 22420
rect 3752 22380 3758 22392
rect 4065 22389 4077 22392
rect 4111 22420 4123 22423
rect 5074 22420 5080 22432
rect 4111 22392 5080 22420
rect 4111 22389 4123 22392
rect 4065 22383 4123 22389
rect 5074 22380 5080 22392
rect 5132 22380 5138 22432
rect 5629 22423 5687 22429
rect 5629 22389 5641 22423
rect 5675 22420 5687 22423
rect 6181 22423 6239 22429
rect 6181 22420 6193 22423
rect 5675 22392 6193 22420
rect 5675 22389 5687 22392
rect 5629 22383 5687 22389
rect 6181 22389 6193 22392
rect 6227 22420 6239 22423
rect 6454 22420 6460 22432
rect 6227 22392 6460 22420
rect 6227 22389 6239 22392
rect 6181 22383 6239 22389
rect 6454 22380 6460 22392
rect 6512 22380 6518 22432
rect 8202 22380 8208 22432
rect 8260 22420 8266 22432
rect 8312 22429 8340 22460
rect 10410 22448 10416 22460
rect 10468 22448 10474 22500
rect 8297 22423 8355 22429
rect 8297 22420 8309 22423
rect 8260 22392 8309 22420
rect 8260 22380 8266 22392
rect 8297 22389 8309 22392
rect 8343 22389 8355 22423
rect 9122 22420 9128 22432
rect 9083 22392 9128 22420
rect 8297 22383 8355 22389
rect 9122 22380 9128 22392
rect 9180 22380 9186 22432
rect 9950 22380 9956 22432
rect 10008 22420 10014 22432
rect 10796 22429 10824 22596
rect 12253 22593 12265 22627
rect 12299 22624 12311 22627
rect 15381 22627 15439 22633
rect 12299 22596 12572 22624
rect 12299 22593 12311 22596
rect 12253 22587 12311 22593
rect 11241 22559 11299 22565
rect 11241 22525 11253 22559
rect 11287 22556 11299 22559
rect 12434 22556 12440 22568
rect 11287 22528 11928 22556
rect 12395 22528 12440 22556
rect 11287 22525 11299 22528
rect 11241 22519 11299 22525
rect 11900 22432 11928 22528
rect 12434 22516 12440 22528
rect 12492 22516 12498 22568
rect 12544 22556 12572 22596
rect 15381 22593 15393 22627
rect 15427 22593 15439 22627
rect 15381 22587 15439 22593
rect 15473 22627 15531 22633
rect 15473 22593 15485 22627
rect 15519 22593 15531 22627
rect 16850 22624 16856 22636
rect 16811 22596 16856 22624
rect 15473 22587 15531 22593
rect 12704 22559 12762 22565
rect 12704 22556 12716 22559
rect 12544 22528 12716 22556
rect 12704 22525 12716 22528
rect 12750 22556 12762 22559
rect 13998 22556 14004 22568
rect 12750 22528 14004 22556
rect 12750 22525 12762 22528
rect 12704 22519 12762 22525
rect 13998 22516 14004 22528
rect 14056 22516 14062 22568
rect 14090 22516 14096 22568
rect 14148 22556 14154 22568
rect 15286 22556 15292 22568
rect 14148 22528 15292 22556
rect 14148 22516 14154 22528
rect 15286 22516 15292 22528
rect 15344 22556 15350 22568
rect 15488 22556 15516 22587
rect 16850 22584 16856 22596
rect 16908 22584 16914 22636
rect 15344 22528 15516 22556
rect 16669 22559 16727 22565
rect 15344 22516 15350 22528
rect 16669 22525 16681 22559
rect 16715 22556 16727 22559
rect 17512 22556 17540 22723
rect 17770 22720 17776 22732
rect 17828 22720 17834 22772
rect 19150 22760 19156 22772
rect 19111 22732 19156 22760
rect 19150 22720 19156 22732
rect 19208 22760 19214 22772
rect 19610 22760 19616 22772
rect 19208 22732 19616 22760
rect 19208 22720 19214 22732
rect 19610 22720 19616 22732
rect 19668 22760 19674 22772
rect 19978 22760 19984 22772
rect 19668 22732 19984 22760
rect 19668 22720 19674 22732
rect 19978 22720 19984 22732
rect 20036 22720 20042 22772
rect 20530 22720 20536 22772
rect 20588 22760 20594 22772
rect 20717 22763 20775 22769
rect 20717 22760 20729 22763
rect 20588 22732 20729 22760
rect 20588 22720 20594 22732
rect 20717 22729 20729 22732
rect 20763 22729 20775 22763
rect 22002 22760 22008 22772
rect 21963 22732 22008 22760
rect 20717 22723 20775 22729
rect 22002 22720 22008 22732
rect 22060 22720 22066 22772
rect 22094 22720 22100 22772
rect 22152 22760 22158 22772
rect 23017 22763 23075 22769
rect 23017 22760 23029 22763
rect 22152 22732 23029 22760
rect 22152 22720 22158 22732
rect 23017 22729 23029 22732
rect 23063 22729 23075 22763
rect 23017 22723 23075 22729
rect 24762 22720 24768 22772
rect 24820 22760 24826 22772
rect 25593 22763 25651 22769
rect 25593 22760 25605 22763
rect 24820 22732 25605 22760
rect 24820 22720 24826 22732
rect 25593 22729 25605 22732
rect 25639 22729 25651 22763
rect 25593 22723 25651 22729
rect 25866 22720 25872 22772
rect 25924 22760 25930 22772
rect 25961 22763 26019 22769
rect 25961 22760 25973 22763
rect 25924 22732 25973 22760
rect 25924 22720 25930 22732
rect 25961 22729 25973 22732
rect 26007 22729 26019 22763
rect 25961 22723 26019 22729
rect 18322 22584 18328 22636
rect 18380 22624 18386 22636
rect 19150 22624 19156 22636
rect 18380 22596 19156 22624
rect 18380 22584 18386 22596
rect 19150 22584 19156 22596
rect 19208 22584 19214 22636
rect 22649 22627 22707 22633
rect 22649 22593 22661 22627
rect 22695 22624 22707 22627
rect 23014 22624 23020 22636
rect 22695 22596 23020 22624
rect 22695 22593 22707 22596
rect 22649 22587 22707 22593
rect 23014 22584 23020 22596
rect 23072 22624 23078 22636
rect 23072 22596 23796 22624
rect 23072 22584 23078 22596
rect 16715 22528 17540 22556
rect 17865 22559 17923 22565
rect 16715 22525 16727 22528
rect 16669 22519 16727 22525
rect 17865 22525 17877 22559
rect 17911 22556 17923 22559
rect 18046 22556 18052 22568
rect 17911 22528 18052 22556
rect 17911 22525 17923 22528
rect 17865 22519 17923 22525
rect 18046 22516 18052 22528
rect 18104 22516 18110 22568
rect 18690 22516 18696 22568
rect 18748 22556 18754 22568
rect 19334 22556 19340 22568
rect 18748 22528 19340 22556
rect 18748 22516 18754 22528
rect 19334 22516 19340 22528
rect 19392 22516 19398 22568
rect 21450 22516 21456 22568
rect 21508 22556 21514 22568
rect 21729 22559 21787 22565
rect 21729 22556 21741 22559
rect 21508 22528 21741 22556
rect 21508 22516 21514 22528
rect 21729 22525 21741 22528
rect 21775 22556 21787 22559
rect 21821 22559 21879 22565
rect 21821 22556 21833 22559
rect 21775 22528 21833 22556
rect 21775 22525 21787 22528
rect 21729 22519 21787 22525
rect 21821 22525 21833 22528
rect 21867 22525 21879 22559
rect 21821 22519 21879 22525
rect 23566 22516 23572 22568
rect 23624 22556 23630 22568
rect 23661 22559 23719 22565
rect 23661 22556 23673 22559
rect 23624 22528 23673 22556
rect 23624 22516 23630 22528
rect 23661 22525 23673 22528
rect 23707 22525 23719 22559
rect 23768 22556 23796 22596
rect 23928 22559 23986 22565
rect 23928 22556 23940 22559
rect 23768 22528 23940 22556
rect 23661 22519 23719 22525
rect 23928 22525 23940 22528
rect 23974 22556 23986 22559
rect 24210 22556 24216 22568
rect 23974 22528 24216 22556
rect 23974 22525 23986 22528
rect 23928 22519 23986 22525
rect 15562 22448 15568 22500
rect 15620 22488 15626 22500
rect 15746 22488 15752 22500
rect 15620 22460 15752 22488
rect 15620 22448 15626 22460
rect 15746 22448 15752 22460
rect 15804 22448 15810 22500
rect 18322 22488 18328 22500
rect 18283 22460 18328 22488
rect 18322 22448 18328 22460
rect 18380 22448 18386 22500
rect 19518 22448 19524 22500
rect 19576 22497 19582 22500
rect 19576 22491 19640 22497
rect 19576 22457 19594 22491
rect 19628 22457 19640 22491
rect 19576 22451 19640 22457
rect 19576 22448 19582 22451
rect 19702 22448 19708 22500
rect 19760 22448 19766 22500
rect 22465 22491 22523 22497
rect 22465 22488 22477 22491
rect 21468 22460 22477 22488
rect 10045 22423 10103 22429
rect 10045 22420 10057 22423
rect 10008 22392 10057 22420
rect 10008 22380 10014 22392
rect 10045 22389 10057 22392
rect 10091 22389 10103 22423
rect 10045 22383 10103 22389
rect 10781 22423 10839 22429
rect 10781 22389 10793 22423
rect 10827 22420 10839 22423
rect 11149 22423 11207 22429
rect 11149 22420 11161 22423
rect 10827 22392 11161 22420
rect 10827 22389 10839 22392
rect 10781 22383 10839 22389
rect 11149 22389 11161 22392
rect 11195 22420 11207 22423
rect 11606 22420 11612 22432
rect 11195 22392 11612 22420
rect 11195 22389 11207 22392
rect 11149 22383 11207 22389
rect 11606 22380 11612 22392
rect 11664 22380 11670 22432
rect 11882 22420 11888 22432
rect 11843 22392 11888 22420
rect 11882 22380 11888 22392
rect 11940 22380 11946 22432
rect 13817 22423 13875 22429
rect 13817 22389 13829 22423
rect 13863 22420 13875 22423
rect 13906 22420 13912 22432
rect 13863 22392 13912 22420
rect 13863 22389 13875 22392
rect 13817 22383 13875 22389
rect 13906 22380 13912 22392
rect 13964 22380 13970 22432
rect 14918 22420 14924 22432
rect 14879 22392 14924 22420
rect 14918 22380 14924 22392
rect 14976 22380 14982 22432
rect 15102 22380 15108 22432
rect 15160 22420 15166 22432
rect 15289 22423 15347 22429
rect 15289 22420 15301 22423
rect 15160 22392 15301 22420
rect 15160 22380 15166 22392
rect 15289 22389 15301 22392
rect 15335 22389 15347 22423
rect 16022 22420 16028 22432
rect 15983 22392 16028 22420
rect 15289 22383 15347 22389
rect 16022 22380 16028 22392
rect 16080 22380 16086 22432
rect 18690 22380 18696 22432
rect 18748 22420 18754 22432
rect 18785 22423 18843 22429
rect 18785 22420 18797 22423
rect 18748 22392 18797 22420
rect 18748 22380 18754 22392
rect 18785 22389 18797 22392
rect 18831 22420 18843 22423
rect 19720 22420 19748 22448
rect 18831 22392 19748 22420
rect 18831 22389 18843 22392
rect 18785 22383 18843 22389
rect 20990 22380 20996 22432
rect 21048 22420 21054 22432
rect 21468 22429 21496 22460
rect 22465 22457 22477 22460
rect 22511 22457 22523 22491
rect 23676 22488 23704 22519
rect 24210 22516 24216 22528
rect 24268 22516 24274 22568
rect 23750 22488 23756 22500
rect 23676 22460 23756 22488
rect 22465 22451 22523 22457
rect 23750 22448 23756 22460
rect 23808 22448 23814 22500
rect 21453 22423 21511 22429
rect 21453 22420 21465 22423
rect 21048 22392 21465 22420
rect 21048 22380 21054 22392
rect 21453 22389 21465 22392
rect 21499 22389 21511 22423
rect 21453 22383 21511 22389
rect 21729 22423 21787 22429
rect 21729 22389 21741 22423
rect 21775 22420 21787 22423
rect 22373 22423 22431 22429
rect 22373 22420 22385 22423
rect 21775 22392 22385 22420
rect 21775 22389 21787 22392
rect 21729 22383 21787 22389
rect 22373 22389 22385 22392
rect 22419 22389 22431 22423
rect 23474 22420 23480 22432
rect 23435 22392 23480 22420
rect 22373 22383 22431 22389
rect 23474 22380 23480 22392
rect 23532 22380 23538 22432
rect 24762 22380 24768 22432
rect 24820 22420 24826 22432
rect 25041 22423 25099 22429
rect 25041 22420 25053 22423
rect 24820 22392 25053 22420
rect 24820 22380 24826 22392
rect 25041 22389 25053 22392
rect 25087 22389 25099 22423
rect 26326 22420 26332 22432
rect 26287 22392 26332 22420
rect 25041 22383 25099 22389
rect 26326 22380 26332 22392
rect 26384 22380 26390 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 2774 22176 2780 22228
rect 2832 22216 2838 22228
rect 2958 22216 2964 22228
rect 2832 22188 2964 22216
rect 2832 22176 2838 22188
rect 2958 22176 2964 22188
rect 3016 22176 3022 22228
rect 3697 22219 3755 22225
rect 3697 22185 3709 22219
rect 3743 22216 3755 22219
rect 4154 22216 4160 22228
rect 3743 22188 4160 22216
rect 3743 22185 3755 22188
rect 3697 22179 3755 22185
rect 4154 22176 4160 22188
rect 4212 22176 4218 22228
rect 5442 22216 5448 22228
rect 5403 22188 5448 22216
rect 5442 22176 5448 22188
rect 5500 22176 5506 22228
rect 5994 22216 6000 22228
rect 5955 22188 6000 22216
rect 5994 22176 6000 22188
rect 6052 22176 6058 22228
rect 6454 22176 6460 22228
rect 6512 22216 6518 22228
rect 6549 22219 6607 22225
rect 6549 22216 6561 22219
rect 6512 22188 6561 22216
rect 6512 22176 6518 22188
rect 6549 22185 6561 22188
rect 6595 22185 6607 22219
rect 6914 22216 6920 22228
rect 6875 22188 6920 22216
rect 6549 22179 6607 22185
rect 6914 22176 6920 22188
rect 6972 22176 6978 22228
rect 7009 22219 7067 22225
rect 7009 22185 7021 22219
rect 7055 22216 7067 22219
rect 7098 22216 7104 22228
rect 7055 22188 7104 22216
rect 7055 22185 7067 22188
rect 7009 22179 7067 22185
rect 7098 22176 7104 22188
rect 7156 22216 7162 22228
rect 7466 22216 7472 22228
rect 7156 22188 7472 22216
rect 7156 22176 7162 22188
rect 7466 22176 7472 22188
rect 7524 22176 7530 22228
rect 7926 22216 7932 22228
rect 7887 22188 7932 22216
rect 7926 22176 7932 22188
rect 7984 22176 7990 22228
rect 9674 22176 9680 22228
rect 9732 22216 9738 22228
rect 10045 22219 10103 22225
rect 10045 22216 10057 22219
rect 9732 22188 10057 22216
rect 9732 22176 9738 22188
rect 10045 22185 10057 22188
rect 10091 22185 10103 22219
rect 10045 22179 10103 22185
rect 12345 22219 12403 22225
rect 12345 22185 12357 22219
rect 12391 22216 12403 22219
rect 13262 22216 13268 22228
rect 12391 22188 13268 22216
rect 12391 22185 12403 22188
rect 12345 22179 12403 22185
rect 13262 22176 13268 22188
rect 13320 22176 13326 22228
rect 13541 22219 13599 22225
rect 13541 22185 13553 22219
rect 13587 22216 13599 22219
rect 13998 22216 14004 22228
rect 13587 22188 14004 22216
rect 13587 22185 13599 22188
rect 13541 22179 13599 22185
rect 13998 22176 14004 22188
rect 14056 22176 14062 22228
rect 16022 22176 16028 22228
rect 16080 22216 16086 22228
rect 17129 22219 17187 22225
rect 17129 22216 17141 22219
rect 16080 22188 17141 22216
rect 16080 22176 16086 22188
rect 17129 22185 17141 22188
rect 17175 22185 17187 22219
rect 17129 22179 17187 22185
rect 19429 22219 19487 22225
rect 19429 22185 19441 22219
rect 19475 22216 19487 22219
rect 19518 22216 19524 22228
rect 19475 22188 19524 22216
rect 19475 22185 19487 22188
rect 19429 22179 19487 22185
rect 19518 22176 19524 22188
rect 19576 22176 19582 22228
rect 19797 22219 19855 22225
rect 19797 22185 19809 22219
rect 19843 22216 19855 22219
rect 20070 22216 20076 22228
rect 19843 22188 20076 22216
rect 19843 22185 19855 22188
rect 19797 22179 19855 22185
rect 20070 22176 20076 22188
rect 20128 22176 20134 22228
rect 20530 22216 20536 22228
rect 20491 22188 20536 22216
rect 20530 22176 20536 22188
rect 20588 22216 20594 22228
rect 20714 22216 20720 22228
rect 20588 22188 20720 22216
rect 20588 22176 20594 22188
rect 20714 22176 20720 22188
rect 20772 22176 20778 22228
rect 22094 22176 22100 22228
rect 22152 22216 22158 22228
rect 22281 22219 22339 22225
rect 22281 22216 22293 22219
rect 22152 22188 22293 22216
rect 22152 22176 22158 22188
rect 22281 22185 22293 22188
rect 22327 22185 22339 22219
rect 22281 22179 22339 22185
rect 22925 22219 22983 22225
rect 22925 22185 22937 22219
rect 22971 22216 22983 22219
rect 23014 22216 23020 22228
rect 22971 22188 23020 22216
rect 22971 22185 22983 22188
rect 22925 22179 22983 22185
rect 23014 22176 23020 22188
rect 23072 22176 23078 22228
rect 1397 22151 1455 22157
rect 1397 22117 1409 22151
rect 1443 22148 1455 22151
rect 2222 22148 2228 22160
rect 1443 22120 2228 22148
rect 1443 22117 1455 22120
rect 1397 22111 1455 22117
rect 2222 22108 2228 22120
rect 2280 22108 2286 22160
rect 2866 22108 2872 22160
rect 2924 22148 2930 22160
rect 2924 22120 2969 22148
rect 2924 22108 2930 22120
rect 3602 22108 3608 22160
rect 3660 22148 3666 22160
rect 3878 22148 3884 22160
rect 3660 22120 3884 22148
rect 3660 22108 3666 22120
rect 3878 22108 3884 22120
rect 3936 22108 3942 22160
rect 3970 22108 3976 22160
rect 4028 22148 4034 22160
rect 4172 22148 4200 22176
rect 5534 22148 5540 22160
rect 4028 22120 4108 22148
rect 4172 22120 5540 22148
rect 4028 22108 4034 22120
rect 1949 22083 2007 22089
rect 1949 22049 1961 22083
rect 1995 22080 2007 22083
rect 2314 22080 2320 22092
rect 1995 22052 2320 22080
rect 1995 22049 2007 22052
rect 1949 22043 2007 22049
rect 2314 22040 2320 22052
rect 2372 22080 2378 22092
rect 3142 22080 3148 22092
rect 2372 22052 3148 22080
rect 2372 22040 2378 22052
rect 3142 22040 3148 22052
rect 3200 22080 3206 22092
rect 4080 22089 4108 22120
rect 5534 22108 5540 22120
rect 5592 22108 5598 22160
rect 7653 22151 7711 22157
rect 7653 22117 7665 22151
rect 7699 22148 7711 22151
rect 8018 22148 8024 22160
rect 7699 22120 8024 22148
rect 7699 22117 7711 22120
rect 7653 22111 7711 22117
rect 8018 22108 8024 22120
rect 8076 22108 8082 22160
rect 12713 22151 12771 22157
rect 12713 22148 12725 22151
rect 12452 22120 12725 22148
rect 4338 22089 4344 22092
rect 4065 22083 4123 22089
rect 4065 22080 4077 22083
rect 3200 22052 4077 22080
rect 3200 22040 3206 22052
rect 4065 22049 4077 22052
rect 4111 22080 4123 22083
rect 4332 22080 4344 22089
rect 4111 22052 4145 22080
rect 4299 22052 4344 22080
rect 4111 22049 4123 22052
rect 4065 22043 4123 22049
rect 4332 22043 4344 22052
rect 4338 22040 4344 22043
rect 4396 22040 4402 22092
rect 8110 22080 8116 22092
rect 8071 22052 8116 22080
rect 8110 22040 8116 22052
rect 8168 22040 8174 22092
rect 9493 22083 9551 22089
rect 9493 22049 9505 22083
rect 9539 22080 9551 22083
rect 9582 22080 9588 22092
rect 9539 22052 9588 22080
rect 9539 22049 9551 22052
rect 9493 22043 9551 22049
rect 9582 22040 9588 22052
rect 9640 22040 9646 22092
rect 9950 22040 9956 22092
rect 10008 22080 10014 22092
rect 11238 22080 11244 22092
rect 10008 22052 10272 22080
rect 11199 22052 11244 22080
rect 10008 22040 10014 22052
rect 3053 22015 3111 22021
rect 3053 21981 3065 22015
rect 3099 22012 3111 22015
rect 3234 22012 3240 22024
rect 3099 21984 3240 22012
rect 3099 21981 3111 21984
rect 3053 21975 3111 21981
rect 3234 21972 3240 21984
rect 3292 22012 3298 22024
rect 3786 22012 3792 22024
rect 3292 21984 3792 22012
rect 3292 21972 3298 21984
rect 3786 21972 3792 21984
rect 3844 21972 3850 22024
rect 6546 21972 6552 22024
rect 6604 22012 6610 22024
rect 7101 22015 7159 22021
rect 7101 22012 7113 22015
rect 6604 21984 7113 22012
rect 6604 21972 6610 21984
rect 7101 21981 7113 21984
rect 7147 21981 7159 22015
rect 7101 21975 7159 21981
rect 10042 21972 10048 22024
rect 10100 22012 10106 22024
rect 10244 22021 10272 22052
rect 11238 22040 11244 22052
rect 11296 22040 11302 22092
rect 12253 22083 12311 22089
rect 12253 22049 12265 22083
rect 12299 22080 12311 22083
rect 12452 22080 12480 22120
rect 12713 22117 12725 22120
rect 12759 22148 12771 22151
rect 13354 22148 13360 22160
rect 12759 22120 13360 22148
rect 12759 22117 12771 22120
rect 12713 22111 12771 22117
rect 13354 22108 13360 22120
rect 13412 22108 13418 22160
rect 16574 22148 16580 22160
rect 15764 22120 16580 22148
rect 12299 22052 12480 22080
rect 13909 22083 13967 22089
rect 12299 22049 12311 22052
rect 12253 22043 12311 22049
rect 13909 22049 13921 22083
rect 13955 22080 13967 22083
rect 13998 22080 14004 22092
rect 13955 22052 14004 22080
rect 13955 22049 13967 22052
rect 13909 22043 13967 22049
rect 13998 22040 14004 22052
rect 14056 22040 14062 22092
rect 14185 22083 14243 22089
rect 14185 22049 14197 22083
rect 14231 22080 14243 22083
rect 14826 22080 14832 22092
rect 14231 22052 14832 22080
rect 14231 22049 14243 22052
rect 14185 22043 14243 22049
rect 14826 22040 14832 22052
rect 14884 22040 14890 22092
rect 15013 22083 15071 22089
rect 15013 22049 15025 22083
rect 15059 22080 15071 22083
rect 15102 22080 15108 22092
rect 15059 22052 15108 22080
rect 15059 22049 15071 22052
rect 15013 22043 15071 22049
rect 10137 22015 10195 22021
rect 10137 22012 10149 22015
rect 10100 21984 10149 22012
rect 10100 21972 10106 21984
rect 10137 21981 10149 21984
rect 10183 21981 10195 22015
rect 10137 21975 10195 21981
rect 10229 22015 10287 22021
rect 10229 21981 10241 22015
rect 10275 21981 10287 22015
rect 12802 22012 12808 22024
rect 12763 21984 12808 22012
rect 10229 21975 10287 21981
rect 12802 21972 12808 21984
rect 12860 21972 12866 22024
rect 12986 22012 12992 22024
rect 12947 21984 12992 22012
rect 12986 21972 12992 21984
rect 13044 21972 13050 22024
rect 14274 21972 14280 22024
rect 14332 22012 14338 22024
rect 15028 22012 15056 22043
rect 15102 22040 15108 22052
rect 15160 22040 15166 22092
rect 15764 22021 15792 22120
rect 16574 22108 16580 22120
rect 16632 22108 16638 22160
rect 17954 22108 17960 22160
rect 18012 22148 18018 22160
rect 18601 22151 18659 22157
rect 18601 22148 18613 22151
rect 18012 22120 18613 22148
rect 18012 22108 18018 22120
rect 18601 22117 18613 22120
rect 18647 22117 18659 22151
rect 18601 22111 18659 22117
rect 19334 22108 19340 22160
rect 19392 22148 19398 22160
rect 20732 22148 20760 22176
rect 21146 22151 21204 22157
rect 21146 22148 21158 22151
rect 19392 22120 20668 22148
rect 20732 22120 21158 22148
rect 19392 22108 19398 22120
rect 16016 22083 16074 22089
rect 16016 22049 16028 22083
rect 16062 22080 16074 22083
rect 16390 22080 16396 22092
rect 16062 22052 16396 22080
rect 16062 22049 16074 22052
rect 16016 22043 16074 22049
rect 16390 22040 16396 22052
rect 16448 22040 16454 22092
rect 18414 22040 18420 22092
rect 18472 22080 18478 22092
rect 18693 22083 18751 22089
rect 18693 22080 18705 22083
rect 18472 22052 18705 22080
rect 18472 22040 18478 22052
rect 18693 22049 18705 22052
rect 18739 22049 18751 22083
rect 20640 22080 20668 22120
rect 21146 22117 21158 22120
rect 21192 22117 21204 22151
rect 22554 22148 22560 22160
rect 21146 22111 21204 22117
rect 22480 22120 22560 22148
rect 21634 22080 21640 22092
rect 20640 22052 21640 22080
rect 18693 22043 18751 22049
rect 15749 22015 15807 22021
rect 15749 22012 15761 22015
rect 14332 21984 15056 22012
rect 15488 21984 15761 22012
rect 14332 21972 14338 21984
rect 2317 21947 2375 21953
rect 2317 21913 2329 21947
rect 2363 21944 2375 21947
rect 2590 21944 2596 21956
rect 2363 21916 2596 21944
rect 2363 21913 2375 21916
rect 2317 21907 2375 21913
rect 2590 21904 2596 21916
rect 2648 21904 2654 21956
rect 8297 21947 8355 21953
rect 8297 21913 8309 21947
rect 8343 21944 8355 21947
rect 8386 21944 8392 21956
rect 8343 21916 8392 21944
rect 8343 21913 8355 21916
rect 8297 21907 8355 21913
rect 8386 21904 8392 21916
rect 8444 21904 8450 21956
rect 9677 21947 9735 21953
rect 9677 21913 9689 21947
rect 9723 21944 9735 21947
rect 10962 21944 10968 21956
rect 9723 21916 10968 21944
rect 9723 21913 9735 21916
rect 9677 21907 9735 21913
rect 10962 21904 10968 21916
rect 11020 21944 11026 21956
rect 11057 21947 11115 21953
rect 11057 21944 11069 21947
rect 11020 21916 11069 21944
rect 11020 21904 11026 21916
rect 11057 21913 11069 21916
rect 11103 21913 11115 21947
rect 11422 21944 11428 21956
rect 11383 21916 11428 21944
rect 11057 21907 11115 21913
rect 11422 21904 11428 21916
rect 11480 21904 11486 21956
rect 2406 21876 2412 21888
rect 2367 21848 2412 21876
rect 2406 21836 2412 21848
rect 2464 21836 2470 21888
rect 6454 21876 6460 21888
rect 6415 21848 6460 21876
rect 6454 21836 6460 21848
rect 6512 21836 6518 21888
rect 7650 21836 7656 21888
rect 7708 21876 7714 21888
rect 8757 21879 8815 21885
rect 8757 21876 8769 21879
rect 7708 21848 8769 21876
rect 7708 21836 7714 21848
rect 8757 21845 8769 21848
rect 8803 21876 8815 21879
rect 9030 21876 9036 21888
rect 8803 21848 9036 21876
rect 8803 21845 8815 21848
rect 8757 21839 8815 21845
rect 9030 21836 9036 21848
rect 9088 21836 9094 21888
rect 9125 21879 9183 21885
rect 9125 21845 9137 21879
rect 9171 21876 9183 21879
rect 9306 21876 9312 21888
rect 9171 21848 9312 21876
rect 9171 21845 9183 21848
rect 9125 21839 9183 21845
rect 9306 21836 9312 21848
rect 9364 21836 9370 21888
rect 10781 21879 10839 21885
rect 10781 21845 10793 21879
rect 10827 21876 10839 21879
rect 11238 21876 11244 21888
rect 10827 21848 11244 21876
rect 10827 21845 10839 21848
rect 10781 21839 10839 21845
rect 11238 21836 11244 21848
rect 11296 21836 11302 21888
rect 11885 21879 11943 21885
rect 11885 21845 11897 21879
rect 11931 21876 11943 21879
rect 12250 21876 12256 21888
rect 11931 21848 12256 21876
rect 11931 21845 11943 21848
rect 11885 21839 11943 21845
rect 12250 21836 12256 21848
rect 12308 21836 12314 21888
rect 15286 21836 15292 21888
rect 15344 21876 15350 21888
rect 15488 21885 15516 21984
rect 15749 21981 15761 21984
rect 15795 21981 15807 22015
rect 18782 22012 18788 22024
rect 18743 21984 18788 22012
rect 15749 21975 15807 21981
rect 18782 21972 18788 21984
rect 18840 21972 18846 22024
rect 19886 21972 19892 22024
rect 19944 22012 19950 22024
rect 20070 22012 20076 22024
rect 19944 21984 20076 22012
rect 19944 21972 19950 21984
rect 20070 21972 20076 21984
rect 20128 21972 20134 22024
rect 20254 21972 20260 22024
rect 20312 21972 20318 22024
rect 20916 22021 20944 22052
rect 21634 22040 21640 22052
rect 21692 22080 21698 22092
rect 22480 22080 22508 22120
rect 22554 22108 22560 22120
rect 22612 22108 22618 22160
rect 23474 22108 23480 22160
rect 23532 22148 23538 22160
rect 23998 22151 24056 22157
rect 23998 22148 24010 22151
rect 23532 22120 24010 22148
rect 23532 22108 23538 22120
rect 23998 22117 24010 22120
rect 24044 22148 24056 22151
rect 24762 22148 24768 22160
rect 24044 22120 24768 22148
rect 24044 22117 24056 22120
rect 23998 22111 24056 22117
rect 24762 22108 24768 22120
rect 24820 22108 24826 22160
rect 23382 22080 23388 22092
rect 21692 22052 21956 22080
rect 22480 22052 23388 22080
rect 21692 22040 21698 22052
rect 20901 22015 20959 22021
rect 20901 22012 20913 22015
rect 20824 21984 20913 22012
rect 18233 21947 18291 21953
rect 18233 21913 18245 21947
rect 18279 21944 18291 21947
rect 19058 21944 19064 21956
rect 18279 21916 19064 21944
rect 18279 21913 18291 21916
rect 18233 21907 18291 21913
rect 19058 21904 19064 21916
rect 19116 21904 19122 21956
rect 19978 21904 19984 21956
rect 20036 21944 20042 21956
rect 20272 21944 20300 21972
rect 20036 21916 20300 21944
rect 20036 21904 20042 21916
rect 20824 21888 20852 21984
rect 20901 21981 20913 21984
rect 20947 21981 20959 22015
rect 21928 22012 21956 22052
rect 23382 22040 23388 22052
rect 23440 22040 23446 22092
rect 23293 22015 23351 22021
rect 23293 22012 23305 22015
rect 21928 21984 23305 22012
rect 20901 21975 20959 21981
rect 23293 21981 23305 21984
rect 23339 22012 23351 22015
rect 23661 22015 23719 22021
rect 23661 22012 23673 22015
rect 23339 21984 23673 22012
rect 23339 21981 23351 21984
rect 23293 21975 23351 21981
rect 23661 21981 23673 21984
rect 23707 22012 23719 22015
rect 23750 22012 23756 22024
rect 23707 21984 23756 22012
rect 23707 21981 23719 21984
rect 23661 21975 23719 21981
rect 23750 21972 23756 21984
rect 23808 21972 23814 22024
rect 15473 21879 15531 21885
rect 15473 21876 15485 21879
rect 15344 21848 15485 21876
rect 15344 21836 15350 21848
rect 15473 21845 15485 21848
rect 15519 21845 15531 21879
rect 15473 21839 15531 21845
rect 17494 21836 17500 21888
rect 17552 21876 17558 21888
rect 17681 21879 17739 21885
rect 17681 21876 17693 21879
rect 17552 21848 17693 21876
rect 17552 21836 17558 21848
rect 17681 21845 17693 21848
rect 17727 21845 17739 21879
rect 18138 21876 18144 21888
rect 18099 21848 18144 21876
rect 17681 21839 17739 21845
rect 18138 21836 18144 21848
rect 18196 21836 18202 21888
rect 20254 21836 20260 21888
rect 20312 21876 20318 21888
rect 20530 21876 20536 21888
rect 20312 21848 20536 21876
rect 20312 21836 20318 21848
rect 20530 21836 20536 21848
rect 20588 21836 20594 21888
rect 20806 21836 20812 21888
rect 20864 21836 20870 21888
rect 25130 21876 25136 21888
rect 25091 21848 25136 21876
rect 25130 21836 25136 21848
rect 25188 21836 25194 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1854 21672 1860 21684
rect 1815 21644 1860 21672
rect 1854 21632 1860 21644
rect 1912 21632 1918 21684
rect 2225 21675 2283 21681
rect 2225 21641 2237 21675
rect 2271 21672 2283 21675
rect 2682 21672 2688 21684
rect 2271 21644 2688 21672
rect 2271 21641 2283 21644
rect 2225 21635 2283 21641
rect 2682 21632 2688 21644
rect 2740 21632 2746 21684
rect 5074 21672 5080 21684
rect 5035 21644 5080 21672
rect 5074 21632 5080 21644
rect 5132 21632 5138 21684
rect 6273 21675 6331 21681
rect 6273 21641 6285 21675
rect 6319 21672 6331 21675
rect 6822 21672 6828 21684
rect 6319 21644 6828 21672
rect 6319 21641 6331 21644
rect 6273 21635 6331 21641
rect 6822 21632 6828 21644
rect 6880 21632 6886 21684
rect 7098 21672 7104 21684
rect 7059 21644 7104 21672
rect 7098 21632 7104 21644
rect 7156 21632 7162 21684
rect 9674 21672 9680 21684
rect 9635 21644 9680 21672
rect 9674 21632 9680 21644
rect 9732 21632 9738 21684
rect 10505 21675 10563 21681
rect 10505 21641 10517 21675
rect 10551 21672 10563 21675
rect 10778 21672 10784 21684
rect 10551 21644 10784 21672
rect 10551 21641 10563 21644
rect 10505 21635 10563 21641
rect 10778 21632 10784 21644
rect 10836 21632 10842 21684
rect 11606 21632 11612 21684
rect 11664 21672 11670 21684
rect 11793 21675 11851 21681
rect 11793 21672 11805 21675
rect 11664 21644 11805 21672
rect 11664 21632 11670 21644
rect 11793 21641 11805 21644
rect 11839 21641 11851 21675
rect 11793 21635 11851 21641
rect 5534 21564 5540 21616
rect 5592 21604 5598 21616
rect 6546 21604 6552 21616
rect 5592 21576 6552 21604
rect 5592 21564 5598 21576
rect 6546 21564 6552 21576
rect 6604 21564 6610 21616
rect 2314 21536 2320 21548
rect 2275 21508 2320 21536
rect 2314 21496 2320 21508
rect 2372 21496 2378 21548
rect 5442 21496 5448 21548
rect 5500 21536 5506 21548
rect 5629 21539 5687 21545
rect 5629 21536 5641 21539
rect 5500 21508 5641 21536
rect 5500 21496 5506 21508
rect 5629 21505 5641 21508
rect 5675 21505 5687 21539
rect 7558 21536 7564 21548
rect 7519 21508 7564 21536
rect 5629 21499 5687 21505
rect 7558 21496 7564 21508
rect 7616 21496 7622 21548
rect 10962 21536 10968 21548
rect 10923 21508 10968 21536
rect 10962 21496 10968 21508
rect 11020 21496 11026 21548
rect 11149 21539 11207 21545
rect 11149 21505 11161 21539
rect 11195 21536 11207 21539
rect 11238 21536 11244 21548
rect 11195 21508 11244 21536
rect 11195 21505 11207 21508
rect 11149 21499 11207 21505
rect 11238 21496 11244 21508
rect 11296 21496 11302 21548
rect 11808 21536 11836 21635
rect 12066 21632 12072 21684
rect 12124 21672 12130 21684
rect 12437 21675 12495 21681
rect 12437 21672 12449 21675
rect 12124 21644 12449 21672
rect 12124 21632 12130 21644
rect 12437 21641 12449 21644
rect 12483 21641 12495 21675
rect 12437 21635 12495 21641
rect 12986 21632 12992 21684
rect 13044 21672 13050 21684
rect 13449 21675 13507 21681
rect 13449 21672 13461 21675
rect 13044 21644 13461 21672
rect 13044 21632 13050 21644
rect 13449 21641 13461 21644
rect 13495 21641 13507 21675
rect 17034 21672 17040 21684
rect 16995 21644 17040 21672
rect 13449 21635 13507 21641
rect 17034 21632 17040 21644
rect 17092 21632 17098 21684
rect 17770 21672 17776 21684
rect 17731 21644 17776 21672
rect 17770 21632 17776 21644
rect 17828 21632 17834 21684
rect 20441 21675 20499 21681
rect 20441 21641 20453 21675
rect 20487 21672 20499 21675
rect 20622 21672 20628 21684
rect 20487 21644 20628 21672
rect 20487 21641 20499 21644
rect 20441 21635 20499 21641
rect 20622 21632 20628 21644
rect 20680 21632 20686 21684
rect 22002 21672 22008 21684
rect 21963 21644 22008 21672
rect 22002 21632 22008 21644
rect 22060 21632 22066 21684
rect 24762 21672 24768 21684
rect 24723 21644 24768 21672
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 25130 21672 25136 21684
rect 25091 21644 25136 21672
rect 25130 21632 25136 21644
rect 25188 21632 25194 21684
rect 12802 21564 12808 21616
rect 12860 21604 12866 21616
rect 13817 21607 13875 21613
rect 13817 21604 13829 21607
rect 12860 21576 13829 21604
rect 12860 21564 12866 21576
rect 13817 21573 13829 21576
rect 13863 21573 13875 21607
rect 13817 21567 13875 21573
rect 17497 21607 17555 21613
rect 17497 21573 17509 21607
rect 17543 21604 17555 21607
rect 18782 21604 18788 21616
rect 17543 21576 18788 21604
rect 17543 21573 17555 21576
rect 17497 21567 17555 21573
rect 18782 21564 18788 21576
rect 18840 21564 18846 21616
rect 22094 21564 22100 21616
rect 22152 21604 22158 21616
rect 22152 21576 22692 21604
rect 22152 21564 22158 21576
rect 12989 21539 13047 21545
rect 12989 21536 13001 21539
rect 11808 21508 13001 21536
rect 12989 21505 13001 21508
rect 13035 21536 13047 21539
rect 13722 21536 13728 21548
rect 13035 21508 13728 21536
rect 13035 21505 13047 21508
rect 12989 21499 13047 21505
rect 13722 21496 13728 21508
rect 13780 21496 13786 21548
rect 14274 21496 14280 21548
rect 14332 21536 14338 21548
rect 14369 21539 14427 21545
rect 14369 21536 14381 21539
rect 14332 21508 14381 21536
rect 14332 21496 14338 21508
rect 14369 21505 14381 21508
rect 14415 21505 14427 21539
rect 14369 21499 14427 21505
rect 18138 21496 18144 21548
rect 18196 21536 18202 21548
rect 18601 21539 18659 21545
rect 18601 21536 18613 21539
rect 18196 21508 18613 21536
rect 18196 21496 18202 21508
rect 18601 21505 18613 21508
rect 18647 21505 18659 21539
rect 18601 21499 18659 21505
rect 19521 21539 19579 21545
rect 19521 21505 19533 21539
rect 19567 21536 19579 21539
rect 20714 21536 20720 21548
rect 19567 21508 20720 21536
rect 19567 21505 19579 21508
rect 19521 21499 19579 21505
rect 20714 21496 20720 21508
rect 20772 21536 20778 21548
rect 20993 21539 21051 21545
rect 20993 21536 21005 21539
rect 20772 21508 21005 21536
rect 20772 21496 20778 21508
rect 20993 21505 21005 21508
rect 21039 21536 21051 21539
rect 21453 21539 21511 21545
rect 21453 21536 21465 21539
rect 21039 21508 21465 21536
rect 21039 21505 21051 21508
rect 20993 21499 21051 21505
rect 21453 21505 21465 21508
rect 21499 21505 21511 21539
rect 21453 21499 21511 21505
rect 21913 21539 21971 21545
rect 21913 21505 21925 21539
rect 21959 21536 21971 21539
rect 22002 21536 22008 21548
rect 21959 21508 22008 21536
rect 21959 21505 21971 21508
rect 21913 21499 21971 21505
rect 22002 21496 22008 21508
rect 22060 21496 22066 21548
rect 22664 21545 22692 21576
rect 22649 21539 22707 21545
rect 22649 21505 22661 21539
rect 22695 21505 22707 21539
rect 24302 21536 24308 21548
rect 24215 21508 24308 21536
rect 22649 21499 22707 21505
rect 24302 21496 24308 21508
rect 24360 21536 24366 21548
rect 25148 21536 25176 21632
rect 25406 21536 25412 21548
rect 24360 21508 25176 21536
rect 25367 21508 25412 21536
rect 24360 21496 24366 21508
rect 25406 21496 25412 21508
rect 25464 21496 25470 21548
rect 2590 21477 2596 21480
rect 2584 21468 2596 21477
rect 2551 21440 2596 21468
rect 2584 21431 2596 21440
rect 2648 21468 2654 21480
rect 3602 21468 3608 21480
rect 2648 21440 3608 21468
rect 2590 21428 2596 21431
rect 2648 21428 2654 21440
rect 3602 21428 3608 21440
rect 3660 21428 3666 21480
rect 7650 21428 7656 21480
rect 7708 21468 7714 21480
rect 7828 21471 7886 21477
rect 7828 21468 7840 21471
rect 7708 21440 7840 21468
rect 7708 21428 7714 21440
rect 7828 21437 7840 21440
rect 7874 21468 7886 21471
rect 8202 21468 8208 21480
rect 7874 21440 8208 21468
rect 7874 21437 7886 21440
rect 7828 21431 7886 21437
rect 8202 21428 8208 21440
rect 8260 21428 8266 21480
rect 12253 21471 12311 21477
rect 12253 21437 12265 21471
rect 12299 21468 12311 21471
rect 12897 21471 12955 21477
rect 12897 21468 12909 21471
rect 12299 21440 12909 21468
rect 12299 21437 12311 21440
rect 12253 21431 12311 21437
rect 12897 21437 12909 21440
rect 12943 21468 12955 21471
rect 13078 21468 13084 21480
rect 12943 21440 13084 21468
rect 12943 21437 12955 21440
rect 12897 21431 12955 21437
rect 13078 21428 13084 21440
rect 13136 21428 13142 21480
rect 13170 21428 13176 21480
rect 13228 21468 13234 21480
rect 15930 21468 15936 21480
rect 13228 21440 15936 21468
rect 13228 21428 13234 21440
rect 15930 21428 15936 21440
rect 15988 21428 15994 21480
rect 16853 21471 16911 21477
rect 16853 21437 16865 21471
rect 16899 21437 16911 21471
rect 18506 21468 18512 21480
rect 18419 21440 18512 21468
rect 16853 21431 16911 21437
rect 4985 21403 5043 21409
rect 4985 21369 4997 21403
rect 5031 21400 5043 21403
rect 5537 21403 5595 21409
rect 5537 21400 5549 21403
rect 5031 21372 5549 21400
rect 5031 21369 5043 21372
rect 4985 21363 5043 21369
rect 5537 21369 5549 21372
rect 5583 21400 5595 21403
rect 7469 21403 7527 21409
rect 7469 21400 7481 21403
rect 5583 21372 7481 21400
rect 5583 21369 5595 21372
rect 5537 21363 5595 21369
rect 7469 21369 7481 21372
rect 7515 21400 7527 21403
rect 8110 21400 8116 21412
rect 7515 21372 8116 21400
rect 7515 21369 7527 21372
rect 7469 21363 7527 21369
rect 8110 21360 8116 21372
rect 8168 21360 8174 21412
rect 10226 21360 10232 21412
rect 10284 21400 10290 21412
rect 10778 21400 10784 21412
rect 10284 21372 10784 21400
rect 10284 21360 10290 21372
rect 10778 21360 10784 21372
rect 10836 21360 10842 21412
rect 14277 21403 14335 21409
rect 14277 21369 14289 21403
rect 14323 21400 14335 21403
rect 14636 21403 14694 21409
rect 14636 21400 14648 21403
rect 14323 21372 14648 21400
rect 14323 21369 14335 21372
rect 14277 21363 14335 21369
rect 14636 21369 14648 21372
rect 14682 21400 14694 21403
rect 14734 21400 14740 21412
rect 14682 21372 14740 21400
rect 14682 21369 14694 21372
rect 14636 21363 14694 21369
rect 14734 21360 14740 21372
rect 14792 21360 14798 21412
rect 2682 21292 2688 21344
rect 2740 21332 2746 21344
rect 3697 21335 3755 21341
rect 3697 21332 3709 21335
rect 2740 21304 3709 21332
rect 2740 21292 2746 21304
rect 3697 21301 3709 21304
rect 3743 21332 3755 21335
rect 4249 21335 4307 21341
rect 4249 21332 4261 21335
rect 3743 21304 4261 21332
rect 3743 21301 3755 21304
rect 3697 21295 3755 21301
rect 4249 21301 4261 21304
rect 4295 21332 4307 21335
rect 4338 21332 4344 21344
rect 4295 21304 4344 21332
rect 4295 21301 4307 21304
rect 4249 21295 4307 21301
rect 4338 21292 4344 21304
rect 4396 21292 4402 21344
rect 5166 21292 5172 21344
rect 5224 21332 5230 21344
rect 5445 21335 5503 21341
rect 5445 21332 5457 21335
rect 5224 21304 5457 21332
rect 5224 21292 5230 21304
rect 5445 21301 5457 21304
rect 5491 21301 5503 21335
rect 5445 21295 5503 21301
rect 8294 21292 8300 21344
rect 8352 21332 8358 21344
rect 8941 21335 8999 21341
rect 8941 21332 8953 21335
rect 8352 21304 8953 21332
rect 8352 21292 8358 21304
rect 8941 21301 8953 21304
rect 8987 21301 8999 21335
rect 10042 21332 10048 21344
rect 10003 21304 10048 21332
rect 8941 21295 8999 21301
rect 10042 21292 10048 21304
rect 10100 21292 10106 21344
rect 10873 21335 10931 21341
rect 10873 21301 10885 21335
rect 10919 21332 10931 21335
rect 12250 21332 12256 21344
rect 10919 21304 12256 21332
rect 10919 21301 10931 21304
rect 10873 21295 10931 21301
rect 12250 21292 12256 21304
rect 12308 21292 12314 21344
rect 12434 21292 12440 21344
rect 12492 21332 12498 21344
rect 12805 21335 12863 21341
rect 12805 21332 12817 21335
rect 12492 21304 12817 21332
rect 12492 21292 12498 21304
rect 12805 21301 12817 21304
rect 12851 21301 12863 21335
rect 15746 21332 15752 21344
rect 15707 21304 15752 21332
rect 12805 21295 12863 21301
rect 15746 21292 15752 21304
rect 15804 21292 15810 21344
rect 16390 21332 16396 21344
rect 16351 21304 16396 21332
rect 16390 21292 16396 21304
rect 16448 21292 16454 21344
rect 16761 21335 16819 21341
rect 16761 21301 16773 21335
rect 16807 21332 16819 21335
rect 16868 21332 16896 21431
rect 18506 21428 18512 21440
rect 18564 21468 18570 21480
rect 19797 21471 19855 21477
rect 19797 21468 19809 21471
rect 18564 21440 19809 21468
rect 18564 21428 18570 21440
rect 19797 21437 19809 21440
rect 19843 21437 19855 21471
rect 22462 21468 22468 21480
rect 22423 21440 22468 21468
rect 19797 21431 19855 21437
rect 22462 21428 22468 21440
rect 22520 21428 22526 21480
rect 23474 21428 23480 21480
rect 23532 21468 23538 21480
rect 24029 21471 24087 21477
rect 24029 21468 24041 21471
rect 23532 21440 24041 21468
rect 23532 21428 23538 21440
rect 24029 21437 24041 21440
rect 24075 21437 24087 21471
rect 25222 21468 25228 21480
rect 25183 21440 25228 21468
rect 24029 21431 24087 21437
rect 25222 21428 25228 21440
rect 25280 21468 25286 21480
rect 25961 21471 26019 21477
rect 25961 21468 25973 21471
rect 25280 21440 25973 21468
rect 25280 21428 25286 21440
rect 25961 21437 25973 21440
rect 26007 21437 26019 21471
rect 25961 21431 26019 21437
rect 17494 21360 17500 21412
rect 17552 21400 17558 21412
rect 18417 21403 18475 21409
rect 18417 21400 18429 21403
rect 17552 21372 18429 21400
rect 17552 21360 17558 21372
rect 18417 21369 18429 21372
rect 18463 21369 18475 21403
rect 18417 21363 18475 21369
rect 20438 21360 20444 21412
rect 20496 21400 20502 21412
rect 20809 21403 20867 21409
rect 20809 21400 20821 21403
rect 20496 21372 20821 21400
rect 20496 21360 20502 21372
rect 20809 21369 20821 21372
rect 20855 21369 20867 21403
rect 20809 21363 20867 21369
rect 22094 21360 22100 21412
rect 22152 21400 22158 21412
rect 23109 21403 23167 21409
rect 23109 21400 23121 21403
rect 22152 21372 23121 21400
rect 22152 21360 22158 21372
rect 23109 21369 23121 21372
rect 23155 21400 23167 21403
rect 24121 21403 24179 21409
rect 24121 21400 24133 21403
rect 23155 21372 24133 21400
rect 23155 21369 23167 21372
rect 23109 21363 23167 21369
rect 24121 21369 24133 21372
rect 24167 21369 24179 21403
rect 24121 21363 24179 21369
rect 16942 21332 16948 21344
rect 16807 21304 16948 21332
rect 16807 21301 16819 21304
rect 16761 21295 16819 21301
rect 16942 21292 16948 21304
rect 17000 21292 17006 21344
rect 17862 21292 17868 21344
rect 17920 21332 17926 21344
rect 18049 21335 18107 21341
rect 18049 21332 18061 21335
rect 17920 21304 18061 21332
rect 17920 21292 17926 21304
rect 18049 21301 18061 21304
rect 18095 21301 18107 21335
rect 18049 21295 18107 21301
rect 18322 21292 18328 21344
rect 18380 21332 18386 21344
rect 19061 21335 19119 21341
rect 19061 21332 19073 21335
rect 18380 21304 19073 21332
rect 18380 21292 18386 21304
rect 19061 21301 19073 21304
rect 19107 21301 19119 21335
rect 19061 21295 19119 21301
rect 20349 21335 20407 21341
rect 20349 21301 20361 21335
rect 20395 21332 20407 21335
rect 20901 21335 20959 21341
rect 20901 21332 20913 21335
rect 20395 21304 20913 21332
rect 20395 21301 20407 21304
rect 20349 21295 20407 21301
rect 20901 21301 20913 21304
rect 20947 21332 20959 21335
rect 21634 21332 21640 21344
rect 20947 21304 21640 21332
rect 20947 21301 20959 21304
rect 20901 21295 20959 21301
rect 21634 21292 21640 21304
rect 21692 21292 21698 21344
rect 22373 21335 22431 21341
rect 22373 21301 22385 21335
rect 22419 21332 22431 21335
rect 22554 21332 22560 21344
rect 22419 21304 22560 21332
rect 22419 21301 22431 21304
rect 22373 21295 22431 21301
rect 22554 21292 22560 21304
rect 22612 21292 22618 21344
rect 23474 21332 23480 21344
rect 23435 21304 23480 21332
rect 23474 21292 23480 21304
rect 23532 21292 23538 21344
rect 23658 21332 23664 21344
rect 23619 21304 23664 21332
rect 23658 21292 23664 21304
rect 23716 21292 23722 21344
rect 26326 21332 26332 21344
rect 26287 21304 26332 21332
rect 26326 21292 26332 21304
rect 26384 21292 26390 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 2038 21128 2044 21140
rect 1999 21100 2044 21128
rect 2038 21088 2044 21100
rect 2096 21088 2102 21140
rect 2501 21131 2559 21137
rect 2501 21097 2513 21131
rect 2547 21128 2559 21131
rect 2958 21128 2964 21140
rect 2547 21100 2964 21128
rect 2547 21097 2559 21100
rect 2501 21091 2559 21097
rect 2958 21088 2964 21100
rect 3016 21128 3022 21140
rect 4065 21131 4123 21137
rect 4065 21128 4077 21131
rect 3016 21100 4077 21128
rect 3016 21088 3022 21100
rect 4065 21097 4077 21100
rect 4111 21097 4123 21131
rect 4522 21128 4528 21140
rect 4483 21100 4528 21128
rect 4065 21091 4123 21097
rect 4522 21088 4528 21100
rect 4580 21088 4586 21140
rect 5166 21128 5172 21140
rect 5127 21100 5172 21128
rect 5166 21088 5172 21100
rect 5224 21088 5230 21140
rect 5442 21128 5448 21140
rect 5403 21100 5448 21128
rect 5442 21088 5448 21100
rect 5500 21088 5506 21140
rect 6454 21128 6460 21140
rect 6415 21100 6460 21128
rect 6454 21088 6460 21100
rect 6512 21088 6518 21140
rect 7650 21128 7656 21140
rect 7611 21100 7656 21128
rect 7650 21088 7656 21100
rect 7708 21088 7714 21140
rect 8202 21088 8208 21140
rect 8260 21128 8266 21140
rect 8481 21131 8539 21137
rect 8481 21128 8493 21131
rect 8260 21100 8493 21128
rect 8260 21088 8266 21100
rect 8481 21097 8493 21100
rect 8527 21128 8539 21131
rect 8570 21128 8576 21140
rect 8527 21100 8576 21128
rect 8527 21097 8539 21100
rect 8481 21091 8539 21097
rect 8570 21088 8576 21100
rect 8628 21088 8634 21140
rect 9030 21128 9036 21140
rect 8991 21100 9036 21128
rect 9030 21088 9036 21100
rect 9088 21088 9094 21140
rect 9398 21128 9404 21140
rect 9359 21100 9404 21128
rect 9398 21088 9404 21100
rect 9456 21088 9462 21140
rect 14550 21128 14556 21140
rect 14511 21100 14556 21128
rect 14550 21088 14556 21100
rect 14608 21128 14614 21140
rect 14829 21131 14887 21137
rect 14829 21128 14841 21131
rect 14608 21100 14841 21128
rect 14608 21088 14614 21100
rect 14829 21097 14841 21100
rect 14875 21097 14887 21131
rect 16666 21128 16672 21140
rect 16627 21100 16672 21128
rect 14829 21091 14887 21097
rect 16666 21088 16672 21100
rect 16724 21088 16730 21140
rect 19150 21128 19156 21140
rect 19111 21100 19156 21128
rect 19150 21088 19156 21100
rect 19208 21088 19214 21140
rect 20438 21128 20444 21140
rect 20399 21100 20444 21128
rect 20438 21088 20444 21100
rect 20496 21088 20502 21140
rect 20530 21088 20536 21140
rect 20588 21128 20594 21140
rect 22002 21128 22008 21140
rect 20588 21100 22008 21128
rect 20588 21088 20594 21100
rect 22002 21088 22008 21100
rect 22060 21088 22066 21140
rect 22186 21128 22192 21140
rect 22147 21100 22192 21128
rect 22186 21088 22192 21100
rect 22244 21088 22250 21140
rect 22649 21131 22707 21137
rect 22649 21097 22661 21131
rect 22695 21128 22707 21131
rect 23658 21128 23664 21140
rect 22695 21100 23664 21128
rect 22695 21097 22707 21100
rect 22649 21091 22707 21097
rect 23658 21088 23664 21100
rect 23716 21088 23722 21140
rect 3145 21063 3203 21069
rect 3145 21029 3157 21063
rect 3191 21060 3203 21063
rect 3234 21060 3240 21072
rect 3191 21032 3240 21060
rect 3191 21029 3203 21032
rect 3145 21023 3203 21029
rect 3234 21020 3240 21032
rect 3292 21020 3298 21072
rect 4430 21060 4436 21072
rect 4391 21032 4436 21060
rect 4430 21020 4436 21032
rect 4488 21020 4494 21072
rect 8110 21020 8116 21072
rect 8168 21060 8174 21072
rect 8389 21063 8447 21069
rect 8389 21060 8401 21063
rect 8168 21032 8401 21060
rect 8168 21020 8174 21032
rect 8389 21029 8401 21032
rect 8435 21060 8447 21063
rect 9490 21060 9496 21072
rect 8435 21032 9496 21060
rect 8435 21029 8447 21032
rect 8389 21023 8447 21029
rect 9490 21020 9496 21032
rect 9548 21020 9554 21072
rect 13081 21063 13139 21069
rect 13081 21029 13093 21063
rect 13127 21060 13139 21063
rect 13262 21060 13268 21072
rect 13127 21032 13268 21060
rect 13127 21029 13139 21032
rect 13081 21023 13139 21029
rect 13262 21020 13268 21032
rect 13320 21020 13326 21072
rect 15556 21063 15614 21069
rect 15556 21029 15568 21063
rect 15602 21060 15614 21063
rect 15746 21060 15752 21072
rect 15602 21032 15752 21060
rect 15602 21029 15614 21032
rect 15556 21023 15614 21029
rect 15746 21020 15752 21032
rect 15804 21020 15810 21072
rect 19705 21063 19763 21069
rect 19705 21060 19717 21063
rect 17788 21032 19717 21060
rect 1854 20952 1860 21004
rect 1912 20992 1918 21004
rect 2409 20995 2467 21001
rect 2409 20992 2421 20995
rect 1912 20964 2421 20992
rect 1912 20952 1918 20964
rect 2409 20961 2421 20964
rect 2455 20961 2467 20995
rect 7006 20992 7012 21004
rect 2409 20955 2467 20961
rect 6564 20964 7012 20992
rect 2590 20924 2596 20936
rect 2551 20896 2596 20924
rect 2590 20884 2596 20896
rect 2648 20884 2654 20936
rect 3602 20884 3608 20936
rect 3660 20924 3666 20936
rect 4617 20927 4675 20933
rect 4617 20924 4629 20927
rect 3660 20896 4629 20924
rect 3660 20884 3666 20896
rect 4617 20893 4629 20896
rect 4663 20893 4675 20927
rect 4617 20887 4675 20893
rect 6086 20884 6092 20936
rect 6144 20924 6150 20936
rect 6564 20933 6592 20964
rect 7006 20952 7012 20964
rect 7064 20952 7070 21004
rect 9950 20952 9956 21004
rect 10008 20992 10014 21004
rect 10485 20995 10543 21001
rect 10485 20992 10497 20995
rect 10008 20964 10497 20992
rect 10008 20952 10014 20964
rect 10485 20961 10497 20964
rect 10531 20961 10543 20995
rect 17221 20995 17279 21001
rect 17221 20992 17233 20995
rect 10485 20955 10543 20961
rect 15304 20964 17233 20992
rect 15304 20936 15332 20964
rect 17221 20961 17233 20964
rect 17267 20992 17279 20995
rect 17586 20992 17592 21004
rect 17267 20964 17592 20992
rect 17267 20961 17279 20964
rect 17221 20955 17279 20961
rect 17586 20952 17592 20964
rect 17644 20992 17650 21004
rect 17788 21001 17816 21032
rect 19705 21029 19717 21032
rect 19751 21060 19763 21063
rect 20162 21060 20168 21072
rect 19751 21032 20168 21060
rect 19751 21029 19763 21032
rect 19705 21023 19763 21029
rect 20162 21020 20168 21032
rect 20220 21020 20226 21072
rect 21174 21060 21180 21072
rect 20916 21032 21180 21060
rect 18046 21001 18052 21004
rect 17773 20995 17831 21001
rect 17773 20992 17785 20995
rect 17644 20964 17785 20992
rect 17644 20952 17650 20964
rect 17773 20961 17785 20964
rect 17819 20961 17831 20995
rect 18040 20992 18052 21001
rect 17959 20964 18052 20992
rect 17773 20955 17831 20961
rect 18040 20955 18052 20964
rect 18104 20992 18110 21004
rect 20916 21001 20944 21032
rect 21174 21020 21180 21032
rect 21232 21060 21238 21072
rect 22370 21060 22376 21072
rect 21232 21032 22376 21060
rect 21232 21020 21238 21032
rect 22370 21020 22376 21032
rect 22428 21020 22434 21072
rect 23474 21020 23480 21072
rect 23532 21060 23538 21072
rect 23842 21060 23848 21072
rect 23532 21032 23848 21060
rect 23532 21020 23538 21032
rect 23842 21020 23848 21032
rect 23900 21020 23906 21072
rect 24020 21063 24078 21069
rect 24020 21029 24032 21063
rect 24066 21060 24078 21063
rect 24302 21060 24308 21072
rect 24066 21032 24308 21060
rect 24066 21029 24078 21032
rect 24020 21023 24078 21029
rect 24302 21020 24308 21032
rect 24360 21060 24366 21072
rect 24670 21060 24676 21072
rect 24360 21032 24676 21060
rect 24360 21020 24366 21032
rect 24670 21020 24676 21032
rect 24728 21020 24734 21072
rect 20901 20995 20959 21001
rect 18104 20964 19288 20992
rect 18046 20952 18052 20955
rect 18104 20952 18110 20964
rect 19260 20936 19288 20964
rect 20901 20961 20913 20995
rect 20947 20961 20959 20995
rect 20901 20955 20959 20961
rect 22002 20952 22008 21004
rect 22060 20992 22066 21004
rect 22557 20995 22615 21001
rect 22557 20992 22569 20995
rect 22060 20964 22569 20992
rect 22060 20952 22066 20964
rect 22557 20961 22569 20964
rect 22603 20992 22615 20995
rect 23382 20992 23388 21004
rect 22603 20964 23388 20992
rect 22603 20961 22615 20964
rect 22557 20955 22615 20961
rect 23382 20952 23388 20964
rect 23440 20952 23446 21004
rect 23750 20992 23756 21004
rect 23663 20964 23756 20992
rect 23750 20952 23756 20964
rect 23808 20992 23814 21004
rect 24762 20992 24768 21004
rect 23808 20964 24768 20992
rect 23808 20952 23814 20964
rect 24762 20952 24768 20964
rect 24820 20952 24826 21004
rect 6549 20927 6607 20933
rect 6549 20924 6561 20927
rect 6144 20896 6561 20924
rect 6144 20884 6150 20896
rect 6549 20893 6561 20896
rect 6595 20893 6607 20927
rect 6549 20887 6607 20893
rect 6638 20884 6644 20936
rect 6696 20924 6702 20936
rect 7285 20927 7343 20933
rect 6696 20896 6741 20924
rect 6696 20884 6702 20896
rect 7285 20893 7297 20927
rect 7331 20924 7343 20927
rect 8573 20927 8631 20933
rect 8573 20924 8585 20927
rect 7331 20896 8585 20924
rect 7331 20893 7343 20896
rect 7285 20887 7343 20893
rect 8573 20893 8585 20896
rect 8619 20924 8631 20927
rect 9858 20924 9864 20936
rect 8619 20896 9864 20924
rect 8619 20893 8631 20896
rect 8573 20887 8631 20893
rect 9858 20884 9864 20896
rect 9916 20884 9922 20936
rect 10042 20884 10048 20936
rect 10100 20924 10106 20936
rect 10229 20927 10287 20933
rect 10229 20924 10241 20927
rect 10100 20896 10241 20924
rect 10100 20884 10106 20896
rect 10229 20893 10241 20896
rect 10275 20893 10287 20927
rect 10229 20887 10287 20893
rect 12434 20884 12440 20936
rect 12492 20924 12498 20936
rect 13170 20924 13176 20936
rect 12492 20896 12537 20924
rect 13131 20896 13176 20924
rect 12492 20884 12498 20896
rect 13170 20884 13176 20896
rect 13228 20884 13234 20936
rect 13354 20924 13360 20936
rect 13267 20896 13360 20924
rect 13354 20884 13360 20896
rect 13412 20924 13418 20936
rect 13906 20924 13912 20936
rect 13412 20896 13912 20924
rect 13412 20884 13418 20896
rect 13906 20884 13912 20896
rect 13964 20884 13970 20936
rect 14274 20884 14280 20936
rect 14332 20924 14338 20936
rect 15286 20924 15292 20936
rect 14332 20896 15292 20924
rect 14332 20884 14338 20896
rect 15286 20884 15292 20896
rect 15344 20884 15350 20936
rect 19242 20884 19248 20936
rect 19300 20884 19306 20936
rect 20714 20884 20720 20936
rect 20772 20924 20778 20936
rect 21085 20927 21143 20933
rect 21085 20924 21097 20927
rect 20772 20896 21097 20924
rect 20772 20884 20778 20896
rect 21085 20893 21097 20896
rect 21131 20893 21143 20927
rect 21085 20887 21143 20893
rect 22097 20927 22155 20933
rect 22097 20893 22109 20927
rect 22143 20924 22155 20927
rect 22462 20924 22468 20936
rect 22143 20896 22468 20924
rect 22143 20893 22155 20896
rect 22097 20887 22155 20893
rect 22462 20884 22468 20896
rect 22520 20884 22526 20936
rect 22833 20927 22891 20933
rect 22833 20893 22845 20927
rect 22879 20893 22891 20927
rect 22833 20887 22891 20893
rect 11974 20816 11980 20868
rect 12032 20856 12038 20868
rect 12526 20856 12532 20868
rect 12032 20828 12532 20856
rect 12032 20816 12038 20828
rect 12526 20816 12532 20828
rect 12584 20816 12590 20868
rect 14090 20856 14096 20868
rect 13924 20828 14096 20856
rect 13924 20800 13952 20828
rect 14090 20816 14096 20828
rect 14148 20816 14154 20868
rect 22848 20856 22876 20887
rect 23014 20856 23020 20868
rect 22848 20828 23020 20856
rect 23014 20816 23020 20828
rect 23072 20856 23078 20868
rect 23072 20828 23612 20856
rect 23072 20816 23078 20828
rect 1854 20788 1860 20800
rect 1815 20760 1860 20788
rect 1854 20748 1860 20760
rect 1912 20748 1918 20800
rect 3510 20788 3516 20800
rect 3471 20760 3516 20788
rect 3510 20748 3516 20760
rect 3568 20748 3574 20800
rect 3881 20791 3939 20797
rect 3881 20757 3893 20791
rect 3927 20788 3939 20791
rect 3970 20788 3976 20800
rect 3927 20760 3976 20788
rect 3927 20757 3939 20760
rect 3881 20751 3939 20757
rect 3970 20748 3976 20760
rect 4028 20748 4034 20800
rect 5534 20748 5540 20800
rect 5592 20788 5598 20800
rect 5813 20791 5871 20797
rect 5813 20788 5825 20791
rect 5592 20760 5825 20788
rect 5592 20748 5598 20760
rect 5813 20757 5825 20760
rect 5859 20757 5871 20791
rect 5813 20751 5871 20757
rect 6089 20791 6147 20797
rect 6089 20757 6101 20791
rect 6135 20788 6147 20791
rect 6178 20788 6184 20800
rect 6135 20760 6184 20788
rect 6135 20757 6147 20760
rect 6089 20751 6147 20757
rect 6178 20748 6184 20760
rect 6236 20748 6242 20800
rect 8018 20788 8024 20800
rect 7979 20760 8024 20788
rect 8018 20748 8024 20760
rect 8076 20748 8082 20800
rect 9950 20788 9956 20800
rect 9911 20760 9956 20788
rect 9950 20748 9956 20760
rect 10008 20748 10014 20800
rect 11606 20788 11612 20800
rect 11567 20760 11612 20788
rect 11606 20748 11612 20760
rect 11664 20748 11670 20800
rect 12710 20788 12716 20800
rect 12671 20760 12716 20788
rect 12710 20748 12716 20760
rect 12768 20748 12774 20800
rect 13817 20791 13875 20797
rect 13817 20757 13829 20791
rect 13863 20788 13875 20791
rect 13906 20788 13912 20800
rect 13863 20760 13912 20788
rect 13863 20757 13875 20760
rect 13817 20751 13875 20757
rect 13906 20748 13912 20760
rect 13964 20748 13970 20800
rect 13998 20748 14004 20800
rect 14056 20788 14062 20800
rect 14185 20791 14243 20797
rect 14185 20788 14197 20791
rect 14056 20760 14197 20788
rect 14056 20748 14062 20760
rect 14185 20757 14197 20760
rect 14231 20788 14243 20791
rect 14642 20788 14648 20800
rect 14231 20760 14648 20788
rect 14231 20757 14243 20760
rect 14185 20751 14243 20757
rect 14642 20748 14648 20760
rect 14700 20748 14706 20800
rect 19242 20748 19248 20800
rect 19300 20788 19306 20800
rect 20073 20791 20131 20797
rect 20073 20788 20085 20791
rect 19300 20760 20085 20788
rect 19300 20748 19306 20760
rect 20073 20757 20085 20760
rect 20119 20788 20131 20791
rect 20806 20788 20812 20800
rect 20119 20760 20812 20788
rect 20119 20757 20131 20760
rect 20073 20751 20131 20757
rect 20806 20748 20812 20760
rect 20864 20748 20870 20800
rect 21729 20791 21787 20797
rect 21729 20757 21741 20791
rect 21775 20788 21787 20791
rect 21818 20788 21824 20800
rect 21775 20760 21824 20788
rect 21775 20757 21787 20760
rect 21729 20751 21787 20757
rect 21818 20748 21824 20760
rect 21876 20748 21882 20800
rect 22094 20748 22100 20800
rect 22152 20788 22158 20800
rect 22370 20788 22376 20800
rect 22152 20760 22376 20788
rect 22152 20748 22158 20760
rect 22370 20748 22376 20760
rect 22428 20748 22434 20800
rect 22554 20748 22560 20800
rect 22612 20788 22618 20800
rect 23293 20791 23351 20797
rect 23293 20788 23305 20791
rect 22612 20760 23305 20788
rect 22612 20748 22618 20760
rect 23293 20757 23305 20760
rect 23339 20788 23351 20791
rect 23474 20788 23480 20800
rect 23339 20760 23480 20788
rect 23339 20757 23351 20760
rect 23293 20751 23351 20757
rect 23474 20748 23480 20760
rect 23532 20748 23538 20800
rect 23584 20788 23612 20828
rect 25133 20791 25191 20797
rect 25133 20788 25145 20791
rect 23584 20760 25145 20788
rect 25133 20757 25145 20760
rect 25179 20757 25191 20791
rect 25133 20751 25191 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 2133 20587 2191 20593
rect 2133 20553 2145 20587
rect 2179 20584 2191 20587
rect 2590 20584 2596 20596
rect 2179 20556 2596 20584
rect 2179 20553 2191 20556
rect 2133 20547 2191 20553
rect 2590 20544 2596 20556
rect 2648 20544 2654 20596
rect 3602 20584 3608 20596
rect 3563 20556 3608 20584
rect 3602 20544 3608 20556
rect 3660 20584 3666 20596
rect 4157 20587 4215 20593
rect 4157 20584 4169 20587
rect 3660 20556 4169 20584
rect 3660 20544 3666 20556
rect 4157 20553 4169 20556
rect 4203 20553 4215 20587
rect 4157 20547 4215 20553
rect 5813 20587 5871 20593
rect 5813 20553 5825 20587
rect 5859 20584 5871 20587
rect 6086 20584 6092 20596
rect 5859 20556 6092 20584
rect 5859 20553 5871 20556
rect 5813 20547 5871 20553
rect 6086 20544 6092 20556
rect 6144 20544 6150 20596
rect 6181 20587 6239 20593
rect 6181 20553 6193 20587
rect 6227 20584 6239 20587
rect 6454 20584 6460 20596
rect 6227 20556 6460 20584
rect 6227 20553 6239 20556
rect 6181 20547 6239 20553
rect 6454 20544 6460 20556
rect 6512 20544 6518 20596
rect 7745 20587 7803 20593
rect 7745 20553 7757 20587
rect 7791 20584 7803 20587
rect 8202 20584 8208 20596
rect 7791 20556 8208 20584
rect 7791 20553 7803 20556
rect 7745 20547 7803 20553
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 10597 20587 10655 20593
rect 10597 20553 10609 20587
rect 10643 20584 10655 20587
rect 10686 20584 10692 20596
rect 10643 20556 10692 20584
rect 10643 20553 10655 20556
rect 10597 20547 10655 20553
rect 10686 20544 10692 20556
rect 10744 20544 10750 20596
rect 12253 20587 12311 20593
rect 12253 20553 12265 20587
rect 12299 20584 12311 20587
rect 13354 20584 13360 20596
rect 12299 20556 13360 20584
rect 12299 20553 12311 20556
rect 12253 20547 12311 20553
rect 6273 20519 6331 20525
rect 6273 20485 6285 20519
rect 6319 20485 6331 20519
rect 6273 20479 6331 20485
rect 4522 20408 4528 20460
rect 4580 20448 4586 20460
rect 5261 20451 5319 20457
rect 5261 20448 5273 20451
rect 4580 20420 5273 20448
rect 4580 20408 4586 20420
rect 5261 20417 5273 20420
rect 5307 20417 5319 20451
rect 6288 20448 6316 20479
rect 9950 20476 9956 20528
rect 10008 20516 10014 20528
rect 10137 20519 10195 20525
rect 10137 20516 10149 20519
rect 10008 20488 10149 20516
rect 10008 20476 10014 20488
rect 10137 20485 10149 20488
rect 10183 20516 10195 20519
rect 12268 20516 12296 20547
rect 13354 20544 13360 20556
rect 13412 20544 13418 20596
rect 14734 20544 14740 20596
rect 14792 20584 14798 20596
rect 15105 20587 15163 20593
rect 15105 20584 15117 20587
rect 14792 20556 15117 20584
rect 14792 20544 14798 20556
rect 15105 20553 15117 20556
rect 15151 20553 15163 20587
rect 15746 20584 15752 20596
rect 15707 20556 15752 20584
rect 15105 20547 15163 20553
rect 15746 20544 15752 20556
rect 15804 20584 15810 20596
rect 16025 20587 16083 20593
rect 16025 20584 16037 20587
rect 15804 20556 16037 20584
rect 15804 20544 15810 20556
rect 16025 20553 16037 20556
rect 16071 20553 16083 20587
rect 16025 20547 16083 20553
rect 17865 20587 17923 20593
rect 17865 20553 17877 20587
rect 17911 20584 17923 20587
rect 18046 20584 18052 20596
rect 17911 20556 18052 20584
rect 17911 20553 17923 20556
rect 17865 20547 17923 20553
rect 10183 20488 12296 20516
rect 10183 20485 10195 20488
rect 10137 20479 10195 20485
rect 12342 20476 12348 20528
rect 12400 20516 12406 20528
rect 13262 20516 13268 20528
rect 12400 20488 13268 20516
rect 12400 20476 12406 20488
rect 13262 20476 13268 20488
rect 13320 20476 13326 20528
rect 6362 20448 6368 20460
rect 6275 20420 6368 20448
rect 5261 20411 5319 20417
rect 6362 20408 6368 20420
rect 6420 20448 6426 20460
rect 7558 20448 7564 20460
rect 6420 20420 7564 20448
rect 6420 20408 6426 20420
rect 7558 20408 7564 20420
rect 7616 20448 7622 20460
rect 7837 20451 7895 20457
rect 7837 20448 7849 20451
rect 7616 20420 7849 20448
rect 7616 20408 7622 20420
rect 7837 20417 7849 20420
rect 7883 20417 7895 20451
rect 7837 20411 7895 20417
rect 10962 20408 10968 20460
rect 11020 20448 11026 20460
rect 11057 20451 11115 20457
rect 11057 20448 11069 20451
rect 11020 20420 11069 20448
rect 11020 20408 11026 20420
rect 11057 20417 11069 20420
rect 11103 20417 11115 20451
rect 11238 20448 11244 20460
rect 11199 20420 11244 20448
rect 11057 20411 11115 20417
rect 11238 20408 11244 20420
rect 11296 20448 11302 20460
rect 11606 20448 11612 20460
rect 11296 20420 11612 20448
rect 11296 20408 11302 20420
rect 11606 20408 11612 20420
rect 11664 20408 11670 20460
rect 12713 20451 12771 20457
rect 12713 20417 12725 20451
rect 12759 20448 12771 20451
rect 12986 20448 12992 20460
rect 12759 20420 12992 20448
rect 12759 20417 12771 20420
rect 12713 20411 12771 20417
rect 12986 20408 12992 20420
rect 13044 20408 13050 20460
rect 16040 20448 16068 20547
rect 18046 20544 18052 20556
rect 18104 20544 18110 20596
rect 19334 20544 19340 20596
rect 19392 20584 19398 20596
rect 20346 20584 20352 20596
rect 19392 20556 20352 20584
rect 19392 20544 19398 20556
rect 20346 20544 20352 20556
rect 20404 20584 20410 20596
rect 20533 20587 20591 20593
rect 20533 20584 20545 20587
rect 20404 20556 20545 20584
rect 20404 20544 20410 20556
rect 20533 20553 20545 20556
rect 20579 20553 20591 20587
rect 21174 20584 21180 20596
rect 21135 20556 21180 20584
rect 20533 20547 20591 20553
rect 21174 20544 21180 20556
rect 21232 20544 21238 20596
rect 22741 20587 22799 20593
rect 22741 20553 22753 20587
rect 22787 20584 22799 20587
rect 23014 20584 23020 20596
rect 22787 20556 23020 20584
rect 22787 20553 22799 20556
rect 22741 20547 22799 20553
rect 23014 20544 23020 20556
rect 23072 20544 23078 20596
rect 23382 20544 23388 20596
rect 23440 20584 23446 20596
rect 23661 20587 23719 20593
rect 23661 20584 23673 20587
rect 23440 20556 23673 20584
rect 23440 20544 23446 20556
rect 23661 20553 23673 20556
rect 23707 20553 23719 20587
rect 24670 20584 24676 20596
rect 24631 20556 24676 20584
rect 23661 20547 23719 20553
rect 24670 20544 24676 20556
rect 24728 20544 24734 20596
rect 25409 20587 25467 20593
rect 25409 20553 25421 20587
rect 25455 20584 25467 20587
rect 25590 20584 25596 20596
rect 25455 20556 25596 20584
rect 25455 20553 25467 20556
rect 25409 20547 25467 20553
rect 25590 20544 25596 20556
rect 25648 20544 25654 20596
rect 26237 20587 26295 20593
rect 26237 20553 26249 20587
rect 26283 20584 26295 20587
rect 26326 20584 26332 20596
rect 26283 20556 26332 20584
rect 26283 20553 26295 20556
rect 26237 20547 26295 20553
rect 18230 20516 18236 20528
rect 18191 20488 18236 20516
rect 18230 20476 18236 20488
rect 18288 20476 18294 20528
rect 16761 20451 16819 20457
rect 16761 20448 16773 20451
rect 16040 20420 16773 20448
rect 16761 20417 16773 20420
rect 16807 20417 16819 20451
rect 16761 20411 16819 20417
rect 21818 20408 21824 20460
rect 21876 20448 21882 20460
rect 22189 20451 22247 20457
rect 22189 20448 22201 20451
rect 21876 20420 22201 20448
rect 21876 20408 21882 20420
rect 22189 20417 22201 20420
rect 22235 20417 22247 20451
rect 23032 20448 23060 20544
rect 23382 20448 23388 20460
rect 23032 20420 23388 20448
rect 22189 20411 22247 20417
rect 23382 20408 23388 20420
rect 23440 20408 23446 20460
rect 24302 20448 24308 20460
rect 24215 20420 24308 20448
rect 24302 20408 24308 20420
rect 24360 20448 24366 20460
rect 24688 20448 24716 20544
rect 24854 20476 24860 20528
rect 24912 20516 24918 20528
rect 25133 20519 25191 20525
rect 25133 20516 25145 20519
rect 24912 20488 25145 20516
rect 24912 20476 24918 20488
rect 25133 20485 25145 20488
rect 25179 20516 25191 20519
rect 26252 20516 26280 20547
rect 26326 20544 26332 20556
rect 26384 20544 26390 20596
rect 25179 20488 26280 20516
rect 25179 20485 25191 20488
rect 25133 20479 25191 20485
rect 24360 20420 24716 20448
rect 24360 20408 24366 20420
rect 2225 20383 2283 20389
rect 2225 20349 2237 20383
rect 2271 20380 2283 20383
rect 2314 20380 2320 20392
rect 2271 20352 2320 20380
rect 2271 20349 2283 20352
rect 2225 20343 2283 20349
rect 2314 20340 2320 20352
rect 2372 20340 2378 20392
rect 2492 20383 2550 20389
rect 2492 20380 2504 20383
rect 2424 20352 2504 20380
rect 2424 20324 2452 20352
rect 2492 20349 2504 20352
rect 2538 20380 2550 20383
rect 3234 20380 3240 20392
rect 2538 20352 3240 20380
rect 2538 20349 2550 20352
rect 2492 20343 2550 20349
rect 3234 20340 3240 20352
rect 3292 20340 3298 20392
rect 4706 20340 4712 20392
rect 4764 20380 4770 20392
rect 5077 20383 5135 20389
rect 5077 20380 5089 20383
rect 4764 20352 5089 20380
rect 4764 20340 4770 20352
rect 5077 20349 5089 20352
rect 5123 20380 5135 20383
rect 5442 20380 5448 20392
rect 5123 20352 5448 20380
rect 5123 20349 5135 20352
rect 5077 20343 5135 20349
rect 5442 20340 5448 20352
rect 5500 20340 5506 20392
rect 6457 20383 6515 20389
rect 6457 20349 6469 20383
rect 6503 20380 6515 20383
rect 6546 20380 6552 20392
rect 6503 20352 6552 20380
rect 6503 20349 6515 20352
rect 6457 20343 6515 20349
rect 6546 20340 6552 20352
rect 6604 20340 6610 20392
rect 6822 20380 6828 20392
rect 6783 20352 6828 20380
rect 6822 20340 6828 20352
rect 6880 20340 6886 20392
rect 12434 20340 12440 20392
rect 12492 20380 12498 20392
rect 13262 20380 13268 20392
rect 12492 20352 12537 20380
rect 13223 20352 13268 20380
rect 12492 20340 12498 20352
rect 13262 20340 13268 20352
rect 13320 20340 13326 20392
rect 13725 20383 13783 20389
rect 13725 20349 13737 20383
rect 13771 20380 13783 20383
rect 14274 20380 14280 20392
rect 13771 20352 14280 20380
rect 13771 20349 13783 20352
rect 13725 20343 13783 20349
rect 14274 20340 14280 20352
rect 14332 20340 14338 20392
rect 16666 20380 16672 20392
rect 16579 20352 16672 20380
rect 16666 20340 16672 20352
rect 16724 20380 16730 20392
rect 17862 20380 17868 20392
rect 16724 20352 17868 20380
rect 16724 20340 16730 20352
rect 17862 20340 17868 20352
rect 17920 20340 17926 20392
rect 18049 20383 18107 20389
rect 18049 20349 18061 20383
rect 18095 20349 18107 20383
rect 18049 20343 18107 20349
rect 1765 20315 1823 20321
rect 1765 20281 1777 20315
rect 1811 20312 1823 20315
rect 2406 20312 2412 20324
rect 1811 20284 2412 20312
rect 1811 20281 1823 20284
rect 1765 20275 1823 20281
rect 2406 20272 2412 20284
rect 2464 20272 2470 20324
rect 7377 20315 7435 20321
rect 4724 20284 5396 20312
rect 4522 20244 4528 20256
rect 4483 20216 4528 20244
rect 4522 20204 4528 20216
rect 4580 20204 4586 20256
rect 4724 20253 4752 20284
rect 4709 20247 4767 20253
rect 4709 20213 4721 20247
rect 4755 20213 4767 20247
rect 5166 20244 5172 20256
rect 5127 20216 5172 20244
rect 4709 20207 4767 20213
rect 5166 20204 5172 20216
rect 5224 20204 5230 20256
rect 5368 20244 5396 20284
rect 7377 20281 7389 20315
rect 7423 20312 7435 20315
rect 8082 20315 8140 20321
rect 8082 20312 8094 20315
rect 7423 20284 8094 20312
rect 7423 20281 7435 20284
rect 7377 20275 7435 20281
rect 8082 20281 8094 20284
rect 8128 20312 8140 20315
rect 8202 20312 8208 20324
rect 8128 20284 8208 20312
rect 8128 20281 8140 20284
rect 8082 20275 8140 20281
rect 8202 20272 8208 20284
rect 8260 20272 8266 20324
rect 13998 20321 14004 20324
rect 13992 20312 14004 20321
rect 13959 20284 14004 20312
rect 13992 20275 14004 20284
rect 13998 20272 14004 20275
rect 14056 20272 14062 20324
rect 15764 20284 16344 20312
rect 5534 20244 5540 20256
rect 5368 20216 5540 20244
rect 5534 20204 5540 20216
rect 5592 20204 5598 20256
rect 7834 20204 7840 20256
rect 7892 20244 7898 20256
rect 9122 20244 9128 20256
rect 7892 20216 9128 20244
rect 7892 20204 7898 20216
rect 9122 20204 9128 20216
rect 9180 20244 9186 20256
rect 9217 20247 9275 20253
rect 9217 20244 9229 20247
rect 9180 20216 9229 20244
rect 9180 20204 9186 20216
rect 9217 20213 9229 20216
rect 9263 20213 9275 20247
rect 9217 20207 9275 20213
rect 9766 20204 9772 20256
rect 9824 20244 9830 20256
rect 10413 20247 10471 20253
rect 10413 20244 10425 20247
rect 9824 20216 10425 20244
rect 9824 20204 9830 20216
rect 10413 20213 10425 20216
rect 10459 20244 10471 20247
rect 10965 20247 11023 20253
rect 10965 20244 10977 20247
rect 10459 20216 10977 20244
rect 10459 20213 10471 20216
rect 10413 20207 10471 20213
rect 10965 20213 10977 20216
rect 11011 20213 11023 20247
rect 10965 20207 11023 20213
rect 12986 20204 12992 20256
rect 13044 20244 13050 20256
rect 13170 20244 13176 20256
rect 13044 20216 13176 20244
rect 13044 20204 13050 20216
rect 13170 20204 13176 20216
rect 13228 20244 13234 20256
rect 13541 20247 13599 20253
rect 13541 20244 13553 20247
rect 13228 20216 13553 20244
rect 13228 20204 13234 20216
rect 13541 20213 13553 20216
rect 13587 20244 13599 20247
rect 15764 20244 15792 20284
rect 16206 20244 16212 20256
rect 13587 20216 15792 20244
rect 16167 20216 16212 20244
rect 13587 20213 13599 20216
rect 13541 20207 13599 20213
rect 16206 20204 16212 20216
rect 16264 20204 16270 20256
rect 16316 20244 16344 20284
rect 16390 20272 16396 20324
rect 16448 20312 16454 20324
rect 16577 20315 16635 20321
rect 16577 20312 16589 20315
rect 16448 20284 16589 20312
rect 16448 20272 16454 20284
rect 16577 20281 16589 20284
rect 16623 20312 16635 20315
rect 17221 20315 17279 20321
rect 17221 20312 17233 20315
rect 16623 20284 17233 20312
rect 16623 20281 16635 20284
rect 16577 20275 16635 20281
rect 17221 20281 17233 20284
rect 17267 20281 17279 20315
rect 17221 20275 17279 20281
rect 18064 20244 18092 20343
rect 18138 20340 18144 20392
rect 18196 20380 18202 20392
rect 19153 20383 19211 20389
rect 19153 20380 19165 20383
rect 18196 20352 19165 20380
rect 18196 20340 18202 20352
rect 19153 20349 19165 20352
rect 19199 20380 19211 20383
rect 19242 20380 19248 20392
rect 19199 20352 19248 20380
rect 19199 20349 19211 20352
rect 19153 20343 19211 20349
rect 19242 20340 19248 20352
rect 19300 20340 19306 20392
rect 21545 20383 21603 20389
rect 21545 20380 21557 20383
rect 20640 20352 21557 20380
rect 19061 20315 19119 20321
rect 19061 20281 19073 20315
rect 19107 20312 19119 20315
rect 19420 20315 19478 20321
rect 19420 20312 19432 20315
rect 19107 20284 19432 20312
rect 19107 20281 19119 20284
rect 19061 20275 19119 20281
rect 19420 20281 19432 20284
rect 19466 20312 19478 20315
rect 19518 20312 19524 20324
rect 19466 20284 19524 20312
rect 19466 20281 19478 20284
rect 19420 20275 19478 20281
rect 19518 20272 19524 20284
rect 19576 20312 19582 20324
rect 20530 20312 20536 20324
rect 19576 20284 20536 20312
rect 19576 20272 19582 20284
rect 20530 20272 20536 20284
rect 20588 20272 20594 20324
rect 18601 20247 18659 20253
rect 18601 20244 18613 20247
rect 16316 20216 18613 20244
rect 18601 20213 18613 20216
rect 18647 20213 18659 20247
rect 18601 20207 18659 20213
rect 19334 20204 19340 20256
rect 19392 20244 19398 20256
rect 20640 20244 20668 20352
rect 21545 20349 21557 20352
rect 21591 20380 21603 20383
rect 21634 20380 21640 20392
rect 21591 20352 21640 20380
rect 21591 20349 21603 20352
rect 21545 20343 21603 20349
rect 21634 20340 21640 20352
rect 21692 20380 21698 20392
rect 23477 20383 23535 20389
rect 21692 20352 22140 20380
rect 21692 20340 21698 20352
rect 21358 20272 21364 20324
rect 21416 20312 21422 20324
rect 22112 20321 22140 20352
rect 23477 20349 23489 20383
rect 23523 20380 23535 20383
rect 23566 20380 23572 20392
rect 23523 20352 23572 20380
rect 23523 20349 23535 20352
rect 23477 20343 23535 20349
rect 23566 20340 23572 20352
rect 23624 20380 23630 20392
rect 23934 20380 23940 20392
rect 23624 20352 23940 20380
rect 23624 20340 23630 20352
rect 23934 20340 23940 20352
rect 23992 20380 23998 20392
rect 24121 20383 24179 20389
rect 24121 20380 24133 20383
rect 23992 20352 24133 20380
rect 23992 20340 23998 20352
rect 24121 20349 24133 20352
rect 24167 20349 24179 20383
rect 25222 20380 25228 20392
rect 25183 20352 25228 20380
rect 24121 20343 24179 20349
rect 25222 20340 25228 20352
rect 25280 20380 25286 20392
rect 25777 20383 25835 20389
rect 25777 20380 25789 20383
rect 25280 20352 25789 20380
rect 25280 20340 25286 20352
rect 25777 20349 25789 20352
rect 25823 20349 25835 20383
rect 25777 20343 25835 20349
rect 22005 20315 22063 20321
rect 22005 20312 22017 20315
rect 21416 20284 22017 20312
rect 21416 20272 21422 20284
rect 22005 20281 22017 20284
rect 22051 20281 22063 20315
rect 22005 20275 22063 20281
rect 22097 20315 22155 20321
rect 22097 20281 22109 20315
rect 22143 20312 22155 20315
rect 22186 20312 22192 20324
rect 22143 20284 22192 20312
rect 22143 20281 22155 20284
rect 22097 20275 22155 20281
rect 22186 20272 22192 20284
rect 22244 20272 22250 20324
rect 24029 20315 24087 20321
rect 24029 20312 24041 20315
rect 23032 20284 24041 20312
rect 23032 20256 23060 20284
rect 24029 20281 24041 20284
rect 24075 20281 24087 20315
rect 24029 20275 24087 20281
rect 21634 20244 21640 20256
rect 19392 20216 20668 20244
rect 21595 20216 21640 20244
rect 19392 20204 19398 20216
rect 21634 20204 21640 20216
rect 21692 20204 21698 20256
rect 23014 20244 23020 20256
rect 22975 20216 23020 20244
rect 23014 20204 23020 20216
rect 23072 20204 23078 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 2222 20040 2228 20052
rect 2183 20012 2228 20040
rect 2222 20000 2228 20012
rect 2280 20000 2286 20052
rect 2958 20040 2964 20052
rect 2919 20012 2964 20040
rect 2958 20000 2964 20012
rect 3016 20000 3022 20052
rect 4341 20043 4399 20049
rect 4341 20009 4353 20043
rect 4387 20040 4399 20043
rect 4430 20040 4436 20052
rect 4387 20012 4436 20040
rect 4387 20009 4399 20012
rect 4341 20003 4399 20009
rect 4430 20000 4436 20012
rect 4488 20000 4494 20052
rect 8110 20040 8116 20052
rect 8071 20012 8116 20040
rect 8110 20000 8116 20012
rect 8168 20000 8174 20052
rect 10137 20043 10195 20049
rect 10137 20009 10149 20043
rect 10183 20040 10195 20043
rect 10962 20040 10968 20052
rect 10183 20012 10968 20040
rect 10183 20009 10195 20012
rect 10137 20003 10195 20009
rect 10962 20000 10968 20012
rect 11020 20000 11026 20052
rect 12250 20000 12256 20052
rect 12308 20040 12314 20052
rect 12713 20043 12771 20049
rect 12713 20040 12725 20043
rect 12308 20012 12725 20040
rect 12308 20000 12314 20012
rect 12713 20009 12725 20012
rect 12759 20009 12771 20043
rect 12713 20003 12771 20009
rect 13446 20000 13452 20052
rect 13504 20040 13510 20052
rect 13722 20040 13728 20052
rect 13504 20012 13728 20040
rect 13504 20000 13510 20012
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 13814 20000 13820 20052
rect 13872 20040 13878 20052
rect 14458 20040 14464 20052
rect 13872 20012 14464 20040
rect 13872 20000 13878 20012
rect 14458 20000 14464 20012
rect 14516 20000 14522 20052
rect 15289 20043 15347 20049
rect 15289 20009 15301 20043
rect 15335 20040 15347 20043
rect 15378 20040 15384 20052
rect 15335 20012 15384 20040
rect 15335 20009 15347 20012
rect 15289 20003 15347 20009
rect 15378 20000 15384 20012
rect 15436 20000 15442 20052
rect 15749 20043 15807 20049
rect 15749 20009 15761 20043
rect 15795 20040 15807 20043
rect 15930 20040 15936 20052
rect 15795 20012 15936 20040
rect 15795 20009 15807 20012
rect 15749 20003 15807 20009
rect 15930 20000 15936 20012
rect 15988 20000 15994 20052
rect 16666 20040 16672 20052
rect 16627 20012 16672 20040
rect 16666 20000 16672 20012
rect 16724 20000 16730 20052
rect 17586 20040 17592 20052
rect 17547 20012 17592 20040
rect 17586 20000 17592 20012
rect 17644 20000 17650 20052
rect 19518 20000 19524 20052
rect 19576 20040 19582 20052
rect 19705 20043 19763 20049
rect 19705 20040 19717 20043
rect 19576 20012 19717 20040
rect 19576 20000 19582 20012
rect 19705 20009 19717 20012
rect 19751 20009 19763 20043
rect 19705 20003 19763 20009
rect 20162 20000 20168 20052
rect 20220 20040 20226 20052
rect 20257 20043 20315 20049
rect 20257 20040 20269 20043
rect 20220 20012 20269 20040
rect 20220 20000 20226 20012
rect 20257 20009 20269 20012
rect 20303 20009 20315 20043
rect 20257 20003 20315 20009
rect 20901 20043 20959 20049
rect 20901 20009 20913 20043
rect 20947 20040 20959 20043
rect 23014 20040 23020 20052
rect 20947 20012 23020 20040
rect 20947 20009 20959 20012
rect 20901 20003 20959 20009
rect 23014 20000 23020 20012
rect 23072 20000 23078 20052
rect 24302 20040 24308 20052
rect 24263 20012 24308 20040
rect 24302 20000 24308 20012
rect 24360 20000 24366 20052
rect 4522 19932 4528 19984
rect 4580 19972 4586 19984
rect 4862 19975 4920 19981
rect 4862 19972 4874 19975
rect 4580 19944 4874 19972
rect 4580 19932 4586 19944
rect 4862 19941 4874 19944
rect 4908 19941 4920 19975
rect 4862 19935 4920 19941
rect 7469 19975 7527 19981
rect 7469 19941 7481 19975
rect 7515 19972 7527 19975
rect 7650 19972 7656 19984
rect 7515 19944 7656 19972
rect 7515 19941 7527 19944
rect 7469 19935 7527 19941
rect 7650 19932 7656 19944
rect 7708 19932 7714 19984
rect 12434 19932 12440 19984
rect 12492 19972 12498 19984
rect 13173 19975 13231 19981
rect 13173 19972 13185 19975
rect 12492 19944 12537 19972
rect 12636 19944 13185 19972
rect 12492 19932 12498 19944
rect 1762 19864 1768 19916
rect 1820 19904 1826 19916
rect 2317 19907 2375 19913
rect 2317 19904 2329 19907
rect 1820 19876 2329 19904
rect 1820 19864 1826 19876
rect 2317 19873 2329 19876
rect 2363 19873 2375 19907
rect 2317 19867 2375 19873
rect 3329 19907 3387 19913
rect 3329 19873 3341 19907
rect 3375 19904 3387 19907
rect 3510 19904 3516 19916
rect 3375 19876 3516 19904
rect 3375 19873 3387 19876
rect 3329 19867 3387 19873
rect 3510 19864 3516 19876
rect 3568 19904 3574 19916
rect 4617 19907 4675 19913
rect 4617 19904 4629 19907
rect 3568 19876 4629 19904
rect 3568 19864 3574 19876
rect 4617 19873 4629 19876
rect 4663 19904 4675 19907
rect 6362 19904 6368 19916
rect 4663 19876 6368 19904
rect 4663 19873 4675 19876
rect 4617 19867 4675 19873
rect 6362 19864 6368 19876
rect 6420 19864 6426 19916
rect 6546 19864 6552 19916
rect 6604 19904 6610 19916
rect 9214 19904 9220 19916
rect 6604 19876 9220 19904
rect 6604 19864 6610 19876
rect 9214 19864 9220 19876
rect 9272 19904 9278 19916
rect 9493 19907 9551 19913
rect 9493 19904 9505 19907
rect 9272 19876 9505 19904
rect 9272 19864 9278 19876
rect 9493 19873 9505 19876
rect 9539 19873 9551 19907
rect 9493 19867 9551 19873
rect 9674 19864 9680 19916
rect 9732 19904 9738 19916
rect 10485 19907 10543 19913
rect 10485 19904 10497 19907
rect 9732 19876 10497 19904
rect 9732 19864 9738 19876
rect 10485 19873 10497 19876
rect 10531 19904 10543 19907
rect 11238 19904 11244 19916
rect 10531 19876 11244 19904
rect 10531 19873 10543 19876
rect 10485 19867 10543 19873
rect 11238 19864 11244 19876
rect 11296 19864 11302 19916
rect 12250 19864 12256 19916
rect 12308 19904 12314 19916
rect 12636 19904 12664 19944
rect 13173 19941 13185 19944
rect 13219 19972 13231 19975
rect 14550 19972 14556 19984
rect 13219 19944 14556 19972
rect 13219 19941 13231 19944
rect 13173 19935 13231 19941
rect 14550 19932 14556 19944
rect 14608 19932 14614 19984
rect 15470 19932 15476 19984
rect 15528 19972 15534 19984
rect 16301 19975 16359 19981
rect 16301 19972 16313 19975
rect 15528 19944 16313 19972
rect 15528 19932 15534 19944
rect 16301 19941 16313 19944
rect 16347 19972 16359 19975
rect 16482 19972 16488 19984
rect 16347 19944 16488 19972
rect 16347 19941 16359 19944
rect 16301 19935 16359 19941
rect 16482 19932 16488 19944
rect 16540 19932 16546 19984
rect 20717 19975 20775 19981
rect 20717 19941 20729 19975
rect 20763 19972 20775 19975
rect 22002 19972 22008 19984
rect 20763 19944 22008 19972
rect 20763 19941 20775 19944
rect 20717 19935 20775 19941
rect 22002 19932 22008 19944
rect 22060 19932 22066 19984
rect 22094 19932 22100 19984
rect 22152 19981 22158 19984
rect 22152 19975 22216 19981
rect 22152 19941 22170 19975
rect 22204 19941 22216 19975
rect 22152 19935 22216 19941
rect 22152 19932 22158 19935
rect 12308 19876 12664 19904
rect 13081 19907 13139 19913
rect 12308 19864 12314 19876
rect 13081 19873 13093 19907
rect 13127 19873 13139 19907
rect 13081 19867 13139 19873
rect 2406 19836 2412 19848
rect 2367 19808 2412 19836
rect 2406 19796 2412 19808
rect 2464 19796 2470 19848
rect 3881 19839 3939 19845
rect 3881 19805 3893 19839
rect 3927 19836 3939 19839
rect 4338 19836 4344 19848
rect 3927 19808 4344 19836
rect 3927 19805 3939 19808
rect 3881 19799 3939 19805
rect 4338 19796 4344 19808
rect 4396 19796 4402 19848
rect 6638 19836 6644 19848
rect 6551 19808 6644 19836
rect 6564 19712 6592 19808
rect 6638 19796 6644 19808
rect 6696 19836 6702 19848
rect 7558 19836 7564 19848
rect 6696 19808 7328 19836
rect 7519 19808 7564 19836
rect 6696 19796 6702 19808
rect 7006 19768 7012 19780
rect 6967 19740 7012 19768
rect 7006 19728 7012 19740
rect 7064 19728 7070 19780
rect 7300 19768 7328 19808
rect 7558 19796 7564 19808
rect 7616 19796 7622 19848
rect 7653 19839 7711 19845
rect 7653 19805 7665 19839
rect 7699 19805 7711 19839
rect 7653 19799 7711 19805
rect 8665 19839 8723 19845
rect 8665 19805 8677 19839
rect 8711 19836 8723 19839
rect 8938 19836 8944 19848
rect 8711 19808 8944 19836
rect 8711 19805 8723 19808
rect 8665 19799 8723 19805
rect 7668 19768 7696 19799
rect 8938 19796 8944 19808
rect 8996 19796 9002 19848
rect 10042 19836 10048 19848
rect 9324 19808 10048 19836
rect 7300 19740 7696 19768
rect 9324 19712 9352 19808
rect 10042 19796 10048 19808
rect 10100 19836 10106 19848
rect 10229 19839 10287 19845
rect 10229 19836 10241 19839
rect 10100 19808 10241 19836
rect 10100 19796 10106 19808
rect 10229 19805 10241 19808
rect 10275 19805 10287 19839
rect 10229 19799 10287 19805
rect 12066 19796 12072 19848
rect 12124 19836 12130 19848
rect 13096 19836 13124 19867
rect 14090 19864 14096 19916
rect 14148 19904 14154 19916
rect 15105 19907 15163 19913
rect 15105 19904 15117 19907
rect 14148 19876 15117 19904
rect 14148 19864 14154 19876
rect 15105 19873 15117 19876
rect 15151 19873 15163 19907
rect 15105 19867 15163 19873
rect 15657 19907 15715 19913
rect 15657 19873 15669 19907
rect 15703 19904 15715 19907
rect 15746 19904 15752 19916
rect 15703 19876 15752 19904
rect 15703 19873 15715 19876
rect 15657 19867 15715 19873
rect 15746 19864 15752 19876
rect 15804 19864 15810 19916
rect 16206 19864 16212 19916
rect 16264 19904 16270 19916
rect 16853 19907 16911 19913
rect 16853 19904 16865 19907
rect 16264 19876 16865 19904
rect 16264 19864 16270 19876
rect 16853 19873 16865 19876
rect 16899 19904 16911 19907
rect 17402 19904 17408 19916
rect 16899 19876 17408 19904
rect 16899 19873 16911 19876
rect 16853 19867 16911 19873
rect 17402 19864 17408 19876
rect 17460 19864 17466 19916
rect 18592 19907 18650 19913
rect 18592 19873 18604 19907
rect 18638 19904 18650 19907
rect 19150 19904 19156 19916
rect 18638 19876 19156 19904
rect 18638 19873 18650 19876
rect 18592 19867 18650 19873
rect 19150 19864 19156 19876
rect 19208 19864 19214 19916
rect 24762 19904 24768 19916
rect 24723 19876 24768 19904
rect 24762 19864 24768 19876
rect 24820 19864 24826 19916
rect 13354 19836 13360 19848
rect 12124 19808 13124 19836
rect 13315 19808 13360 19836
rect 12124 19796 12130 19808
rect 13354 19796 13360 19808
rect 13412 19796 13418 19848
rect 13998 19796 14004 19848
rect 14056 19836 14062 19848
rect 15933 19839 15991 19845
rect 15933 19836 15945 19839
rect 14056 19808 15945 19836
rect 14056 19796 14062 19808
rect 15933 19805 15945 19808
rect 15979 19836 15991 19839
rect 16666 19836 16672 19848
rect 15979 19808 16672 19836
rect 15979 19805 15991 19808
rect 15933 19799 15991 19805
rect 16666 19796 16672 19808
rect 16724 19796 16730 19848
rect 17129 19839 17187 19845
rect 17129 19805 17141 19839
rect 17175 19836 17187 19839
rect 17310 19836 17316 19848
rect 17175 19808 17316 19836
rect 17175 19805 17187 19808
rect 17129 19799 17187 19805
rect 17310 19796 17316 19808
rect 17368 19796 17374 19848
rect 18138 19796 18144 19848
rect 18196 19836 18202 19848
rect 18325 19839 18383 19845
rect 18325 19836 18337 19839
rect 18196 19808 18337 19836
rect 18196 19796 18202 19808
rect 18325 19805 18337 19808
rect 18371 19805 18383 19839
rect 18325 19799 18383 19805
rect 21082 19796 21088 19848
rect 21140 19836 21146 19848
rect 21913 19839 21971 19845
rect 21913 19836 21925 19839
rect 21140 19808 21925 19836
rect 21140 19796 21146 19808
rect 21913 19805 21925 19808
rect 21959 19805 21971 19839
rect 24854 19836 24860 19848
rect 24815 19808 24860 19836
rect 21913 19799 21971 19805
rect 24854 19796 24860 19808
rect 24912 19796 24918 19848
rect 24949 19839 25007 19845
rect 24949 19805 24961 19839
rect 24995 19805 25007 19839
rect 24949 19799 25007 19805
rect 22922 19728 22928 19780
rect 22980 19768 22986 19780
rect 23293 19771 23351 19777
rect 23293 19768 23305 19771
rect 22980 19740 23305 19768
rect 22980 19728 22986 19740
rect 23293 19737 23305 19740
rect 23339 19737 23351 19771
rect 23293 19731 23351 19737
rect 23474 19728 23480 19780
rect 23532 19768 23538 19780
rect 24397 19771 24455 19777
rect 24397 19768 24409 19771
rect 23532 19740 24409 19768
rect 23532 19728 23538 19740
rect 24397 19737 24409 19740
rect 24443 19737 24455 19771
rect 24397 19731 24455 19737
rect 24670 19728 24676 19780
rect 24728 19768 24734 19780
rect 24964 19768 24992 19799
rect 24728 19740 24992 19768
rect 24728 19728 24734 19740
rect 1765 19703 1823 19709
rect 1765 19669 1777 19703
rect 1811 19700 1823 19703
rect 1857 19703 1915 19709
rect 1857 19700 1869 19703
rect 1811 19672 1869 19700
rect 1811 19669 1823 19672
rect 1765 19663 1823 19669
rect 1857 19669 1869 19672
rect 1903 19700 1915 19703
rect 2222 19700 2228 19712
rect 1903 19672 2228 19700
rect 1903 19669 1915 19672
rect 1857 19663 1915 19669
rect 2222 19660 2228 19672
rect 2280 19660 2286 19712
rect 5994 19700 6000 19712
rect 5955 19672 6000 19700
rect 5994 19660 6000 19672
rect 6052 19660 6058 19712
rect 6546 19700 6552 19712
rect 6507 19672 6552 19700
rect 6546 19660 6552 19672
rect 6604 19660 6610 19712
rect 7098 19700 7104 19712
rect 7059 19672 7104 19700
rect 7098 19660 7104 19672
rect 7156 19660 7162 19712
rect 9030 19700 9036 19712
rect 8991 19672 9036 19700
rect 9030 19660 9036 19672
rect 9088 19660 9094 19712
rect 9306 19700 9312 19712
rect 9267 19672 9312 19700
rect 9306 19660 9312 19672
rect 9364 19660 9370 19712
rect 10134 19660 10140 19712
rect 10192 19700 10198 19712
rect 11330 19700 11336 19712
rect 10192 19672 11336 19700
rect 10192 19660 10198 19672
rect 11330 19660 11336 19672
rect 11388 19700 11394 19712
rect 11609 19703 11667 19709
rect 11609 19700 11621 19703
rect 11388 19672 11621 19700
rect 11388 19660 11394 19672
rect 11609 19669 11621 19672
rect 11655 19669 11667 19703
rect 14090 19700 14096 19712
rect 14051 19672 14096 19700
rect 11609 19663 11667 19669
rect 14090 19660 14096 19672
rect 14148 19660 14154 19712
rect 14274 19660 14280 19712
rect 14332 19700 14338 19712
rect 14921 19703 14979 19709
rect 14921 19700 14933 19703
rect 14332 19672 14933 19700
rect 14332 19660 14338 19672
rect 14921 19669 14933 19672
rect 14967 19669 14979 19703
rect 14921 19663 14979 19669
rect 18141 19703 18199 19709
rect 18141 19669 18153 19703
rect 18187 19700 18199 19703
rect 18966 19700 18972 19712
rect 18187 19672 18972 19700
rect 18187 19669 18199 19672
rect 18141 19663 18199 19669
rect 18966 19660 18972 19672
rect 19024 19660 19030 19712
rect 20714 19660 20720 19712
rect 20772 19700 20778 19712
rect 21358 19700 21364 19712
rect 20772 19672 21364 19700
rect 20772 19660 20778 19672
rect 21358 19660 21364 19672
rect 21416 19700 21422 19712
rect 21637 19703 21695 19709
rect 21637 19700 21649 19703
rect 21416 19672 21649 19700
rect 21416 19660 21422 19672
rect 21637 19669 21649 19672
rect 21683 19669 21695 19703
rect 23934 19700 23940 19712
rect 23895 19672 23940 19700
rect 21637 19663 21695 19669
rect 23934 19660 23940 19672
rect 23992 19660 23998 19712
rect 25222 19660 25228 19712
rect 25280 19700 25286 19712
rect 25409 19703 25467 19709
rect 25409 19700 25421 19703
rect 25280 19672 25421 19700
rect 25280 19660 25286 19672
rect 25409 19669 25421 19672
rect 25455 19669 25467 19703
rect 25409 19663 25467 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1854 19496 1860 19508
rect 1815 19468 1860 19496
rect 1854 19456 1860 19468
rect 1912 19456 1918 19508
rect 4157 19499 4215 19505
rect 4157 19465 4169 19499
rect 4203 19496 4215 19499
rect 4522 19496 4528 19508
rect 4203 19468 4528 19496
rect 4203 19465 4215 19468
rect 4157 19459 4215 19465
rect 4522 19456 4528 19468
rect 4580 19496 4586 19508
rect 5629 19499 5687 19505
rect 5629 19496 5641 19499
rect 4580 19468 5641 19496
rect 4580 19456 4586 19468
rect 5629 19465 5641 19468
rect 5675 19465 5687 19499
rect 5629 19459 5687 19465
rect 6086 19456 6092 19508
rect 6144 19496 6150 19508
rect 9398 19496 9404 19508
rect 6144 19468 9404 19496
rect 6144 19456 6150 19468
rect 9398 19456 9404 19468
rect 9456 19456 9462 19508
rect 9674 19496 9680 19508
rect 9635 19468 9680 19496
rect 9674 19456 9680 19468
rect 9732 19456 9738 19508
rect 11790 19456 11796 19508
rect 11848 19496 11854 19508
rect 11885 19499 11943 19505
rect 11885 19496 11897 19499
rect 11848 19468 11897 19496
rect 11848 19456 11854 19468
rect 11885 19465 11897 19468
rect 11931 19496 11943 19499
rect 12066 19496 12072 19508
rect 11931 19468 12072 19496
rect 11931 19465 11943 19468
rect 11885 19459 11943 19465
rect 12066 19456 12072 19468
rect 12124 19456 12130 19508
rect 15565 19499 15623 19505
rect 15565 19465 15577 19499
rect 15611 19496 15623 19499
rect 15930 19496 15936 19508
rect 15611 19468 15936 19496
rect 15611 19465 15623 19468
rect 15565 19459 15623 19465
rect 15930 19456 15936 19468
rect 15988 19456 15994 19508
rect 17402 19496 17408 19508
rect 17363 19468 17408 19496
rect 17402 19456 17408 19468
rect 17460 19456 17466 19508
rect 3329 19431 3387 19437
rect 3329 19428 3341 19431
rect 2516 19400 3341 19428
rect 2516 19369 2544 19400
rect 3329 19397 3341 19400
rect 3375 19428 3387 19431
rect 3602 19428 3608 19440
rect 3375 19400 3608 19428
rect 3375 19397 3387 19400
rect 3329 19391 3387 19397
rect 3602 19388 3608 19400
rect 3660 19388 3666 19440
rect 7282 19388 7288 19440
rect 7340 19428 7346 19440
rect 7340 19400 7512 19428
rect 7340 19388 7346 19400
rect 7484 19372 7512 19400
rect 9214 19388 9220 19440
rect 9272 19428 9278 19440
rect 9490 19428 9496 19440
rect 9272 19400 9496 19428
rect 9272 19388 9278 19400
rect 9490 19388 9496 19400
rect 9548 19388 9554 19440
rect 12250 19388 12256 19440
rect 12308 19388 12314 19440
rect 13354 19388 13360 19440
rect 13412 19428 13418 19440
rect 13412 19400 13584 19428
rect 13412 19388 13418 19400
rect 2501 19363 2559 19369
rect 2501 19329 2513 19363
rect 2547 19329 2559 19363
rect 2501 19323 2559 19329
rect 7006 19320 7012 19372
rect 7064 19360 7070 19372
rect 7377 19363 7435 19369
rect 7377 19360 7389 19363
rect 7064 19332 7389 19360
rect 7064 19320 7070 19332
rect 7377 19329 7389 19332
rect 7423 19329 7435 19363
rect 7377 19323 7435 19329
rect 7466 19320 7472 19372
rect 7524 19320 7530 19372
rect 8754 19320 8760 19372
rect 8812 19360 8818 19372
rect 8846 19360 8852 19372
rect 8812 19332 8852 19360
rect 8812 19320 8818 19332
rect 8846 19320 8852 19332
rect 8904 19320 8910 19372
rect 9030 19320 9036 19372
rect 9088 19360 9094 19372
rect 9125 19363 9183 19369
rect 9125 19360 9137 19363
rect 9088 19332 9137 19360
rect 9088 19320 9094 19332
rect 9125 19329 9137 19332
rect 9171 19360 9183 19363
rect 9582 19360 9588 19372
rect 9171 19332 9588 19360
rect 9171 19329 9183 19332
rect 9125 19323 9183 19329
rect 9582 19320 9588 19332
rect 9640 19320 9646 19372
rect 9950 19320 9956 19372
rect 10008 19360 10014 19372
rect 10045 19363 10103 19369
rect 10045 19360 10057 19363
rect 10008 19332 10057 19360
rect 10008 19320 10014 19332
rect 10045 19329 10057 19332
rect 10091 19360 10103 19363
rect 10689 19363 10747 19369
rect 10689 19360 10701 19363
rect 10091 19332 10701 19360
rect 10091 19329 10103 19332
rect 10045 19323 10103 19329
rect 10689 19329 10701 19332
rect 10735 19329 10747 19363
rect 10689 19323 10747 19329
rect 2314 19292 2320 19304
rect 2275 19264 2320 19292
rect 2314 19252 2320 19264
rect 2372 19252 2378 19304
rect 2406 19252 2412 19304
rect 2464 19292 2470 19304
rect 2590 19292 2596 19304
rect 2464 19264 2596 19292
rect 2464 19252 2470 19264
rect 2590 19252 2596 19264
rect 2648 19292 2654 19304
rect 2869 19295 2927 19301
rect 2869 19292 2881 19295
rect 2648 19264 2881 19292
rect 2648 19252 2654 19264
rect 2869 19261 2881 19264
rect 2915 19261 2927 19295
rect 2869 19255 2927 19261
rect 4154 19252 4160 19304
rect 4212 19292 4218 19304
rect 4249 19295 4307 19301
rect 4249 19292 4261 19295
rect 4212 19264 4261 19292
rect 4212 19252 4218 19264
rect 4249 19261 4261 19264
rect 4295 19261 4307 19295
rect 6178 19292 6184 19304
rect 6139 19264 6184 19292
rect 4249 19255 4307 19261
rect 6178 19252 6184 19264
rect 6236 19252 6242 19304
rect 7098 19252 7104 19304
rect 7156 19292 7162 19304
rect 7193 19295 7251 19301
rect 7193 19292 7205 19295
rect 7156 19264 7205 19292
rect 7156 19252 7162 19264
rect 7193 19261 7205 19264
rect 7239 19261 7251 19295
rect 7193 19255 7251 19261
rect 12066 19252 12072 19304
rect 12124 19292 12130 19304
rect 12161 19295 12219 19301
rect 12161 19292 12173 19295
rect 12124 19264 12173 19292
rect 12124 19252 12130 19264
rect 12161 19261 12173 19264
rect 12207 19292 12219 19295
rect 12268 19292 12296 19388
rect 13446 19360 13452 19372
rect 13407 19332 13452 19360
rect 13446 19320 13452 19332
rect 13504 19320 13510 19372
rect 13556 19360 13584 19400
rect 16114 19388 16120 19440
rect 16172 19428 16178 19440
rect 19150 19428 19156 19440
rect 16172 19400 16620 19428
rect 19111 19400 19156 19428
rect 16172 19388 16178 19400
rect 13556 19332 13768 19360
rect 12207 19264 12296 19292
rect 13740 19292 13768 19332
rect 14550 19320 14556 19372
rect 14608 19360 14614 19372
rect 15013 19363 15071 19369
rect 15013 19360 15025 19363
rect 14608 19332 15025 19360
rect 14608 19320 14614 19332
rect 15013 19329 15025 19332
rect 15059 19329 15071 19363
rect 16482 19360 16488 19372
rect 16443 19332 16488 19360
rect 15013 19323 15071 19329
rect 16482 19320 16488 19332
rect 16540 19320 16546 19372
rect 16592 19369 16620 19400
rect 19150 19388 19156 19400
rect 19208 19388 19214 19440
rect 24578 19388 24584 19440
rect 24636 19428 24642 19440
rect 24854 19428 24860 19440
rect 24636 19400 24860 19428
rect 24636 19388 24642 19400
rect 24854 19388 24860 19400
rect 24912 19388 24918 19440
rect 16577 19363 16635 19369
rect 16577 19329 16589 19363
rect 16623 19329 16635 19363
rect 16577 19323 16635 19329
rect 18693 19363 18751 19369
rect 18693 19329 18705 19363
rect 18739 19360 18751 19363
rect 18966 19360 18972 19372
rect 18739 19332 18972 19360
rect 18739 19329 18751 19332
rect 18693 19323 18751 19329
rect 18966 19320 18972 19332
rect 19024 19320 19030 19372
rect 22922 19360 22928 19372
rect 22112 19332 22928 19360
rect 14277 19295 14335 19301
rect 14277 19292 14289 19295
rect 13740 19264 14289 19292
rect 12207 19261 12219 19264
rect 12161 19255 12219 19261
rect 14277 19261 14289 19264
rect 14323 19261 14335 19295
rect 14277 19255 14335 19261
rect 14458 19252 14464 19304
rect 14516 19292 14522 19304
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 14516 19264 14933 19292
rect 14516 19252 14522 19264
rect 14921 19261 14933 19264
rect 14967 19261 14979 19295
rect 17126 19292 17132 19304
rect 17087 19264 17132 19292
rect 14921 19255 14979 19261
rect 17126 19252 17132 19264
rect 17184 19252 17190 19304
rect 19426 19252 19432 19304
rect 19484 19252 19490 19304
rect 19610 19292 19616 19304
rect 19571 19264 19616 19292
rect 19610 19252 19616 19264
rect 19668 19292 19674 19304
rect 20349 19295 20407 19301
rect 20349 19292 20361 19295
rect 19668 19264 20361 19292
rect 19668 19252 19674 19264
rect 20349 19261 20361 19264
rect 20395 19261 20407 19295
rect 21082 19292 21088 19304
rect 21043 19264 21088 19292
rect 20349 19255 20407 19261
rect 21082 19252 21088 19264
rect 21140 19252 21146 19304
rect 22112 19292 22140 19332
rect 22922 19320 22928 19332
rect 22980 19320 22986 19372
rect 23934 19320 23940 19372
rect 23992 19360 23998 19372
rect 24213 19363 24271 19369
rect 24213 19360 24225 19363
rect 23992 19332 24225 19360
rect 23992 19320 23998 19332
rect 24213 19329 24225 19332
rect 24259 19329 24271 19363
rect 24213 19323 24271 19329
rect 24670 19320 24676 19372
rect 24728 19360 24734 19372
rect 24728 19332 24808 19360
rect 24728 19320 24734 19332
rect 23474 19292 23480 19304
rect 21468 19264 22140 19292
rect 23387 19264 23480 19292
rect 2222 19224 2228 19236
rect 2183 19196 2228 19224
rect 2222 19184 2228 19196
rect 2280 19184 2286 19236
rect 2332 19224 2360 19252
rect 4522 19233 4528 19236
rect 3605 19227 3663 19233
rect 3605 19224 3617 19227
rect 2332 19196 3617 19224
rect 3605 19193 3617 19196
rect 3651 19193 3663 19227
rect 4516 19224 4528 19233
rect 4483 19196 4528 19224
rect 3605 19187 3663 19193
rect 4516 19187 4528 19196
rect 4522 19184 4528 19187
rect 4580 19184 4586 19236
rect 6196 19224 6224 19252
rect 7285 19227 7343 19233
rect 7285 19224 7297 19227
rect 6196 19196 7297 19224
rect 7285 19193 7297 19196
rect 7331 19193 7343 19227
rect 7285 19187 7343 19193
rect 8481 19227 8539 19233
rect 8481 19193 8493 19227
rect 8527 19224 8539 19227
rect 10505 19227 10563 19233
rect 8527 19196 9076 19224
rect 8527 19193 8539 19196
rect 8481 19187 8539 19193
rect 9048 19168 9076 19196
rect 10505 19193 10517 19227
rect 10551 19224 10563 19227
rect 11241 19227 11299 19233
rect 11241 19224 11253 19227
rect 10551 19196 11253 19224
rect 10551 19193 10563 19196
rect 10505 19187 10563 19193
rect 11241 19193 11253 19196
rect 11287 19224 11299 19227
rect 12434 19224 12440 19236
rect 11287 19196 12440 19224
rect 11287 19193 11299 19196
rect 11241 19187 11299 19193
rect 12434 19184 12440 19196
rect 12492 19184 12498 19236
rect 12713 19227 12771 19233
rect 12713 19193 12725 19227
rect 12759 19224 12771 19227
rect 13265 19227 13323 19233
rect 13265 19224 13277 19227
rect 12759 19196 13277 19224
rect 12759 19193 12771 19196
rect 12713 19187 12771 19193
rect 13265 19193 13277 19196
rect 13311 19224 13323 19227
rect 13538 19224 13544 19236
rect 13311 19196 13544 19224
rect 13311 19193 13323 19196
rect 13265 19187 13323 19193
rect 13538 19184 13544 19196
rect 13596 19184 13602 19236
rect 17678 19184 17684 19236
rect 17736 19224 17742 19236
rect 17773 19227 17831 19233
rect 17773 19224 17785 19227
rect 17736 19196 17785 19224
rect 17736 19184 17742 19196
rect 17773 19193 17785 19196
rect 17819 19224 17831 19227
rect 18506 19224 18512 19236
rect 17819 19196 18512 19224
rect 17819 19193 17831 19196
rect 17773 19187 17831 19193
rect 18506 19184 18512 19196
rect 18564 19184 18570 19236
rect 19444 19224 19472 19252
rect 19889 19227 19947 19233
rect 19889 19224 19901 19227
rect 19444 19196 19901 19224
rect 19889 19193 19901 19196
rect 19935 19193 19947 19227
rect 19889 19187 19947 19193
rect 20993 19227 21051 19233
rect 20993 19193 21005 19227
rect 21039 19224 21051 19227
rect 21330 19227 21388 19233
rect 21330 19224 21342 19227
rect 21039 19196 21342 19224
rect 21039 19193 21051 19196
rect 20993 19187 21051 19193
rect 21330 19193 21342 19196
rect 21376 19224 21388 19227
rect 21468 19224 21496 19264
rect 23474 19252 23480 19264
rect 23532 19292 23538 19304
rect 24780 19292 24808 19332
rect 25222 19292 25228 19304
rect 23532 19264 24256 19292
rect 24780 19264 24900 19292
rect 25183 19264 25228 19292
rect 23532 19252 23538 19264
rect 21376 19196 21496 19224
rect 21376 19193 21388 19196
rect 21330 19187 21388 19193
rect 21726 19184 21732 19236
rect 21784 19224 21790 19236
rect 23109 19227 23167 19233
rect 23109 19224 23121 19227
rect 21784 19196 23121 19224
rect 21784 19184 21790 19196
rect 23109 19193 23121 19196
rect 23155 19224 23167 19227
rect 24121 19227 24179 19233
rect 24121 19224 24133 19227
rect 23155 19196 24133 19224
rect 23155 19193 23167 19196
rect 23109 19187 23167 19193
rect 24121 19193 24133 19196
rect 24167 19193 24179 19227
rect 24121 19187 24179 19193
rect 1765 19159 1823 19165
rect 1765 19125 1777 19159
rect 1811 19156 1823 19159
rect 1854 19156 1860 19168
rect 1811 19128 1860 19156
rect 1811 19125 1823 19128
rect 1765 19119 1823 19125
rect 1854 19116 1860 19128
rect 1912 19116 1918 19168
rect 6546 19156 6552 19168
rect 6507 19128 6552 19156
rect 6546 19116 6552 19128
rect 6604 19116 6610 19168
rect 6730 19116 6736 19168
rect 6788 19156 6794 19168
rect 6825 19159 6883 19165
rect 6825 19156 6837 19159
rect 6788 19128 6837 19156
rect 6788 19116 6794 19128
rect 6825 19125 6837 19128
rect 6871 19125 6883 19159
rect 6825 19119 6883 19125
rect 7742 19116 7748 19168
rect 7800 19156 7806 19168
rect 7837 19159 7895 19165
rect 7837 19156 7849 19159
rect 7800 19128 7849 19156
rect 7800 19116 7806 19128
rect 7837 19125 7849 19128
rect 7883 19125 7895 19159
rect 8570 19156 8576 19168
rect 8531 19128 8576 19156
rect 7837 19119 7895 19125
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 8938 19156 8944 19168
rect 8899 19128 8944 19156
rect 8938 19116 8944 19128
rect 8996 19116 9002 19168
rect 9030 19116 9036 19168
rect 9088 19156 9094 19168
rect 9088 19128 9133 19156
rect 9088 19116 9094 19128
rect 10042 19116 10048 19168
rect 10100 19156 10106 19168
rect 10137 19159 10195 19165
rect 10137 19156 10149 19159
rect 10100 19128 10149 19156
rect 10100 19116 10106 19128
rect 10137 19125 10149 19128
rect 10183 19125 10195 19159
rect 10137 19119 10195 19125
rect 10597 19159 10655 19165
rect 10597 19125 10609 19159
rect 10643 19156 10655 19159
rect 10962 19156 10968 19168
rect 10643 19128 10968 19156
rect 10643 19125 10655 19128
rect 10597 19119 10655 19125
rect 10962 19116 10968 19128
rect 11020 19116 11026 19168
rect 12802 19116 12808 19168
rect 12860 19156 12866 19168
rect 12897 19159 12955 19165
rect 12897 19156 12909 19159
rect 12860 19128 12909 19156
rect 12860 19116 12866 19128
rect 12897 19125 12909 19128
rect 12943 19125 12955 19159
rect 12897 19119 12955 19125
rect 13357 19159 13415 19165
rect 13357 19125 13369 19159
rect 13403 19156 13415 19159
rect 13906 19156 13912 19168
rect 13403 19128 13912 19156
rect 13403 19125 13415 19128
rect 13357 19119 13415 19125
rect 13906 19116 13912 19128
rect 13964 19116 13970 19168
rect 14458 19156 14464 19168
rect 14419 19128 14464 19156
rect 14458 19116 14464 19128
rect 14516 19116 14522 19168
rect 14826 19156 14832 19168
rect 14787 19128 14832 19156
rect 14826 19116 14832 19128
rect 14884 19116 14890 19168
rect 15746 19116 15752 19168
rect 15804 19156 15810 19168
rect 15841 19159 15899 19165
rect 15841 19156 15853 19159
rect 15804 19128 15853 19156
rect 15804 19116 15810 19128
rect 15841 19125 15853 19128
rect 15887 19125 15899 19159
rect 15841 19119 15899 19125
rect 16025 19159 16083 19165
rect 16025 19125 16037 19159
rect 16071 19156 16083 19159
rect 16298 19156 16304 19168
rect 16071 19128 16304 19156
rect 16071 19125 16083 19128
rect 16025 19119 16083 19125
rect 16298 19116 16304 19128
rect 16356 19116 16362 19168
rect 16393 19159 16451 19165
rect 16393 19125 16405 19159
rect 16439 19156 16451 19159
rect 16850 19156 16856 19168
rect 16439 19128 16856 19156
rect 16439 19125 16451 19128
rect 16393 19119 16451 19125
rect 16850 19116 16856 19128
rect 16908 19116 16914 19168
rect 18046 19156 18052 19168
rect 18007 19128 18052 19156
rect 18046 19116 18052 19128
rect 18104 19116 18110 19168
rect 18414 19156 18420 19168
rect 18375 19128 18420 19156
rect 18414 19116 18420 19128
rect 18472 19116 18478 19168
rect 19521 19159 19579 19165
rect 19521 19125 19533 19159
rect 19567 19156 19579 19159
rect 20162 19156 20168 19168
rect 19567 19128 20168 19156
rect 19567 19125 19579 19128
rect 19521 19119 19579 19125
rect 20162 19116 20168 19128
rect 20220 19116 20226 19168
rect 22462 19156 22468 19168
rect 22423 19128 22468 19156
rect 22462 19116 22468 19128
rect 22520 19116 22526 19168
rect 23658 19156 23664 19168
rect 23619 19128 23664 19156
rect 23658 19116 23664 19128
rect 23716 19116 23722 19168
rect 24029 19159 24087 19165
rect 24029 19125 24041 19159
rect 24075 19156 24087 19159
rect 24228 19156 24256 19264
rect 24872 19224 24900 19264
rect 25222 19252 25228 19264
rect 25280 19252 25286 19304
rect 25777 19227 25835 19233
rect 25777 19224 25789 19227
rect 24872 19196 25789 19224
rect 25777 19193 25789 19196
rect 25823 19193 25835 19227
rect 25777 19187 25835 19193
rect 24302 19156 24308 19168
rect 24075 19128 24308 19156
rect 24075 19125 24087 19128
rect 24029 19119 24087 19125
rect 24302 19116 24308 19128
rect 24360 19116 24366 19168
rect 24578 19116 24584 19168
rect 24636 19156 24642 19168
rect 24673 19159 24731 19165
rect 24673 19156 24685 19159
rect 24636 19128 24685 19156
rect 24636 19116 24642 19128
rect 24673 19125 24685 19128
rect 24719 19125 24731 19159
rect 24673 19119 24731 19125
rect 24762 19116 24768 19168
rect 24820 19156 24826 19168
rect 25133 19159 25191 19165
rect 25133 19156 25145 19159
rect 24820 19128 25145 19156
rect 24820 19116 24826 19128
rect 25133 19125 25145 19128
rect 25179 19156 25191 19159
rect 25222 19156 25228 19168
rect 25179 19128 25228 19156
rect 25179 19125 25191 19128
rect 25133 19119 25191 19125
rect 25222 19116 25228 19128
rect 25280 19116 25286 19168
rect 25409 19159 25467 19165
rect 25409 19125 25421 19159
rect 25455 19156 25467 19159
rect 25498 19156 25504 19168
rect 25455 19128 25504 19156
rect 25455 19125 25467 19128
rect 25409 19119 25467 19125
rect 25498 19116 25504 19128
rect 25556 19116 25562 19168
rect 26142 19156 26148 19168
rect 26103 19128 26148 19156
rect 26142 19116 26148 19128
rect 26200 19116 26206 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 2041 18955 2099 18961
rect 2041 18921 2053 18955
rect 2087 18952 2099 18955
rect 2314 18952 2320 18964
rect 2087 18924 2320 18952
rect 2087 18921 2099 18924
rect 2041 18915 2099 18921
rect 2314 18912 2320 18924
rect 2372 18912 2378 18964
rect 2498 18952 2504 18964
rect 2459 18924 2504 18952
rect 2498 18912 2504 18924
rect 2556 18912 2562 18964
rect 4341 18955 4399 18961
rect 4341 18921 4353 18955
rect 4387 18952 4399 18955
rect 4522 18952 4528 18964
rect 4387 18924 4528 18952
rect 4387 18921 4399 18924
rect 4341 18915 4399 18921
rect 4522 18912 4528 18924
rect 4580 18952 4586 18964
rect 5350 18952 5356 18964
rect 4580 18924 5356 18952
rect 4580 18912 4586 18924
rect 5350 18912 5356 18924
rect 5408 18952 5414 18964
rect 6089 18955 6147 18961
rect 6089 18952 6101 18955
rect 5408 18924 6101 18952
rect 5408 18912 5414 18924
rect 6089 18921 6101 18924
rect 6135 18952 6147 18955
rect 6822 18952 6828 18964
rect 6135 18924 6828 18952
rect 6135 18921 6147 18924
rect 6089 18915 6147 18921
rect 6822 18912 6828 18924
rect 6880 18912 6886 18964
rect 7098 18912 7104 18964
rect 7156 18952 7162 18964
rect 7469 18955 7527 18961
rect 7469 18952 7481 18955
rect 7156 18924 7481 18952
rect 7156 18912 7162 18924
rect 7469 18921 7481 18924
rect 7515 18921 7527 18955
rect 8478 18952 8484 18964
rect 8439 18924 8484 18952
rect 7469 18915 7527 18921
rect 8478 18912 8484 18924
rect 8536 18912 8542 18964
rect 8662 18912 8668 18964
rect 8720 18952 8726 18964
rect 9582 18952 9588 18964
rect 8720 18924 9588 18952
rect 8720 18912 8726 18924
rect 9582 18912 9588 18924
rect 9640 18912 9646 18964
rect 9674 18912 9680 18964
rect 9732 18952 9738 18964
rect 11238 18952 11244 18964
rect 9732 18924 11244 18952
rect 9732 18912 9738 18924
rect 11238 18912 11244 18924
rect 11296 18912 11302 18964
rect 11790 18912 11796 18964
rect 11848 18952 11854 18964
rect 12066 18952 12072 18964
rect 11848 18924 12072 18952
rect 11848 18912 11854 18924
rect 12066 18912 12072 18924
rect 12124 18912 12130 18964
rect 12894 18912 12900 18964
rect 12952 18952 12958 18964
rect 13265 18955 13323 18961
rect 13265 18952 13277 18955
rect 12952 18924 13277 18952
rect 12952 18912 12958 18924
rect 13265 18921 13277 18924
rect 13311 18921 13323 18955
rect 13265 18915 13323 18921
rect 15289 18955 15347 18961
rect 15289 18921 15301 18955
rect 15335 18952 15347 18955
rect 15562 18952 15568 18964
rect 15335 18924 15568 18952
rect 15335 18921 15347 18924
rect 15289 18915 15347 18921
rect 15562 18912 15568 18924
rect 15620 18912 15626 18964
rect 16114 18912 16120 18964
rect 16172 18952 16178 18964
rect 16301 18955 16359 18961
rect 16301 18952 16313 18955
rect 16172 18924 16313 18952
rect 16172 18912 16178 18924
rect 16301 18921 16313 18924
rect 16347 18921 16359 18955
rect 16301 18915 16359 18921
rect 16945 18955 17003 18961
rect 16945 18921 16957 18955
rect 16991 18952 17003 18955
rect 17862 18952 17868 18964
rect 16991 18924 17868 18952
rect 16991 18921 17003 18924
rect 16945 18915 17003 18921
rect 17862 18912 17868 18924
rect 17920 18912 17926 18964
rect 18141 18955 18199 18961
rect 18141 18921 18153 18955
rect 18187 18952 18199 18955
rect 18414 18952 18420 18964
rect 18187 18924 18420 18952
rect 18187 18921 18199 18924
rect 18141 18915 18199 18921
rect 18414 18912 18420 18924
rect 18472 18912 18478 18964
rect 18598 18912 18604 18964
rect 18656 18952 18662 18964
rect 18969 18955 19027 18961
rect 18969 18952 18981 18955
rect 18656 18924 18981 18952
rect 18656 18912 18662 18924
rect 18969 18921 18981 18924
rect 19015 18952 19027 18955
rect 19058 18952 19064 18964
rect 19015 18924 19064 18952
rect 19015 18921 19027 18924
rect 18969 18915 19027 18921
rect 19058 18912 19064 18924
rect 19116 18912 19122 18964
rect 19334 18912 19340 18964
rect 19392 18952 19398 18964
rect 20073 18955 20131 18961
rect 20073 18952 20085 18955
rect 19392 18924 20085 18952
rect 19392 18912 19398 18924
rect 20073 18921 20085 18924
rect 20119 18952 20131 18955
rect 21082 18952 21088 18964
rect 20119 18924 21088 18952
rect 20119 18921 20131 18924
rect 20073 18915 20131 18921
rect 21082 18912 21088 18924
rect 21140 18912 21146 18964
rect 21174 18912 21180 18964
rect 21232 18952 21238 18964
rect 21269 18955 21327 18961
rect 21269 18952 21281 18955
rect 21232 18924 21281 18952
rect 21232 18912 21238 18924
rect 21269 18921 21281 18924
rect 21315 18921 21327 18955
rect 22002 18952 22008 18964
rect 21963 18924 22008 18952
rect 21269 18915 21327 18921
rect 22002 18912 22008 18924
rect 22060 18912 22066 18964
rect 22741 18955 22799 18961
rect 22741 18921 22753 18955
rect 22787 18952 22799 18955
rect 23290 18952 23296 18964
rect 22787 18924 23296 18952
rect 22787 18921 22799 18924
rect 22741 18915 22799 18921
rect 23290 18912 23296 18924
rect 23348 18912 23354 18964
rect 25041 18955 25099 18961
rect 25041 18921 25053 18955
rect 25087 18952 25099 18955
rect 25130 18952 25136 18964
rect 25087 18924 25136 18952
rect 25087 18921 25099 18924
rect 25041 18915 25099 18921
rect 25130 18912 25136 18924
rect 25188 18912 25194 18964
rect 1949 18887 2007 18893
rect 1949 18853 1961 18887
rect 1995 18884 2007 18887
rect 2130 18884 2136 18896
rect 1995 18856 2136 18884
rect 1995 18853 2007 18856
rect 1949 18847 2007 18853
rect 2130 18844 2136 18856
rect 2188 18844 2194 18896
rect 3513 18887 3571 18893
rect 3513 18853 3525 18887
rect 3559 18884 3571 18887
rect 3602 18884 3608 18896
rect 3559 18856 3608 18884
rect 3559 18853 3571 18856
rect 3513 18847 3571 18853
rect 3602 18844 3608 18856
rect 3660 18884 3666 18896
rect 3881 18887 3939 18893
rect 3881 18884 3893 18887
rect 3660 18856 3893 18884
rect 3660 18844 3666 18856
rect 3881 18853 3893 18856
rect 3927 18884 3939 18887
rect 4154 18884 4160 18896
rect 3927 18856 4160 18884
rect 3927 18853 3939 18856
rect 3881 18847 3939 18853
rect 4154 18844 4160 18856
rect 4212 18884 4218 18896
rect 6362 18884 6368 18896
rect 4212 18856 6368 18884
rect 4212 18844 4218 18856
rect 2406 18816 2412 18828
rect 2367 18788 2412 18816
rect 2406 18776 2412 18788
rect 2464 18776 2470 18828
rect 4724 18825 4752 18856
rect 6362 18844 6368 18856
rect 6420 18884 6426 18896
rect 6641 18887 6699 18893
rect 6641 18884 6653 18887
rect 6420 18856 6653 18884
rect 6420 18844 6426 18856
rect 6641 18853 6653 18856
rect 6687 18853 6699 18887
rect 6641 18847 6699 18853
rect 7193 18887 7251 18893
rect 7193 18853 7205 18887
rect 7239 18884 7251 18887
rect 7558 18884 7564 18896
rect 7239 18856 7564 18884
rect 7239 18853 7251 18856
rect 7193 18847 7251 18853
rect 4709 18819 4767 18825
rect 4709 18785 4721 18819
rect 4755 18785 4767 18819
rect 4709 18779 4767 18785
rect 4976 18819 5034 18825
rect 4976 18785 4988 18819
rect 5022 18816 5034 18819
rect 5258 18816 5264 18828
rect 5022 18788 5264 18816
rect 5022 18785 5034 18788
rect 4976 18779 5034 18785
rect 5258 18776 5264 18788
rect 5316 18816 5322 18828
rect 6546 18816 6552 18828
rect 5316 18788 6552 18816
rect 5316 18776 5322 18788
rect 6546 18776 6552 18788
rect 6604 18776 6610 18828
rect 6656 18816 6684 18847
rect 7558 18844 7564 18856
rect 7616 18844 7622 18896
rect 8110 18844 8116 18896
rect 8168 18884 8174 18896
rect 8389 18887 8447 18893
rect 8389 18884 8401 18887
rect 8168 18856 8401 18884
rect 8168 18844 8174 18856
rect 8389 18853 8401 18856
rect 8435 18884 8447 18887
rect 9398 18884 9404 18896
rect 8435 18856 9404 18884
rect 8435 18853 8447 18856
rect 8389 18847 8447 18853
rect 9398 18844 9404 18856
rect 9456 18844 9462 18896
rect 10134 18844 10140 18896
rect 10192 18884 10198 18896
rect 10566 18887 10624 18893
rect 10566 18884 10578 18887
rect 10192 18856 10578 18884
rect 10192 18844 10198 18856
rect 10566 18853 10578 18856
rect 10612 18853 10624 18887
rect 10566 18847 10624 18853
rect 12250 18844 12256 18896
rect 12308 18884 12314 18896
rect 13173 18887 13231 18893
rect 13173 18884 13185 18887
rect 12308 18856 13185 18884
rect 12308 18844 12314 18856
rect 13173 18853 13185 18856
rect 13219 18853 13231 18887
rect 13173 18847 13231 18853
rect 7837 18819 7895 18825
rect 7837 18816 7849 18819
rect 6656 18788 7849 18816
rect 7837 18785 7849 18788
rect 7883 18785 7895 18819
rect 7837 18779 7895 18785
rect 8846 18776 8852 18828
rect 8904 18816 8910 18828
rect 9306 18816 9312 18828
rect 8904 18788 9312 18816
rect 8904 18776 8910 18788
rect 9306 18776 9312 18788
rect 9364 18816 9370 18828
rect 10321 18819 10379 18825
rect 10321 18816 10333 18819
rect 9364 18788 10333 18816
rect 9364 18776 9370 18788
rect 10321 18785 10333 18788
rect 10367 18785 10379 18819
rect 10321 18779 10379 18785
rect 13188 18760 13216 18847
rect 14734 18844 14740 18896
rect 14792 18884 14798 18896
rect 15749 18887 15807 18893
rect 15749 18884 15761 18887
rect 14792 18856 15761 18884
rect 14792 18844 14798 18856
rect 15749 18853 15761 18856
rect 15795 18853 15807 18887
rect 15749 18847 15807 18853
rect 16761 18887 16819 18893
rect 16761 18853 16773 18887
rect 16807 18884 16819 18887
rect 16850 18884 16856 18896
rect 16807 18856 16856 18884
rect 16807 18853 16819 18856
rect 16761 18847 16819 18853
rect 16850 18844 16856 18856
rect 16908 18844 16914 18896
rect 18506 18844 18512 18896
rect 18564 18884 18570 18896
rect 21100 18884 21128 18912
rect 23477 18887 23535 18893
rect 23477 18884 23489 18887
rect 18564 18856 20852 18884
rect 21100 18856 23489 18884
rect 18564 18844 18570 18856
rect 15657 18819 15715 18825
rect 15657 18785 15669 18819
rect 15703 18785 15715 18819
rect 15657 18779 15715 18785
rect 2590 18748 2596 18760
rect 2551 18720 2596 18748
rect 2590 18708 2596 18720
rect 2648 18748 2654 18760
rect 2774 18748 2780 18760
rect 2648 18720 2780 18748
rect 2648 18708 2654 18720
rect 2774 18708 2780 18720
rect 2832 18708 2838 18760
rect 8665 18751 8723 18757
rect 8665 18717 8677 18751
rect 8711 18748 8723 18751
rect 9214 18748 9220 18760
rect 8711 18720 9220 18748
rect 8711 18717 8723 18720
rect 8665 18711 8723 18717
rect 9214 18708 9220 18720
rect 9272 18708 9278 18760
rect 13170 18708 13176 18760
rect 13228 18708 13234 18760
rect 13262 18708 13268 18760
rect 13320 18748 13326 18760
rect 13357 18751 13415 18757
rect 13357 18748 13369 18751
rect 13320 18720 13369 18748
rect 13320 18708 13326 18720
rect 13357 18717 13369 18720
rect 13403 18717 13415 18751
rect 13357 18711 13415 18717
rect 14185 18751 14243 18757
rect 14185 18717 14197 18751
rect 14231 18748 14243 18751
rect 14826 18748 14832 18760
rect 14231 18720 14832 18748
rect 14231 18717 14243 18720
rect 14185 18711 14243 18717
rect 14826 18708 14832 18720
rect 14884 18708 14890 18760
rect 2130 18640 2136 18692
rect 2188 18680 2194 18692
rect 3602 18680 3608 18692
rect 2188 18652 3608 18680
rect 2188 18640 2194 18652
rect 3602 18640 3608 18652
rect 3660 18640 3666 18692
rect 12805 18683 12863 18689
rect 12805 18649 12817 18683
rect 12851 18680 12863 18683
rect 15013 18683 15071 18689
rect 15013 18680 15025 18683
rect 12851 18652 15025 18680
rect 12851 18649 12863 18652
rect 12805 18643 12863 18649
rect 15013 18649 15025 18652
rect 15059 18680 15071 18683
rect 15672 18680 15700 18779
rect 16574 18776 16580 18828
rect 16632 18816 16638 18828
rect 17313 18819 17371 18825
rect 17313 18816 17325 18819
rect 16632 18788 17325 18816
rect 16632 18776 16638 18788
rect 17313 18785 17325 18788
rect 17359 18785 17371 18819
rect 17313 18779 17371 18785
rect 17405 18819 17463 18825
rect 17405 18785 17417 18819
rect 17451 18816 17463 18819
rect 17862 18816 17868 18828
rect 17451 18788 17868 18816
rect 17451 18785 17463 18788
rect 17405 18779 17463 18785
rect 17862 18776 17868 18788
rect 17920 18776 17926 18828
rect 18877 18819 18935 18825
rect 18877 18785 18889 18819
rect 18923 18816 18935 18819
rect 19886 18816 19892 18828
rect 18923 18788 19892 18816
rect 18923 18785 18935 18788
rect 18877 18779 18935 18785
rect 15933 18751 15991 18757
rect 15933 18717 15945 18751
rect 15979 18748 15991 18751
rect 16022 18748 16028 18760
rect 15979 18720 16028 18748
rect 15979 18717 15991 18720
rect 15933 18711 15991 18717
rect 16022 18708 16028 18720
rect 16080 18708 16086 18760
rect 17494 18748 17500 18760
rect 17455 18720 17500 18748
rect 17494 18708 17500 18720
rect 17552 18708 17558 18760
rect 17770 18708 17776 18760
rect 17828 18748 17834 18760
rect 18892 18748 18920 18779
rect 19886 18776 19892 18788
rect 19944 18776 19950 18828
rect 20162 18776 20168 18828
rect 20220 18816 20226 18828
rect 20257 18819 20315 18825
rect 20257 18816 20269 18819
rect 20220 18788 20269 18816
rect 20220 18776 20226 18788
rect 20257 18785 20269 18788
rect 20303 18785 20315 18819
rect 20824 18816 20852 18856
rect 23477 18853 23489 18856
rect 23523 18884 23535 18887
rect 23566 18884 23572 18896
rect 23523 18856 23572 18884
rect 23523 18853 23535 18856
rect 23477 18847 23535 18853
rect 23566 18844 23572 18856
rect 23624 18884 23630 18896
rect 23624 18856 23704 18884
rect 23624 18844 23630 18856
rect 21358 18816 21364 18828
rect 20824 18788 21364 18816
rect 20257 18779 20315 18785
rect 17828 18720 18920 18748
rect 17828 18708 17834 18720
rect 18966 18708 18972 18760
rect 19024 18748 19030 18760
rect 19061 18751 19119 18757
rect 19061 18748 19073 18751
rect 19024 18720 19073 18748
rect 19024 18708 19030 18720
rect 19061 18717 19073 18720
rect 19107 18717 19119 18751
rect 19904 18748 19932 18776
rect 21008 18760 21036 18788
rect 21358 18776 21364 18788
rect 21416 18816 21422 18828
rect 21726 18816 21732 18828
rect 21416 18788 21732 18816
rect 21416 18776 21422 18788
rect 21726 18776 21732 18788
rect 21784 18776 21790 18828
rect 22554 18816 22560 18828
rect 22515 18788 22560 18816
rect 22554 18776 22560 18788
rect 22612 18776 22618 18828
rect 23676 18825 23704 18856
rect 23661 18819 23719 18825
rect 23661 18785 23673 18819
rect 23707 18785 23719 18819
rect 23661 18779 23719 18785
rect 23750 18776 23756 18828
rect 23808 18776 23814 18828
rect 23934 18825 23940 18828
rect 23928 18816 23940 18825
rect 23895 18788 23940 18816
rect 23928 18779 23940 18788
rect 23934 18776 23940 18779
rect 23992 18776 23998 18828
rect 20898 18748 20904 18760
rect 19904 18720 20904 18748
rect 19061 18711 19119 18717
rect 20898 18708 20904 18720
rect 20956 18708 20962 18760
rect 20990 18708 20996 18760
rect 21048 18708 21054 18760
rect 21453 18751 21511 18757
rect 21453 18717 21465 18751
rect 21499 18717 21511 18751
rect 21453 18711 21511 18717
rect 15059 18652 15700 18680
rect 15059 18649 15071 18652
rect 15013 18643 15071 18649
rect 20806 18640 20812 18692
rect 20864 18680 20870 18692
rect 21468 18680 21496 18711
rect 23290 18708 23296 18760
rect 23348 18748 23354 18760
rect 23768 18748 23796 18776
rect 23348 18720 23796 18748
rect 23348 18708 23354 18720
rect 20864 18652 21496 18680
rect 20864 18640 20870 18652
rect 2682 18572 2688 18624
rect 2740 18612 2746 18624
rect 3053 18615 3111 18621
rect 3053 18612 3065 18615
rect 2740 18584 3065 18612
rect 2740 18572 2746 18584
rect 3053 18581 3065 18584
rect 3099 18581 3111 18615
rect 8018 18612 8024 18624
rect 7979 18584 8024 18612
rect 3053 18575 3111 18581
rect 8018 18572 8024 18584
rect 8076 18572 8082 18624
rect 9306 18612 9312 18624
rect 9267 18584 9312 18612
rect 9306 18572 9312 18584
rect 9364 18612 9370 18624
rect 9490 18612 9496 18624
rect 9364 18584 9496 18612
rect 9364 18572 9370 18584
rect 9490 18572 9496 18584
rect 9548 18572 9554 18624
rect 10229 18615 10287 18621
rect 10229 18581 10241 18615
rect 10275 18612 10287 18615
rect 10962 18612 10968 18624
rect 10275 18584 10968 18612
rect 10275 18581 10287 18584
rect 10229 18575 10287 18581
rect 10962 18572 10968 18584
rect 11020 18572 11026 18624
rect 11330 18572 11336 18624
rect 11388 18612 11394 18624
rect 11701 18615 11759 18621
rect 11701 18612 11713 18615
rect 11388 18584 11713 18612
rect 11388 18572 11394 18584
rect 11701 18581 11713 18584
rect 11747 18581 11759 18615
rect 11701 18575 11759 18581
rect 12529 18615 12587 18621
rect 12529 18581 12541 18615
rect 12575 18612 12587 18615
rect 12710 18612 12716 18624
rect 12575 18584 12716 18612
rect 12575 18581 12587 18584
rect 12529 18575 12587 18581
rect 12710 18572 12716 18584
rect 12768 18572 12774 18624
rect 14550 18612 14556 18624
rect 14511 18584 14556 18612
rect 14550 18572 14556 18584
rect 14608 18572 14614 18624
rect 18414 18572 18420 18624
rect 18472 18612 18478 18624
rect 18509 18615 18567 18621
rect 18509 18612 18521 18615
rect 18472 18584 18521 18612
rect 18472 18572 18478 18584
rect 18509 18581 18521 18584
rect 18555 18612 18567 18615
rect 19521 18615 19579 18621
rect 19521 18612 19533 18615
rect 18555 18584 19533 18612
rect 18555 18581 18567 18584
rect 18509 18575 18567 18581
rect 19521 18581 19533 18584
rect 19567 18581 19579 18615
rect 19521 18575 19579 18581
rect 20717 18615 20775 18621
rect 20717 18581 20729 18615
rect 20763 18612 20775 18615
rect 20898 18612 20904 18624
rect 20763 18584 20904 18612
rect 20763 18581 20775 18584
rect 20717 18575 20775 18581
rect 20898 18572 20904 18584
rect 20956 18572 20962 18624
rect 22094 18572 22100 18624
rect 22152 18612 22158 18624
rect 22281 18615 22339 18621
rect 22281 18612 22293 18615
rect 22152 18584 22293 18612
rect 22152 18572 22158 18584
rect 22281 18581 22293 18584
rect 22327 18581 22339 18615
rect 22281 18575 22339 18581
rect 23014 18572 23020 18624
rect 23072 18612 23078 18624
rect 23109 18615 23167 18621
rect 23109 18612 23121 18615
rect 23072 18584 23121 18612
rect 23072 18572 23078 18584
rect 23109 18581 23121 18584
rect 23155 18581 23167 18615
rect 23109 18575 23167 18581
rect 24762 18572 24768 18624
rect 24820 18612 24826 18624
rect 25593 18615 25651 18621
rect 25593 18612 25605 18615
rect 24820 18584 25605 18612
rect 24820 18572 24826 18584
rect 25593 18581 25605 18584
rect 25639 18612 25651 18615
rect 26142 18612 26148 18624
rect 25639 18584 26148 18612
rect 25639 18581 25651 18584
rect 25593 18575 25651 18581
rect 26142 18572 26148 18584
rect 26200 18572 26206 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 2041 18411 2099 18417
rect 2041 18377 2053 18411
rect 2087 18408 2099 18411
rect 2498 18408 2504 18420
rect 2087 18380 2504 18408
rect 2087 18377 2099 18380
rect 2041 18371 2099 18377
rect 2498 18368 2504 18380
rect 2556 18368 2562 18420
rect 4706 18408 4712 18420
rect 4667 18380 4712 18408
rect 4706 18368 4712 18380
rect 4764 18368 4770 18420
rect 5534 18368 5540 18420
rect 5592 18408 5598 18420
rect 6549 18411 6607 18417
rect 6549 18408 6561 18411
rect 5592 18380 6561 18408
rect 5592 18368 5598 18380
rect 6549 18377 6561 18380
rect 6595 18377 6607 18411
rect 6549 18371 6607 18377
rect 2130 18272 2136 18284
rect 2091 18244 2136 18272
rect 2130 18232 2136 18244
rect 2188 18232 2194 18284
rect 4249 18275 4307 18281
rect 4249 18241 4261 18275
rect 4295 18272 4307 18275
rect 5350 18272 5356 18284
rect 4295 18244 5356 18272
rect 4295 18241 4307 18244
rect 4249 18235 4307 18241
rect 5350 18232 5356 18244
rect 5408 18232 5414 18284
rect 4617 18207 4675 18213
rect 4617 18173 4629 18207
rect 4663 18204 4675 18207
rect 5258 18204 5264 18216
rect 4663 18176 5264 18204
rect 4663 18173 4675 18176
rect 4617 18167 4675 18173
rect 5258 18164 5264 18176
rect 5316 18164 5322 18216
rect 6564 18204 6592 18371
rect 7190 18368 7196 18420
rect 7248 18408 7254 18420
rect 7745 18411 7803 18417
rect 7745 18408 7757 18411
rect 7248 18380 7757 18408
rect 7248 18368 7254 18380
rect 7745 18377 7757 18380
rect 7791 18408 7803 18411
rect 8478 18408 8484 18420
rect 7791 18380 8484 18408
rect 7791 18377 7803 18380
rect 7745 18371 7803 18377
rect 8478 18368 8484 18380
rect 8536 18368 8542 18420
rect 8662 18368 8668 18420
rect 8720 18408 8726 18420
rect 9582 18408 9588 18420
rect 8720 18380 9588 18408
rect 8720 18368 8726 18380
rect 9582 18368 9588 18380
rect 9640 18408 9646 18420
rect 9674 18408 9680 18420
rect 9640 18380 9680 18408
rect 9640 18368 9646 18380
rect 9674 18368 9680 18380
rect 9732 18368 9738 18420
rect 10134 18368 10140 18420
rect 10192 18408 10198 18420
rect 10229 18411 10287 18417
rect 10229 18408 10241 18411
rect 10192 18380 10241 18408
rect 10192 18368 10198 18380
rect 10229 18377 10241 18380
rect 10275 18377 10287 18411
rect 12250 18408 12256 18420
rect 12211 18380 12256 18408
rect 10229 18371 10287 18377
rect 12250 18368 12256 18380
rect 12308 18368 12314 18420
rect 13814 18408 13820 18420
rect 12360 18380 13400 18408
rect 13775 18380 13820 18408
rect 8110 18340 8116 18352
rect 8071 18312 8116 18340
rect 8110 18300 8116 18312
rect 8168 18300 8174 18352
rect 12360 18340 12388 18380
rect 9324 18312 12388 18340
rect 13372 18340 13400 18380
rect 13814 18368 13820 18380
rect 13872 18368 13878 18420
rect 15562 18408 15568 18420
rect 14384 18380 15568 18408
rect 14384 18340 14412 18380
rect 15562 18368 15568 18380
rect 15620 18368 15626 18420
rect 16301 18411 16359 18417
rect 16301 18377 16313 18411
rect 16347 18408 16359 18411
rect 16666 18408 16672 18420
rect 16347 18380 16672 18408
rect 16347 18377 16359 18380
rect 16301 18371 16359 18377
rect 16666 18368 16672 18380
rect 16724 18368 16730 18420
rect 17037 18411 17095 18417
rect 17037 18377 17049 18411
rect 17083 18408 17095 18411
rect 17494 18408 17500 18420
rect 17083 18380 17500 18408
rect 17083 18377 17095 18380
rect 17037 18371 17095 18377
rect 17494 18368 17500 18380
rect 17552 18368 17558 18420
rect 19058 18408 19064 18420
rect 19019 18380 19064 18408
rect 19058 18368 19064 18380
rect 19116 18408 19122 18420
rect 19705 18411 19763 18417
rect 19705 18408 19717 18411
rect 19116 18380 19717 18408
rect 19116 18368 19122 18380
rect 19705 18377 19717 18380
rect 19751 18408 19763 18411
rect 20990 18408 20996 18420
rect 19751 18380 20392 18408
rect 20951 18380 20996 18408
rect 19751 18377 19763 18380
rect 19705 18371 19763 18377
rect 13372 18312 14412 18340
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 6564 18176 6837 18204
rect 6825 18173 6837 18176
rect 6871 18173 6883 18207
rect 6825 18167 6883 18173
rect 8297 18207 8355 18213
rect 8297 18173 8309 18207
rect 8343 18204 8355 18207
rect 8846 18204 8852 18216
rect 8343 18176 8852 18204
rect 8343 18173 8355 18176
rect 8297 18167 8355 18173
rect 8846 18164 8852 18176
rect 8904 18164 8910 18216
rect 9030 18164 9036 18216
rect 9088 18204 9094 18216
rect 9324 18204 9352 18312
rect 11054 18232 11060 18284
rect 11112 18272 11118 18284
rect 11333 18275 11391 18281
rect 11333 18272 11345 18275
rect 11112 18244 11345 18272
rect 11112 18232 11118 18244
rect 11333 18241 11345 18244
rect 11379 18241 11391 18275
rect 14734 18272 14740 18284
rect 11333 18235 11391 18241
rect 14200 18244 14740 18272
rect 10686 18204 10692 18216
rect 9088 18176 9352 18204
rect 10599 18176 10692 18204
rect 9088 18164 9094 18176
rect 10686 18164 10692 18176
rect 10744 18204 10750 18216
rect 11149 18207 11207 18213
rect 11149 18204 11161 18207
rect 10744 18176 11161 18204
rect 10744 18164 10750 18176
rect 11149 18173 11161 18176
rect 11195 18204 11207 18207
rect 11974 18204 11980 18216
rect 11195 18176 11980 18204
rect 11195 18173 11207 18176
rect 11149 18167 11207 18173
rect 11974 18164 11980 18176
rect 12032 18164 12038 18216
rect 12250 18164 12256 18216
rect 12308 18204 12314 18216
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 12308 18176 12449 18204
rect 12308 18164 12314 18176
rect 12437 18173 12449 18176
rect 12483 18173 12495 18207
rect 14200 18204 14228 18244
rect 14734 18232 14740 18244
rect 14792 18232 14798 18284
rect 18046 18232 18052 18284
rect 18104 18272 18110 18284
rect 18509 18275 18567 18281
rect 18509 18272 18521 18275
rect 18104 18244 18521 18272
rect 18104 18232 18110 18244
rect 18509 18241 18521 18244
rect 18555 18241 18567 18275
rect 18509 18235 18567 18241
rect 12437 18167 12495 18173
rect 12544 18176 14228 18204
rect 2038 18096 2044 18148
rect 2096 18136 2102 18148
rect 2378 18139 2436 18145
rect 2378 18136 2390 18139
rect 2096 18108 2390 18136
rect 2096 18096 2102 18108
rect 2378 18105 2390 18108
rect 2424 18105 2436 18139
rect 5074 18136 5080 18148
rect 4987 18108 5080 18136
rect 2378 18099 2436 18105
rect 5074 18096 5080 18108
rect 5132 18136 5138 18148
rect 6089 18139 6147 18145
rect 6089 18136 6101 18139
rect 5132 18108 6101 18136
rect 5132 18096 5138 18108
rect 6089 18105 6101 18108
rect 6135 18105 6147 18139
rect 6089 18099 6147 18105
rect 7101 18139 7159 18145
rect 7101 18105 7113 18139
rect 7147 18105 7159 18139
rect 7101 18099 7159 18105
rect 8564 18139 8622 18145
rect 8564 18105 8576 18139
rect 8610 18136 8622 18139
rect 9214 18136 9220 18148
rect 8610 18108 9220 18136
rect 8610 18105 8622 18108
rect 8564 18099 8622 18105
rect 1673 18071 1731 18077
rect 1673 18037 1685 18071
rect 1719 18068 1731 18071
rect 2590 18068 2596 18080
rect 1719 18040 2596 18068
rect 1719 18037 1731 18040
rect 1673 18031 1731 18037
rect 2590 18028 2596 18040
rect 2648 18028 2654 18080
rect 2866 18028 2872 18080
rect 2924 18068 2930 18080
rect 3513 18071 3571 18077
rect 3513 18068 3525 18071
rect 2924 18040 3525 18068
rect 2924 18028 2930 18040
rect 3513 18037 3525 18040
rect 3559 18068 3571 18071
rect 4062 18068 4068 18080
rect 3559 18040 4068 18068
rect 3559 18037 3571 18040
rect 3513 18031 3571 18037
rect 4062 18028 4068 18040
rect 4120 18028 4126 18080
rect 4982 18028 4988 18080
rect 5040 18068 5046 18080
rect 5169 18071 5227 18077
rect 5169 18068 5181 18071
rect 5040 18040 5181 18068
rect 5040 18028 5046 18040
rect 5169 18037 5181 18040
rect 5215 18068 5227 18071
rect 5721 18071 5779 18077
rect 5721 18068 5733 18071
rect 5215 18040 5733 18068
rect 5215 18037 5227 18040
rect 5169 18031 5227 18037
rect 5721 18037 5733 18040
rect 5767 18037 5779 18071
rect 5721 18031 5779 18037
rect 6822 18028 6828 18080
rect 6880 18068 6886 18080
rect 7116 18068 7144 18099
rect 9214 18096 9220 18108
rect 9272 18096 9278 18148
rect 11238 18136 11244 18148
rect 10612 18108 11100 18136
rect 11199 18108 11244 18136
rect 6880 18040 7144 18068
rect 6880 18028 6886 18040
rect 8386 18028 8392 18080
rect 8444 18068 8450 18080
rect 10612 18068 10640 18108
rect 10778 18068 10784 18080
rect 8444 18040 10640 18068
rect 10739 18040 10784 18068
rect 8444 18028 8450 18040
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 11072 18068 11100 18108
rect 11238 18096 11244 18108
rect 11296 18136 11302 18148
rect 11793 18139 11851 18145
rect 11793 18136 11805 18139
rect 11296 18108 11805 18136
rect 11296 18096 11302 18108
rect 11793 18105 11805 18108
rect 11839 18105 11851 18139
rect 11793 18099 11851 18105
rect 12544 18068 12572 18176
rect 14274 18164 14280 18216
rect 14332 18204 14338 18216
rect 14918 18204 14924 18216
rect 14332 18176 14924 18204
rect 14332 18164 14338 18176
rect 14918 18164 14924 18176
rect 14976 18164 14982 18216
rect 17770 18204 17776 18216
rect 17731 18176 17776 18204
rect 17770 18164 17776 18176
rect 17828 18164 17834 18216
rect 18414 18204 18420 18216
rect 18375 18176 18420 18204
rect 18414 18164 18420 18176
rect 18472 18164 18478 18216
rect 18524 18204 18552 18235
rect 18598 18232 18604 18284
rect 18656 18272 18662 18284
rect 20364 18281 20392 18380
rect 20990 18368 20996 18380
rect 21048 18368 21054 18420
rect 21174 18368 21180 18420
rect 21232 18408 21238 18420
rect 21269 18411 21327 18417
rect 21269 18408 21281 18411
rect 21232 18380 21281 18408
rect 21232 18368 21238 18380
rect 21269 18377 21281 18380
rect 21315 18377 21327 18411
rect 22554 18408 22560 18420
rect 22515 18380 22560 18408
rect 21269 18371 21327 18377
rect 22554 18368 22560 18380
rect 22612 18368 22618 18420
rect 23109 18411 23167 18417
rect 23109 18377 23121 18411
rect 23155 18408 23167 18411
rect 23934 18408 23940 18420
rect 23155 18380 23940 18408
rect 23155 18377 23167 18380
rect 23109 18371 23167 18377
rect 23934 18368 23940 18380
rect 23992 18408 23998 18420
rect 25041 18411 25099 18417
rect 25041 18408 25053 18411
rect 23992 18380 25053 18408
rect 23992 18368 23998 18380
rect 25041 18377 25053 18380
rect 25087 18377 25099 18411
rect 25041 18371 25099 18377
rect 20714 18300 20720 18352
rect 20772 18340 20778 18352
rect 21453 18343 21511 18349
rect 21453 18340 21465 18343
rect 20772 18312 21465 18340
rect 20772 18300 20778 18312
rect 21453 18309 21465 18312
rect 21499 18309 21511 18343
rect 21453 18303 21511 18309
rect 20349 18275 20407 18281
rect 18656 18244 18701 18272
rect 18656 18232 18662 18244
rect 20349 18241 20361 18275
rect 20395 18241 20407 18275
rect 20349 18235 20407 18241
rect 20533 18275 20591 18281
rect 20533 18241 20545 18275
rect 20579 18272 20591 18275
rect 20806 18272 20812 18284
rect 20579 18244 20812 18272
rect 20579 18241 20591 18244
rect 20533 18235 20591 18241
rect 20806 18232 20812 18244
rect 20864 18232 20870 18284
rect 20898 18232 20904 18284
rect 20956 18272 20962 18284
rect 21913 18275 21971 18281
rect 21913 18272 21925 18275
rect 20956 18244 21925 18272
rect 20956 18232 20962 18244
rect 21913 18241 21925 18244
rect 21959 18241 21971 18275
rect 22094 18272 22100 18284
rect 22055 18244 22100 18272
rect 21913 18235 21971 18241
rect 22094 18232 22100 18244
rect 22152 18232 22158 18284
rect 23566 18232 23572 18284
rect 23624 18272 23630 18284
rect 23661 18275 23719 18281
rect 23661 18272 23673 18275
rect 23624 18244 23673 18272
rect 23624 18232 23630 18244
rect 23661 18241 23673 18244
rect 23707 18241 23719 18275
rect 23661 18235 23719 18241
rect 19242 18204 19248 18216
rect 18524 18176 19248 18204
rect 19242 18164 19248 18176
rect 19300 18164 19306 18216
rect 19886 18164 19892 18216
rect 19944 18204 19950 18216
rect 20257 18207 20315 18213
rect 20257 18204 20269 18207
rect 19944 18176 20269 18204
rect 19944 18164 19950 18176
rect 20257 18173 20269 18176
rect 20303 18173 20315 18207
rect 20257 18167 20315 18173
rect 21450 18164 21456 18216
rect 21508 18204 21514 18216
rect 22554 18204 22560 18216
rect 21508 18176 22560 18204
rect 21508 18164 21514 18176
rect 22554 18164 22560 18176
rect 22612 18164 22618 18216
rect 23676 18204 23704 18235
rect 24762 18204 24768 18216
rect 23676 18176 24768 18204
rect 24762 18164 24768 18176
rect 24820 18164 24826 18216
rect 12710 18145 12716 18148
rect 12704 18136 12716 18145
rect 12671 18108 12716 18136
rect 12704 18099 12716 18108
rect 12768 18136 12774 18148
rect 14369 18139 14427 18145
rect 14369 18136 14381 18139
rect 12768 18108 14381 18136
rect 12710 18096 12716 18099
rect 12768 18096 12774 18108
rect 14369 18105 14381 18108
rect 14415 18105 14427 18139
rect 14369 18099 14427 18105
rect 11072 18040 12572 18068
rect 14384 18068 14412 18099
rect 14550 18096 14556 18148
rect 14608 18136 14614 18148
rect 14829 18139 14887 18145
rect 14829 18136 14841 18139
rect 14608 18108 14841 18136
rect 14608 18096 14614 18108
rect 14829 18105 14841 18108
rect 14875 18136 14887 18139
rect 15188 18139 15246 18145
rect 15188 18136 15200 18139
rect 14875 18108 15200 18136
rect 14875 18105 14887 18108
rect 14829 18099 14887 18105
rect 15188 18105 15200 18108
rect 15234 18136 15246 18139
rect 15378 18136 15384 18148
rect 15234 18108 15384 18136
rect 15234 18105 15246 18108
rect 15188 18099 15246 18105
rect 15378 18096 15384 18108
rect 15436 18096 15442 18148
rect 21821 18139 21879 18145
rect 21821 18136 21833 18139
rect 19904 18108 21833 18136
rect 16022 18068 16028 18080
rect 14384 18040 16028 18068
rect 16022 18028 16028 18040
rect 16080 18028 16086 18080
rect 17497 18071 17555 18077
rect 17497 18037 17509 18071
rect 17543 18068 17555 18071
rect 17678 18068 17684 18080
rect 17543 18040 17684 18068
rect 17543 18037 17555 18040
rect 17497 18031 17555 18037
rect 17678 18028 17684 18040
rect 17736 18028 17742 18080
rect 17862 18028 17868 18080
rect 17920 18068 17926 18080
rect 19904 18077 19932 18108
rect 21821 18105 21833 18108
rect 21867 18136 21879 18139
rect 22094 18136 22100 18148
rect 21867 18108 22100 18136
rect 21867 18105 21879 18108
rect 21821 18099 21879 18105
rect 22094 18096 22100 18108
rect 22152 18096 22158 18148
rect 23934 18145 23940 18148
rect 23477 18139 23535 18145
rect 23477 18105 23489 18139
rect 23523 18136 23535 18139
rect 23928 18136 23940 18145
rect 23523 18108 23940 18136
rect 23523 18105 23535 18108
rect 23477 18099 23535 18105
rect 23928 18099 23940 18108
rect 23934 18096 23940 18099
rect 23992 18096 23998 18148
rect 18049 18071 18107 18077
rect 18049 18068 18061 18071
rect 17920 18040 18061 18068
rect 17920 18028 17926 18040
rect 18049 18037 18061 18040
rect 18095 18037 18107 18071
rect 18049 18031 18107 18037
rect 19889 18071 19947 18077
rect 19889 18037 19901 18071
rect 19935 18037 19947 18071
rect 19889 18031 19947 18037
rect 24026 18028 24032 18080
rect 24084 18068 24090 18080
rect 25406 18068 25412 18080
rect 24084 18040 25412 18068
rect 24084 18028 24090 18040
rect 25406 18028 25412 18040
rect 25464 18028 25470 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1670 17824 1676 17876
rect 1728 17864 1734 17876
rect 2133 17867 2191 17873
rect 2133 17864 2145 17867
rect 1728 17836 2145 17864
rect 1728 17824 1734 17836
rect 2133 17833 2145 17836
rect 2179 17864 2191 17867
rect 2682 17864 2688 17876
rect 2179 17836 2688 17864
rect 2179 17833 2191 17836
rect 2133 17827 2191 17833
rect 2682 17824 2688 17836
rect 2740 17824 2746 17876
rect 2774 17824 2780 17876
rect 2832 17864 2838 17876
rect 6089 17867 6147 17873
rect 2832 17836 2877 17864
rect 2832 17824 2838 17836
rect 6089 17833 6101 17867
rect 6135 17864 6147 17867
rect 6362 17864 6368 17876
rect 6135 17836 6368 17864
rect 6135 17833 6147 17836
rect 6089 17827 6147 17833
rect 6362 17824 6368 17836
rect 6420 17824 6426 17876
rect 6730 17864 6736 17876
rect 6691 17836 6736 17864
rect 6730 17824 6736 17836
rect 6788 17824 6794 17876
rect 7561 17867 7619 17873
rect 7561 17833 7573 17867
rect 7607 17864 7619 17867
rect 8018 17864 8024 17876
rect 7607 17836 8024 17864
rect 7607 17833 7619 17836
rect 7561 17827 7619 17833
rect 8018 17824 8024 17836
rect 8076 17864 8082 17876
rect 8481 17867 8539 17873
rect 8481 17864 8493 17867
rect 8076 17836 8493 17864
rect 8076 17824 8082 17836
rect 8481 17833 8493 17836
rect 8527 17833 8539 17867
rect 8481 17827 8539 17833
rect 9858 17824 9864 17876
rect 9916 17864 9922 17876
rect 10505 17867 10563 17873
rect 10505 17864 10517 17867
rect 9916 17836 10517 17864
rect 9916 17824 9922 17836
rect 10505 17833 10517 17836
rect 10551 17864 10563 17867
rect 12894 17864 12900 17876
rect 10551 17836 11008 17864
rect 12855 17836 12900 17864
rect 10551 17833 10563 17836
rect 10505 17827 10563 17833
rect 1302 17756 1308 17808
rect 1360 17796 1366 17808
rect 9030 17796 9036 17808
rect 1360 17768 9036 17796
rect 1360 17756 1366 17768
rect 9030 17756 9036 17768
rect 9088 17756 9094 17808
rect 10980 17796 11008 17836
rect 12894 17824 12900 17836
rect 12952 17824 12958 17876
rect 13814 17824 13820 17876
rect 13872 17864 13878 17876
rect 14274 17864 14280 17876
rect 13872 17836 14280 17864
rect 13872 17824 13878 17836
rect 14274 17824 14280 17836
rect 14332 17864 14338 17876
rect 14461 17867 14519 17873
rect 14461 17864 14473 17867
rect 14332 17836 14473 17864
rect 14332 17824 14338 17836
rect 14461 17833 14473 17836
rect 14507 17833 14519 17867
rect 14461 17827 14519 17833
rect 14734 17824 14740 17876
rect 14792 17864 14798 17876
rect 15013 17867 15071 17873
rect 15013 17864 15025 17867
rect 14792 17836 15025 17864
rect 14792 17824 14798 17836
rect 15013 17833 15025 17836
rect 15059 17833 15071 17867
rect 15286 17864 15292 17876
rect 15247 17836 15292 17864
rect 15013 17827 15071 17833
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 15654 17824 15660 17876
rect 15712 17824 15718 17876
rect 16574 17864 16580 17876
rect 16535 17836 16580 17864
rect 16574 17824 16580 17836
rect 16632 17824 16638 17876
rect 16945 17867 17003 17873
rect 16945 17833 16957 17867
rect 16991 17864 17003 17867
rect 17862 17864 17868 17876
rect 16991 17836 17868 17864
rect 16991 17833 17003 17836
rect 16945 17827 17003 17833
rect 17862 17824 17868 17836
rect 17920 17824 17926 17876
rect 19334 17864 19340 17876
rect 19295 17836 19340 17864
rect 19334 17824 19340 17836
rect 19392 17824 19398 17876
rect 20070 17824 20076 17876
rect 20128 17864 20134 17876
rect 20438 17864 20444 17876
rect 20128 17836 20444 17864
rect 20128 17824 20134 17836
rect 20438 17824 20444 17836
rect 20496 17824 20502 17876
rect 22094 17824 22100 17876
rect 22152 17864 22158 17876
rect 22833 17867 22891 17873
rect 22833 17864 22845 17867
rect 22152 17836 22845 17864
rect 22152 17824 22158 17836
rect 22833 17833 22845 17836
rect 22879 17833 22891 17867
rect 24854 17864 24860 17876
rect 24815 17836 24860 17864
rect 22833 17827 22891 17833
rect 24854 17824 24860 17836
rect 24912 17824 24918 17876
rect 11232 17799 11290 17805
rect 11232 17796 11244 17799
rect 10980 17768 11244 17796
rect 11232 17765 11244 17768
rect 11278 17796 11290 17799
rect 12342 17796 12348 17808
rect 11278 17768 12348 17796
rect 11278 17765 11290 17768
rect 11232 17759 11290 17765
rect 12342 17756 12348 17768
rect 12400 17756 12406 17808
rect 13909 17799 13967 17805
rect 13909 17765 13921 17799
rect 13955 17796 13967 17799
rect 13998 17796 14004 17808
rect 13955 17768 14004 17796
rect 13955 17765 13967 17768
rect 13909 17759 13967 17765
rect 13998 17756 14004 17768
rect 14056 17796 14062 17808
rect 15672 17796 15700 17824
rect 14056 17768 15700 17796
rect 17304 17799 17362 17805
rect 14056 17756 14062 17768
rect 17304 17765 17316 17799
rect 17350 17796 17362 17799
rect 17402 17796 17408 17808
rect 17350 17768 17408 17796
rect 17350 17765 17362 17768
rect 17304 17759 17362 17765
rect 17402 17756 17408 17768
rect 17460 17796 17466 17808
rect 18966 17796 18972 17808
rect 17460 17768 18972 17796
rect 17460 17756 17466 17768
rect 18966 17756 18972 17768
rect 19024 17756 19030 17808
rect 19797 17799 19855 17805
rect 19797 17765 19809 17799
rect 19843 17796 19855 17799
rect 19978 17796 19984 17808
rect 19843 17768 19984 17796
rect 19843 17765 19855 17768
rect 19797 17759 19855 17765
rect 19978 17756 19984 17768
rect 20036 17756 20042 17808
rect 20530 17756 20536 17808
rect 20588 17756 20594 17808
rect 25038 17756 25044 17808
rect 25096 17796 25102 17808
rect 25225 17799 25283 17805
rect 25225 17796 25237 17799
rect 25096 17768 25237 17796
rect 25096 17756 25102 17768
rect 25225 17765 25237 17768
rect 25271 17765 25283 17799
rect 25225 17759 25283 17765
rect 1673 17731 1731 17737
rect 1673 17697 1685 17731
rect 1719 17728 1731 17731
rect 2038 17728 2044 17740
rect 1719 17700 2044 17728
rect 1719 17697 1731 17700
rect 1673 17691 1731 17697
rect 2038 17688 2044 17700
rect 2096 17688 2102 17740
rect 2225 17731 2283 17737
rect 2225 17697 2237 17731
rect 2271 17728 2283 17731
rect 2682 17728 2688 17740
rect 2271 17700 2688 17728
rect 2271 17697 2283 17700
rect 2225 17691 2283 17697
rect 2682 17688 2688 17700
rect 2740 17728 2746 17740
rect 3513 17731 3571 17737
rect 3513 17728 3525 17731
rect 2740 17700 3525 17728
rect 2740 17688 2746 17700
rect 3513 17697 3525 17700
rect 3559 17697 3571 17731
rect 3513 17691 3571 17697
rect 3602 17688 3608 17740
rect 3660 17728 3666 17740
rect 4065 17731 4123 17737
rect 4065 17728 4077 17731
rect 3660 17700 4077 17728
rect 3660 17688 3666 17700
rect 4065 17697 4077 17700
rect 4111 17697 4123 17731
rect 4065 17691 4123 17697
rect 4154 17688 4160 17740
rect 4212 17728 4218 17740
rect 4321 17731 4379 17737
rect 4321 17728 4333 17731
rect 4212 17700 4333 17728
rect 4212 17688 4218 17700
rect 4321 17697 4333 17700
rect 4367 17697 4379 17731
rect 4321 17691 4379 17697
rect 6549 17731 6607 17737
rect 6549 17697 6561 17731
rect 6595 17728 6607 17731
rect 6638 17728 6644 17740
rect 6595 17700 6644 17728
rect 6595 17697 6607 17700
rect 6549 17691 6607 17697
rect 6638 17688 6644 17700
rect 6696 17688 6702 17740
rect 7193 17731 7251 17737
rect 7193 17697 7205 17731
rect 7239 17728 7251 17731
rect 8386 17728 8392 17740
rect 7239 17700 8392 17728
rect 7239 17697 7251 17700
rect 7193 17691 7251 17697
rect 8386 17688 8392 17700
rect 8444 17688 8450 17740
rect 9490 17688 9496 17740
rect 9548 17728 9554 17740
rect 9677 17731 9735 17737
rect 9677 17728 9689 17731
rect 9548 17700 9689 17728
rect 9548 17688 9554 17700
rect 9677 17697 9689 17700
rect 9723 17728 9735 17731
rect 10686 17728 10692 17740
rect 9723 17700 10692 17728
rect 9723 17697 9735 17700
rect 9677 17691 9735 17697
rect 10686 17688 10692 17700
rect 10744 17688 10750 17740
rect 10873 17731 10931 17737
rect 10873 17697 10885 17731
rect 10919 17728 10931 17731
rect 11054 17728 11060 17740
rect 10919 17700 11060 17728
rect 10919 17697 10931 17700
rect 10873 17691 10931 17697
rect 2314 17620 2320 17672
rect 2372 17660 2378 17672
rect 2866 17660 2872 17672
rect 2372 17632 2872 17660
rect 2372 17620 2378 17632
rect 2866 17620 2872 17632
rect 2924 17620 2930 17672
rect 8202 17620 8208 17672
rect 8260 17660 8266 17672
rect 8662 17660 8668 17672
rect 8260 17632 8668 17660
rect 8260 17620 8266 17632
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 9950 17660 9956 17672
rect 9911 17632 9956 17660
rect 9950 17620 9956 17632
rect 10008 17620 10014 17672
rect 10594 17620 10600 17672
rect 10652 17660 10658 17672
rect 10888 17660 10916 17691
rect 11054 17688 11060 17700
rect 11112 17688 11118 17740
rect 13722 17688 13728 17740
rect 13780 17728 13786 17740
rect 13817 17731 13875 17737
rect 13817 17728 13829 17731
rect 13780 17700 13829 17728
rect 13780 17688 13786 17700
rect 13817 17697 13829 17700
rect 13863 17697 13875 17731
rect 13817 17691 13875 17697
rect 14550 17688 14556 17740
rect 14608 17728 14614 17740
rect 15657 17731 15715 17737
rect 15657 17728 15669 17731
rect 14608 17700 15669 17728
rect 14608 17688 14614 17700
rect 15657 17697 15669 17700
rect 15703 17697 15715 17731
rect 15657 17691 15715 17697
rect 15746 17688 15752 17740
rect 15804 17728 15810 17740
rect 19518 17728 19524 17740
rect 15804 17700 15849 17728
rect 19479 17700 19524 17728
rect 15804 17688 15810 17700
rect 19518 17688 19524 17700
rect 19576 17688 19582 17740
rect 20548 17728 20576 17756
rect 19996 17700 20576 17728
rect 19996 17672 20024 17700
rect 20806 17688 20812 17740
rect 20864 17728 20870 17740
rect 21157 17731 21215 17737
rect 21157 17728 21169 17731
rect 20864 17700 21169 17728
rect 20864 17688 20870 17700
rect 21157 17697 21169 17700
rect 21203 17697 21215 17731
rect 21157 17691 21215 17697
rect 23753 17731 23811 17737
rect 23753 17697 23765 17731
rect 23799 17728 23811 17731
rect 24026 17728 24032 17740
rect 23799 17700 24032 17728
rect 23799 17697 23811 17700
rect 23753 17691 23811 17697
rect 24026 17688 24032 17700
rect 24084 17688 24090 17740
rect 24949 17731 25007 17737
rect 24949 17697 24961 17731
rect 24995 17697 25007 17731
rect 24949 17691 25007 17697
rect 10652 17632 10916 17660
rect 10965 17663 11023 17669
rect 10652 17620 10658 17632
rect 10965 17629 10977 17663
rect 11011 17629 11023 17663
rect 10965 17623 11023 17629
rect 8018 17592 8024 17604
rect 7979 17564 8024 17592
rect 8018 17552 8024 17564
rect 8076 17552 8082 17604
rect 8846 17552 8852 17604
rect 8904 17592 8910 17604
rect 9401 17595 9459 17601
rect 9401 17592 9413 17595
rect 8904 17564 9413 17592
rect 8904 17552 8910 17564
rect 9401 17561 9413 17564
rect 9447 17592 9459 17595
rect 10980 17592 11008 17623
rect 12434 17620 12440 17672
rect 12492 17660 12498 17672
rect 14093 17663 14151 17669
rect 12492 17632 13492 17660
rect 12492 17620 12498 17632
rect 9447 17564 11008 17592
rect 9447 17561 9459 17564
rect 9401 17555 9459 17561
rect 10980 17536 11008 17564
rect 12345 17595 12403 17601
rect 12345 17561 12357 17595
rect 12391 17592 12403 17595
rect 12710 17592 12716 17604
rect 12391 17564 12716 17592
rect 12391 17561 12403 17564
rect 12345 17555 12403 17561
rect 12710 17552 12716 17564
rect 12768 17592 12774 17604
rect 13354 17592 13360 17604
rect 12768 17564 13360 17592
rect 12768 17552 12774 17564
rect 13354 17552 13360 17564
rect 13412 17552 13418 17604
rect 13464 17601 13492 17632
rect 14093 17629 14105 17663
rect 14139 17660 14151 17663
rect 14182 17660 14188 17672
rect 14139 17632 14188 17660
rect 14139 17629 14151 17632
rect 14093 17623 14151 17629
rect 14182 17620 14188 17632
rect 14240 17620 14246 17672
rect 14734 17620 14740 17672
rect 14792 17660 14798 17672
rect 14918 17660 14924 17672
rect 14792 17632 14924 17660
rect 14792 17620 14798 17632
rect 14918 17620 14924 17632
rect 14976 17620 14982 17672
rect 15930 17660 15936 17672
rect 15891 17632 15936 17660
rect 15930 17620 15936 17632
rect 15988 17620 15994 17672
rect 17037 17663 17095 17669
rect 17037 17629 17049 17663
rect 17083 17629 17095 17663
rect 17037 17623 17095 17629
rect 13449 17595 13507 17601
rect 13449 17561 13461 17595
rect 13495 17561 13507 17595
rect 14936 17592 14964 17620
rect 17052 17592 17080 17623
rect 19978 17620 19984 17672
rect 20036 17620 20042 17672
rect 20901 17663 20959 17669
rect 20901 17629 20913 17663
rect 20947 17629 20959 17663
rect 20901 17623 20959 17629
rect 14936 17564 17080 17592
rect 13449 17555 13507 17561
rect 20530 17552 20536 17604
rect 20588 17592 20594 17604
rect 20916 17592 20944 17623
rect 22738 17620 22744 17672
rect 22796 17660 22802 17672
rect 23566 17660 23572 17672
rect 22796 17632 23572 17660
rect 22796 17620 22802 17632
rect 23566 17620 23572 17632
rect 23624 17660 23630 17672
rect 23845 17663 23903 17669
rect 23845 17660 23857 17663
rect 23624 17632 23857 17660
rect 23624 17620 23630 17632
rect 23845 17629 23857 17632
rect 23891 17629 23903 17663
rect 23845 17623 23903 17629
rect 23934 17620 23940 17672
rect 23992 17660 23998 17672
rect 23992 17632 24037 17660
rect 23992 17620 23998 17632
rect 20588 17564 20944 17592
rect 20588 17552 20594 17564
rect 1762 17524 1768 17536
rect 1723 17496 1768 17524
rect 1762 17484 1768 17496
rect 1820 17484 1826 17536
rect 3142 17524 3148 17536
rect 3103 17496 3148 17524
rect 3142 17484 3148 17496
rect 3200 17484 3206 17536
rect 5258 17484 5264 17536
rect 5316 17524 5322 17536
rect 5445 17527 5503 17533
rect 5445 17524 5457 17527
rect 5316 17496 5457 17524
rect 5316 17484 5322 17496
rect 5445 17493 5457 17496
rect 5491 17493 5503 17527
rect 5445 17487 5503 17493
rect 7929 17527 7987 17533
rect 7929 17493 7941 17527
rect 7975 17524 7987 17527
rect 9125 17527 9183 17533
rect 9125 17524 9137 17527
rect 7975 17496 9137 17524
rect 7975 17493 7987 17496
rect 7929 17487 7987 17493
rect 9125 17493 9137 17496
rect 9171 17524 9183 17527
rect 9214 17524 9220 17536
rect 9171 17496 9220 17524
rect 9171 17493 9183 17496
rect 9125 17487 9183 17493
rect 9214 17484 9220 17496
rect 9272 17484 9278 17536
rect 10962 17484 10968 17536
rect 11020 17524 11026 17536
rect 12250 17524 12256 17536
rect 11020 17496 12256 17524
rect 11020 17484 11026 17496
rect 12250 17484 12256 17496
rect 12308 17484 12314 17536
rect 12434 17484 12440 17536
rect 12492 17524 12498 17536
rect 13262 17524 13268 17536
rect 12492 17496 13268 17524
rect 12492 17484 12498 17496
rect 13262 17484 13268 17496
rect 13320 17484 13326 17536
rect 16114 17484 16120 17536
rect 16172 17524 16178 17536
rect 17034 17524 17040 17536
rect 16172 17496 17040 17524
rect 16172 17484 16178 17496
rect 17034 17484 17040 17496
rect 17092 17484 17098 17536
rect 18414 17524 18420 17536
rect 18375 17496 18420 17524
rect 18414 17484 18420 17496
rect 18472 17484 18478 17536
rect 20349 17527 20407 17533
rect 20349 17493 20361 17527
rect 20395 17524 20407 17527
rect 20717 17527 20775 17533
rect 20717 17524 20729 17527
rect 20395 17496 20729 17524
rect 20395 17493 20407 17496
rect 20349 17487 20407 17493
rect 20717 17493 20729 17496
rect 20763 17524 20775 17527
rect 20806 17524 20812 17536
rect 20763 17496 20812 17524
rect 20763 17493 20775 17496
rect 20717 17487 20775 17493
rect 20806 17484 20812 17496
rect 20864 17484 20870 17536
rect 20916 17524 20944 17564
rect 23385 17595 23443 17601
rect 23385 17561 23397 17595
rect 23431 17592 23443 17595
rect 24964 17592 24992 17691
rect 25682 17592 25688 17604
rect 23431 17564 25688 17592
rect 23431 17561 23443 17564
rect 23385 17555 23443 17561
rect 25682 17552 25688 17564
rect 25740 17552 25746 17604
rect 21634 17524 21640 17536
rect 20916 17496 21640 17524
rect 21634 17484 21640 17496
rect 21692 17484 21698 17536
rect 22186 17484 22192 17536
rect 22244 17524 22250 17536
rect 22281 17527 22339 17533
rect 22281 17524 22293 17527
rect 22244 17496 22293 17524
rect 22244 17484 22250 17496
rect 22281 17493 22293 17496
rect 22327 17493 22339 17527
rect 22281 17487 22339 17493
rect 23014 17484 23020 17536
rect 23072 17524 23078 17536
rect 23293 17527 23351 17533
rect 23293 17524 23305 17527
rect 23072 17496 23305 17524
rect 23072 17484 23078 17496
rect 23293 17493 23305 17496
rect 23339 17524 23351 17527
rect 24489 17527 24547 17533
rect 24489 17524 24501 17527
rect 23339 17496 24501 17524
rect 23339 17493 23351 17496
rect 23293 17487 23351 17493
rect 24489 17493 24501 17496
rect 24535 17524 24547 17527
rect 24670 17524 24676 17536
rect 24535 17496 24676 17524
rect 24535 17493 24547 17496
rect 24489 17487 24547 17493
rect 24670 17484 24676 17496
rect 24728 17484 24734 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1857 17323 1915 17329
rect 1857 17289 1869 17323
rect 1903 17320 1915 17323
rect 2314 17320 2320 17332
rect 1903 17292 2320 17320
rect 1903 17289 1915 17292
rect 1857 17283 1915 17289
rect 2314 17280 2320 17292
rect 2372 17280 2378 17332
rect 4154 17320 4160 17332
rect 4115 17292 4160 17320
rect 4154 17280 4160 17292
rect 4212 17280 4218 17332
rect 5074 17320 5080 17332
rect 5035 17292 5080 17320
rect 5074 17280 5080 17292
rect 5132 17280 5138 17332
rect 7745 17323 7803 17329
rect 7745 17289 7757 17323
rect 7791 17320 7803 17323
rect 8113 17323 8171 17329
rect 8113 17320 8125 17323
rect 7791 17292 8125 17320
rect 7791 17289 7803 17292
rect 7745 17283 7803 17289
rect 8113 17289 8125 17292
rect 8159 17320 8171 17323
rect 8202 17320 8208 17332
rect 8159 17292 8208 17320
rect 8159 17289 8171 17292
rect 8113 17283 8171 17289
rect 8202 17280 8208 17292
rect 8260 17280 8266 17332
rect 8386 17280 8392 17332
rect 8444 17320 8450 17332
rect 10689 17323 10747 17329
rect 10689 17320 10701 17323
rect 8444 17292 10701 17320
rect 8444 17280 8450 17292
rect 10689 17289 10701 17292
rect 10735 17289 10747 17323
rect 10689 17283 10747 17289
rect 13909 17323 13967 17329
rect 13909 17289 13921 17323
rect 13955 17320 13967 17323
rect 13998 17320 14004 17332
rect 13955 17292 14004 17320
rect 13955 17289 13967 17292
rect 13909 17283 13967 17289
rect 5258 17144 5264 17196
rect 5316 17184 5322 17196
rect 5629 17187 5687 17193
rect 5629 17184 5641 17187
rect 5316 17156 5641 17184
rect 5316 17144 5322 17156
rect 5629 17153 5641 17156
rect 5675 17184 5687 17187
rect 6089 17187 6147 17193
rect 6089 17184 6101 17187
rect 5675 17156 6101 17184
rect 5675 17153 5687 17156
rect 5629 17147 5687 17153
rect 6089 17153 6101 17156
rect 6135 17153 6147 17187
rect 8220 17184 8248 17280
rect 9582 17252 9588 17264
rect 9543 17224 9588 17252
rect 9582 17212 9588 17224
rect 9640 17212 9646 17264
rect 13924 17252 13952 17283
rect 13998 17280 14004 17292
rect 14056 17280 14062 17332
rect 15378 17320 15384 17332
rect 15339 17292 15384 17320
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 15746 17280 15752 17332
rect 15804 17320 15810 17332
rect 16301 17323 16359 17329
rect 16301 17320 16313 17323
rect 15804 17292 16313 17320
rect 15804 17280 15810 17292
rect 16301 17289 16313 17292
rect 16347 17289 16359 17323
rect 19426 17320 19432 17332
rect 19387 17292 19432 17320
rect 16301 17283 16359 17289
rect 19426 17280 19432 17292
rect 19484 17280 19490 17332
rect 20073 17323 20131 17329
rect 20073 17289 20085 17323
rect 20119 17320 20131 17323
rect 20622 17320 20628 17332
rect 20119 17292 20628 17320
rect 20119 17289 20131 17292
rect 20073 17283 20131 17289
rect 20622 17280 20628 17292
rect 20680 17280 20686 17332
rect 22738 17320 22744 17332
rect 22699 17292 22744 17320
rect 22738 17280 22744 17292
rect 22796 17280 22802 17332
rect 23477 17323 23535 17329
rect 23477 17289 23489 17323
rect 23523 17320 23535 17323
rect 23934 17320 23940 17332
rect 23523 17292 23940 17320
rect 23523 17289 23535 17292
rect 23477 17283 23535 17289
rect 23934 17280 23940 17292
rect 23992 17320 23998 17332
rect 25133 17323 25191 17329
rect 25133 17320 25145 17323
rect 23992 17292 25145 17320
rect 23992 17280 23998 17292
rect 25133 17289 25145 17292
rect 25179 17289 25191 17323
rect 25682 17320 25688 17332
rect 25643 17292 25688 17320
rect 25133 17283 25191 17289
rect 25682 17280 25688 17292
rect 25740 17280 25746 17332
rect 26142 17320 26148 17332
rect 26103 17292 26148 17320
rect 26142 17280 26148 17292
rect 26200 17280 26206 17332
rect 15930 17252 15936 17264
rect 12176 17224 13952 17252
rect 15891 17224 15936 17252
rect 8220 17156 8340 17184
rect 6089 17147 6147 17153
rect 1949 17119 2007 17125
rect 1949 17085 1961 17119
rect 1995 17116 2007 17119
rect 2038 17116 2044 17128
rect 1995 17088 2044 17116
rect 1995 17085 2007 17088
rect 1949 17079 2007 17085
rect 2038 17076 2044 17088
rect 2096 17076 2102 17128
rect 4430 17076 4436 17128
rect 4488 17116 4494 17128
rect 4985 17119 5043 17125
rect 4985 17116 4997 17119
rect 4488 17088 4997 17116
rect 4488 17076 4494 17088
rect 4985 17085 4997 17088
rect 5031 17116 5043 17119
rect 5537 17119 5595 17125
rect 5537 17116 5549 17119
rect 5031 17088 5549 17116
rect 5031 17085 5043 17088
rect 4985 17079 5043 17085
rect 5537 17085 5549 17088
rect 5583 17085 5595 17119
rect 5537 17079 5595 17085
rect 6730 17076 6736 17128
rect 6788 17116 6794 17128
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 6788 17088 6837 17116
rect 6788 17076 6794 17088
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 8202 17116 8208 17128
rect 8163 17088 8208 17116
rect 6825 17079 6883 17085
rect 8202 17076 8208 17088
rect 8260 17076 8266 17128
rect 8312 17116 8340 17156
rect 9214 17144 9220 17196
rect 9272 17184 9278 17196
rect 10229 17187 10287 17193
rect 10229 17184 10241 17187
rect 9272 17156 10241 17184
rect 9272 17144 9278 17156
rect 10229 17153 10241 17156
rect 10275 17184 10287 17187
rect 11330 17184 11336 17196
rect 10275 17156 11336 17184
rect 10275 17153 10287 17156
rect 10229 17147 10287 17153
rect 11330 17144 11336 17156
rect 11388 17144 11394 17196
rect 12176 17184 12204 17224
rect 15930 17212 15936 17224
rect 15988 17212 15994 17264
rect 11808 17156 12204 17184
rect 12253 17187 12311 17193
rect 8472 17119 8530 17125
rect 8472 17116 8484 17119
rect 8312 17088 8484 17116
rect 8472 17085 8484 17088
rect 8518 17085 8530 17119
rect 8472 17079 8530 17085
rect 10597 17119 10655 17125
rect 10597 17085 10609 17119
rect 10643 17116 10655 17119
rect 11149 17119 11207 17125
rect 11149 17116 11161 17119
rect 10643 17088 11161 17116
rect 10643 17085 10655 17088
rect 10597 17079 10655 17085
rect 11149 17085 11161 17088
rect 11195 17116 11207 17119
rect 11808 17116 11836 17156
rect 12253 17153 12265 17187
rect 12299 17184 12311 17187
rect 12526 17184 12532 17196
rect 12299 17156 12532 17184
rect 12299 17153 12311 17156
rect 12253 17147 12311 17153
rect 12526 17144 12532 17156
rect 12584 17184 12590 17196
rect 12894 17184 12900 17196
rect 12584 17156 12900 17184
rect 12584 17144 12590 17156
rect 12894 17144 12900 17156
rect 12952 17144 12958 17196
rect 13081 17187 13139 17193
rect 13081 17153 13093 17187
rect 13127 17184 13139 17187
rect 13262 17184 13268 17196
rect 13127 17156 13268 17184
rect 13127 17153 13139 17156
rect 13081 17147 13139 17153
rect 13262 17144 13268 17156
rect 13320 17144 13326 17196
rect 20530 17144 20536 17196
rect 20588 17184 20594 17196
rect 20625 17187 20683 17193
rect 20625 17184 20637 17187
rect 20588 17156 20637 17184
rect 20588 17144 20594 17156
rect 20625 17153 20637 17156
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 23661 17187 23719 17193
rect 23661 17153 23673 17187
rect 23707 17184 23719 17187
rect 23753 17187 23811 17193
rect 23753 17184 23765 17187
rect 23707 17156 23765 17184
rect 23707 17153 23719 17156
rect 23661 17147 23719 17153
rect 23753 17153 23765 17156
rect 23799 17153 23811 17187
rect 23753 17147 23811 17153
rect 11195 17088 11836 17116
rect 11885 17119 11943 17125
rect 11195 17085 11207 17088
rect 11149 17079 11207 17085
rect 11885 17085 11897 17119
rect 11931 17116 11943 17119
rect 12066 17116 12072 17128
rect 11931 17088 12072 17116
rect 11931 17085 11943 17088
rect 11885 17079 11943 17085
rect 12066 17076 12072 17088
rect 12124 17116 12130 17128
rect 14274 17125 14280 17128
rect 12805 17119 12863 17125
rect 12805 17116 12817 17119
rect 12124 17088 12817 17116
rect 12124 17076 12130 17088
rect 12805 17085 12817 17088
rect 12851 17085 12863 17119
rect 12805 17079 12863 17085
rect 14001 17119 14059 17125
rect 14001 17085 14013 17119
rect 14047 17085 14059 17119
rect 14268 17116 14280 17125
rect 14235 17088 14280 17116
rect 14001 17079 14059 17085
rect 14268 17079 14280 17088
rect 14332 17116 14338 17128
rect 15194 17116 15200 17128
rect 14332 17088 15200 17116
rect 2216 17051 2274 17057
rect 2216 17017 2228 17051
rect 2262 17048 2274 17051
rect 2774 17048 2780 17060
rect 2262 17020 2780 17048
rect 2262 17017 2274 17020
rect 2216 17011 2274 17017
rect 2774 17008 2780 17020
rect 2832 17008 2838 17060
rect 7098 17048 7104 17060
rect 7059 17020 7104 17048
rect 7098 17008 7104 17020
rect 7156 17008 7162 17060
rect 14016 17048 14044 17079
rect 14274 17076 14280 17079
rect 14332 17076 14338 17088
rect 15194 17076 15200 17088
rect 15252 17076 15258 17128
rect 16482 17116 16488 17128
rect 16443 17088 16488 17116
rect 16482 17076 16488 17088
rect 16540 17076 16546 17128
rect 18049 17119 18107 17125
rect 18049 17085 18061 17119
rect 18095 17116 18107 17119
rect 18138 17116 18144 17128
rect 18095 17088 18144 17116
rect 18095 17085 18107 17088
rect 18049 17079 18107 17085
rect 18138 17076 18144 17088
rect 18196 17076 18202 17128
rect 20714 17076 20720 17128
rect 20772 17116 20778 17128
rect 20892 17119 20950 17125
rect 20892 17116 20904 17119
rect 20772 17088 20904 17116
rect 20772 17076 20778 17088
rect 20892 17085 20904 17088
rect 20938 17116 20950 17119
rect 22186 17116 22192 17128
rect 20938 17088 22192 17116
rect 20938 17085 20950 17088
rect 20892 17079 20950 17085
rect 22186 17076 22192 17088
rect 22244 17076 22250 17128
rect 25222 17116 25228 17128
rect 23032 17088 25228 17116
rect 14734 17048 14740 17060
rect 14016 17020 14740 17048
rect 14734 17008 14740 17020
rect 14792 17008 14798 17060
rect 16761 17051 16819 17057
rect 16761 17017 16773 17051
rect 16807 17048 16819 17051
rect 17586 17048 17592 17060
rect 16807 17020 17592 17048
rect 16807 17017 16819 17020
rect 16761 17011 16819 17017
rect 17586 17008 17592 17020
rect 17644 17008 17650 17060
rect 18294 17051 18352 17057
rect 18294 17048 18306 17051
rect 17788 17020 18306 17048
rect 3326 16980 3332 16992
rect 3287 16952 3332 16980
rect 3326 16940 3332 16952
rect 3384 16940 3390 16992
rect 4617 16983 4675 16989
rect 4617 16949 4629 16983
rect 4663 16980 4675 16983
rect 5445 16983 5503 16989
rect 5445 16980 5457 16983
rect 4663 16952 5457 16980
rect 4663 16949 4675 16952
rect 4617 16943 4675 16949
rect 5445 16949 5457 16952
rect 5491 16980 5503 16983
rect 6178 16980 6184 16992
rect 5491 16952 6184 16980
rect 5491 16949 5503 16952
rect 5445 16943 5503 16949
rect 6178 16940 6184 16952
rect 6236 16940 6242 16992
rect 6638 16980 6644 16992
rect 6599 16952 6644 16980
rect 6638 16940 6644 16952
rect 6696 16940 6702 16992
rect 11054 16980 11060 16992
rect 11015 16952 11060 16980
rect 11054 16940 11060 16952
rect 11112 16940 11118 16992
rect 12437 16983 12495 16989
rect 12437 16949 12449 16983
rect 12483 16980 12495 16983
rect 12710 16980 12716 16992
rect 12483 16952 12716 16980
rect 12483 16949 12495 16952
rect 12437 16943 12495 16949
rect 12710 16940 12716 16952
rect 12768 16940 12774 16992
rect 12894 16980 12900 16992
rect 12855 16952 12900 16980
rect 12894 16940 12900 16952
rect 12952 16940 12958 16992
rect 13541 16983 13599 16989
rect 13541 16949 13553 16983
rect 13587 16980 13599 16983
rect 13722 16980 13728 16992
rect 13587 16952 13728 16980
rect 13587 16949 13599 16952
rect 13541 16943 13599 16949
rect 13722 16940 13728 16952
rect 13780 16940 13786 16992
rect 17313 16983 17371 16989
rect 17313 16949 17325 16983
rect 17359 16980 17371 16983
rect 17402 16980 17408 16992
rect 17359 16952 17408 16980
rect 17359 16949 17371 16952
rect 17313 16943 17371 16949
rect 17402 16940 17408 16952
rect 17460 16940 17466 16992
rect 17678 16940 17684 16992
rect 17736 16980 17742 16992
rect 17788 16989 17816 17020
rect 18294 17017 18306 17020
rect 18340 17048 18352 17051
rect 18414 17048 18420 17060
rect 18340 17020 18420 17048
rect 18340 17017 18352 17020
rect 18294 17011 18352 17017
rect 18414 17008 18420 17020
rect 18472 17008 18478 17060
rect 20346 17008 20352 17060
rect 20404 17048 20410 17060
rect 23032 17048 23060 17088
rect 25222 17076 25228 17088
rect 25280 17076 25286 17128
rect 20404 17020 23060 17048
rect 23109 17051 23167 17057
rect 20404 17008 20410 17020
rect 23109 17017 23121 17051
rect 23155 17048 23167 17051
rect 23998 17051 24056 17057
rect 23998 17048 24010 17051
rect 23155 17020 24010 17048
rect 23155 17017 23167 17020
rect 23109 17011 23167 17017
rect 23998 17017 24010 17020
rect 24044 17048 24056 17051
rect 24302 17048 24308 17060
rect 24044 17020 24308 17048
rect 24044 17017 24056 17020
rect 23998 17011 24056 17017
rect 24302 17008 24308 17020
rect 24360 17008 24366 17060
rect 17773 16983 17831 16989
rect 17773 16980 17785 16983
rect 17736 16952 17785 16980
rect 17736 16940 17742 16952
rect 17773 16949 17785 16952
rect 17819 16949 17831 16983
rect 17773 16943 17831 16949
rect 20533 16983 20591 16989
rect 20533 16949 20545 16983
rect 20579 16980 20591 16983
rect 20806 16980 20812 16992
rect 20579 16952 20812 16980
rect 20579 16949 20591 16952
rect 20533 16943 20591 16949
rect 20806 16940 20812 16952
rect 20864 16980 20870 16992
rect 21174 16980 21180 16992
rect 20864 16952 21180 16980
rect 20864 16940 20870 16952
rect 21174 16940 21180 16952
rect 21232 16940 21238 16992
rect 22002 16980 22008 16992
rect 21963 16952 22008 16980
rect 22002 16940 22008 16952
rect 22060 16940 22066 16992
rect 23661 16983 23719 16989
rect 23661 16949 23673 16983
rect 23707 16980 23719 16983
rect 24670 16980 24676 16992
rect 23707 16952 24676 16980
rect 23707 16949 23719 16952
rect 23661 16943 23719 16949
rect 24670 16940 24676 16952
rect 24728 16980 24734 16992
rect 25222 16980 25228 16992
rect 24728 16952 25228 16980
rect 24728 16940 24734 16952
rect 25222 16940 25228 16952
rect 25280 16940 25286 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1670 16776 1676 16788
rect 1631 16748 1676 16776
rect 1670 16736 1676 16748
rect 1728 16736 1734 16788
rect 3142 16776 3148 16788
rect 2056 16748 3148 16776
rect 2056 16652 2084 16748
rect 3142 16736 3148 16748
rect 3200 16736 3206 16788
rect 3510 16776 3516 16788
rect 3471 16748 3516 16776
rect 3510 16736 3516 16748
rect 3568 16736 3574 16788
rect 3878 16736 3884 16788
rect 3936 16776 3942 16788
rect 4065 16779 4123 16785
rect 4065 16776 4077 16779
rect 3936 16748 4077 16776
rect 3936 16736 3942 16748
rect 4065 16745 4077 16748
rect 4111 16745 4123 16779
rect 4065 16739 4123 16745
rect 6730 16736 6736 16788
rect 6788 16776 6794 16788
rect 7009 16779 7067 16785
rect 7009 16776 7021 16779
rect 6788 16748 7021 16776
rect 6788 16736 6794 16748
rect 7009 16745 7021 16748
rect 7055 16745 7067 16779
rect 7558 16776 7564 16788
rect 7519 16748 7564 16776
rect 7009 16739 7067 16745
rect 7558 16736 7564 16748
rect 7616 16736 7622 16788
rect 8662 16776 8668 16788
rect 8575 16748 8668 16776
rect 8662 16736 8668 16748
rect 8720 16776 8726 16788
rect 9582 16776 9588 16788
rect 8720 16748 9588 16776
rect 8720 16736 8726 16748
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 9858 16776 9864 16788
rect 9819 16748 9864 16776
rect 9858 16736 9864 16748
rect 9916 16736 9922 16788
rect 10413 16779 10471 16785
rect 10413 16745 10425 16779
rect 10459 16776 10471 16779
rect 10778 16776 10784 16788
rect 10459 16748 10784 16776
rect 10459 16745 10471 16748
rect 10413 16739 10471 16745
rect 10778 16736 10784 16748
rect 10836 16736 10842 16788
rect 13630 16776 13636 16788
rect 13591 16748 13636 16776
rect 13630 16736 13636 16748
rect 13688 16736 13694 16788
rect 13998 16776 14004 16788
rect 13959 16748 14004 16776
rect 13998 16736 14004 16748
rect 14056 16736 14062 16788
rect 14090 16736 14096 16788
rect 14148 16776 14154 16788
rect 14148 16748 14193 16776
rect 14148 16736 14154 16748
rect 14826 16736 14832 16788
rect 14884 16776 14890 16788
rect 15289 16779 15347 16785
rect 15289 16776 15301 16779
rect 14884 16748 15301 16776
rect 14884 16736 14890 16748
rect 15289 16745 15301 16748
rect 15335 16745 15347 16779
rect 16482 16776 16488 16788
rect 16443 16748 16488 16776
rect 15289 16739 15347 16745
rect 16482 16736 16488 16748
rect 16540 16736 16546 16788
rect 17313 16779 17371 16785
rect 17313 16745 17325 16779
rect 17359 16776 17371 16779
rect 17865 16779 17923 16785
rect 17865 16776 17877 16779
rect 17359 16748 17877 16776
rect 17359 16745 17371 16748
rect 17313 16739 17371 16745
rect 17865 16745 17877 16748
rect 17911 16776 17923 16779
rect 18969 16779 19027 16785
rect 18969 16776 18981 16779
rect 17911 16748 18981 16776
rect 17911 16745 17923 16748
rect 17865 16739 17923 16745
rect 18969 16745 18981 16748
rect 19015 16745 19027 16779
rect 20714 16776 20720 16788
rect 20675 16748 20720 16776
rect 18969 16739 19027 16745
rect 20714 16736 20720 16748
rect 20772 16736 20778 16788
rect 24026 16776 24032 16788
rect 23987 16748 24032 16776
rect 24026 16736 24032 16748
rect 24084 16776 24090 16788
rect 24213 16779 24271 16785
rect 24213 16776 24225 16779
rect 24084 16748 24225 16776
rect 24084 16736 24090 16748
rect 24213 16745 24225 16748
rect 24259 16745 24271 16779
rect 24213 16739 24271 16745
rect 3789 16711 3847 16717
rect 3789 16708 3801 16711
rect 2148 16680 3801 16708
rect 2148 16652 2176 16680
rect 3789 16677 3801 16680
rect 3835 16677 3847 16711
rect 9490 16708 9496 16720
rect 3789 16671 3847 16677
rect 3896 16680 6500 16708
rect 9451 16680 9496 16708
rect 2038 16640 2044 16652
rect 1999 16612 2044 16640
rect 2038 16600 2044 16612
rect 2096 16600 2102 16652
rect 2130 16600 2136 16652
rect 2188 16640 2194 16652
rect 2498 16640 2504 16652
rect 2188 16612 2233 16640
rect 2332 16612 2504 16640
rect 2188 16600 2194 16612
rect 1946 16532 1952 16584
rect 2004 16572 2010 16584
rect 2225 16575 2283 16581
rect 2225 16572 2237 16575
rect 2004 16544 2237 16572
rect 2004 16532 2010 16544
rect 2225 16541 2237 16544
rect 2271 16572 2283 16575
rect 2332 16572 2360 16612
rect 2498 16600 2504 16612
rect 2556 16640 2562 16652
rect 3145 16643 3203 16649
rect 3145 16640 3157 16643
rect 2556 16612 3157 16640
rect 2556 16600 2562 16612
rect 3145 16609 3157 16612
rect 3191 16640 3203 16643
rect 3326 16640 3332 16652
rect 3191 16612 3332 16640
rect 3191 16609 3203 16612
rect 3145 16603 3203 16609
rect 3326 16600 3332 16612
rect 3384 16600 3390 16652
rect 3896 16584 3924 16680
rect 5350 16649 5356 16652
rect 5344 16640 5356 16649
rect 5263 16612 5356 16640
rect 5344 16603 5356 16612
rect 5408 16640 5414 16652
rect 5408 16612 6132 16640
rect 5350 16600 5356 16603
rect 5408 16600 5414 16612
rect 6104 16584 6132 16612
rect 2774 16572 2780 16584
rect 2271 16544 2360 16572
rect 2687 16544 2780 16572
rect 2271 16541 2283 16544
rect 2225 16535 2283 16541
rect 2774 16532 2780 16544
rect 2832 16572 2838 16584
rect 3878 16572 3884 16584
rect 2832 16544 3884 16572
rect 2832 16532 2838 16544
rect 3878 16532 3884 16544
rect 3936 16532 3942 16584
rect 5077 16575 5135 16581
rect 5077 16572 5089 16575
rect 4908 16544 5089 16572
rect 4617 16439 4675 16445
rect 4617 16405 4629 16439
rect 4663 16436 4675 16439
rect 4706 16436 4712 16448
rect 4663 16408 4712 16436
rect 4663 16405 4675 16408
rect 4617 16399 4675 16405
rect 4706 16396 4712 16408
rect 4764 16436 4770 16448
rect 4908 16445 4936 16544
rect 5077 16541 5089 16544
rect 5123 16541 5135 16575
rect 5077 16535 5135 16541
rect 6086 16532 6092 16584
rect 6144 16532 6150 16584
rect 6472 16513 6500 16680
rect 9490 16668 9496 16680
rect 9548 16668 9554 16720
rect 10689 16711 10747 16717
rect 10689 16677 10701 16711
rect 10735 16708 10747 16711
rect 11054 16708 11060 16720
rect 10735 16680 11060 16708
rect 10735 16677 10747 16680
rect 10689 16671 10747 16677
rect 11054 16668 11060 16680
rect 11112 16708 11118 16720
rect 12158 16708 12164 16720
rect 11112 16680 12164 16708
rect 11112 16668 11118 16680
rect 12158 16668 12164 16680
rect 12216 16668 12222 16720
rect 14550 16668 14556 16720
rect 14608 16708 14614 16720
rect 15013 16711 15071 16717
rect 15013 16708 15025 16711
rect 14608 16680 15025 16708
rect 14608 16668 14614 16680
rect 15013 16677 15025 16680
rect 15059 16677 15071 16711
rect 15013 16671 15071 16677
rect 19337 16711 19395 16717
rect 19337 16677 19349 16711
rect 19383 16708 19395 16711
rect 19426 16708 19432 16720
rect 19383 16680 19432 16708
rect 19383 16677 19395 16680
rect 19337 16671 19395 16677
rect 19426 16668 19432 16680
rect 19484 16668 19490 16720
rect 19518 16668 19524 16720
rect 19576 16708 19582 16720
rect 22002 16717 22008 16720
rect 21453 16711 21511 16717
rect 21453 16708 21465 16711
rect 19576 16680 21465 16708
rect 19576 16668 19582 16680
rect 21453 16677 21465 16680
rect 21499 16677 21511 16711
rect 21996 16708 22008 16717
rect 21963 16680 22008 16708
rect 21453 16671 21511 16677
rect 21996 16671 22008 16680
rect 22002 16668 22008 16671
rect 22060 16668 22066 16720
rect 24581 16711 24639 16717
rect 24581 16677 24593 16711
rect 24627 16708 24639 16711
rect 24670 16708 24676 16720
rect 24627 16680 24676 16708
rect 24627 16677 24639 16680
rect 24581 16671 24639 16677
rect 24670 16668 24676 16680
rect 24728 16668 24734 16720
rect 7650 16600 7656 16652
rect 7708 16640 7714 16652
rect 7929 16643 7987 16649
rect 7929 16640 7941 16643
rect 7708 16612 7941 16640
rect 7708 16600 7714 16612
rect 7929 16609 7941 16612
rect 7975 16640 7987 16643
rect 9398 16640 9404 16652
rect 7975 16612 9404 16640
rect 7975 16609 7987 16612
rect 7929 16603 7987 16609
rect 9398 16600 9404 16612
rect 9456 16600 9462 16652
rect 9674 16640 9680 16652
rect 9635 16612 9680 16640
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 10962 16600 10968 16652
rect 11020 16640 11026 16652
rect 11422 16649 11428 16652
rect 11149 16643 11207 16649
rect 11149 16640 11161 16643
rect 11020 16612 11161 16640
rect 11020 16600 11026 16612
rect 11149 16609 11161 16612
rect 11195 16609 11207 16643
rect 11416 16640 11428 16649
rect 11383 16612 11428 16640
rect 11149 16603 11207 16609
rect 11416 16603 11428 16612
rect 11422 16600 11428 16603
rect 11480 16600 11486 16652
rect 14737 16643 14795 16649
rect 14737 16609 14749 16643
rect 14783 16640 14795 16643
rect 14783 16612 15148 16640
rect 14783 16609 14795 16612
rect 14737 16603 14795 16609
rect 7469 16575 7527 16581
rect 7469 16541 7481 16575
rect 7515 16572 7527 16575
rect 7834 16572 7840 16584
rect 7515 16544 7840 16572
rect 7515 16541 7527 16544
rect 7469 16535 7527 16541
rect 7834 16532 7840 16544
rect 7892 16572 7898 16584
rect 8021 16575 8079 16581
rect 8021 16572 8033 16575
rect 7892 16544 8033 16572
rect 7892 16532 7898 16544
rect 8021 16541 8033 16544
rect 8067 16541 8079 16575
rect 8021 16535 8079 16541
rect 8110 16532 8116 16584
rect 8168 16572 8174 16584
rect 14277 16575 14335 16581
rect 8168 16544 8213 16572
rect 8168 16532 8174 16544
rect 14277 16541 14289 16575
rect 14323 16541 14335 16575
rect 15120 16572 15148 16612
rect 15470 16600 15476 16652
rect 15528 16640 15534 16652
rect 15657 16643 15715 16649
rect 15657 16640 15669 16643
rect 15528 16612 15669 16640
rect 15528 16600 15534 16612
rect 15657 16609 15669 16612
rect 15703 16609 15715 16643
rect 15657 16603 15715 16609
rect 16574 16600 16580 16652
rect 16632 16640 16638 16652
rect 17773 16643 17831 16649
rect 16632 16612 17448 16640
rect 16632 16600 16638 16612
rect 15378 16572 15384 16584
rect 15120 16544 15384 16572
rect 14277 16535 14335 16541
rect 6457 16507 6515 16513
rect 6457 16473 6469 16507
rect 6503 16504 6515 16507
rect 6914 16504 6920 16516
rect 6503 16476 6920 16504
rect 6503 16473 6515 16476
rect 6457 16467 6515 16473
rect 6914 16464 6920 16476
rect 6972 16464 6978 16516
rect 4893 16439 4951 16445
rect 4893 16436 4905 16439
rect 4764 16408 4905 16436
rect 4764 16396 4770 16408
rect 4893 16405 4905 16408
rect 4939 16405 4951 16439
rect 9030 16436 9036 16448
rect 8991 16408 9036 16436
rect 4893 16399 4951 16405
rect 9030 16396 9036 16408
rect 9088 16396 9094 16448
rect 12529 16439 12587 16445
rect 12529 16405 12541 16439
rect 12575 16436 12587 16439
rect 12618 16436 12624 16448
rect 12575 16408 12624 16436
rect 12575 16405 12587 16408
rect 12529 16399 12587 16405
rect 12618 16396 12624 16408
rect 12676 16396 12682 16448
rect 13173 16439 13231 16445
rect 13173 16405 13185 16439
rect 13219 16436 13231 16439
rect 13262 16436 13268 16448
rect 13219 16408 13268 16436
rect 13219 16405 13231 16408
rect 13173 16399 13231 16405
rect 13262 16396 13268 16408
rect 13320 16396 13326 16448
rect 13446 16436 13452 16448
rect 13407 16408 13452 16436
rect 13446 16396 13452 16408
rect 13504 16436 13510 16448
rect 14182 16436 14188 16448
rect 13504 16408 14188 16436
rect 13504 16396 13510 16408
rect 14182 16396 14188 16408
rect 14240 16436 14246 16448
rect 14292 16436 14320 16535
rect 15378 16532 15384 16544
rect 15436 16532 15442 16584
rect 15562 16532 15568 16584
rect 15620 16572 15626 16584
rect 15749 16575 15807 16581
rect 15749 16572 15761 16575
rect 15620 16544 15761 16572
rect 15620 16532 15626 16544
rect 15749 16541 15761 16544
rect 15795 16541 15807 16575
rect 15749 16535 15807 16541
rect 15841 16575 15899 16581
rect 15841 16541 15853 16575
rect 15887 16541 15899 16575
rect 15841 16535 15899 16541
rect 15194 16464 15200 16516
rect 15252 16504 15258 16516
rect 15856 16504 15884 16535
rect 15930 16504 15936 16516
rect 15252 16476 15936 16504
rect 15252 16464 15258 16476
rect 15930 16464 15936 16476
rect 15988 16464 15994 16516
rect 17420 16513 17448 16612
rect 17773 16609 17785 16643
rect 17819 16640 17831 16643
rect 17862 16640 17868 16652
rect 17819 16612 17868 16640
rect 17819 16609 17831 16612
rect 17773 16603 17831 16609
rect 17862 16600 17868 16612
rect 17920 16600 17926 16652
rect 18506 16640 18512 16652
rect 18467 16612 18512 16640
rect 18506 16600 18512 16612
rect 18564 16600 18570 16652
rect 23198 16600 23204 16652
rect 23256 16640 23262 16652
rect 24854 16640 24860 16652
rect 23256 16612 24860 16640
rect 23256 16600 23262 16612
rect 24854 16600 24860 16612
rect 24912 16600 24918 16652
rect 17678 16532 17684 16584
rect 17736 16572 17742 16584
rect 17957 16575 18015 16581
rect 17957 16572 17969 16575
rect 17736 16544 17969 16572
rect 17736 16532 17742 16544
rect 17957 16541 17969 16544
rect 18003 16541 18015 16575
rect 17957 16535 18015 16541
rect 19150 16532 19156 16584
rect 19208 16572 19214 16584
rect 19429 16575 19487 16581
rect 19429 16572 19441 16575
rect 19208 16544 19441 16572
rect 19208 16532 19214 16544
rect 19429 16541 19441 16544
rect 19475 16541 19487 16575
rect 19429 16535 19487 16541
rect 19521 16575 19579 16581
rect 19521 16541 19533 16575
rect 19567 16541 19579 16575
rect 19521 16535 19579 16541
rect 17405 16507 17463 16513
rect 17405 16473 17417 16507
rect 17451 16473 17463 16507
rect 19536 16504 19564 16535
rect 20806 16532 20812 16584
rect 20864 16572 20870 16584
rect 21082 16572 21088 16584
rect 20864 16544 21088 16572
rect 20864 16532 20870 16544
rect 21082 16532 21088 16544
rect 21140 16532 21146 16584
rect 21726 16572 21732 16584
rect 21687 16544 21732 16572
rect 21726 16532 21732 16544
rect 21784 16532 21790 16584
rect 24026 16532 24032 16584
rect 24084 16572 24090 16584
rect 24673 16575 24731 16581
rect 24673 16572 24685 16575
rect 24084 16544 24685 16572
rect 24084 16532 24090 16544
rect 24673 16541 24685 16544
rect 24719 16541 24731 16575
rect 24673 16535 24731 16541
rect 24765 16575 24823 16581
rect 24765 16541 24777 16575
rect 24811 16541 24823 16575
rect 24765 16535 24823 16541
rect 17405 16467 17463 16473
rect 18800 16476 19564 16504
rect 18800 16448 18828 16476
rect 20162 16464 20168 16516
rect 20220 16504 20226 16516
rect 20530 16504 20536 16516
rect 20220 16476 20536 16504
rect 20220 16464 20226 16476
rect 20530 16464 20536 16476
rect 20588 16464 20594 16516
rect 24302 16464 24308 16516
rect 24360 16504 24366 16516
rect 24780 16504 24808 16535
rect 24946 16504 24952 16516
rect 24360 16476 24952 16504
rect 24360 16464 24366 16476
rect 24946 16464 24952 16476
rect 25004 16464 25010 16516
rect 14734 16436 14740 16448
rect 14240 16408 14740 16436
rect 14240 16396 14246 16408
rect 14734 16396 14740 16408
rect 14792 16396 14798 16448
rect 16850 16436 16856 16448
rect 16811 16408 16856 16436
rect 16850 16396 16856 16408
rect 16908 16396 16914 16448
rect 18782 16436 18788 16448
rect 18743 16408 18788 16436
rect 18782 16396 18788 16408
rect 18840 16396 18846 16448
rect 20070 16436 20076 16448
rect 20031 16408 20076 16436
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 21082 16436 21088 16448
rect 21043 16408 21088 16436
rect 21082 16396 21088 16408
rect 21140 16396 21146 16448
rect 23106 16436 23112 16448
rect 23019 16408 23112 16436
rect 23106 16396 23112 16408
rect 23164 16436 23170 16448
rect 23661 16439 23719 16445
rect 23661 16436 23673 16439
rect 23164 16408 23673 16436
rect 23164 16396 23170 16408
rect 23661 16405 23673 16408
rect 23707 16436 23719 16439
rect 23750 16436 23756 16448
rect 23707 16408 23756 16436
rect 23707 16405 23719 16408
rect 23661 16399 23719 16405
rect 23750 16396 23756 16408
rect 23808 16396 23814 16448
rect 24210 16396 24216 16448
rect 24268 16436 24274 16448
rect 24762 16436 24768 16448
rect 24268 16408 24768 16436
rect 24268 16396 24274 16408
rect 24762 16396 24768 16408
rect 24820 16396 24826 16448
rect 25222 16436 25228 16448
rect 25183 16408 25228 16436
rect 25222 16396 25228 16408
rect 25280 16396 25286 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2498 16232 2504 16244
rect 2459 16204 2504 16232
rect 2498 16192 2504 16204
rect 2556 16192 2562 16244
rect 2682 16232 2688 16244
rect 2643 16204 2688 16232
rect 2682 16192 2688 16204
rect 2740 16192 2746 16244
rect 4614 16192 4620 16244
rect 4672 16232 4678 16244
rect 4801 16235 4859 16241
rect 4801 16232 4813 16235
rect 4672 16204 4813 16232
rect 4672 16192 4678 16204
rect 4801 16201 4813 16204
rect 4847 16201 4859 16235
rect 4982 16232 4988 16244
rect 4943 16204 4988 16232
rect 4801 16195 4859 16201
rect 2225 16167 2283 16173
rect 2225 16133 2237 16167
rect 2271 16164 2283 16167
rect 2774 16164 2780 16176
rect 2271 16136 2780 16164
rect 2271 16133 2283 16136
rect 2225 16127 2283 16133
rect 2774 16124 2780 16136
rect 2832 16124 2838 16176
rect 3510 16164 3516 16176
rect 3160 16136 3516 16164
rect 3160 16105 3188 16136
rect 3510 16124 3516 16136
rect 3568 16124 3574 16176
rect 3145 16099 3203 16105
rect 3145 16065 3157 16099
rect 3191 16065 3203 16099
rect 3326 16096 3332 16108
rect 3287 16068 3332 16096
rect 3145 16059 3203 16065
rect 3326 16056 3332 16068
rect 3384 16056 3390 16108
rect 4816 16096 4844 16195
rect 4982 16192 4988 16204
rect 5040 16192 5046 16244
rect 7650 16232 7656 16244
rect 7611 16204 7656 16232
rect 7650 16192 7656 16204
rect 7708 16192 7714 16244
rect 9674 16192 9680 16244
rect 9732 16232 9738 16244
rect 9953 16235 10011 16241
rect 9953 16232 9965 16235
rect 9732 16204 9965 16232
rect 9732 16192 9738 16204
rect 9953 16201 9965 16204
rect 9999 16201 10011 16235
rect 9953 16195 10011 16201
rect 13998 16192 14004 16244
rect 14056 16232 14062 16244
rect 14369 16235 14427 16241
rect 14369 16232 14381 16235
rect 14056 16204 14381 16232
rect 14056 16192 14062 16204
rect 14369 16201 14381 16204
rect 14415 16201 14427 16235
rect 14369 16195 14427 16201
rect 14642 16192 14648 16244
rect 14700 16232 14706 16244
rect 14921 16235 14979 16241
rect 14921 16232 14933 16235
rect 14700 16204 14933 16232
rect 14700 16192 14706 16204
rect 14921 16201 14933 16204
rect 14967 16201 14979 16235
rect 15930 16232 15936 16244
rect 15891 16204 15936 16232
rect 14921 16195 14979 16201
rect 15930 16192 15936 16204
rect 15988 16192 15994 16244
rect 19518 16192 19524 16244
rect 19576 16232 19582 16244
rect 19889 16235 19947 16241
rect 19889 16232 19901 16235
rect 19576 16204 19901 16232
rect 19576 16192 19582 16204
rect 19889 16201 19901 16204
rect 19935 16201 19947 16235
rect 19889 16195 19947 16201
rect 21269 16235 21327 16241
rect 21269 16201 21281 16235
rect 21315 16232 21327 16235
rect 22002 16232 22008 16244
rect 21315 16204 22008 16232
rect 21315 16201 21327 16204
rect 21269 16195 21327 16201
rect 7006 16164 7012 16176
rect 6967 16136 7012 16164
rect 7006 16124 7012 16136
rect 7064 16124 7070 16176
rect 10689 16167 10747 16173
rect 10689 16133 10701 16167
rect 10735 16164 10747 16167
rect 14734 16164 14740 16176
rect 10735 16136 11468 16164
rect 14695 16136 14740 16164
rect 10735 16133 10747 16136
rect 10689 16127 10747 16133
rect 11440 16108 11468 16136
rect 14734 16124 14740 16136
rect 14792 16124 14798 16176
rect 5445 16099 5503 16105
rect 5445 16096 5457 16099
rect 4816 16068 5457 16096
rect 5445 16065 5457 16068
rect 5491 16065 5503 16099
rect 5445 16059 5503 16065
rect 5537 16099 5595 16105
rect 5537 16065 5549 16099
rect 5583 16065 5595 16099
rect 6086 16096 6092 16108
rect 5999 16068 6092 16096
rect 5537 16059 5595 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 4157 16031 4215 16037
rect 1443 16000 3832 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 1670 15960 1676 15972
rect 1631 15932 1676 15960
rect 1670 15920 1676 15932
rect 1728 15920 1734 15972
rect 3053 15963 3111 15969
rect 3053 15929 3065 15963
rect 3099 15960 3111 15963
rect 3326 15960 3332 15972
rect 3099 15932 3332 15960
rect 3099 15929 3111 15932
rect 3053 15923 3111 15929
rect 3326 15920 3332 15932
rect 3384 15920 3390 15972
rect 3804 15904 3832 16000
rect 4157 15997 4169 16031
rect 4203 16028 4215 16031
rect 5258 16028 5264 16040
rect 4203 16000 5264 16028
rect 4203 15997 4215 16000
rect 4157 15991 4215 15997
rect 5258 15988 5264 16000
rect 5316 16028 5322 16040
rect 5552 16028 5580 16059
rect 6086 16056 6092 16068
rect 6144 16096 6150 16108
rect 7190 16096 7196 16108
rect 6144 16068 7196 16096
rect 6144 16056 6150 16068
rect 7190 16056 7196 16068
rect 7248 16056 7254 16108
rect 10778 16056 10784 16108
rect 10836 16096 10842 16108
rect 11241 16099 11299 16105
rect 11241 16096 11253 16099
rect 10836 16068 11253 16096
rect 10836 16056 10842 16068
rect 11241 16065 11253 16068
rect 11287 16065 11299 16099
rect 11422 16096 11428 16108
rect 11335 16068 11428 16096
rect 11241 16059 11299 16065
rect 11422 16056 11428 16068
rect 11480 16096 11486 16108
rect 11882 16096 11888 16108
rect 11480 16068 11888 16096
rect 11480 16056 11486 16068
rect 11882 16056 11888 16068
rect 11940 16056 11946 16108
rect 15565 16099 15623 16105
rect 15565 16065 15577 16099
rect 15611 16096 15623 16099
rect 16022 16096 16028 16108
rect 15611 16068 16028 16096
rect 15611 16065 15623 16068
rect 15565 16059 15623 16065
rect 16022 16056 16028 16068
rect 16080 16056 16086 16108
rect 16942 16096 16948 16108
rect 16903 16068 16948 16096
rect 16942 16056 16948 16068
rect 17000 16056 17006 16108
rect 17402 16056 17408 16108
rect 17460 16096 17466 16108
rect 18601 16099 18659 16105
rect 18601 16096 18613 16099
rect 17460 16068 18613 16096
rect 17460 16056 17466 16068
rect 18601 16065 18613 16068
rect 18647 16096 18659 16099
rect 18782 16096 18788 16108
rect 18647 16068 18788 16096
rect 18647 16065 18659 16068
rect 18601 16059 18659 16065
rect 18782 16056 18788 16068
rect 18840 16056 18846 16108
rect 20070 16056 20076 16108
rect 20128 16096 20134 16108
rect 20533 16099 20591 16105
rect 20533 16096 20545 16099
rect 20128 16068 20545 16096
rect 20128 16056 20134 16068
rect 20533 16065 20545 16068
rect 20579 16096 20591 16099
rect 21284 16096 21312 16195
rect 22002 16192 22008 16204
rect 22060 16192 22066 16244
rect 23106 16232 23112 16244
rect 22664 16204 23112 16232
rect 21726 16164 21732 16176
rect 21639 16136 21732 16164
rect 21726 16124 21732 16136
rect 21784 16164 21790 16176
rect 21784 16136 22039 16164
rect 21784 16124 21790 16136
rect 20579 16068 21312 16096
rect 20579 16065 20591 16068
rect 20533 16059 20591 16065
rect 5316 16000 5580 16028
rect 6641 16031 6699 16037
rect 5316 15988 5322 16000
rect 6641 15997 6653 16031
rect 6687 16028 6699 16031
rect 6822 16028 6828 16040
rect 6687 16000 6828 16028
rect 6687 15997 6699 16000
rect 6641 15991 6699 15997
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 8021 16031 8079 16037
rect 8021 15997 8033 16031
rect 8067 15997 8079 16031
rect 8021 15991 8079 15997
rect 8288 16031 8346 16037
rect 8288 15997 8300 16031
rect 8334 16028 8346 16031
rect 8662 16028 8668 16040
rect 8334 16000 8668 16028
rect 8334 15997 8346 16000
rect 8288 15991 8346 15997
rect 5353 15963 5411 15969
rect 5353 15960 5365 15963
rect 4448 15932 5365 15960
rect 3786 15892 3792 15904
rect 3747 15864 3792 15892
rect 3786 15852 3792 15864
rect 3844 15852 3850 15904
rect 4246 15852 4252 15904
rect 4304 15892 4310 15904
rect 4448 15901 4476 15932
rect 5353 15929 5365 15932
rect 5399 15929 5411 15963
rect 5353 15923 5411 15929
rect 7926 15920 7932 15972
rect 7984 15960 7990 15972
rect 8036 15960 8064 15991
rect 8662 15988 8668 16000
rect 8720 15988 8726 16040
rect 10042 15988 10048 16040
rect 10100 16028 10106 16040
rect 11149 16031 11207 16037
rect 11149 16028 11161 16031
rect 10100 16000 11161 16028
rect 10100 15988 10106 16000
rect 11149 15997 11161 16000
rect 11195 16028 11207 16031
rect 12342 16028 12348 16040
rect 11195 16000 12348 16028
rect 11195 15997 11207 16000
rect 11149 15991 11207 15997
rect 12342 15988 12348 16000
rect 12400 15988 12406 16040
rect 12437 16031 12495 16037
rect 12437 15997 12449 16031
rect 12483 16028 12495 16031
rect 12526 16028 12532 16040
rect 12483 16000 12532 16028
rect 12483 15997 12495 16000
rect 12437 15991 12495 15997
rect 12526 15988 12532 16000
rect 12584 15988 12590 16040
rect 12704 16031 12762 16037
rect 12704 16028 12716 16031
rect 12636 16000 12716 16028
rect 12636 15972 12664 16000
rect 12704 15997 12716 16000
rect 12750 16028 12762 16031
rect 13538 16028 13544 16040
rect 12750 16000 13544 16028
rect 12750 15997 12762 16000
rect 12704 15991 12762 15997
rect 13538 15988 13544 16000
rect 13596 15988 13602 16040
rect 16669 16031 16727 16037
rect 16669 15997 16681 16031
rect 16715 16028 16727 16031
rect 16850 16028 16856 16040
rect 16715 16000 16856 16028
rect 16715 15997 16727 16000
rect 16669 15991 16727 15997
rect 16850 15988 16856 16000
rect 16908 15988 16914 16040
rect 18046 15988 18052 16040
rect 18104 16028 18110 16040
rect 18417 16031 18475 16037
rect 18417 16028 18429 16031
rect 18104 16000 18429 16028
rect 18104 15988 18110 16000
rect 18417 15997 18429 16000
rect 18463 15997 18475 16031
rect 18417 15991 18475 15997
rect 20349 16031 20407 16037
rect 20349 15997 20361 16031
rect 20395 16028 20407 16031
rect 20622 16028 20628 16040
rect 20395 16000 20628 16028
rect 20395 15997 20407 16000
rect 20349 15991 20407 15997
rect 20622 15988 20628 16000
rect 20680 15988 20686 16040
rect 21726 15988 21732 16040
rect 21784 16028 21790 16040
rect 21913 16031 21971 16037
rect 21913 16028 21925 16031
rect 21784 16000 21925 16028
rect 21784 15988 21790 16000
rect 21913 15997 21925 16000
rect 21959 15997 21971 16031
rect 22011 16028 22039 16136
rect 22370 16056 22376 16108
rect 22428 16096 22434 16108
rect 22664 16105 22692 16204
rect 23106 16192 23112 16204
rect 23164 16192 23170 16244
rect 23477 16235 23535 16241
rect 23477 16201 23489 16235
rect 23523 16232 23535 16235
rect 24026 16232 24032 16244
rect 23523 16204 24032 16232
rect 23523 16201 23535 16204
rect 23477 16195 23535 16201
rect 24026 16192 24032 16204
rect 24084 16192 24090 16244
rect 24946 16192 24952 16244
rect 25004 16232 25010 16244
rect 25041 16235 25099 16241
rect 25041 16232 25053 16235
rect 25004 16204 25053 16232
rect 25004 16192 25010 16204
rect 25041 16201 25053 16204
rect 25087 16201 25099 16235
rect 25041 16195 25099 16201
rect 22465 16099 22523 16105
rect 22465 16096 22477 16099
rect 22428 16068 22477 16096
rect 22428 16056 22434 16068
rect 22465 16065 22477 16068
rect 22511 16065 22523 16099
rect 22465 16059 22523 16065
rect 22649 16099 22707 16105
rect 22649 16065 22661 16099
rect 22695 16065 22707 16099
rect 22649 16059 22707 16065
rect 23661 16031 23719 16037
rect 23661 16028 23673 16031
rect 22011 16000 23673 16028
rect 21913 15991 21971 15997
rect 23661 15997 23673 16000
rect 23707 15997 23719 16031
rect 23661 15991 23719 15997
rect 8202 15960 8208 15972
rect 7984 15932 8208 15960
rect 7984 15920 7990 15932
rect 8202 15920 8208 15932
rect 8260 15960 8266 15972
rect 9030 15960 9036 15972
rect 8260 15932 9036 15960
rect 8260 15920 8266 15932
rect 9030 15920 9036 15932
rect 9088 15920 9094 15972
rect 12253 15963 12311 15969
rect 12253 15929 12265 15963
rect 12299 15960 12311 15963
rect 12618 15960 12624 15972
rect 12299 15932 12624 15960
rect 12299 15929 12311 15932
rect 12253 15923 12311 15929
rect 12618 15920 12624 15932
rect 12676 15920 12682 15972
rect 14642 15920 14648 15972
rect 14700 15960 14706 15972
rect 15289 15963 15347 15969
rect 15289 15960 15301 15963
rect 14700 15932 15301 15960
rect 14700 15920 14706 15932
rect 15289 15929 15301 15932
rect 15335 15929 15347 15963
rect 15289 15923 15347 15929
rect 15470 15920 15476 15972
rect 15528 15960 15534 15972
rect 16301 15963 16359 15969
rect 16301 15960 16313 15963
rect 15528 15932 16313 15960
rect 15528 15920 15534 15932
rect 16301 15929 16313 15932
rect 16347 15929 16359 15963
rect 18509 15963 18567 15969
rect 18509 15960 18521 15963
rect 16301 15923 16359 15929
rect 17788 15932 18521 15960
rect 17788 15904 17816 15932
rect 18509 15929 18521 15932
rect 18555 15929 18567 15963
rect 18509 15923 18567 15929
rect 20257 15963 20315 15969
rect 20257 15929 20269 15963
rect 20303 15960 20315 15963
rect 21082 15960 21088 15972
rect 20303 15932 21088 15960
rect 20303 15929 20315 15932
rect 20257 15923 20315 15929
rect 21082 15920 21088 15932
rect 21140 15920 21146 15972
rect 21450 15920 21456 15972
rect 21508 15960 21514 15972
rect 21545 15963 21603 15969
rect 21545 15960 21557 15963
rect 21508 15932 21557 15960
rect 21508 15920 21514 15932
rect 21545 15929 21557 15932
rect 21591 15960 21603 15963
rect 21818 15960 21824 15972
rect 21591 15932 21824 15960
rect 21591 15929 21603 15932
rect 21545 15923 21603 15929
rect 21818 15920 21824 15932
rect 21876 15960 21882 15972
rect 22373 15963 22431 15969
rect 22373 15960 22385 15963
rect 21876 15932 22385 15960
rect 21876 15920 21882 15932
rect 22373 15929 22385 15932
rect 22419 15929 22431 15963
rect 22373 15923 22431 15929
rect 4433 15895 4491 15901
rect 4433 15892 4445 15895
rect 4304 15864 4445 15892
rect 4304 15852 4310 15864
rect 4433 15861 4445 15864
rect 4479 15861 4491 15895
rect 4433 15855 4491 15861
rect 8570 15852 8576 15904
rect 8628 15892 8634 15904
rect 9401 15895 9459 15901
rect 9401 15892 9413 15895
rect 8628 15864 9413 15892
rect 8628 15852 8634 15864
rect 9401 15861 9413 15864
rect 9447 15861 9459 15895
rect 10778 15892 10784 15904
rect 10739 15864 10784 15892
rect 9401 15855 9459 15861
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 11882 15892 11888 15904
rect 11843 15864 11888 15892
rect 11882 15852 11888 15864
rect 11940 15852 11946 15904
rect 13262 15852 13268 15904
rect 13320 15892 13326 15904
rect 13817 15895 13875 15901
rect 13817 15892 13829 15895
rect 13320 15864 13829 15892
rect 13320 15852 13326 15864
rect 13817 15861 13829 15864
rect 13863 15861 13875 15895
rect 13817 15855 13875 15861
rect 15378 15852 15384 15904
rect 15436 15892 15442 15904
rect 17402 15892 17408 15904
rect 15436 15864 15481 15892
rect 17363 15864 17408 15892
rect 15436 15852 15442 15864
rect 17402 15852 17408 15864
rect 17460 15852 17466 15904
rect 17770 15892 17776 15904
rect 17731 15864 17776 15892
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 17954 15852 17960 15904
rect 18012 15892 18018 15904
rect 18049 15895 18107 15901
rect 18049 15892 18061 15895
rect 18012 15864 18061 15892
rect 18012 15852 18018 15864
rect 18049 15861 18061 15864
rect 18095 15861 18107 15895
rect 19150 15892 19156 15904
rect 19111 15864 19156 15892
rect 18049 15855 18107 15861
rect 19150 15852 19156 15864
rect 19208 15852 19214 15904
rect 19426 15892 19432 15904
rect 19387 15864 19432 15892
rect 19426 15852 19432 15864
rect 19484 15852 19490 15904
rect 22002 15892 22008 15904
rect 21963 15864 22008 15892
rect 22002 15852 22008 15864
rect 22060 15852 22066 15904
rect 23676 15892 23704 15991
rect 23750 15988 23756 16040
rect 23808 16028 23814 16040
rect 23917 16031 23975 16037
rect 23917 16028 23929 16031
rect 23808 16000 23929 16028
rect 23808 15988 23814 16000
rect 23917 15997 23929 16000
rect 23963 15997 23975 16031
rect 23917 15991 23975 15997
rect 23934 15892 23940 15904
rect 23676 15864 23940 15892
rect 23934 15852 23940 15864
rect 23992 15892 23998 15904
rect 25222 15892 25228 15904
rect 23992 15864 25228 15892
rect 23992 15852 23998 15864
rect 25222 15852 25228 15864
rect 25280 15892 25286 15904
rect 25593 15895 25651 15901
rect 25593 15892 25605 15895
rect 25280 15864 25605 15892
rect 25280 15852 25286 15864
rect 25593 15861 25605 15864
rect 25639 15861 25651 15895
rect 25593 15855 25651 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1765 15691 1823 15697
rect 1765 15657 1777 15691
rect 1811 15688 1823 15691
rect 2038 15688 2044 15700
rect 1811 15660 2044 15688
rect 1811 15657 1823 15660
rect 1765 15651 1823 15657
rect 2038 15648 2044 15660
rect 2096 15648 2102 15700
rect 2406 15648 2412 15700
rect 2464 15688 2470 15700
rect 2774 15688 2780 15700
rect 2464 15660 2780 15688
rect 2464 15648 2470 15660
rect 2774 15648 2780 15660
rect 2832 15648 2838 15700
rect 3234 15648 3240 15700
rect 3292 15688 3298 15700
rect 6825 15691 6883 15697
rect 6825 15688 6837 15691
rect 3292 15660 6837 15688
rect 3292 15648 3298 15660
rect 6825 15657 6837 15660
rect 6871 15657 6883 15691
rect 6825 15651 6883 15657
rect 7834 15648 7840 15700
rect 7892 15688 7898 15700
rect 7929 15691 7987 15697
rect 7929 15688 7941 15691
rect 7892 15660 7941 15688
rect 7892 15648 7898 15660
rect 7929 15657 7941 15660
rect 7975 15657 7987 15691
rect 8294 15688 8300 15700
rect 8207 15660 8300 15688
rect 7929 15651 7987 15657
rect 8294 15648 8300 15660
rect 8352 15688 8358 15700
rect 8754 15688 8760 15700
rect 8352 15660 8760 15688
rect 8352 15648 8358 15660
rect 8754 15648 8760 15660
rect 8812 15648 8818 15700
rect 10042 15688 10048 15700
rect 10003 15660 10048 15688
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 10962 15688 10968 15700
rect 10336 15660 10968 15688
rect 4985 15623 5043 15629
rect 4985 15589 4997 15623
rect 5031 15620 5043 15623
rect 6086 15620 6092 15632
rect 5031 15592 6092 15620
rect 5031 15589 5043 15592
rect 4985 15583 5043 15589
rect 6086 15580 6092 15592
rect 6144 15580 6150 15632
rect 6181 15623 6239 15629
rect 6181 15589 6193 15623
rect 6227 15620 6239 15623
rect 6457 15623 6515 15629
rect 6457 15620 6469 15623
rect 6227 15592 6469 15620
rect 6227 15589 6239 15592
rect 6181 15583 6239 15589
rect 6457 15589 6469 15592
rect 6503 15589 6515 15623
rect 6457 15583 6515 15589
rect 7469 15623 7527 15629
rect 7469 15589 7481 15623
rect 7515 15620 7527 15623
rect 8110 15620 8116 15632
rect 7515 15592 8116 15620
rect 7515 15589 7527 15592
rect 7469 15583 7527 15589
rect 1673 15555 1731 15561
rect 1673 15521 1685 15555
rect 1719 15552 1731 15555
rect 1762 15552 1768 15564
rect 1719 15524 1768 15552
rect 1719 15521 1731 15524
rect 1673 15515 1731 15521
rect 1762 15512 1768 15524
rect 1820 15512 1826 15564
rect 1854 15512 1860 15564
rect 1912 15552 1918 15564
rect 2133 15555 2191 15561
rect 2133 15552 2145 15555
rect 1912 15524 2145 15552
rect 1912 15512 1918 15524
rect 2133 15521 2145 15524
rect 2179 15552 2191 15555
rect 4065 15555 4123 15561
rect 4065 15552 4077 15555
rect 2179 15524 4077 15552
rect 2179 15521 2191 15524
rect 2133 15515 2191 15521
rect 4065 15521 4077 15524
rect 4111 15521 4123 15555
rect 5442 15552 5448 15564
rect 5403 15524 5448 15552
rect 4065 15515 4123 15521
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 1946 15444 1952 15496
rect 2004 15484 2010 15496
rect 2222 15484 2228 15496
rect 2004 15456 2228 15484
rect 2004 15444 2010 15456
rect 2222 15444 2228 15456
rect 2280 15444 2286 15496
rect 2406 15444 2412 15496
rect 2464 15484 2470 15496
rect 2464 15456 2509 15484
rect 2464 15444 2470 15456
rect 5166 15444 5172 15496
rect 5224 15484 5230 15496
rect 5537 15487 5595 15493
rect 5537 15484 5549 15487
rect 5224 15456 5549 15484
rect 5224 15444 5230 15456
rect 5537 15453 5549 15456
rect 5583 15453 5595 15487
rect 5537 15447 5595 15453
rect 5626 15444 5632 15496
rect 5684 15484 5690 15496
rect 5684 15456 5729 15484
rect 5684 15444 5690 15456
rect 4617 15419 4675 15425
rect 4617 15385 4629 15419
rect 4663 15416 4675 15419
rect 4706 15416 4712 15428
rect 4663 15388 4712 15416
rect 4663 15385 4675 15388
rect 4617 15379 4675 15385
rect 4706 15376 4712 15388
rect 4764 15416 4770 15428
rect 5258 15416 5264 15428
rect 4764 15388 5264 15416
rect 4764 15376 4770 15388
rect 5258 15376 5264 15388
rect 5316 15376 5322 15428
rect 3234 15348 3240 15360
rect 3195 15320 3240 15348
rect 3234 15308 3240 15320
rect 3292 15308 3298 15360
rect 3326 15308 3332 15360
rect 3384 15348 3390 15360
rect 3513 15351 3571 15357
rect 3513 15348 3525 15351
rect 3384 15320 3525 15348
rect 3384 15308 3390 15320
rect 3513 15317 3525 15320
rect 3559 15317 3571 15351
rect 5074 15348 5080 15360
rect 5035 15320 5080 15348
rect 3513 15311 3571 15317
rect 5074 15308 5080 15320
rect 5132 15308 5138 15360
rect 6472 15348 6500 15583
rect 8110 15580 8116 15592
rect 8168 15580 8174 15632
rect 6638 15552 6644 15564
rect 6599 15524 6644 15552
rect 6638 15512 6644 15524
rect 6696 15512 6702 15564
rect 7650 15512 7656 15564
rect 7708 15552 7714 15564
rect 8389 15555 8447 15561
rect 8389 15552 8401 15555
rect 7708 15524 8401 15552
rect 7708 15512 7714 15524
rect 8389 15521 8401 15524
rect 8435 15552 8447 15555
rect 8662 15552 8668 15564
rect 8435 15524 8668 15552
rect 8435 15521 8447 15524
rect 8389 15515 8447 15521
rect 8662 15512 8668 15524
rect 8720 15512 8726 15564
rect 9030 15552 9036 15564
rect 8943 15524 9036 15552
rect 9030 15512 9036 15524
rect 9088 15552 9094 15564
rect 9398 15552 9404 15564
rect 9088 15524 9404 15552
rect 9088 15512 9094 15524
rect 9398 15512 9404 15524
rect 9456 15552 9462 15564
rect 9493 15555 9551 15561
rect 9493 15552 9505 15555
rect 9456 15524 9505 15552
rect 9456 15512 9462 15524
rect 9493 15521 9505 15524
rect 9539 15552 9551 15555
rect 10336 15552 10364 15660
rect 10962 15648 10968 15660
rect 11020 15648 11026 15700
rect 13446 15688 13452 15700
rect 13407 15660 13452 15688
rect 13446 15648 13452 15660
rect 13504 15688 13510 15700
rect 13906 15688 13912 15700
rect 13504 15660 13912 15688
rect 13504 15648 13510 15660
rect 13906 15648 13912 15660
rect 13964 15648 13970 15700
rect 14090 15688 14096 15700
rect 14051 15660 14096 15688
rect 14090 15648 14096 15660
rect 14148 15648 14154 15700
rect 17129 15691 17187 15697
rect 17129 15657 17141 15691
rect 17175 15688 17187 15691
rect 17402 15688 17408 15700
rect 17175 15660 17408 15688
rect 17175 15657 17187 15660
rect 17129 15651 17187 15657
rect 17402 15648 17408 15660
rect 17460 15648 17466 15700
rect 17678 15688 17684 15700
rect 17639 15660 17684 15688
rect 17678 15648 17684 15660
rect 17736 15648 17742 15700
rect 20901 15691 20959 15697
rect 20901 15657 20913 15691
rect 20947 15688 20959 15691
rect 21082 15688 21088 15700
rect 20947 15660 21088 15688
rect 20947 15657 20959 15660
rect 20901 15651 20959 15657
rect 21082 15648 21088 15660
rect 21140 15648 21146 15700
rect 22094 15648 22100 15700
rect 22152 15688 22158 15700
rect 22649 15691 22707 15697
rect 22649 15688 22661 15691
rect 22152 15660 22661 15688
rect 22152 15648 22158 15660
rect 22649 15657 22661 15660
rect 22695 15657 22707 15691
rect 23474 15688 23480 15700
rect 23435 15660 23480 15688
rect 22649 15651 22707 15657
rect 23474 15648 23480 15660
rect 23532 15688 23538 15700
rect 24029 15691 24087 15697
rect 24029 15688 24041 15691
rect 23532 15660 24041 15688
rect 23532 15648 23538 15660
rect 24029 15657 24041 15660
rect 24075 15657 24087 15691
rect 24946 15688 24952 15700
rect 24907 15660 24952 15688
rect 24029 15651 24087 15657
rect 24946 15648 24952 15660
rect 25004 15648 25010 15700
rect 10413 15623 10471 15629
rect 10413 15589 10425 15623
rect 10459 15620 10471 15623
rect 10686 15620 10692 15632
rect 10459 15592 10692 15620
rect 10459 15589 10471 15592
rect 10413 15583 10471 15589
rect 10686 15580 10692 15592
rect 10744 15629 10750 15632
rect 10744 15623 10808 15629
rect 10744 15589 10762 15623
rect 10796 15620 10808 15623
rect 12805 15623 12863 15629
rect 12805 15620 12817 15623
rect 10796 15592 12817 15620
rect 10796 15589 10808 15592
rect 10744 15583 10808 15589
rect 12805 15589 12817 15592
rect 12851 15620 12863 15623
rect 13078 15620 13084 15632
rect 12851 15592 13084 15620
rect 12851 15589 12863 15592
rect 12805 15583 12863 15589
rect 10744 15580 10750 15583
rect 13078 15580 13084 15592
rect 13136 15580 13142 15632
rect 18500 15623 18558 15629
rect 18500 15589 18512 15623
rect 18546 15620 18558 15623
rect 18598 15620 18604 15632
rect 18546 15592 18604 15620
rect 18546 15589 18558 15592
rect 18500 15583 18558 15589
rect 18598 15580 18604 15592
rect 18656 15580 18662 15632
rect 21358 15580 21364 15632
rect 21416 15580 21422 15632
rect 21450 15580 21456 15632
rect 21508 15620 21514 15632
rect 21726 15620 21732 15632
rect 21508 15592 21732 15620
rect 21508 15580 21514 15592
rect 21726 15580 21732 15592
rect 21784 15620 21790 15632
rect 23017 15623 23075 15629
rect 23017 15620 23029 15623
rect 21784 15592 23029 15620
rect 21784 15580 21790 15592
rect 23017 15589 23029 15592
rect 23063 15589 23075 15623
rect 24578 15620 24584 15632
rect 24539 15592 24584 15620
rect 23017 15583 23075 15589
rect 24578 15580 24584 15592
rect 24636 15580 24642 15632
rect 10505 15555 10563 15561
rect 10505 15552 10517 15555
rect 9539 15524 10517 15552
rect 9539 15521 9551 15524
rect 9493 15515 9551 15521
rect 10505 15521 10517 15524
rect 10551 15521 10563 15555
rect 10505 15515 10563 15521
rect 12526 15512 12532 15564
rect 12584 15552 12590 15564
rect 13357 15555 13415 15561
rect 13357 15552 13369 15555
rect 12584 15524 13369 15552
rect 12584 15512 12590 15524
rect 13357 15521 13369 15524
rect 13403 15552 13415 15555
rect 13722 15552 13728 15564
rect 13403 15524 13728 15552
rect 13403 15521 13415 15524
rect 13357 15515 13415 15521
rect 13722 15512 13728 15524
rect 13780 15512 13786 15564
rect 16022 15561 16028 15564
rect 15013 15555 15071 15561
rect 15013 15521 15025 15555
rect 15059 15552 15071 15555
rect 16016 15552 16028 15561
rect 15059 15524 16028 15552
rect 15059 15521 15071 15524
rect 15013 15515 15071 15521
rect 16016 15515 16028 15524
rect 16022 15512 16028 15515
rect 16080 15512 16086 15564
rect 20717 15555 20775 15561
rect 20717 15521 20729 15555
rect 20763 15552 20775 15555
rect 20898 15552 20904 15564
rect 20763 15524 20904 15552
rect 20763 15521 20775 15524
rect 20717 15515 20775 15521
rect 20898 15512 20904 15524
rect 20956 15552 20962 15564
rect 21269 15555 21327 15561
rect 21269 15552 21281 15555
rect 20956 15524 21281 15552
rect 20956 15512 20962 15524
rect 21269 15521 21281 15524
rect 21315 15521 21327 15555
rect 21376 15552 21404 15580
rect 22094 15552 22100 15564
rect 21376 15524 22100 15552
rect 21269 15515 21327 15521
rect 22094 15512 22100 15524
rect 22152 15512 22158 15564
rect 22462 15552 22468 15564
rect 22423 15524 22468 15552
rect 22462 15512 22468 15524
rect 22520 15512 22526 15564
rect 23750 15512 23756 15564
rect 23808 15552 23814 15564
rect 23937 15555 23995 15561
rect 23937 15552 23949 15555
rect 23808 15524 23949 15552
rect 23808 15512 23814 15524
rect 23937 15521 23949 15524
rect 23983 15521 23995 15555
rect 25130 15552 25136 15564
rect 25091 15524 25136 15552
rect 23937 15515 23995 15521
rect 25130 15512 25136 15524
rect 25188 15512 25194 15564
rect 8570 15484 8576 15496
rect 8531 15456 8576 15484
rect 8570 15444 8576 15456
rect 8628 15444 8634 15496
rect 13538 15484 13544 15496
rect 13499 15456 13544 15484
rect 13538 15444 13544 15456
rect 13596 15444 13602 15496
rect 15286 15444 15292 15496
rect 15344 15484 15350 15496
rect 15749 15487 15807 15493
rect 15749 15484 15761 15487
rect 15344 15456 15761 15484
rect 15344 15444 15350 15456
rect 15749 15453 15761 15456
rect 15795 15453 15807 15487
rect 15749 15447 15807 15453
rect 18138 15444 18144 15496
rect 18196 15484 18202 15496
rect 18233 15487 18291 15493
rect 18233 15484 18245 15487
rect 18196 15456 18245 15484
rect 18196 15444 18202 15456
rect 18233 15453 18245 15456
rect 18279 15453 18291 15487
rect 21358 15484 21364 15496
rect 21319 15456 21364 15484
rect 18233 15447 18291 15453
rect 21358 15444 21364 15456
rect 21416 15444 21422 15496
rect 21545 15487 21603 15493
rect 21545 15453 21557 15487
rect 21591 15453 21603 15487
rect 21545 15447 21603 15453
rect 24213 15487 24271 15493
rect 24213 15453 24225 15487
rect 24259 15484 24271 15487
rect 24670 15484 24676 15496
rect 24259 15456 24676 15484
rect 24259 15453 24271 15456
rect 24213 15447 24271 15453
rect 7837 15419 7895 15425
rect 7837 15385 7849 15419
rect 7883 15416 7895 15419
rect 8110 15416 8116 15428
rect 7883 15388 8116 15416
rect 7883 15385 7895 15388
rect 7837 15379 7895 15385
rect 8110 15376 8116 15388
rect 8168 15416 8174 15428
rect 8588 15416 8616 15444
rect 8168 15388 8616 15416
rect 8168 15376 8174 15388
rect 19334 15376 19340 15428
rect 19392 15416 19398 15428
rect 20165 15419 20223 15425
rect 20165 15416 20177 15419
rect 19392 15388 20177 15416
rect 19392 15376 19398 15388
rect 20165 15385 20177 15388
rect 20211 15385 20223 15419
rect 20165 15379 20223 15385
rect 20714 15376 20720 15428
rect 20772 15416 20778 15428
rect 21450 15416 21456 15428
rect 20772 15388 21456 15416
rect 20772 15376 20778 15388
rect 21450 15376 21456 15388
rect 21508 15416 21514 15428
rect 21560 15416 21588 15447
rect 24670 15444 24676 15456
rect 24728 15484 24734 15496
rect 24946 15484 24952 15496
rect 24728 15456 24952 15484
rect 24728 15444 24734 15456
rect 24946 15444 24952 15456
rect 25004 15444 25010 15496
rect 23566 15416 23572 15428
rect 21508 15388 21588 15416
rect 23527 15388 23572 15416
rect 21508 15376 21514 15388
rect 23566 15376 23572 15388
rect 23624 15376 23630 15428
rect 24854 15376 24860 15428
rect 24912 15416 24918 15428
rect 25317 15419 25375 15425
rect 25317 15416 25329 15419
rect 24912 15388 25329 15416
rect 24912 15376 24918 15388
rect 25317 15385 25329 15388
rect 25363 15385 25375 15419
rect 25317 15379 25375 15385
rect 8570 15348 8576 15360
rect 6472 15320 8576 15348
rect 8570 15308 8576 15320
rect 8628 15348 8634 15360
rect 8846 15348 8852 15360
rect 8628 15320 8852 15348
rect 8628 15308 8634 15320
rect 8846 15308 8852 15320
rect 8904 15308 8910 15360
rect 11882 15348 11888 15360
rect 11843 15320 11888 15348
rect 11882 15308 11888 15320
rect 11940 15308 11946 15360
rect 12158 15308 12164 15360
rect 12216 15348 12222 15360
rect 12529 15351 12587 15357
rect 12529 15348 12541 15351
rect 12216 15320 12541 15348
rect 12216 15308 12222 15320
rect 12529 15317 12541 15320
rect 12575 15348 12587 15351
rect 12618 15348 12624 15360
rect 12575 15320 12624 15348
rect 12575 15317 12587 15320
rect 12529 15311 12587 15317
rect 12618 15308 12624 15320
rect 12676 15308 12682 15360
rect 12989 15351 13047 15357
rect 12989 15317 13001 15351
rect 13035 15348 13047 15351
rect 13814 15348 13820 15360
rect 13035 15320 13820 15348
rect 13035 15317 13047 15320
rect 12989 15311 13047 15317
rect 13814 15308 13820 15320
rect 13872 15308 13878 15360
rect 14090 15308 14096 15360
rect 14148 15348 14154 15360
rect 14553 15351 14611 15357
rect 14553 15348 14565 15351
rect 14148 15320 14565 15348
rect 14148 15308 14154 15320
rect 14553 15317 14565 15320
rect 14599 15348 14611 15351
rect 14642 15348 14648 15360
rect 14599 15320 14648 15348
rect 14599 15317 14611 15320
rect 14553 15311 14611 15317
rect 14642 15308 14648 15320
rect 14700 15308 14706 15360
rect 14734 15308 14740 15360
rect 14792 15348 14798 15360
rect 15473 15351 15531 15357
rect 15473 15348 15485 15351
rect 14792 15320 15485 15348
rect 14792 15308 14798 15320
rect 15473 15317 15485 15320
rect 15519 15348 15531 15351
rect 15562 15348 15568 15360
rect 15519 15320 15568 15348
rect 15519 15317 15531 15320
rect 15473 15311 15531 15317
rect 15562 15308 15568 15320
rect 15620 15308 15626 15360
rect 18046 15348 18052 15360
rect 18007 15320 18052 15348
rect 18046 15308 18052 15320
rect 18104 15308 18110 15360
rect 19613 15351 19671 15357
rect 19613 15317 19625 15351
rect 19659 15348 19671 15351
rect 19978 15348 19984 15360
rect 19659 15320 19984 15348
rect 19659 15317 19671 15320
rect 19613 15311 19671 15317
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 20622 15308 20628 15360
rect 20680 15348 20686 15360
rect 22005 15351 22063 15357
rect 22005 15348 22017 15351
rect 20680 15320 22017 15348
rect 20680 15308 20686 15320
rect 22005 15317 22017 15320
rect 22051 15348 22063 15351
rect 22370 15348 22376 15360
rect 22051 15320 22376 15348
rect 22051 15317 22063 15320
rect 22005 15311 22063 15317
rect 22370 15308 22376 15320
rect 22428 15308 22434 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1581 15147 1639 15153
rect 1581 15113 1593 15147
rect 1627 15144 1639 15147
rect 2130 15144 2136 15156
rect 1627 15116 2136 15144
rect 1627 15113 1639 15116
rect 1581 15107 1639 15113
rect 2130 15104 2136 15116
rect 2188 15104 2194 15156
rect 2869 15147 2927 15153
rect 2869 15113 2881 15147
rect 2915 15144 2927 15147
rect 3053 15147 3111 15153
rect 3053 15144 3065 15147
rect 2915 15116 3065 15144
rect 2915 15113 2927 15116
rect 2869 15107 2927 15113
rect 3053 15113 3065 15116
rect 3099 15144 3111 15147
rect 4430 15144 4436 15156
rect 3099 15116 4436 15144
rect 3099 15113 3111 15116
rect 3053 15107 3111 15113
rect 4430 15104 4436 15116
rect 4488 15144 4494 15156
rect 4706 15144 4712 15156
rect 4488 15116 4712 15144
rect 4488 15104 4494 15116
rect 4706 15104 4712 15116
rect 4764 15104 4770 15156
rect 7650 15144 7656 15156
rect 7611 15116 7656 15144
rect 7650 15104 7656 15116
rect 7708 15104 7714 15156
rect 7834 15104 7840 15156
rect 7892 15144 7898 15156
rect 8202 15144 8208 15156
rect 7892 15116 8208 15144
rect 7892 15104 7898 15116
rect 8202 15104 8208 15116
rect 8260 15144 8266 15156
rect 9217 15147 9275 15153
rect 9217 15144 9229 15147
rect 8260 15116 9229 15144
rect 8260 15104 8266 15116
rect 9217 15113 9229 15116
rect 9263 15113 9275 15147
rect 9217 15107 9275 15113
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 13538 15144 13544 15156
rect 12492 15116 12537 15144
rect 13499 15116 13544 15144
rect 12492 15104 12498 15116
rect 13538 15104 13544 15116
rect 13596 15104 13602 15156
rect 13906 15144 13912 15156
rect 13867 15116 13912 15144
rect 13906 15104 13912 15116
rect 13964 15104 13970 15156
rect 16022 15104 16028 15156
rect 16080 15144 16086 15156
rect 16209 15147 16267 15153
rect 16209 15144 16221 15147
rect 16080 15116 16221 15144
rect 16080 15104 16086 15116
rect 16209 15113 16221 15116
rect 16255 15144 16267 15147
rect 16761 15147 16819 15153
rect 16761 15144 16773 15147
rect 16255 15116 16773 15144
rect 16255 15113 16267 15116
rect 16209 15107 16267 15113
rect 16761 15113 16773 15116
rect 16807 15113 16819 15147
rect 16761 15107 16819 15113
rect 17497 15147 17555 15153
rect 17497 15113 17509 15147
rect 17543 15144 17555 15147
rect 17862 15144 17868 15156
rect 17543 15116 17868 15144
rect 17543 15113 17555 15116
rect 17497 15107 17555 15113
rect 17862 15104 17868 15116
rect 17920 15104 17926 15156
rect 18598 15104 18604 15156
rect 18656 15144 18662 15156
rect 19061 15147 19119 15153
rect 19061 15144 19073 15147
rect 18656 15116 19073 15144
rect 18656 15104 18662 15116
rect 19061 15113 19073 15116
rect 19107 15113 19119 15147
rect 19061 15107 19119 15113
rect 21450 15104 21456 15156
rect 21508 15144 21514 15156
rect 21729 15147 21787 15153
rect 21729 15144 21741 15147
rect 21508 15116 21741 15144
rect 21508 15104 21514 15116
rect 21729 15113 21741 15116
rect 21775 15113 21787 15147
rect 21729 15107 21787 15113
rect 22189 15147 22247 15153
rect 22189 15113 22201 15147
rect 22235 15144 22247 15147
rect 22462 15144 22468 15156
rect 22235 15116 22468 15144
rect 22235 15113 22247 15116
rect 22189 15107 22247 15113
rect 22462 15104 22468 15116
rect 22520 15104 22526 15156
rect 22922 15104 22928 15156
rect 22980 15144 22986 15156
rect 23017 15147 23075 15153
rect 23017 15144 23029 15147
rect 22980 15116 23029 15144
rect 22980 15104 22986 15116
rect 23017 15113 23029 15116
rect 23063 15113 23075 15147
rect 23017 15107 23075 15113
rect 23661 15147 23719 15153
rect 23661 15113 23673 15147
rect 23707 15144 23719 15147
rect 23842 15144 23848 15156
rect 23707 15116 23848 15144
rect 23707 15113 23719 15116
rect 23661 15107 23719 15113
rect 2406 15076 2412 15088
rect 2240 15048 2412 15076
rect 1762 14968 1768 15020
rect 1820 15008 1826 15020
rect 2240 15017 2268 15048
rect 2406 15036 2412 15048
rect 2464 15036 2470 15088
rect 4525 15079 4583 15085
rect 4525 15045 4537 15079
rect 4571 15076 4583 15079
rect 5350 15076 5356 15088
rect 4571 15048 5356 15076
rect 4571 15045 4583 15048
rect 4525 15039 4583 15045
rect 5350 15036 5356 15048
rect 5408 15036 5414 15088
rect 10042 15076 10048 15088
rect 10003 15048 10048 15076
rect 10042 15036 10048 15048
rect 10100 15036 10106 15088
rect 13722 15036 13728 15088
rect 13780 15076 13786 15088
rect 14185 15079 14243 15085
rect 14185 15076 14197 15079
rect 13780 15048 14197 15076
rect 13780 15036 13786 15048
rect 14185 15045 14197 15048
rect 14231 15045 14243 15079
rect 14185 15039 14243 15045
rect 17218 15036 17224 15088
rect 17276 15076 17282 15088
rect 18049 15079 18107 15085
rect 18049 15076 18061 15079
rect 17276 15048 18061 15076
rect 17276 15036 17282 15048
rect 18049 15045 18061 15048
rect 18095 15045 18107 15079
rect 23032 15076 23060 15107
rect 23842 15104 23848 15116
rect 23900 15104 23906 15156
rect 24670 15144 24676 15156
rect 24631 15116 24676 15144
rect 24670 15104 24676 15116
rect 24728 15104 24734 15156
rect 25314 15104 25320 15156
rect 25372 15144 25378 15156
rect 25409 15147 25467 15153
rect 25409 15144 25421 15147
rect 25372 15116 25421 15144
rect 25372 15104 25378 15116
rect 25409 15113 25421 15116
rect 25455 15113 25467 15147
rect 25409 15107 25467 15113
rect 23106 15076 23112 15088
rect 23019 15048 23112 15076
rect 18049 15039 18107 15045
rect 23106 15036 23112 15048
rect 23164 15076 23170 15088
rect 25041 15079 25099 15085
rect 25041 15076 25053 15079
rect 23164 15048 23612 15076
rect 23164 15036 23170 15048
rect 2041 15011 2099 15017
rect 2041 15008 2053 15011
rect 1820 14980 2053 15008
rect 1820 14968 1826 14980
rect 2041 14977 2053 14980
rect 2087 14977 2099 15011
rect 2041 14971 2099 14977
rect 2225 15011 2283 15017
rect 2225 14977 2237 15011
rect 2271 14977 2283 15011
rect 2225 14971 2283 14977
rect 5258 14968 5264 15020
rect 5316 15008 5322 15020
rect 6549 15011 6607 15017
rect 6549 15008 6561 15011
rect 5316 14980 6561 15008
rect 5316 14968 5322 14980
rect 6549 14977 6561 14980
rect 6595 14977 6607 15011
rect 10060 15008 10088 15036
rect 11057 15011 11115 15017
rect 11057 15008 11069 15011
rect 10060 14980 11069 15008
rect 6549 14971 6607 14977
rect 11057 14977 11069 14980
rect 11103 14977 11115 15011
rect 11057 14971 11115 14977
rect 11241 15011 11299 15017
rect 11241 14977 11253 15011
rect 11287 15008 11299 15011
rect 11330 15008 11336 15020
rect 11287 14980 11336 15008
rect 11287 14977 11299 14980
rect 11241 14971 11299 14977
rect 11330 14968 11336 14980
rect 11388 14968 11394 15020
rect 13078 15008 13084 15020
rect 13039 14980 13084 15008
rect 13078 14968 13084 14980
rect 13136 14968 13142 15020
rect 18598 15008 18604 15020
rect 18559 14980 18604 15008
rect 18598 14968 18604 14980
rect 18656 14968 18662 15020
rect 19242 14968 19248 15020
rect 19300 14968 19306 15020
rect 3145 14943 3203 14949
rect 3145 14909 3157 14943
rect 3191 14909 3203 14943
rect 3145 14903 3203 14909
rect 1949 14875 2007 14881
rect 1949 14841 1961 14875
rect 1995 14872 2007 14875
rect 3160 14872 3188 14903
rect 3234 14900 3240 14952
rect 3292 14940 3298 14952
rect 3401 14943 3459 14949
rect 3401 14940 3413 14943
rect 3292 14912 3413 14940
rect 3292 14900 3298 14912
rect 3401 14909 3413 14912
rect 3447 14909 3459 14943
rect 3401 14903 3459 14909
rect 5169 14943 5227 14949
rect 5169 14909 5181 14943
rect 5215 14940 5227 14943
rect 5534 14940 5540 14952
rect 5215 14912 5540 14940
rect 5215 14909 5227 14912
rect 5169 14903 5227 14909
rect 5534 14900 5540 14912
rect 5592 14900 5598 14952
rect 5629 14943 5687 14949
rect 5629 14909 5641 14943
rect 5675 14940 5687 14943
rect 7837 14943 7895 14949
rect 5675 14912 6040 14940
rect 5675 14909 5687 14912
rect 5629 14903 5687 14909
rect 5258 14872 5264 14884
rect 1995 14844 2728 14872
rect 3160 14844 5264 14872
rect 1995 14841 2007 14844
rect 1949 14835 2007 14841
rect 2314 14764 2320 14816
rect 2372 14804 2378 14816
rect 2593 14807 2651 14813
rect 2593 14804 2605 14807
rect 2372 14776 2605 14804
rect 2372 14764 2378 14776
rect 2593 14773 2605 14776
rect 2639 14773 2651 14807
rect 2700 14804 2728 14844
rect 5258 14832 5264 14844
rect 5316 14832 5322 14884
rect 6012 14816 6040 14912
rect 7837 14909 7849 14943
rect 7883 14940 7895 14943
rect 7926 14940 7932 14952
rect 7883 14912 7932 14940
rect 7883 14909 7895 14912
rect 7837 14903 7895 14909
rect 7926 14900 7932 14912
rect 7984 14900 7990 14952
rect 8110 14949 8116 14952
rect 8104 14940 8116 14949
rect 8071 14912 8116 14940
rect 8104 14903 8116 14912
rect 8110 14900 8116 14903
rect 8168 14900 8174 14952
rect 10502 14940 10508 14952
rect 10415 14912 10508 14940
rect 10502 14900 10508 14912
rect 10560 14940 10566 14952
rect 10965 14943 11023 14949
rect 10965 14940 10977 14943
rect 10560 14912 10977 14940
rect 10560 14900 10566 14912
rect 10965 14909 10977 14912
rect 11011 14940 11023 14943
rect 11514 14940 11520 14952
rect 11011 14912 11520 14940
rect 11011 14909 11023 14912
rect 10965 14903 11023 14909
rect 11514 14900 11520 14912
rect 11572 14900 11578 14952
rect 14826 14940 14832 14952
rect 14787 14912 14832 14940
rect 14826 14900 14832 14912
rect 14884 14940 14890 14952
rect 17862 14940 17868 14952
rect 14884 14912 15332 14940
rect 17823 14912 17868 14940
rect 14884 14900 14890 14912
rect 15304 14884 15332 14912
rect 17862 14900 17868 14912
rect 17920 14900 17926 14952
rect 18414 14940 18420 14952
rect 18327 14912 18420 14940
rect 18414 14900 18420 14912
rect 18472 14940 18478 14952
rect 19260 14940 19288 14968
rect 18472 14912 19288 14940
rect 19797 14943 19855 14949
rect 18472 14900 18478 14912
rect 19797 14909 19809 14943
rect 19843 14940 19855 14943
rect 21082 14940 21088 14952
rect 19843 14912 21088 14940
rect 19843 14909 19855 14912
rect 19797 14903 19855 14909
rect 20180 14884 20208 14912
rect 21082 14900 21088 14912
rect 21140 14900 21146 14952
rect 22278 14940 22284 14952
rect 22239 14912 22284 14940
rect 22278 14900 22284 14912
rect 22336 14900 22342 14952
rect 23014 14900 23020 14952
rect 23072 14900 23078 14952
rect 23584 14940 23612 15048
rect 24136 15048 25053 15076
rect 23658 14968 23664 15020
rect 23716 15008 23722 15020
rect 24136 15017 24164 15048
rect 25041 15045 25053 15048
rect 25087 15045 25099 15079
rect 25041 15039 25099 15045
rect 24121 15011 24179 15017
rect 24121 15008 24133 15011
rect 23716 14980 24133 15008
rect 23716 14968 23722 14980
rect 24121 14977 24133 14980
rect 24167 14977 24179 15011
rect 24121 14971 24179 14977
rect 24213 15011 24271 15017
rect 24213 14977 24225 15011
rect 24259 14977 24271 15011
rect 24213 14971 24271 14977
rect 24026 14940 24032 14952
rect 23584 14912 23888 14940
rect 23987 14912 24032 14940
rect 6638 14832 6644 14884
rect 6696 14872 6702 14884
rect 6696 14844 7328 14872
rect 6696 14832 6702 14844
rect 7300 14816 7328 14844
rect 9490 14832 9496 14884
rect 9548 14872 9554 14884
rect 12434 14872 12440 14884
rect 9548 14844 12440 14872
rect 9548 14832 9554 14844
rect 12434 14832 12440 14844
rect 12492 14832 12498 14884
rect 12618 14832 12624 14884
rect 12676 14872 12682 14884
rect 12805 14875 12863 14881
rect 12805 14872 12817 14875
rect 12676 14844 12817 14872
rect 12676 14832 12682 14844
rect 12805 14841 12817 14844
rect 12851 14872 12863 14875
rect 12986 14872 12992 14884
rect 12851 14844 12992 14872
rect 12851 14841 12863 14844
rect 12805 14835 12863 14841
rect 12986 14832 12992 14844
rect 13044 14832 13050 14884
rect 15074 14875 15132 14881
rect 15074 14872 15086 14875
rect 14660 14844 15086 14872
rect 14660 14816 14688 14844
rect 15074 14841 15086 14844
rect 15120 14841 15132 14875
rect 15074 14835 15132 14841
rect 15286 14832 15292 14884
rect 15344 14872 15350 14884
rect 18506 14872 18512 14884
rect 15344 14844 17724 14872
rect 18419 14844 18512 14872
rect 15344 14832 15350 14844
rect 2869 14807 2927 14813
rect 2869 14804 2881 14807
rect 2700 14776 2881 14804
rect 2593 14767 2651 14773
rect 2869 14773 2881 14776
rect 2915 14804 2927 14807
rect 3142 14804 3148 14816
rect 2915 14776 3148 14804
rect 2915 14773 2927 14776
rect 2869 14767 2927 14773
rect 3142 14764 3148 14776
rect 3200 14764 3206 14816
rect 5166 14764 5172 14816
rect 5224 14804 5230 14816
rect 5537 14807 5595 14813
rect 5537 14804 5549 14807
rect 5224 14776 5549 14804
rect 5224 14764 5230 14776
rect 5537 14773 5549 14776
rect 5583 14773 5595 14807
rect 5810 14804 5816 14816
rect 5771 14776 5816 14804
rect 5537 14767 5595 14773
rect 5810 14764 5816 14776
rect 5868 14764 5874 14816
rect 5994 14764 6000 14816
rect 6052 14804 6058 14816
rect 6181 14807 6239 14813
rect 6181 14804 6193 14807
rect 6052 14776 6193 14804
rect 6052 14764 6058 14776
rect 6181 14773 6193 14776
rect 6227 14773 6239 14807
rect 6822 14804 6828 14816
rect 6783 14776 6828 14804
rect 6181 14767 6239 14773
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7282 14804 7288 14816
rect 7243 14776 7288 14804
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 10597 14807 10655 14813
rect 10597 14773 10609 14807
rect 10643 14804 10655 14807
rect 10686 14804 10692 14816
rect 10643 14776 10692 14804
rect 10643 14773 10655 14776
rect 10597 14767 10655 14773
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 11330 14764 11336 14816
rect 11388 14804 11394 14816
rect 11609 14807 11667 14813
rect 11609 14804 11621 14807
rect 11388 14776 11621 14804
rect 11388 14764 11394 14776
rect 11609 14773 11621 14776
rect 11655 14773 11667 14807
rect 11609 14767 11667 14773
rect 12253 14807 12311 14813
rect 12253 14773 12265 14807
rect 12299 14804 12311 14807
rect 12894 14804 12900 14816
rect 12299 14776 12900 14804
rect 12299 14773 12311 14776
rect 12253 14767 12311 14773
rect 12894 14764 12900 14776
rect 12952 14804 12958 14816
rect 13446 14804 13452 14816
rect 12952 14776 13452 14804
rect 12952 14764 12958 14776
rect 13446 14764 13452 14776
rect 13504 14764 13510 14816
rect 14642 14804 14648 14816
rect 14603 14776 14648 14804
rect 14642 14764 14648 14776
rect 14700 14764 14706 14816
rect 17696 14813 17724 14844
rect 18506 14832 18512 14844
rect 18564 14872 18570 14884
rect 19242 14872 19248 14884
rect 18564 14844 19248 14872
rect 18564 14832 18570 14844
rect 19242 14832 19248 14844
rect 19300 14832 19306 14884
rect 20042 14875 20100 14881
rect 20042 14872 20054 14875
rect 19628 14844 20054 14872
rect 17681 14807 17739 14813
rect 17681 14773 17693 14807
rect 17727 14804 17739 14807
rect 18046 14804 18052 14816
rect 17727 14776 18052 14804
rect 17727 14773 17739 14776
rect 17681 14767 17739 14773
rect 18046 14764 18052 14776
rect 18104 14764 18110 14816
rect 19518 14764 19524 14816
rect 19576 14804 19582 14816
rect 19628 14813 19656 14844
rect 20042 14841 20054 14844
rect 20088 14841 20100 14875
rect 20042 14835 20100 14841
rect 20162 14832 20168 14884
rect 20220 14832 20226 14884
rect 23032 14872 23060 14900
rect 22480 14844 23060 14872
rect 23477 14875 23535 14881
rect 19613 14807 19671 14813
rect 19613 14804 19625 14807
rect 19576 14776 19625 14804
rect 19576 14764 19582 14776
rect 19613 14773 19625 14776
rect 19659 14773 19671 14807
rect 21174 14804 21180 14816
rect 21087 14776 21180 14804
rect 19613 14767 19671 14773
rect 21174 14764 21180 14776
rect 21232 14804 21238 14816
rect 21450 14804 21456 14816
rect 21232 14776 21456 14804
rect 21232 14764 21238 14776
rect 21450 14764 21456 14776
rect 21508 14764 21514 14816
rect 22480 14813 22508 14844
rect 23477 14841 23489 14875
rect 23523 14872 23535 14875
rect 23750 14872 23756 14884
rect 23523 14844 23756 14872
rect 23523 14841 23535 14844
rect 23477 14835 23535 14841
rect 23750 14832 23756 14844
rect 23808 14832 23814 14884
rect 23860 14872 23888 14912
rect 24026 14900 24032 14912
rect 24084 14900 24090 14952
rect 24228 14940 24256 14971
rect 25222 14940 25228 14952
rect 24136 14912 24256 14940
rect 25183 14912 25228 14940
rect 24136 14872 24164 14912
rect 25222 14900 25228 14912
rect 25280 14940 25286 14952
rect 25777 14943 25835 14949
rect 25777 14940 25789 14943
rect 25280 14912 25789 14940
rect 25280 14900 25286 14912
rect 25777 14909 25789 14912
rect 25823 14909 25835 14943
rect 25777 14903 25835 14909
rect 23860 14844 24164 14872
rect 22465 14807 22523 14813
rect 22465 14773 22477 14807
rect 22511 14773 22523 14807
rect 22465 14767 22523 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 2774 14560 2780 14612
rect 2832 14600 2838 14612
rect 2869 14603 2927 14609
rect 2869 14600 2881 14603
rect 2832 14572 2881 14600
rect 2832 14560 2838 14572
rect 2869 14569 2881 14572
rect 2915 14600 2927 14603
rect 3234 14600 3240 14612
rect 2915 14572 3240 14600
rect 2915 14569 2927 14572
rect 2869 14563 2927 14569
rect 3234 14560 3240 14572
rect 3292 14560 3298 14612
rect 4522 14600 4528 14612
rect 4483 14572 4528 14600
rect 4522 14560 4528 14572
rect 4580 14560 4586 14612
rect 5169 14603 5227 14609
rect 5169 14569 5181 14603
rect 5215 14600 5227 14603
rect 5442 14600 5448 14612
rect 5215 14572 5448 14600
rect 5215 14569 5227 14572
rect 5169 14563 5227 14569
rect 5442 14560 5448 14572
rect 5500 14560 5506 14612
rect 7653 14603 7711 14609
rect 7653 14569 7665 14603
rect 7699 14600 7711 14603
rect 7926 14600 7932 14612
rect 7699 14572 7932 14600
rect 7699 14569 7711 14572
rect 7653 14563 7711 14569
rect 7926 14560 7932 14572
rect 7984 14560 7990 14612
rect 8110 14560 8116 14612
rect 8168 14600 8174 14612
rect 8665 14603 8723 14609
rect 8665 14600 8677 14603
rect 8168 14572 8677 14600
rect 8168 14560 8174 14572
rect 8665 14569 8677 14572
rect 8711 14569 8723 14603
rect 9398 14600 9404 14612
rect 9359 14572 9404 14600
rect 8665 14563 8723 14569
rect 9398 14560 9404 14572
rect 9456 14560 9462 14612
rect 10778 14560 10784 14612
rect 10836 14600 10842 14612
rect 11057 14603 11115 14609
rect 11057 14600 11069 14603
rect 10836 14572 11069 14600
rect 10836 14560 10842 14572
rect 11057 14569 11069 14572
rect 11103 14569 11115 14603
rect 11057 14563 11115 14569
rect 12161 14603 12219 14609
rect 12161 14569 12173 14603
rect 12207 14600 12219 14603
rect 12526 14600 12532 14612
rect 12207 14572 12532 14600
rect 12207 14569 12219 14572
rect 12161 14563 12219 14569
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 15749 14603 15807 14609
rect 15749 14569 15761 14603
rect 15795 14600 15807 14603
rect 16482 14600 16488 14612
rect 15795 14572 16488 14600
rect 15795 14569 15807 14572
rect 15749 14563 15807 14569
rect 16482 14560 16488 14572
rect 16540 14560 16546 14612
rect 16761 14603 16819 14609
rect 16761 14569 16773 14603
rect 16807 14600 16819 14603
rect 16850 14600 16856 14612
rect 16807 14572 16856 14600
rect 16807 14569 16819 14572
rect 16761 14563 16819 14569
rect 16850 14560 16856 14572
rect 16908 14560 16914 14612
rect 17862 14560 17868 14612
rect 17920 14600 17926 14612
rect 20070 14600 20076 14612
rect 17920 14572 20076 14600
rect 17920 14560 17926 14572
rect 20070 14560 20076 14572
rect 20128 14600 20134 14612
rect 20257 14603 20315 14609
rect 20257 14600 20269 14603
rect 20128 14572 20269 14600
rect 20128 14560 20134 14572
rect 20257 14569 20269 14572
rect 20303 14569 20315 14603
rect 20898 14600 20904 14612
rect 20859 14572 20904 14600
rect 20257 14563 20315 14569
rect 20898 14560 20904 14572
rect 20956 14560 20962 14612
rect 21082 14560 21088 14612
rect 21140 14600 21146 14612
rect 21913 14603 21971 14609
rect 21913 14600 21925 14603
rect 21140 14572 21925 14600
rect 21140 14560 21146 14572
rect 21913 14569 21925 14572
rect 21959 14569 21971 14603
rect 22278 14600 22284 14612
rect 22239 14572 22284 14600
rect 21913 14563 21971 14569
rect 22278 14560 22284 14572
rect 22336 14560 22342 14612
rect 22465 14603 22523 14609
rect 22465 14569 22477 14603
rect 22511 14600 22523 14603
rect 22830 14600 22836 14612
rect 22511 14572 22836 14600
rect 22511 14569 22523 14572
rect 22465 14563 22523 14569
rect 22830 14560 22836 14572
rect 22888 14560 22894 14612
rect 23753 14603 23811 14609
rect 23753 14569 23765 14603
rect 23799 14600 23811 14603
rect 24026 14600 24032 14612
rect 23799 14572 24032 14600
rect 23799 14569 23811 14572
rect 23753 14563 23811 14569
rect 24026 14560 24032 14572
rect 24084 14560 24090 14612
rect 24118 14560 24124 14612
rect 24176 14600 24182 14612
rect 25501 14603 25559 14609
rect 25501 14600 25513 14603
rect 24176 14572 25513 14600
rect 24176 14560 24182 14572
rect 25501 14569 25513 14572
rect 25547 14569 25559 14603
rect 25501 14563 25559 14569
rect 1756 14535 1814 14541
rect 1756 14501 1768 14535
rect 1802 14532 1814 14535
rect 1946 14532 1952 14544
rect 1802 14504 1952 14532
rect 1802 14501 1814 14504
rect 1756 14495 1814 14501
rect 1946 14492 1952 14504
rect 2004 14492 2010 14544
rect 8021 14535 8079 14541
rect 8021 14501 8033 14535
rect 8067 14532 8079 14535
rect 8294 14532 8300 14544
rect 8067 14504 8300 14532
rect 8067 14501 8079 14504
rect 8021 14495 8079 14501
rect 8294 14492 8300 14504
rect 8352 14492 8358 14544
rect 8570 14492 8576 14544
rect 8628 14532 8634 14544
rect 9033 14535 9091 14541
rect 9033 14532 9045 14535
rect 8628 14504 9045 14532
rect 8628 14492 8634 14504
rect 9033 14501 9045 14504
rect 9079 14501 9091 14535
rect 9033 14495 9091 14501
rect 9674 14492 9680 14544
rect 9732 14532 9738 14544
rect 9922 14535 9980 14541
rect 9922 14532 9934 14535
rect 9732 14504 9934 14532
rect 9732 14492 9738 14504
rect 9922 14501 9934 14504
rect 9968 14501 9980 14535
rect 12618 14532 12624 14544
rect 12531 14504 12624 14532
rect 9922 14495 9980 14501
rect 12618 14492 12624 14504
rect 12676 14532 12682 14544
rect 13998 14532 14004 14544
rect 12676 14504 14004 14532
rect 12676 14492 12682 14504
rect 13998 14492 14004 14504
rect 14056 14492 14062 14544
rect 20717 14535 20775 14541
rect 20717 14501 20729 14535
rect 20763 14532 20775 14535
rect 20990 14532 20996 14544
rect 20763 14504 20996 14532
rect 20763 14501 20775 14504
rect 20717 14495 20775 14501
rect 20990 14492 20996 14504
rect 21048 14532 21054 14544
rect 21358 14532 21364 14544
rect 21048 14504 21364 14532
rect 21048 14492 21054 14504
rect 21358 14492 21364 14504
rect 21416 14492 21422 14544
rect 22738 14492 22744 14544
rect 22796 14532 22802 14544
rect 22925 14535 22983 14541
rect 22925 14532 22937 14535
rect 22796 14504 22937 14532
rect 22796 14492 22802 14504
rect 22925 14501 22937 14504
rect 22971 14501 22983 14535
rect 22925 14495 22983 14501
rect 23658 14492 23664 14544
rect 23716 14532 23722 14544
rect 24210 14532 24216 14544
rect 23716 14504 24216 14532
rect 23716 14492 23722 14504
rect 24210 14492 24216 14504
rect 24268 14492 24274 14544
rect 25130 14532 25136 14544
rect 25091 14504 25136 14532
rect 25130 14492 25136 14504
rect 25188 14492 25194 14544
rect 4430 14464 4436 14476
rect 4391 14436 4436 14464
rect 4430 14424 4436 14436
rect 4488 14424 4494 14476
rect 5445 14467 5503 14473
rect 5445 14433 5457 14467
rect 5491 14464 5503 14467
rect 5896 14467 5954 14473
rect 5896 14464 5908 14467
rect 5491 14436 5908 14464
rect 5491 14433 5503 14436
rect 5445 14427 5503 14433
rect 5896 14433 5908 14436
rect 5942 14464 5954 14467
rect 6270 14464 6276 14476
rect 5942 14436 6276 14464
rect 5942 14433 5954 14436
rect 5896 14427 5954 14433
rect 6270 14424 6276 14436
rect 6328 14464 6334 14476
rect 7834 14464 7840 14476
rect 6328 14436 7840 14464
rect 6328 14424 6334 14436
rect 7834 14424 7840 14436
rect 7892 14424 7898 14476
rect 8113 14467 8171 14473
rect 8113 14433 8125 14467
rect 8159 14464 8171 14467
rect 8202 14464 8208 14476
rect 8159 14436 8208 14464
rect 8159 14433 8171 14436
rect 8113 14427 8171 14433
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 12434 14424 12440 14476
rect 12492 14464 12498 14476
rect 12529 14467 12587 14473
rect 12529 14464 12541 14467
rect 12492 14436 12541 14464
rect 12492 14424 12498 14436
rect 12529 14433 12541 14436
rect 12575 14464 12587 14467
rect 13541 14467 13599 14473
rect 13541 14464 13553 14467
rect 12575 14436 13553 14464
rect 12575 14433 12587 14436
rect 12529 14427 12587 14433
rect 13541 14433 13553 14436
rect 13587 14433 13599 14467
rect 13541 14427 13599 14433
rect 13814 14424 13820 14476
rect 13872 14464 13878 14476
rect 13909 14467 13967 14473
rect 13909 14464 13921 14467
rect 13872 14436 13921 14464
rect 13872 14424 13878 14436
rect 13909 14433 13921 14436
rect 13955 14464 13967 14467
rect 14645 14467 14703 14473
rect 14645 14464 14657 14467
rect 13955 14436 14657 14464
rect 13955 14433 13967 14436
rect 13909 14427 13967 14433
rect 14645 14433 14657 14436
rect 14691 14433 14703 14467
rect 14645 14427 14703 14433
rect 15657 14467 15715 14473
rect 15657 14433 15669 14467
rect 15703 14464 15715 14467
rect 17129 14467 17187 14473
rect 17129 14464 17141 14467
rect 15703 14436 17141 14464
rect 15703 14433 15715 14436
rect 15657 14427 15715 14433
rect 17129 14433 17141 14436
rect 17175 14464 17187 14467
rect 17954 14464 17960 14476
rect 17175 14436 17960 14464
rect 17175 14433 17187 14436
rect 17129 14427 17187 14433
rect 17954 14424 17960 14436
rect 18012 14424 18018 14476
rect 18598 14473 18604 14476
rect 18141 14467 18199 14473
rect 18141 14433 18153 14467
rect 18187 14464 18199 14467
rect 18592 14464 18604 14473
rect 18187 14436 18604 14464
rect 18187 14433 18199 14436
rect 18141 14427 18199 14433
rect 18592 14427 18604 14436
rect 18656 14464 18662 14476
rect 19058 14464 19064 14476
rect 18656 14436 19064 14464
rect 18598 14424 18604 14427
rect 18656 14424 18662 14436
rect 19058 14424 19064 14436
rect 19116 14424 19122 14476
rect 21269 14467 21327 14473
rect 21269 14433 21281 14467
rect 21315 14464 21327 14467
rect 22002 14464 22008 14476
rect 21315 14436 22008 14464
rect 21315 14433 21327 14436
rect 21269 14427 21327 14433
rect 22002 14424 22008 14436
rect 22060 14424 22066 14476
rect 22370 14424 22376 14476
rect 22428 14464 22434 14476
rect 22833 14467 22891 14473
rect 22833 14464 22845 14467
rect 22428 14436 22845 14464
rect 22428 14424 22434 14436
rect 22833 14433 22845 14436
rect 22879 14433 22891 14467
rect 24026 14464 24032 14476
rect 23987 14436 24032 14464
rect 22833 14427 22891 14433
rect 24026 14424 24032 14436
rect 24084 14464 24090 14476
rect 24765 14467 24823 14473
rect 24765 14464 24777 14467
rect 24084 14436 24777 14464
rect 24084 14424 24090 14436
rect 24765 14433 24777 14436
rect 24811 14433 24823 14467
rect 24765 14427 24823 14433
rect 25317 14467 25375 14473
rect 25317 14433 25329 14467
rect 25363 14464 25375 14467
rect 25498 14464 25504 14476
rect 25363 14436 25504 14464
rect 25363 14433 25375 14436
rect 25317 14427 25375 14433
rect 25498 14424 25504 14436
rect 25556 14424 25562 14476
rect 1394 14356 1400 14408
rect 1452 14396 1458 14408
rect 1489 14399 1547 14405
rect 1489 14396 1501 14399
rect 1452 14368 1501 14396
rect 1452 14356 1458 14368
rect 1489 14365 1501 14368
rect 1535 14365 1547 14399
rect 1489 14359 1547 14365
rect 4614 14356 4620 14408
rect 4672 14396 4678 14408
rect 4709 14399 4767 14405
rect 4709 14396 4721 14399
rect 4672 14368 4721 14396
rect 4672 14356 4678 14368
rect 4709 14365 4721 14368
rect 4755 14396 4767 14399
rect 5534 14396 5540 14408
rect 4755 14368 5540 14396
rect 4755 14365 4767 14368
rect 4709 14359 4767 14365
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 5629 14399 5687 14405
rect 5629 14365 5641 14399
rect 5675 14365 5687 14399
rect 5629 14359 5687 14365
rect 5258 14288 5264 14340
rect 5316 14328 5322 14340
rect 5644 14328 5672 14359
rect 6730 14356 6736 14408
rect 6788 14396 6794 14408
rect 6788 14368 8340 14396
rect 6788 14356 6794 14368
rect 8312 14337 8340 14368
rect 9398 14356 9404 14408
rect 9456 14396 9462 14408
rect 9677 14399 9735 14405
rect 9677 14396 9689 14399
rect 9456 14368 9689 14396
rect 9456 14356 9462 14368
rect 9677 14365 9689 14368
rect 9723 14365 9735 14399
rect 9677 14359 9735 14365
rect 11701 14399 11759 14405
rect 11701 14365 11713 14399
rect 11747 14396 11759 14399
rect 12618 14396 12624 14408
rect 11747 14368 12624 14396
rect 11747 14365 11759 14368
rect 11701 14359 11759 14365
rect 12618 14356 12624 14368
rect 12676 14356 12682 14408
rect 12713 14399 12771 14405
rect 12713 14365 12725 14399
rect 12759 14365 12771 14399
rect 14182 14396 14188 14408
rect 14143 14368 14188 14396
rect 12713 14359 12771 14365
rect 5316 14300 5672 14328
rect 8297 14331 8355 14337
rect 5316 14288 5322 14300
rect 8297 14297 8309 14331
rect 8343 14297 8355 14331
rect 8297 14291 8355 14297
rect 11882 14288 11888 14340
rect 11940 14328 11946 14340
rect 12069 14331 12127 14337
rect 12069 14328 12081 14331
rect 11940 14300 12081 14328
rect 11940 14288 11946 14300
rect 12069 14297 12081 14300
rect 12115 14328 12127 14331
rect 12728 14328 12756 14359
rect 14182 14356 14188 14368
rect 14240 14356 14246 14408
rect 16482 14396 16488 14408
rect 16443 14368 16488 14396
rect 16482 14356 16488 14368
rect 16540 14356 16546 14408
rect 17218 14396 17224 14408
rect 17179 14368 17224 14396
rect 17218 14356 17224 14368
rect 17276 14356 17282 14408
rect 17402 14396 17408 14408
rect 17363 14368 17408 14396
rect 17402 14356 17408 14368
rect 17460 14356 17466 14408
rect 18046 14356 18052 14408
rect 18104 14396 18110 14408
rect 18325 14399 18383 14405
rect 18325 14396 18337 14399
rect 18104 14368 18337 14396
rect 18104 14356 18110 14368
rect 18325 14365 18337 14368
rect 18371 14365 18383 14399
rect 18325 14359 18383 14365
rect 20806 14356 20812 14408
rect 20864 14396 20870 14408
rect 21361 14399 21419 14405
rect 21361 14396 21373 14399
rect 20864 14368 21373 14396
rect 20864 14356 20870 14368
rect 21361 14365 21373 14368
rect 21407 14365 21419 14399
rect 21361 14359 21419 14365
rect 21450 14356 21456 14408
rect 21508 14396 21514 14408
rect 21508 14368 21553 14396
rect 21508 14356 21514 14368
rect 21818 14356 21824 14408
rect 21876 14396 21882 14408
rect 22278 14396 22284 14408
rect 21876 14368 22284 14396
rect 21876 14356 21882 14368
rect 22278 14356 22284 14368
rect 22336 14356 22342 14408
rect 23106 14396 23112 14408
rect 23067 14368 23112 14396
rect 23106 14356 23112 14368
rect 23164 14356 23170 14408
rect 24210 14396 24216 14408
rect 24171 14368 24216 14396
rect 24210 14356 24216 14368
rect 24268 14356 24274 14408
rect 19702 14328 19708 14340
rect 12115 14300 12756 14328
rect 19663 14300 19708 14328
rect 12115 14297 12127 14300
rect 12069 14291 12127 14297
rect 19702 14288 19708 14300
rect 19760 14288 19766 14340
rect 3510 14260 3516 14272
rect 3471 14232 3516 14260
rect 3510 14220 3516 14232
rect 3568 14220 3574 14272
rect 3881 14263 3939 14269
rect 3881 14229 3893 14263
rect 3927 14260 3939 14263
rect 4065 14263 4123 14269
rect 4065 14260 4077 14263
rect 3927 14232 4077 14260
rect 3927 14229 3939 14232
rect 3881 14223 3939 14229
rect 4065 14229 4077 14232
rect 4111 14260 4123 14263
rect 6362 14260 6368 14272
rect 4111 14232 6368 14260
rect 4111 14229 4123 14232
rect 4065 14223 4123 14229
rect 6362 14220 6368 14232
rect 6420 14220 6426 14272
rect 6730 14220 6736 14272
rect 6788 14260 6794 14272
rect 7009 14263 7067 14269
rect 7009 14260 7021 14263
rect 6788 14232 7021 14260
rect 6788 14220 6794 14232
rect 7009 14229 7021 14232
rect 7055 14229 7067 14263
rect 7009 14223 7067 14229
rect 12158 14220 12164 14272
rect 12216 14260 12222 14272
rect 12526 14260 12532 14272
rect 12216 14232 12532 14260
rect 12216 14220 12222 14232
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 12894 14220 12900 14272
rect 12952 14260 12958 14272
rect 13173 14263 13231 14269
rect 13173 14260 13185 14263
rect 12952 14232 13185 14260
rect 12952 14220 12958 14232
rect 13173 14229 13185 14232
rect 13219 14229 13231 14263
rect 13173 14223 13231 14229
rect 14826 14220 14832 14272
rect 14884 14260 14890 14272
rect 15013 14263 15071 14269
rect 15013 14260 15025 14263
rect 14884 14232 15025 14260
rect 14884 14220 14890 14232
rect 15013 14229 15025 14232
rect 15059 14229 15071 14263
rect 15013 14223 15071 14229
rect 22002 14220 22008 14272
rect 22060 14260 22066 14272
rect 22554 14260 22560 14272
rect 22060 14232 22560 14260
rect 22060 14220 22066 14232
rect 22554 14220 22560 14232
rect 22612 14220 22618 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1854 14056 1860 14068
rect 1815 14028 1860 14056
rect 1854 14016 1860 14028
rect 1912 14016 1918 14068
rect 3970 14016 3976 14068
rect 4028 14056 4034 14068
rect 4430 14056 4436 14068
rect 4028 14028 4436 14056
rect 4028 14016 4034 14028
rect 4430 14016 4436 14028
rect 4488 14056 4494 14068
rect 6825 14059 6883 14065
rect 6825 14056 6837 14059
rect 4488 14028 6837 14056
rect 4488 14016 4494 14028
rect 6825 14025 6837 14028
rect 6871 14025 6883 14059
rect 7834 14056 7840 14068
rect 6825 14019 6883 14025
rect 7484 14028 7840 14056
rect 4341 13991 4399 13997
rect 4341 13957 4353 13991
rect 4387 13988 4399 13991
rect 4614 13988 4620 14000
rect 4387 13960 4620 13988
rect 4387 13957 4399 13960
rect 4341 13951 4399 13957
rect 4614 13948 4620 13960
rect 4672 13948 4678 14000
rect 6457 13991 6515 13997
rect 6457 13988 6469 13991
rect 4724 13960 6469 13988
rect 2240 13892 2544 13920
rect 1854 13812 1860 13864
rect 1912 13852 1918 13864
rect 2240 13861 2268 13892
rect 2225 13855 2283 13861
rect 2225 13852 2237 13855
rect 1912 13824 2237 13852
rect 1912 13812 1918 13824
rect 2225 13821 2237 13824
rect 2271 13821 2283 13855
rect 2225 13815 2283 13821
rect 2409 13855 2467 13861
rect 2409 13821 2421 13855
rect 2455 13821 2467 13855
rect 2516 13852 2544 13892
rect 3418 13880 3424 13932
rect 3476 13920 3482 13932
rect 4724 13920 4752 13960
rect 6457 13957 6469 13960
rect 6503 13988 6515 13991
rect 6549 13991 6607 13997
rect 6549 13988 6561 13991
rect 6503 13960 6561 13988
rect 6503 13957 6515 13960
rect 6457 13951 6515 13957
rect 6549 13957 6561 13960
rect 6595 13957 6607 13991
rect 6549 13951 6607 13957
rect 3476 13892 4752 13920
rect 4801 13923 4859 13929
rect 3476 13880 3482 13892
rect 4801 13889 4813 13923
rect 4847 13920 4859 13923
rect 5718 13920 5724 13932
rect 4847 13892 5724 13920
rect 4847 13889 4859 13892
rect 4801 13883 4859 13889
rect 5718 13880 5724 13892
rect 5776 13880 5782 13932
rect 6273 13923 6331 13929
rect 6273 13889 6285 13923
rect 6319 13920 6331 13923
rect 7282 13920 7288 13932
rect 6319 13892 7288 13920
rect 6319 13889 6331 13892
rect 6273 13883 6331 13889
rect 7282 13880 7288 13892
rect 7340 13880 7346 13932
rect 7484 13929 7512 14028
rect 7834 14016 7840 14028
rect 7892 14016 7898 14068
rect 9490 14056 9496 14068
rect 8036 14028 9496 14056
rect 7469 13923 7527 13929
rect 7469 13889 7481 13923
rect 7515 13889 7527 13923
rect 7469 13883 7527 13889
rect 2665 13855 2723 13861
rect 2665 13852 2677 13855
rect 2516 13824 2677 13852
rect 2409 13815 2467 13821
rect 2665 13821 2677 13824
rect 2711 13821 2723 13855
rect 2665 13815 2723 13821
rect 1394 13744 1400 13796
rect 1452 13784 1458 13796
rect 2424 13784 2452 13815
rect 3786 13812 3792 13864
rect 3844 13852 3850 13864
rect 5077 13855 5135 13861
rect 3844 13824 5019 13852
rect 3844 13812 3850 13824
rect 1452 13756 4476 13784
rect 1452 13744 1458 13756
rect 4448 13728 4476 13756
rect 1946 13676 1952 13728
rect 2004 13716 2010 13728
rect 2590 13716 2596 13728
rect 2004 13688 2596 13716
rect 2004 13676 2010 13688
rect 2590 13676 2596 13688
rect 2648 13716 2654 13728
rect 3789 13719 3847 13725
rect 3789 13716 3801 13719
rect 2648 13688 3801 13716
rect 2648 13676 2654 13688
rect 3789 13685 3801 13688
rect 3835 13685 3847 13719
rect 3789 13679 3847 13685
rect 4430 13676 4436 13728
rect 4488 13716 4494 13728
rect 4893 13719 4951 13725
rect 4893 13716 4905 13719
rect 4488 13688 4905 13716
rect 4488 13676 4494 13688
rect 4893 13685 4905 13688
rect 4939 13685 4951 13719
rect 4991 13716 5019 13824
rect 5077 13821 5089 13855
rect 5123 13852 5135 13855
rect 5810 13852 5816 13864
rect 5123 13824 5816 13852
rect 5123 13821 5135 13824
rect 5077 13815 5135 13821
rect 5810 13812 5816 13824
rect 5868 13852 5874 13864
rect 6086 13852 6092 13864
rect 5868 13824 6092 13852
rect 5868 13812 5874 13824
rect 6086 13812 6092 13824
rect 6144 13812 6150 13864
rect 6457 13855 6515 13861
rect 6457 13821 6469 13855
rect 6503 13852 6515 13855
rect 7193 13855 7251 13861
rect 7193 13852 7205 13855
rect 6503 13824 7205 13852
rect 6503 13821 6515 13824
rect 6457 13815 6515 13821
rect 7193 13821 7205 13824
rect 7239 13852 7251 13855
rect 8036 13852 8064 14028
rect 9490 14016 9496 14028
rect 9548 14016 9554 14068
rect 9674 14016 9680 14068
rect 9732 14056 9738 14068
rect 10137 14059 10195 14065
rect 10137 14056 10149 14059
rect 9732 14028 10149 14056
rect 9732 14016 9738 14028
rect 10137 14025 10149 14028
rect 10183 14056 10195 14059
rect 10689 14059 10747 14065
rect 10689 14056 10701 14059
rect 10183 14028 10701 14056
rect 10183 14025 10195 14028
rect 10137 14019 10195 14025
rect 10689 14025 10701 14028
rect 10735 14025 10747 14059
rect 10689 14019 10747 14025
rect 10778 14016 10784 14068
rect 10836 14056 10842 14068
rect 11793 14059 11851 14065
rect 11793 14056 11805 14059
rect 10836 14028 11805 14056
rect 10836 14016 10842 14028
rect 11793 14025 11805 14028
rect 11839 14025 11851 14059
rect 11793 14019 11851 14025
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 13998 14056 14004 14068
rect 12492 14028 12537 14056
rect 13959 14028 14004 14056
rect 12492 14016 12498 14028
rect 13998 14016 14004 14028
rect 14056 14016 14062 14068
rect 15565 14059 15623 14065
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 17218 14056 17224 14068
rect 15611 14028 17224 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 17218 14016 17224 14028
rect 17276 14016 17282 14068
rect 17402 14056 17408 14068
rect 17363 14028 17408 14056
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 20070 14056 20076 14068
rect 20031 14028 20076 14056
rect 20070 14016 20076 14028
rect 20128 14016 20134 14068
rect 20990 14056 20996 14068
rect 20951 14028 20996 14056
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 22738 14016 22744 14068
rect 22796 14056 22802 14068
rect 23017 14059 23075 14065
rect 23017 14056 23029 14059
rect 22796 14028 23029 14056
rect 22796 14016 22802 14028
rect 23017 14025 23029 14028
rect 23063 14025 23075 14059
rect 23017 14019 23075 14025
rect 23290 14016 23296 14068
rect 23348 14056 23354 14068
rect 23477 14059 23535 14065
rect 23477 14056 23489 14059
rect 23348 14028 23489 14056
rect 23348 14016 23354 14028
rect 23477 14025 23489 14028
rect 23523 14025 23535 14059
rect 23477 14019 23535 14025
rect 13541 13991 13599 13997
rect 13541 13957 13553 13991
rect 13587 13988 13599 13991
rect 13906 13988 13912 14000
rect 13587 13960 13912 13988
rect 13587 13957 13599 13960
rect 13541 13951 13599 13957
rect 13906 13948 13912 13960
rect 13964 13948 13970 14000
rect 16390 13988 16396 14000
rect 16351 13960 16396 13988
rect 16390 13948 16396 13960
rect 16448 13948 16454 14000
rect 19058 13948 19064 14000
rect 19116 13988 19122 14000
rect 19429 13991 19487 13997
rect 19429 13988 19441 13991
rect 19116 13960 19441 13988
rect 19116 13948 19122 13960
rect 19429 13957 19441 13960
rect 19475 13957 19487 13991
rect 19429 13951 19487 13957
rect 8665 13923 8723 13929
rect 8665 13889 8677 13923
rect 8711 13920 8723 13923
rect 13078 13920 13084 13932
rect 8711 13892 8892 13920
rect 13039 13892 13084 13920
rect 8711 13889 8723 13892
rect 8665 13883 8723 13889
rect 8202 13852 8208 13864
rect 7239 13824 8064 13852
rect 8163 13824 8208 13852
rect 7239 13821 7251 13824
rect 7193 13815 7251 13821
rect 8202 13812 8208 13824
rect 8260 13812 8266 13864
rect 8757 13855 8815 13861
rect 8757 13821 8769 13855
rect 8803 13821 8815 13855
rect 8864 13852 8892 13892
rect 13078 13880 13084 13892
rect 13136 13920 13142 13932
rect 14553 13923 14611 13929
rect 14553 13920 14565 13923
rect 13136 13892 14565 13920
rect 13136 13880 13142 13892
rect 14553 13889 14565 13892
rect 14599 13920 14611 13923
rect 15013 13923 15071 13929
rect 15013 13920 15025 13923
rect 14599 13892 15025 13920
rect 14599 13889 14611 13892
rect 14553 13883 14611 13889
rect 15013 13889 15025 13892
rect 15059 13889 15071 13923
rect 15013 13883 15071 13889
rect 15933 13923 15991 13929
rect 15933 13889 15945 13923
rect 15979 13920 15991 13923
rect 17037 13923 17095 13929
rect 17037 13920 17049 13923
rect 15979 13892 17049 13920
rect 15979 13889 15991 13892
rect 15933 13883 15991 13889
rect 17037 13889 17049 13892
rect 17083 13920 17095 13923
rect 18046 13920 18052 13932
rect 17083 13892 17908 13920
rect 18007 13892 18052 13920
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 9013 13855 9071 13861
rect 9013 13852 9025 13855
rect 8864 13824 9025 13852
rect 8757 13815 8815 13821
rect 9013 13821 9025 13824
rect 9059 13852 9071 13855
rect 9059 13824 9628 13852
rect 9059 13821 9071 13824
rect 9013 13815 9071 13821
rect 5629 13787 5687 13793
rect 5629 13753 5641 13787
rect 5675 13784 5687 13787
rect 6362 13784 6368 13796
rect 5675 13756 6368 13784
rect 5675 13753 5687 13756
rect 5629 13747 5687 13753
rect 6362 13744 6368 13756
rect 6420 13744 6426 13796
rect 8772 13784 8800 13815
rect 9398 13784 9404 13796
rect 8772 13756 9404 13784
rect 9398 13744 9404 13756
rect 9456 13744 9462 13796
rect 9600 13784 9628 13824
rect 12066 13812 12072 13864
rect 12124 13852 12130 13864
rect 12161 13855 12219 13861
rect 12161 13852 12173 13855
rect 12124 13824 12173 13852
rect 12124 13812 12130 13824
rect 12161 13821 12173 13824
rect 12207 13852 12219 13855
rect 12802 13852 12808 13864
rect 12207 13824 12808 13852
rect 12207 13821 12219 13824
rect 12161 13815 12219 13821
rect 12802 13812 12808 13824
rect 12860 13852 12866 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12860 13824 12909 13852
rect 12860 13812 12866 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 13906 13812 13912 13864
rect 13964 13852 13970 13864
rect 14458 13852 14464 13864
rect 13964 13824 14464 13852
rect 13964 13812 13970 13824
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 16853 13855 16911 13861
rect 16853 13852 16865 13855
rect 16224 13824 16865 13852
rect 10042 13784 10048 13796
rect 9600 13756 10048 13784
rect 10042 13744 10048 13756
rect 10100 13744 10106 13796
rect 11238 13744 11244 13796
rect 11296 13784 11302 13796
rect 11333 13787 11391 13793
rect 11333 13784 11345 13787
rect 11296 13756 11345 13784
rect 11296 13744 11302 13756
rect 11333 13753 11345 13756
rect 11379 13753 11391 13787
rect 11333 13747 11391 13753
rect 14918 13744 14924 13796
rect 14976 13784 14982 13796
rect 15930 13784 15936 13796
rect 14976 13756 15936 13784
rect 14976 13744 14982 13756
rect 15930 13744 15936 13756
rect 15988 13784 15994 13796
rect 16224 13793 16252 13824
rect 16853 13821 16865 13824
rect 16899 13821 16911 13855
rect 16853 13815 16911 13821
rect 16209 13787 16267 13793
rect 16209 13784 16221 13787
rect 15988 13756 16221 13784
rect 15988 13744 15994 13756
rect 16209 13753 16221 13756
rect 16255 13753 16267 13787
rect 16758 13784 16764 13796
rect 16719 13756 16764 13784
rect 16209 13747 16267 13753
rect 16758 13744 16764 13756
rect 16816 13744 16822 13796
rect 17880 13793 17908 13892
rect 18046 13880 18052 13892
rect 18104 13880 18110 13932
rect 20088 13920 20116 14016
rect 22002 13988 22008 14000
rect 21963 13960 22008 13988
rect 22002 13948 22008 13960
rect 22060 13948 22066 14000
rect 20088 13892 20760 13920
rect 20533 13855 20591 13861
rect 20533 13821 20545 13855
rect 20579 13852 20591 13855
rect 20732 13852 20760 13892
rect 21450 13880 21456 13932
rect 21508 13920 21514 13932
rect 21545 13923 21603 13929
rect 21545 13920 21557 13923
rect 21508 13892 21557 13920
rect 21508 13880 21514 13892
rect 21545 13889 21557 13892
rect 21591 13889 21603 13923
rect 23492 13920 23520 14019
rect 25498 14016 25504 14068
rect 25556 14056 25562 14068
rect 25593 14059 25651 14065
rect 25593 14056 25605 14059
rect 25556 14028 25605 14056
rect 25556 14016 25562 14028
rect 25593 14025 25605 14028
rect 25639 14025 25651 14059
rect 25593 14019 25651 14025
rect 24946 13948 24952 14000
rect 25004 13988 25010 14000
rect 25041 13991 25099 13997
rect 25041 13988 25053 13991
rect 25004 13960 25053 13988
rect 25004 13948 25010 13960
rect 25041 13957 25053 13960
rect 25087 13957 25099 13991
rect 25041 13951 25099 13957
rect 23492 13892 23796 13920
rect 21545 13883 21603 13889
rect 21818 13852 21824 13864
rect 20579 13824 20668 13852
rect 20732 13824 21824 13852
rect 20579 13821 20591 13824
rect 20533 13815 20591 13821
rect 17865 13787 17923 13793
rect 17865 13753 17877 13787
rect 17911 13784 17923 13787
rect 18316 13787 18374 13793
rect 18316 13784 18328 13787
rect 17911 13756 18328 13784
rect 17911 13753 17923 13756
rect 17865 13747 17923 13753
rect 18316 13753 18328 13756
rect 18362 13784 18374 13787
rect 19978 13784 19984 13796
rect 18362 13756 19984 13784
rect 18362 13753 18374 13756
rect 18316 13747 18374 13753
rect 19978 13744 19984 13756
rect 20036 13744 20042 13796
rect 20640 13784 20668 13824
rect 21468 13793 21496 13824
rect 21818 13812 21824 13824
rect 21876 13812 21882 13864
rect 22370 13852 22376 13864
rect 22331 13824 22376 13852
rect 22370 13812 22376 13824
rect 22428 13812 22434 13864
rect 22554 13852 22560 13864
rect 22515 13824 22560 13852
rect 22554 13812 22560 13824
rect 22612 13812 22618 13864
rect 23661 13855 23719 13861
rect 23661 13821 23673 13855
rect 23707 13821 23719 13855
rect 23768 13852 23796 13892
rect 23917 13855 23975 13861
rect 23917 13852 23929 13855
rect 23768 13824 23929 13852
rect 23661 13815 23719 13821
rect 23917 13821 23929 13824
rect 23963 13821 23975 13855
rect 23917 13815 23975 13821
rect 21453 13787 21511 13793
rect 20640 13756 21404 13784
rect 21376 13728 21404 13756
rect 21453 13753 21465 13787
rect 21499 13753 21511 13787
rect 21453 13747 21511 13753
rect 5169 13719 5227 13725
rect 5169 13716 5181 13719
rect 4991 13688 5181 13716
rect 4893 13679 4951 13685
rect 5169 13685 5181 13688
rect 5215 13685 5227 13719
rect 5534 13716 5540 13728
rect 5495 13688 5540 13716
rect 5169 13679 5227 13685
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 11054 13716 11060 13728
rect 11015 13688 11060 13716
rect 11054 13676 11060 13688
rect 11112 13676 11118 13728
rect 12526 13676 12532 13728
rect 12584 13716 12590 13728
rect 12805 13719 12863 13725
rect 12805 13716 12817 13719
rect 12584 13688 12817 13716
rect 12584 13676 12590 13688
rect 12805 13685 12817 13688
rect 12851 13685 12863 13719
rect 12805 13679 12863 13685
rect 13722 13676 13728 13728
rect 13780 13716 13786 13728
rect 13817 13719 13875 13725
rect 13817 13716 13829 13719
rect 13780 13688 13829 13716
rect 13780 13676 13786 13688
rect 13817 13685 13829 13688
rect 13863 13716 13875 13719
rect 14369 13719 14427 13725
rect 14369 13716 14381 13719
rect 13863 13688 14381 13716
rect 13863 13685 13875 13688
rect 13817 13679 13875 13685
rect 14369 13685 14381 13688
rect 14415 13716 14427 13719
rect 17770 13716 17776 13728
rect 14415 13688 17776 13716
rect 14415 13685 14427 13688
rect 14369 13679 14427 13685
rect 17770 13676 17776 13688
rect 17828 13676 17834 13728
rect 19334 13676 19340 13728
rect 19392 13716 19398 13728
rect 20806 13716 20812 13728
rect 19392 13688 20812 13716
rect 19392 13676 19398 13688
rect 20806 13676 20812 13688
rect 20864 13676 20870 13728
rect 21358 13716 21364 13728
rect 21319 13688 21364 13716
rect 21358 13676 21364 13688
rect 21416 13676 21422 13728
rect 22186 13676 22192 13728
rect 22244 13716 22250 13728
rect 22738 13716 22744 13728
rect 22244 13688 22744 13716
rect 22244 13676 22250 13688
rect 22738 13676 22744 13688
rect 22796 13676 22802 13728
rect 23676 13716 23704 13815
rect 23842 13716 23848 13728
rect 23676 13688 23848 13716
rect 23842 13676 23848 13688
rect 23900 13676 23906 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1946 13512 1952 13524
rect 1907 13484 1952 13512
rect 1946 13472 1952 13484
rect 2004 13472 2010 13524
rect 2498 13472 2504 13524
rect 2556 13512 2562 13524
rect 2774 13512 2780 13524
rect 2556 13484 2780 13512
rect 2556 13472 2562 13484
rect 2774 13472 2780 13484
rect 2832 13512 2838 13524
rect 2869 13515 2927 13521
rect 2869 13512 2881 13515
rect 2832 13484 2881 13512
rect 2832 13472 2838 13484
rect 2869 13481 2881 13484
rect 2915 13481 2927 13515
rect 2869 13475 2927 13481
rect 3513 13515 3571 13521
rect 3513 13481 3525 13515
rect 3559 13512 3571 13515
rect 3786 13512 3792 13524
rect 3559 13484 3792 13512
rect 3559 13481 3571 13484
rect 3513 13475 3571 13481
rect 3786 13472 3792 13484
rect 3844 13472 3850 13524
rect 3881 13515 3939 13521
rect 3881 13481 3893 13515
rect 3927 13512 3939 13515
rect 3970 13512 3976 13524
rect 3927 13484 3976 13512
rect 3927 13481 3939 13484
rect 3881 13475 3939 13481
rect 3970 13472 3976 13484
rect 4028 13472 4034 13524
rect 4522 13472 4528 13524
rect 4580 13512 4586 13524
rect 4801 13515 4859 13521
rect 4801 13512 4813 13515
rect 4580 13484 4813 13512
rect 4580 13472 4586 13484
rect 4801 13481 4813 13484
rect 4847 13481 4859 13515
rect 4801 13475 4859 13481
rect 5718 13472 5724 13524
rect 5776 13512 5782 13524
rect 6546 13512 6552 13524
rect 5776 13484 6552 13512
rect 5776 13472 5782 13484
rect 6546 13472 6552 13484
rect 6604 13512 6610 13524
rect 6917 13515 6975 13521
rect 6917 13512 6929 13515
rect 6604 13484 6929 13512
rect 6604 13472 6610 13484
rect 6917 13481 6929 13484
rect 6963 13481 6975 13515
rect 8018 13512 8024 13524
rect 7979 13484 8024 13512
rect 6917 13475 6975 13481
rect 8018 13472 8024 13484
rect 8076 13472 8082 13524
rect 8386 13512 8392 13524
rect 8347 13484 8392 13512
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 8481 13515 8539 13521
rect 8481 13481 8493 13515
rect 8527 13512 8539 13515
rect 8662 13512 8668 13524
rect 8527 13484 8668 13512
rect 8527 13481 8539 13484
rect 8481 13475 8539 13481
rect 8662 13472 8668 13484
rect 8720 13472 8726 13524
rect 9125 13515 9183 13521
rect 9125 13481 9137 13515
rect 9171 13512 9183 13515
rect 9398 13512 9404 13524
rect 9171 13484 9404 13512
rect 9171 13481 9183 13484
rect 9125 13475 9183 13481
rect 9398 13472 9404 13484
rect 9456 13472 9462 13524
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 13538 13512 13544 13524
rect 12860 13484 13544 13512
rect 12860 13472 12866 13484
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 17954 13472 17960 13524
rect 18012 13512 18018 13524
rect 18049 13515 18107 13521
rect 18049 13512 18061 13515
rect 18012 13484 18061 13512
rect 18012 13472 18018 13484
rect 18049 13481 18061 13484
rect 18095 13481 18107 13515
rect 18049 13475 18107 13481
rect 19521 13515 19579 13521
rect 19521 13481 19533 13515
rect 19567 13512 19579 13515
rect 20162 13512 20168 13524
rect 19567 13484 20168 13512
rect 19567 13481 19579 13484
rect 19521 13475 19579 13481
rect 20162 13472 20168 13484
rect 20220 13472 20226 13524
rect 20717 13515 20775 13521
rect 20717 13481 20729 13515
rect 20763 13512 20775 13515
rect 21450 13512 21456 13524
rect 20763 13484 21456 13512
rect 20763 13481 20775 13484
rect 20717 13475 20775 13481
rect 21450 13472 21456 13484
rect 21508 13512 21514 13524
rect 21545 13515 21603 13521
rect 21545 13512 21557 13515
rect 21508 13484 21557 13512
rect 21508 13472 21514 13484
rect 21545 13481 21557 13484
rect 21591 13481 21603 13515
rect 21545 13475 21603 13481
rect 22281 13515 22339 13521
rect 22281 13481 22293 13515
rect 22327 13512 22339 13515
rect 22646 13512 22652 13524
rect 22327 13484 22652 13512
rect 22327 13481 22339 13484
rect 22281 13475 22339 13481
rect 22646 13472 22652 13484
rect 22704 13472 22710 13524
rect 22741 13515 22799 13521
rect 22741 13481 22753 13515
rect 22787 13512 22799 13515
rect 23106 13512 23112 13524
rect 22787 13484 23112 13512
rect 22787 13481 22799 13484
rect 22741 13475 22799 13481
rect 23106 13472 23112 13484
rect 23164 13472 23170 13524
rect 4341 13447 4399 13453
rect 4341 13413 4353 13447
rect 4387 13444 4399 13447
rect 4982 13444 4988 13456
rect 4387 13416 4988 13444
rect 4387 13413 4399 13416
rect 4341 13407 4399 13413
rect 4982 13404 4988 13416
rect 5040 13404 5046 13456
rect 5261 13447 5319 13453
rect 5261 13413 5273 13447
rect 5307 13444 5319 13447
rect 5534 13444 5540 13456
rect 5307 13416 5540 13444
rect 5307 13413 5319 13416
rect 5261 13407 5319 13413
rect 5534 13404 5540 13416
rect 5592 13444 5598 13456
rect 6822 13444 6828 13456
rect 5592 13416 6828 13444
rect 5592 13404 5598 13416
rect 6822 13404 6828 13416
rect 6880 13404 6886 13456
rect 2777 13379 2835 13385
rect 2777 13345 2789 13379
rect 2823 13376 2835 13379
rect 3050 13376 3056 13388
rect 2823 13348 3056 13376
rect 2823 13345 2835 13348
rect 2777 13339 2835 13345
rect 3050 13336 3056 13348
rect 3108 13376 3114 13388
rect 3602 13376 3608 13388
rect 3108 13348 3608 13376
rect 3108 13336 3114 13348
rect 3602 13336 3608 13348
rect 3660 13376 3666 13388
rect 3660 13348 3924 13376
rect 3660 13336 3666 13348
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13268 1458 13320
rect 2958 13308 2964 13320
rect 2919 13280 2964 13308
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 3896 13308 3924 13348
rect 3970 13336 3976 13388
rect 4028 13376 4034 13388
rect 4065 13379 4123 13385
rect 4065 13376 4077 13379
rect 4028 13348 4077 13376
rect 4028 13336 4034 13348
rect 4065 13345 4077 13348
rect 4111 13345 4123 13379
rect 4065 13339 4123 13345
rect 5626 13336 5632 13388
rect 5684 13376 5690 13388
rect 5804 13379 5862 13385
rect 5804 13376 5816 13379
rect 5684 13348 5816 13376
rect 5684 13336 5690 13348
rect 5804 13345 5816 13348
rect 5850 13376 5862 13379
rect 6178 13376 6184 13388
rect 5850 13348 6184 13376
rect 5850 13345 5862 13348
rect 5804 13339 5862 13345
rect 6178 13336 6184 13348
rect 6236 13376 6242 13388
rect 6730 13376 6736 13388
rect 6236 13348 6736 13376
rect 6236 13336 6242 13348
rect 6730 13336 6736 13348
rect 6788 13336 6794 13388
rect 9416 13376 9444 13472
rect 9953 13447 10011 13453
rect 9953 13413 9965 13447
rect 9999 13444 10011 13447
rect 12526 13444 12532 13456
rect 9999 13416 12532 13444
rect 9999 13413 10011 13416
rect 9953 13407 10011 13413
rect 12526 13404 12532 13416
rect 12584 13404 12590 13456
rect 21082 13404 21088 13456
rect 21140 13444 21146 13456
rect 21913 13447 21971 13453
rect 21913 13444 21925 13447
rect 21140 13416 21925 13444
rect 21140 13404 21146 13416
rect 21913 13413 21925 13416
rect 21959 13413 21971 13447
rect 21913 13407 21971 13413
rect 10229 13379 10287 13385
rect 10229 13376 10241 13379
rect 9416 13348 10241 13376
rect 10229 13345 10241 13348
rect 10275 13345 10287 13379
rect 10229 13339 10287 13345
rect 10318 13336 10324 13388
rect 10376 13376 10382 13388
rect 10485 13379 10543 13385
rect 10485 13376 10497 13379
rect 10376 13348 10497 13376
rect 10376 13336 10382 13348
rect 10485 13345 10497 13348
rect 10531 13345 10543 13379
rect 10485 13339 10543 13345
rect 12158 13336 12164 13388
rect 12216 13376 12222 13388
rect 15562 13385 15568 13388
rect 12713 13379 12771 13385
rect 12713 13376 12725 13379
rect 12216 13348 12725 13376
rect 12216 13336 12222 13348
rect 12713 13345 12725 13348
rect 12759 13345 12771 13379
rect 12713 13339 12771 13345
rect 15556 13339 15568 13385
rect 15620 13376 15626 13388
rect 17589 13379 17647 13385
rect 15620 13348 15656 13376
rect 15562 13336 15568 13339
rect 15620 13336 15626 13348
rect 17589 13345 17601 13379
rect 17635 13376 17647 13379
rect 18230 13376 18236 13388
rect 17635 13348 18236 13376
rect 17635 13345 17647 13348
rect 17589 13339 17647 13345
rect 18230 13336 18236 13348
rect 18288 13376 18294 13388
rect 18417 13379 18475 13385
rect 18417 13376 18429 13379
rect 18288 13348 18429 13376
rect 18288 13336 18294 13348
rect 18417 13345 18429 13348
rect 18463 13345 18475 13379
rect 20990 13376 20996 13388
rect 20951 13348 20996 13376
rect 18417 13339 18475 13345
rect 20990 13336 20996 13348
rect 21048 13336 21054 13388
rect 22094 13336 22100 13388
rect 22152 13376 22158 13388
rect 22152 13348 22197 13376
rect 22152 13336 22158 13348
rect 23934 13336 23940 13388
rect 23992 13376 23998 13388
rect 24121 13379 24179 13385
rect 24121 13376 24133 13379
rect 23992 13348 24133 13376
rect 23992 13336 23998 13348
rect 24121 13345 24133 13348
rect 24167 13376 24179 13379
rect 24857 13379 24915 13385
rect 24857 13376 24869 13379
rect 24167 13348 24869 13376
rect 24167 13345 24179 13348
rect 24121 13339 24179 13345
rect 24857 13345 24869 13348
rect 24903 13345 24915 13379
rect 24857 13339 24915 13345
rect 4890 13308 4896 13320
rect 3896 13280 4896 13308
rect 4890 13268 4896 13280
rect 4948 13268 4954 13320
rect 5537 13311 5595 13317
rect 5537 13277 5549 13311
rect 5583 13277 5595 13311
rect 5537 13271 5595 13277
rect 4430 13200 4436 13252
rect 4488 13240 4494 13252
rect 5258 13240 5264 13252
rect 4488 13212 5264 13240
rect 4488 13200 4494 13212
rect 5258 13200 5264 13212
rect 5316 13240 5322 13252
rect 5552 13240 5580 13271
rect 8570 13268 8576 13320
rect 8628 13308 8634 13320
rect 9674 13308 9680 13320
rect 8628 13280 9680 13308
rect 8628 13268 8634 13280
rect 9674 13268 9680 13280
rect 9732 13268 9738 13320
rect 14366 13268 14372 13320
rect 14424 13308 14430 13320
rect 14826 13308 14832 13320
rect 14424 13280 14832 13308
rect 14424 13268 14430 13280
rect 14826 13268 14832 13280
rect 14884 13308 14890 13320
rect 15289 13311 15347 13317
rect 15289 13308 15301 13311
rect 14884 13280 15301 13308
rect 14884 13268 14890 13280
rect 15289 13277 15301 13280
rect 15335 13277 15347 13311
rect 15289 13271 15347 13277
rect 17957 13311 18015 13317
rect 17957 13277 17969 13311
rect 18003 13308 18015 13311
rect 18506 13308 18512 13320
rect 18003 13280 18512 13308
rect 18003 13277 18015 13280
rect 17957 13271 18015 13277
rect 18506 13268 18512 13280
rect 18564 13268 18570 13320
rect 18598 13268 18604 13320
rect 18656 13308 18662 13320
rect 19058 13308 19064 13320
rect 18656 13280 19064 13308
rect 18656 13268 18662 13280
rect 19058 13268 19064 13280
rect 19116 13268 19122 13320
rect 19610 13308 19616 13320
rect 19571 13280 19616 13308
rect 19610 13268 19616 13280
rect 19668 13268 19674 13320
rect 23474 13268 23480 13320
rect 23532 13308 23538 13320
rect 24305 13311 24363 13317
rect 24305 13308 24317 13311
rect 23532 13280 24317 13308
rect 23532 13268 23538 13280
rect 24305 13277 24317 13280
rect 24351 13277 24363 13311
rect 25406 13308 25412 13320
rect 25367 13280 25412 13308
rect 24305 13271 24363 13277
rect 25406 13268 25412 13280
rect 25464 13268 25470 13320
rect 21174 13240 21180 13252
rect 5316 13212 5580 13240
rect 21135 13212 21180 13240
rect 5316 13200 5322 13212
rect 2222 13172 2228 13184
rect 2183 13144 2228 13172
rect 2222 13132 2228 13144
rect 2280 13132 2286 13184
rect 2409 13175 2467 13181
rect 2409 13141 2421 13175
rect 2455 13172 2467 13175
rect 3694 13172 3700 13184
rect 2455 13144 3700 13172
rect 2455 13141 2467 13144
rect 2409 13135 2467 13141
rect 3694 13132 3700 13144
rect 3752 13132 3758 13184
rect 5552 13172 5580 13212
rect 21174 13200 21180 13212
rect 21232 13200 21238 13252
rect 23750 13200 23756 13252
rect 23808 13240 23814 13252
rect 23934 13240 23940 13252
rect 23808 13212 23940 13240
rect 23808 13200 23814 13212
rect 23934 13200 23940 13212
rect 23992 13200 23998 13252
rect 6822 13172 6828 13184
rect 5552 13144 6828 13172
rect 6822 13132 6828 13144
rect 6880 13172 6886 13184
rect 7469 13175 7527 13181
rect 7469 13172 7481 13175
rect 6880 13144 7481 13172
rect 6880 13132 6886 13144
rect 7469 13141 7481 13144
rect 7515 13141 7527 13175
rect 11606 13172 11612 13184
rect 11567 13144 11612 13172
rect 7469 13135 7527 13141
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 13998 13172 14004 13184
rect 13959 13144 14004 13172
rect 13998 13132 14004 13144
rect 14056 13132 14062 13184
rect 14274 13132 14280 13184
rect 14332 13172 14338 13184
rect 14737 13175 14795 13181
rect 14737 13172 14749 13175
rect 14332 13144 14749 13172
rect 14332 13132 14338 13144
rect 14737 13141 14749 13144
rect 14783 13141 14795 13175
rect 16666 13172 16672 13184
rect 16627 13144 16672 13172
rect 14737 13135 14795 13141
rect 16666 13132 16672 13144
rect 16724 13132 16730 13184
rect 23661 13175 23719 13181
rect 23661 13141 23673 13175
rect 23707 13172 23719 13175
rect 23842 13172 23848 13184
rect 23707 13144 23848 13172
rect 23707 13141 23719 13144
rect 23661 13135 23719 13141
rect 23842 13132 23848 13144
rect 23900 13132 23906 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 3050 12928 3056 12980
rect 3108 12968 3114 12980
rect 3145 12971 3203 12977
rect 3145 12968 3157 12971
rect 3108 12940 3157 12968
rect 3108 12928 3114 12940
rect 3145 12937 3157 12940
rect 3191 12937 3203 12971
rect 3326 12968 3332 12980
rect 3287 12940 3332 12968
rect 3145 12931 3203 12937
rect 3326 12928 3332 12940
rect 3384 12928 3390 12980
rect 4706 12928 4712 12980
rect 4764 12968 4770 12980
rect 4985 12971 5043 12977
rect 4985 12968 4997 12971
rect 4764 12940 4997 12968
rect 4764 12928 4770 12940
rect 4985 12937 4997 12940
rect 5031 12937 5043 12971
rect 4985 12931 5043 12937
rect 5169 12971 5227 12977
rect 5169 12937 5181 12971
rect 5215 12968 5227 12971
rect 5442 12968 5448 12980
rect 5215 12940 5448 12968
rect 5215 12937 5227 12940
rect 5169 12931 5227 12937
rect 1673 12903 1731 12909
rect 1673 12869 1685 12903
rect 1719 12900 1731 12903
rect 1719 12872 2452 12900
rect 1719 12869 1731 12872
rect 1673 12863 1731 12869
rect 2222 12832 2228 12844
rect 2183 12804 2228 12832
rect 2222 12792 2228 12804
rect 2280 12792 2286 12844
rect 2424 12841 2452 12872
rect 2409 12835 2467 12841
rect 2409 12801 2421 12835
rect 2455 12832 2467 12835
rect 2682 12832 2688 12844
rect 2455 12804 2688 12832
rect 2455 12801 2467 12804
rect 2409 12795 2467 12801
rect 2682 12792 2688 12804
rect 2740 12792 2746 12844
rect 3878 12832 3884 12844
rect 3839 12804 3884 12832
rect 3878 12792 3884 12804
rect 3936 12792 3942 12844
rect 5000 12832 5028 12931
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 6178 12968 6184 12980
rect 6139 12940 6184 12968
rect 6178 12928 6184 12940
rect 6236 12928 6242 12980
rect 6546 12968 6552 12980
rect 6507 12940 6552 12968
rect 6546 12928 6552 12940
rect 6604 12928 6610 12980
rect 8662 12928 8668 12980
rect 8720 12968 8726 12980
rect 8757 12971 8815 12977
rect 8757 12968 8769 12971
rect 8720 12940 8769 12968
rect 8720 12928 8726 12940
rect 8757 12937 8769 12940
rect 8803 12937 8815 12971
rect 8757 12931 8815 12937
rect 9309 12971 9367 12977
rect 9309 12937 9321 12971
rect 9355 12968 9367 12971
rect 9398 12968 9404 12980
rect 9355 12940 9404 12968
rect 9355 12937 9367 12940
rect 9309 12931 9367 12937
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 10042 12928 10048 12980
rect 10100 12968 10106 12980
rect 10597 12971 10655 12977
rect 10597 12968 10609 12971
rect 10100 12940 10609 12968
rect 10100 12928 10106 12940
rect 10597 12937 10609 12940
rect 10643 12937 10655 12971
rect 10597 12931 10655 12937
rect 13541 12971 13599 12977
rect 13541 12937 13553 12971
rect 13587 12968 13599 12971
rect 14090 12968 14096 12980
rect 13587 12940 14096 12968
rect 13587 12937 13599 12940
rect 13541 12931 13599 12937
rect 5629 12835 5687 12841
rect 5629 12832 5641 12835
rect 5000 12804 5641 12832
rect 5629 12801 5641 12804
rect 5675 12801 5687 12835
rect 5629 12795 5687 12801
rect 5718 12792 5724 12844
rect 5776 12832 5782 12844
rect 5813 12835 5871 12841
rect 5813 12832 5825 12835
rect 5776 12804 5825 12832
rect 5776 12792 5782 12804
rect 5813 12801 5825 12804
rect 5859 12832 5871 12835
rect 6270 12832 6276 12844
rect 5859 12804 6276 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 6270 12792 6276 12804
rect 6328 12792 6334 12844
rect 6564 12832 6592 12928
rect 10318 12900 10324 12912
rect 10279 12872 10324 12900
rect 10318 12860 10324 12872
rect 10376 12860 10382 12912
rect 10612 12900 10640 12931
rect 14090 12928 14096 12940
rect 14148 12928 14154 12980
rect 15562 12928 15568 12980
rect 15620 12968 15626 12980
rect 15749 12971 15807 12977
rect 15749 12968 15761 12971
rect 15620 12940 15761 12968
rect 15620 12928 15626 12940
rect 15749 12937 15761 12940
rect 15795 12968 15807 12971
rect 15838 12968 15844 12980
rect 15795 12940 15844 12968
rect 15795 12937 15807 12940
rect 15749 12931 15807 12937
rect 15838 12928 15844 12940
rect 15896 12968 15902 12980
rect 16301 12971 16359 12977
rect 16301 12968 16313 12971
rect 15896 12940 16313 12968
rect 15896 12928 15902 12940
rect 16301 12937 16313 12940
rect 16347 12937 16359 12971
rect 18230 12968 18236 12980
rect 18191 12940 18236 12968
rect 16301 12931 16359 12937
rect 18230 12928 18236 12940
rect 18288 12928 18294 12980
rect 19242 12928 19248 12980
rect 19300 12968 19306 12980
rect 19797 12971 19855 12977
rect 19797 12968 19809 12971
rect 19300 12940 19809 12968
rect 19300 12928 19306 12940
rect 19797 12937 19809 12940
rect 19843 12937 19855 12971
rect 20990 12968 20996 12980
rect 20951 12940 20996 12968
rect 19797 12931 19855 12937
rect 20990 12928 20996 12940
rect 21048 12928 21054 12980
rect 21545 12971 21603 12977
rect 21545 12937 21557 12971
rect 21591 12968 21603 12971
rect 21634 12968 21640 12980
rect 21591 12940 21640 12968
rect 21591 12937 21603 12940
rect 21545 12931 21603 12937
rect 21634 12928 21640 12940
rect 21692 12928 21698 12980
rect 22094 12928 22100 12980
rect 22152 12968 22158 12980
rect 22649 12971 22707 12977
rect 22152 12940 22197 12968
rect 22152 12928 22158 12940
rect 22649 12937 22661 12971
rect 22695 12968 22707 12971
rect 23198 12968 23204 12980
rect 22695 12940 23204 12968
rect 22695 12937 22707 12940
rect 22649 12931 22707 12937
rect 23198 12928 23204 12940
rect 23256 12928 23262 12980
rect 11606 12900 11612 12912
rect 10612 12872 11612 12900
rect 9766 12832 9772 12844
rect 6564 12804 6960 12832
rect 9727 12804 9772 12832
rect 3510 12724 3516 12776
rect 3568 12764 3574 12776
rect 3789 12767 3847 12773
rect 3789 12764 3801 12767
rect 3568 12736 3801 12764
rect 3568 12724 3574 12736
rect 3789 12733 3801 12736
rect 3835 12733 3847 12767
rect 5534 12764 5540 12776
rect 5495 12736 5540 12764
rect 3789 12727 3847 12733
rect 5534 12724 5540 12736
rect 5592 12724 5598 12776
rect 6822 12764 6828 12776
rect 6783 12736 6828 12764
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 6932 12764 6960 12804
rect 9766 12792 9772 12804
rect 9824 12792 9830 12844
rect 7081 12767 7139 12773
rect 7081 12764 7093 12767
rect 6932 12736 7093 12764
rect 7081 12733 7093 12736
rect 7127 12733 7139 12767
rect 7081 12727 7139 12733
rect 9217 12767 9275 12773
rect 9217 12733 9229 12767
rect 9263 12764 9275 12767
rect 9493 12767 9551 12773
rect 9493 12764 9505 12767
rect 9263 12736 9505 12764
rect 9263 12733 9275 12736
rect 9217 12727 9275 12733
rect 9493 12733 9505 12736
rect 9539 12764 9551 12767
rect 9582 12764 9588 12776
rect 9539 12736 9588 12764
rect 9539 12733 9551 12736
rect 9493 12727 9551 12733
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 10336 12764 10364 12860
rect 11054 12792 11060 12844
rect 11112 12832 11118 12844
rect 11238 12832 11244 12844
rect 11112 12804 11244 12832
rect 11112 12792 11118 12804
rect 11238 12792 11244 12804
rect 11296 12792 11302 12844
rect 11348 12841 11376 12872
rect 11606 12860 11612 12872
rect 11664 12860 11670 12912
rect 17497 12903 17555 12909
rect 11808 12872 13032 12900
rect 11333 12835 11391 12841
rect 11333 12801 11345 12835
rect 11379 12801 11391 12835
rect 11333 12795 11391 12801
rect 11698 12764 11704 12776
rect 10336 12736 11704 12764
rect 11698 12724 11704 12736
rect 11756 12764 11762 12776
rect 11808 12773 11836 12872
rect 13004 12844 13032 12872
rect 17497 12869 17509 12903
rect 17543 12900 17555 12903
rect 19337 12903 19395 12909
rect 19337 12900 19349 12903
rect 17543 12872 19349 12900
rect 17543 12869 17555 12872
rect 17497 12863 17555 12869
rect 12894 12832 12900 12844
rect 12855 12804 12900 12832
rect 12894 12792 12900 12804
rect 12952 12792 12958 12844
rect 12986 12792 12992 12844
rect 13044 12832 13050 12844
rect 14090 12832 14096 12844
rect 13044 12804 13089 12832
rect 14051 12804 14096 12832
rect 13044 12792 13050 12804
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 14366 12832 14372 12844
rect 14327 12804 14372 12832
rect 14366 12792 14372 12804
rect 14424 12792 14430 12844
rect 17770 12792 17776 12844
rect 17828 12832 17834 12844
rect 17865 12835 17923 12841
rect 17865 12832 17877 12835
rect 17828 12804 17877 12832
rect 17828 12792 17834 12804
rect 17865 12801 17877 12804
rect 17911 12832 17923 12835
rect 18690 12832 18696 12844
rect 17911 12804 18696 12832
rect 17911 12801 17923 12804
rect 17865 12795 17923 12801
rect 18690 12792 18696 12804
rect 18748 12792 18754 12844
rect 18892 12841 18920 12872
rect 19260 12844 19288 12872
rect 19337 12869 19349 12872
rect 19383 12900 19395 12903
rect 19978 12900 19984 12912
rect 19383 12872 19984 12900
rect 19383 12869 19395 12872
rect 19337 12863 19395 12869
rect 19978 12860 19984 12872
rect 20036 12900 20042 12912
rect 20036 12872 20392 12900
rect 20036 12860 20042 12872
rect 18877 12835 18935 12841
rect 18877 12801 18889 12835
rect 18923 12801 18935 12835
rect 18877 12795 18935 12801
rect 19242 12792 19248 12844
rect 19300 12792 19306 12844
rect 19702 12832 19708 12844
rect 19663 12804 19708 12832
rect 19702 12792 19708 12804
rect 19760 12792 19766 12844
rect 20364 12841 20392 12872
rect 24946 12860 24952 12912
rect 25004 12860 25010 12912
rect 20349 12835 20407 12841
rect 20349 12801 20361 12835
rect 20395 12801 20407 12835
rect 20349 12795 20407 12801
rect 20806 12792 20812 12844
rect 20864 12832 20870 12844
rect 23017 12835 23075 12841
rect 23017 12832 23029 12835
rect 20864 12804 23029 12832
rect 20864 12792 20870 12804
rect 11793 12767 11851 12773
rect 11793 12764 11805 12767
rect 11756 12736 11805 12764
rect 11756 12724 11762 12736
rect 11793 12733 11805 12736
rect 11839 12733 11851 12767
rect 11793 12727 11851 12733
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 12492 12736 12817 12764
rect 12492 12724 12498 12736
rect 12805 12733 12817 12736
rect 12851 12764 12863 12767
rect 14274 12764 14280 12776
rect 12851 12736 14280 12764
rect 12851 12733 12863 12736
rect 12805 12727 12863 12733
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 18322 12724 18328 12776
rect 18380 12764 18386 12776
rect 18601 12767 18659 12773
rect 18601 12764 18613 12767
rect 18380 12736 18613 12764
rect 18380 12724 18386 12736
rect 18601 12733 18613 12736
rect 18647 12764 18659 12767
rect 19610 12764 19616 12776
rect 18647 12736 19616 12764
rect 18647 12733 18659 12736
rect 18601 12727 18659 12733
rect 19610 12724 19616 12736
rect 19668 12724 19674 12776
rect 19720 12764 19748 12792
rect 19978 12764 19984 12776
rect 19720 12736 19984 12764
rect 19978 12724 19984 12736
rect 20036 12724 20042 12776
rect 20165 12767 20223 12773
rect 20165 12733 20177 12767
rect 20211 12764 20223 12767
rect 20254 12764 20260 12776
rect 20211 12736 20260 12764
rect 20211 12733 20223 12736
rect 20165 12727 20223 12733
rect 3970 12696 3976 12708
rect 1780 12668 3976 12696
rect 1780 12637 1808 12668
rect 3970 12656 3976 12668
rect 4028 12656 4034 12708
rect 4709 12699 4767 12705
rect 4709 12665 4721 12699
rect 4755 12696 4767 12699
rect 5718 12696 5724 12708
rect 4755 12668 5724 12696
rect 4755 12665 4767 12668
rect 4709 12659 4767 12665
rect 5718 12656 5724 12668
rect 5776 12656 5782 12708
rect 11164 12668 12480 12696
rect 1765 12631 1823 12637
rect 1765 12597 1777 12631
rect 1811 12597 1823 12631
rect 2130 12628 2136 12640
rect 2091 12600 2136 12628
rect 1765 12591 1823 12597
rect 2130 12588 2136 12600
rect 2188 12588 2194 12640
rect 2774 12588 2780 12640
rect 2832 12628 2838 12640
rect 3694 12628 3700 12640
rect 2832 12600 2877 12628
rect 3655 12600 3700 12628
rect 2832 12588 2838 12600
rect 3694 12588 3700 12600
rect 3752 12588 3758 12640
rect 7834 12588 7840 12640
rect 7892 12628 7898 12640
rect 8205 12631 8263 12637
rect 8205 12628 8217 12631
rect 7892 12600 8217 12628
rect 7892 12588 7898 12600
rect 8205 12597 8217 12600
rect 8251 12597 8263 12631
rect 10778 12628 10784 12640
rect 10739 12600 10784 12628
rect 8205 12591 8263 12597
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 11054 12588 11060 12640
rect 11112 12628 11118 12640
rect 11164 12637 11192 12668
rect 11149 12631 11207 12637
rect 11149 12628 11161 12631
rect 11112 12600 11161 12628
rect 11112 12588 11118 12600
rect 11149 12597 11161 12600
rect 11195 12597 11207 12631
rect 12158 12628 12164 12640
rect 12119 12600 12164 12628
rect 11149 12591 11207 12597
rect 12158 12588 12164 12600
rect 12216 12588 12222 12640
rect 12452 12637 12480 12668
rect 14182 12656 14188 12708
rect 14240 12696 14246 12708
rect 14614 12699 14672 12705
rect 14614 12696 14626 12699
rect 14240 12668 14626 12696
rect 14240 12656 14246 12668
rect 14614 12665 14626 12668
rect 14660 12665 14672 12699
rect 14614 12659 14672 12665
rect 15010 12656 15016 12708
rect 15068 12696 15074 12708
rect 15654 12696 15660 12708
rect 15068 12668 15660 12696
rect 15068 12656 15074 12668
rect 15654 12656 15660 12668
rect 15712 12696 15718 12708
rect 15930 12696 15936 12708
rect 15712 12668 15936 12696
rect 15712 12656 15718 12668
rect 15930 12656 15936 12668
rect 15988 12656 15994 12708
rect 16574 12656 16580 12708
rect 16632 12696 16638 12708
rect 16853 12699 16911 12705
rect 16853 12696 16865 12699
rect 16632 12668 16865 12696
rect 16632 12656 16638 12668
rect 16853 12665 16865 12668
rect 16899 12665 16911 12699
rect 16853 12659 16911 12665
rect 19518 12656 19524 12708
rect 19576 12696 19582 12708
rect 20180 12696 20208 12727
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 21082 12724 21088 12776
rect 21140 12764 21146 12776
rect 22480 12773 22508 12804
rect 23017 12801 23029 12804
rect 23063 12801 23075 12835
rect 23017 12795 23075 12801
rect 23477 12835 23535 12841
rect 23477 12801 23489 12835
rect 23523 12832 23535 12835
rect 23523 12804 23980 12832
rect 23523 12801 23535 12804
rect 23477 12795 23535 12801
rect 21361 12767 21419 12773
rect 21361 12764 21373 12767
rect 21140 12736 21373 12764
rect 21140 12724 21146 12736
rect 21361 12733 21373 12736
rect 21407 12733 21419 12767
rect 21361 12727 21419 12733
rect 22465 12767 22523 12773
rect 22465 12733 22477 12767
rect 22511 12733 22523 12767
rect 23842 12764 23848 12776
rect 23755 12736 23848 12764
rect 22465 12727 22523 12733
rect 23842 12724 23848 12736
rect 23900 12724 23906 12776
rect 23952 12764 23980 12804
rect 24112 12767 24170 12773
rect 24112 12764 24124 12767
rect 23952 12736 24124 12764
rect 24112 12733 24124 12736
rect 24158 12764 24170 12767
rect 24964 12764 24992 12860
rect 24158 12736 24992 12764
rect 24158 12733 24170 12736
rect 24112 12727 24170 12733
rect 19576 12668 20208 12696
rect 23860 12696 23888 12724
rect 24026 12696 24032 12708
rect 23860 12668 24032 12696
rect 19576 12656 19582 12668
rect 24026 12656 24032 12668
rect 24084 12656 24090 12708
rect 25406 12696 25412 12708
rect 24780 12668 25412 12696
rect 24780 12640 24808 12668
rect 25406 12656 25412 12668
rect 25464 12656 25470 12708
rect 12437 12631 12495 12637
rect 12437 12597 12449 12631
rect 12483 12597 12495 12631
rect 13906 12628 13912 12640
rect 13867 12600 13912 12628
rect 12437 12591 12495 12597
rect 13906 12588 13912 12600
rect 13964 12588 13970 12640
rect 14001 12631 14059 12637
rect 14001 12597 14013 12631
rect 14047 12628 14059 12631
rect 15102 12628 15108 12640
rect 14047 12600 15108 12628
rect 14047 12597 14059 12600
rect 14001 12591 14059 12597
rect 15102 12588 15108 12600
rect 15160 12588 15166 12640
rect 16482 12588 16488 12640
rect 16540 12628 16546 12640
rect 16669 12631 16727 12637
rect 16669 12628 16681 12631
rect 16540 12600 16681 12628
rect 16540 12588 16546 12600
rect 16669 12597 16681 12600
rect 16715 12597 16727 12631
rect 16669 12591 16727 12597
rect 19978 12588 19984 12640
rect 20036 12628 20042 12640
rect 20257 12631 20315 12637
rect 20257 12628 20269 12631
rect 20036 12600 20269 12628
rect 20036 12588 20042 12600
rect 20257 12597 20269 12600
rect 20303 12628 20315 12631
rect 20622 12628 20628 12640
rect 20303 12600 20628 12628
rect 20303 12597 20315 12600
rect 20257 12591 20315 12597
rect 20622 12588 20628 12600
rect 20680 12588 20686 12640
rect 24762 12588 24768 12640
rect 24820 12588 24826 12640
rect 24854 12588 24860 12640
rect 24912 12628 24918 12640
rect 25225 12631 25283 12637
rect 25225 12628 25237 12631
rect 24912 12600 25237 12628
rect 24912 12588 24918 12600
rect 25225 12597 25237 12600
rect 25271 12597 25283 12631
rect 25225 12591 25283 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 2041 12427 2099 12433
rect 2041 12393 2053 12427
rect 2087 12424 2099 12427
rect 2130 12424 2136 12436
rect 2087 12396 2136 12424
rect 2087 12393 2099 12396
rect 2041 12387 2099 12393
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 3513 12427 3571 12433
rect 3513 12393 3525 12427
rect 3559 12424 3571 12427
rect 3878 12424 3884 12436
rect 3559 12396 3884 12424
rect 3559 12393 3571 12396
rect 3513 12387 3571 12393
rect 3878 12384 3884 12396
rect 3936 12384 3942 12436
rect 3970 12384 3976 12436
rect 4028 12424 4034 12436
rect 4617 12427 4675 12433
rect 4617 12424 4629 12427
rect 4028 12396 4629 12424
rect 4028 12384 4034 12396
rect 4617 12393 4629 12396
rect 4663 12393 4675 12427
rect 4617 12387 4675 12393
rect 5077 12427 5135 12433
rect 5077 12393 5089 12427
rect 5123 12424 5135 12427
rect 5166 12424 5172 12436
rect 5123 12396 5172 12424
rect 5123 12393 5135 12396
rect 5077 12387 5135 12393
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 6086 12424 6092 12436
rect 6047 12396 6092 12424
rect 6086 12384 6092 12396
rect 6144 12384 6150 12436
rect 6549 12427 6607 12433
rect 6549 12393 6561 12427
rect 6595 12424 6607 12427
rect 6822 12424 6828 12436
rect 6595 12396 6828 12424
rect 6595 12393 6607 12396
rect 6549 12387 6607 12393
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 7374 12384 7380 12436
rect 7432 12424 7438 12436
rect 7561 12427 7619 12433
rect 7561 12424 7573 12427
rect 7432 12396 7573 12424
rect 7432 12384 7438 12396
rect 7561 12393 7573 12396
rect 7607 12393 7619 12427
rect 7561 12387 7619 12393
rect 8205 12427 8263 12433
rect 8205 12393 8217 12427
rect 8251 12424 8263 12427
rect 8386 12424 8392 12436
rect 8251 12396 8392 12424
rect 8251 12393 8263 12396
rect 8205 12387 8263 12393
rect 8386 12384 8392 12396
rect 8444 12384 8450 12436
rect 8570 12424 8576 12436
rect 8531 12396 8576 12424
rect 8570 12384 8576 12396
rect 8628 12384 8634 12436
rect 9953 12427 10011 12433
rect 9953 12393 9965 12427
rect 9999 12424 10011 12427
rect 10870 12424 10876 12436
rect 9999 12396 10876 12424
rect 9999 12393 10011 12396
rect 9953 12387 10011 12393
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 12437 12427 12495 12433
rect 12437 12393 12449 12427
rect 12483 12424 12495 12427
rect 12986 12424 12992 12436
rect 12483 12396 12992 12424
rect 12483 12393 12495 12396
rect 12437 12387 12495 12393
rect 12986 12384 12992 12396
rect 13044 12384 13050 12436
rect 13449 12427 13507 12433
rect 13449 12393 13461 12427
rect 13495 12424 13507 12427
rect 14090 12424 14096 12436
rect 13495 12396 14096 12424
rect 13495 12393 13507 12396
rect 13449 12387 13507 12393
rect 14090 12384 14096 12396
rect 14148 12424 14154 12436
rect 14642 12424 14648 12436
rect 14148 12396 14648 12424
rect 14148 12384 14154 12396
rect 14642 12384 14648 12396
rect 14700 12424 14706 12436
rect 15289 12427 15347 12433
rect 14700 12396 15240 12424
rect 14700 12384 14706 12396
rect 2958 12316 2964 12368
rect 3016 12356 3022 12368
rect 3145 12359 3203 12365
rect 3145 12356 3157 12359
rect 3016 12328 3157 12356
rect 3016 12316 3022 12328
rect 3145 12325 3157 12328
rect 3191 12356 3203 12359
rect 4341 12359 4399 12365
rect 4341 12356 4353 12359
rect 3191 12328 4353 12356
rect 3191 12325 3203 12328
rect 3145 12319 3203 12325
rect 4341 12325 4353 12328
rect 4387 12356 4399 12359
rect 4522 12356 4528 12368
rect 4387 12328 4528 12356
rect 4387 12325 4399 12328
rect 4341 12319 4399 12325
rect 4522 12316 4528 12328
rect 4580 12356 4586 12368
rect 5258 12356 5264 12368
rect 4580 12328 5264 12356
rect 4580 12316 4586 12328
rect 5258 12316 5264 12328
rect 5316 12316 5322 12368
rect 10686 12316 10692 12368
rect 10744 12356 10750 12368
rect 10781 12359 10839 12365
rect 10781 12356 10793 12359
rect 10744 12328 10793 12356
rect 10744 12316 10750 12328
rect 10781 12325 10793 12328
rect 10827 12325 10839 12359
rect 10781 12319 10839 12325
rect 2406 12288 2412 12300
rect 2367 12260 2412 12288
rect 2406 12248 2412 12260
rect 2464 12248 2470 12300
rect 2590 12248 2596 12300
rect 2648 12288 2654 12300
rect 2648 12260 2728 12288
rect 2648 12248 2654 12260
rect 2130 12180 2136 12232
rect 2188 12220 2194 12232
rect 2188 12192 2452 12220
rect 2188 12180 2194 12192
rect 1949 12155 2007 12161
rect 1949 12121 1961 12155
rect 1995 12152 2007 12155
rect 2424 12152 2452 12192
rect 2498 12180 2504 12232
rect 2556 12220 2562 12232
rect 2700 12229 2728 12260
rect 5074 12248 5080 12300
rect 5132 12288 5138 12300
rect 5445 12291 5503 12297
rect 5445 12288 5457 12291
rect 5132 12260 5457 12288
rect 5132 12248 5138 12260
rect 5445 12257 5457 12260
rect 5491 12257 5503 12291
rect 5445 12251 5503 12257
rect 7190 12248 7196 12300
rect 7248 12288 7254 12300
rect 7466 12288 7472 12300
rect 7248 12260 7472 12288
rect 7248 12248 7254 12260
rect 7466 12248 7472 12260
rect 7524 12248 7530 12300
rect 9398 12248 9404 12300
rect 9456 12288 9462 12300
rect 9493 12291 9551 12297
rect 9493 12288 9505 12291
rect 9456 12260 9505 12288
rect 9456 12248 9462 12260
rect 9493 12257 9505 12260
rect 9539 12288 9551 12291
rect 11057 12291 11115 12297
rect 11057 12288 11069 12291
rect 9539 12260 11069 12288
rect 9539 12257 9551 12260
rect 9493 12251 9551 12257
rect 11057 12257 11069 12260
rect 11103 12288 11115 12291
rect 11146 12288 11152 12300
rect 11103 12260 11152 12288
rect 11103 12257 11115 12260
rect 11057 12251 11115 12257
rect 11146 12248 11152 12260
rect 11204 12248 11210 12300
rect 11330 12297 11336 12300
rect 11324 12288 11336 12297
rect 11291 12260 11336 12288
rect 11324 12251 11336 12260
rect 11388 12288 11394 12300
rect 12986 12288 12992 12300
rect 11388 12260 12992 12288
rect 11330 12248 11336 12251
rect 11388 12248 11394 12260
rect 12986 12248 12992 12260
rect 13044 12248 13050 12300
rect 13078 12248 13084 12300
rect 13136 12288 13142 12300
rect 13538 12288 13544 12300
rect 13136 12260 13544 12288
rect 13136 12248 13142 12260
rect 13538 12248 13544 12260
rect 13596 12248 13602 12300
rect 13814 12248 13820 12300
rect 13872 12288 13878 12300
rect 13909 12291 13967 12297
rect 13909 12288 13921 12291
rect 13872 12260 13921 12288
rect 13872 12248 13878 12260
rect 13909 12257 13921 12260
rect 13955 12257 13967 12291
rect 13909 12251 13967 12257
rect 2685 12223 2743 12229
rect 2556 12192 2601 12220
rect 2556 12180 2562 12192
rect 2685 12189 2697 12223
rect 2731 12189 2743 12223
rect 2685 12183 2743 12189
rect 4246 12180 4252 12232
rect 4304 12220 4310 12232
rect 5537 12223 5595 12229
rect 5537 12220 5549 12223
rect 4304 12192 5549 12220
rect 4304 12180 4310 12192
rect 5537 12189 5549 12192
rect 5583 12189 5595 12223
rect 5718 12220 5724 12232
rect 5679 12192 5724 12220
rect 5537 12183 5595 12189
rect 5718 12180 5724 12192
rect 5776 12180 5782 12232
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12220 7803 12223
rect 7834 12220 7840 12232
rect 7791 12192 7840 12220
rect 7791 12189 7803 12192
rect 7745 12183 7803 12189
rect 7834 12180 7840 12192
rect 7892 12180 7898 12232
rect 10045 12223 10103 12229
rect 10045 12189 10057 12223
rect 10091 12189 10103 12223
rect 10045 12183 10103 12189
rect 14001 12223 14059 12229
rect 14001 12189 14013 12223
rect 14047 12220 14059 12223
rect 14090 12220 14096 12232
rect 14047 12192 14096 12220
rect 14047 12189 14059 12192
rect 14001 12183 14059 12189
rect 3789 12155 3847 12161
rect 3789 12152 3801 12155
rect 1995 12124 2360 12152
rect 2424 12124 3801 12152
rect 1995 12121 2007 12124
rect 1949 12115 2007 12121
rect 2332 12084 2360 12124
rect 3789 12121 3801 12124
rect 3835 12121 3847 12155
rect 10060 12152 10088 12183
rect 14090 12180 14096 12192
rect 14148 12180 14154 12232
rect 14185 12223 14243 12229
rect 14185 12189 14197 12223
rect 14231 12220 14243 12223
rect 14366 12220 14372 12232
rect 14231 12192 14372 12220
rect 14231 12189 14243 12192
rect 14185 12183 14243 12189
rect 14366 12180 14372 12192
rect 14424 12180 14430 12232
rect 11054 12152 11060 12164
rect 10060 12124 11060 12152
rect 3789 12115 3847 12121
rect 11054 12112 11060 12124
rect 11112 12112 11118 12164
rect 12894 12112 12900 12164
rect 12952 12152 12958 12164
rect 13541 12155 13599 12161
rect 13541 12152 13553 12155
rect 12952 12124 13553 12152
rect 12952 12112 12958 12124
rect 13541 12121 13553 12124
rect 13587 12121 13599 12155
rect 15212 12152 15240 12396
rect 15289 12393 15301 12427
rect 15335 12424 15347 12427
rect 15378 12424 15384 12436
rect 15335 12396 15384 12424
rect 15335 12393 15347 12396
rect 15289 12387 15347 12393
rect 15378 12384 15384 12396
rect 15436 12384 15442 12436
rect 15562 12384 15568 12436
rect 15620 12424 15626 12436
rect 16114 12424 16120 12436
rect 15620 12396 16120 12424
rect 15620 12384 15626 12396
rect 16114 12384 16120 12396
rect 16172 12384 16178 12436
rect 16758 12384 16764 12436
rect 16816 12424 16822 12436
rect 17313 12427 17371 12433
rect 17313 12424 17325 12427
rect 16816 12396 17325 12424
rect 16816 12384 16822 12396
rect 17313 12393 17325 12396
rect 17359 12424 17371 12427
rect 17402 12424 17408 12436
rect 17359 12396 17408 12424
rect 17359 12393 17371 12396
rect 17313 12387 17371 12393
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 18322 12424 18328 12436
rect 18283 12396 18328 12424
rect 18322 12384 18328 12396
rect 18380 12384 18386 12436
rect 18506 12384 18512 12436
rect 18564 12424 18570 12436
rect 18693 12427 18751 12433
rect 18693 12424 18705 12427
rect 18564 12396 18705 12424
rect 18564 12384 18570 12396
rect 18693 12393 18705 12396
rect 18739 12393 18751 12427
rect 18693 12387 18751 12393
rect 19518 12384 19524 12436
rect 19576 12424 19582 12436
rect 19797 12427 19855 12433
rect 19797 12424 19809 12427
rect 19576 12396 19809 12424
rect 19576 12384 19582 12396
rect 19797 12393 19809 12396
rect 19843 12393 19855 12427
rect 20162 12424 20168 12436
rect 20123 12396 20168 12424
rect 19797 12387 19855 12393
rect 20162 12384 20168 12396
rect 20220 12384 20226 12436
rect 21637 12427 21695 12433
rect 21637 12393 21649 12427
rect 21683 12424 21695 12427
rect 21726 12424 21732 12436
rect 21683 12396 21732 12424
rect 21683 12393 21695 12396
rect 21637 12387 21695 12393
rect 21726 12384 21732 12396
rect 21784 12384 21790 12436
rect 22738 12424 22744 12436
rect 22699 12396 22744 12424
rect 22738 12384 22744 12396
rect 22796 12384 22802 12436
rect 24854 12424 24860 12436
rect 23943 12396 24860 12424
rect 15838 12316 15844 12368
rect 15896 12356 15902 12368
rect 17957 12359 18015 12365
rect 15896 12328 16988 12356
rect 15896 12316 15902 12328
rect 15657 12291 15715 12297
rect 15657 12257 15669 12291
rect 15703 12288 15715 12291
rect 16390 12288 16396 12300
rect 15703 12260 16396 12288
rect 15703 12257 15715 12260
rect 15657 12251 15715 12257
rect 16390 12248 16396 12260
rect 16448 12288 16454 12300
rect 16448 12260 16896 12288
rect 16448 12248 16454 12260
rect 15746 12220 15752 12232
rect 15707 12192 15752 12220
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 15841 12223 15899 12229
rect 15841 12189 15853 12223
rect 15887 12189 15899 12223
rect 15841 12183 15899 12189
rect 15856 12152 15884 12183
rect 15930 12152 15936 12164
rect 15212 12124 15936 12152
rect 13541 12115 13599 12121
rect 15930 12112 15936 12124
rect 15988 12152 15994 12164
rect 16666 12152 16672 12164
rect 15988 12124 16672 12152
rect 15988 12112 15994 12124
rect 16666 12112 16672 12124
rect 16724 12112 16730 12164
rect 16868 12161 16896 12260
rect 16960 12220 16988 12328
rect 17957 12325 17969 12359
rect 18003 12356 18015 12359
rect 18598 12356 18604 12368
rect 18003 12328 18604 12356
rect 18003 12325 18015 12328
rect 17957 12319 18015 12325
rect 18598 12316 18604 12328
rect 18656 12316 18662 12368
rect 19061 12359 19119 12365
rect 19061 12325 19073 12359
rect 19107 12356 19119 12359
rect 19150 12356 19156 12368
rect 19107 12328 19156 12356
rect 19107 12325 19119 12328
rect 19061 12319 19119 12325
rect 19150 12316 19156 12328
rect 19208 12316 19214 12368
rect 23014 12316 23020 12368
rect 23072 12356 23078 12368
rect 23943 12365 23971 12396
rect 24854 12384 24860 12396
rect 24912 12384 24918 12436
rect 23928 12359 23986 12365
rect 23928 12356 23940 12359
rect 23072 12328 23940 12356
rect 23072 12316 23078 12328
rect 23928 12325 23940 12328
rect 23974 12325 23986 12359
rect 23928 12319 23986 12325
rect 24578 12316 24584 12368
rect 24636 12316 24642 12368
rect 17034 12248 17040 12300
rect 17092 12288 17098 12300
rect 17221 12291 17279 12297
rect 17221 12288 17233 12291
rect 17092 12260 17233 12288
rect 17092 12248 17098 12260
rect 17221 12257 17233 12260
rect 17267 12257 17279 12291
rect 21450 12288 21456 12300
rect 21411 12260 21456 12288
rect 17221 12251 17279 12257
rect 21450 12248 21456 12260
rect 21508 12248 21514 12300
rect 22554 12288 22560 12300
rect 22515 12260 22560 12288
rect 22554 12248 22560 12260
rect 22612 12248 22618 12300
rect 23290 12248 23296 12300
rect 23348 12288 23354 12300
rect 23566 12288 23572 12300
rect 23348 12260 23572 12288
rect 23348 12248 23354 12260
rect 23566 12248 23572 12260
rect 23624 12248 23630 12300
rect 24596 12288 24624 12316
rect 24854 12288 24860 12300
rect 24596 12260 24860 12288
rect 24854 12248 24860 12260
rect 24912 12248 24918 12300
rect 17405 12223 17463 12229
rect 17405 12220 17417 12223
rect 16960 12192 17417 12220
rect 17405 12189 17417 12192
rect 17451 12220 17463 12223
rect 17678 12220 17684 12232
rect 17451 12192 17684 12220
rect 17451 12189 17463 12192
rect 17405 12183 17463 12189
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 18782 12180 18788 12232
rect 18840 12220 18846 12232
rect 19153 12223 19211 12229
rect 19153 12220 19165 12223
rect 18840 12192 19165 12220
rect 18840 12180 18846 12192
rect 19153 12189 19165 12192
rect 19199 12189 19211 12223
rect 19153 12183 19211 12189
rect 19242 12180 19248 12232
rect 19300 12220 19306 12232
rect 23661 12223 23719 12229
rect 19300 12192 19345 12220
rect 19300 12180 19306 12192
rect 23661 12189 23673 12223
rect 23707 12189 23719 12223
rect 23661 12183 23719 12189
rect 16853 12155 16911 12161
rect 16853 12121 16865 12155
rect 16899 12121 16911 12155
rect 16853 12115 16911 12121
rect 2774 12084 2780 12096
rect 2332 12056 2780 12084
rect 2774 12044 2780 12056
rect 2832 12044 2838 12096
rect 2958 12044 2964 12096
rect 3016 12084 3022 12096
rect 7101 12087 7159 12093
rect 7101 12084 7113 12087
rect 3016 12056 7113 12084
rect 3016 12044 3022 12056
rect 7101 12053 7113 12056
rect 7147 12053 7159 12087
rect 12986 12084 12992 12096
rect 12947 12056 12992 12084
rect 7101 12047 7159 12053
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 14182 12044 14188 12096
rect 14240 12084 14246 12096
rect 14553 12087 14611 12093
rect 14553 12084 14565 12087
rect 14240 12056 14565 12084
rect 14240 12044 14246 12056
rect 14553 12053 14565 12056
rect 14599 12053 14611 12087
rect 14553 12047 14611 12053
rect 15013 12087 15071 12093
rect 15013 12053 15025 12087
rect 15059 12084 15071 12087
rect 15562 12084 15568 12096
rect 15059 12056 15568 12084
rect 15059 12053 15071 12056
rect 15013 12047 15071 12053
rect 15562 12044 15568 12056
rect 15620 12044 15626 12096
rect 16393 12087 16451 12093
rect 16393 12053 16405 12087
rect 16439 12084 16451 12087
rect 16482 12084 16488 12096
rect 16439 12056 16488 12084
rect 16439 12053 16451 12056
rect 16393 12047 16451 12053
rect 16482 12044 16488 12056
rect 16540 12084 16546 12096
rect 16758 12084 16764 12096
rect 16540 12056 16764 12084
rect 16540 12044 16546 12056
rect 16758 12044 16764 12056
rect 16816 12044 16822 12096
rect 23569 12087 23627 12093
rect 23569 12053 23581 12087
rect 23615 12084 23627 12087
rect 23676 12084 23704 12183
rect 24026 12084 24032 12096
rect 23615 12056 24032 12084
rect 23615 12053 23627 12056
rect 23569 12047 23627 12053
rect 24026 12044 24032 12056
rect 24084 12044 24090 12096
rect 25038 12084 25044 12096
rect 24999 12056 25044 12084
rect 25038 12044 25044 12056
rect 25096 12044 25102 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2222 11840 2228 11892
rect 2280 11880 2286 11892
rect 2409 11883 2467 11889
rect 2409 11880 2421 11883
rect 2280 11852 2421 11880
rect 2280 11840 2286 11852
rect 2409 11849 2421 11852
rect 2455 11849 2467 11883
rect 2409 11843 2467 11849
rect 2590 11840 2596 11892
rect 2648 11880 2654 11892
rect 2648 11852 3096 11880
rect 2648 11840 2654 11852
rect 1765 11747 1823 11753
rect 1765 11713 1777 11747
rect 1811 11744 1823 11747
rect 2133 11747 2191 11753
rect 2133 11744 2145 11747
rect 1811 11716 2145 11744
rect 1811 11713 1823 11716
rect 1765 11707 1823 11713
rect 2133 11713 2145 11716
rect 2179 11744 2191 11747
rect 2590 11744 2596 11756
rect 2179 11716 2596 11744
rect 2179 11713 2191 11716
rect 2133 11707 2191 11713
rect 2590 11704 2596 11716
rect 2648 11704 2654 11756
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11744 2927 11747
rect 2958 11744 2964 11756
rect 2915 11716 2964 11744
rect 2915 11713 2927 11716
rect 2869 11707 2927 11713
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 3068 11753 3096 11852
rect 3510 11840 3516 11892
rect 3568 11880 3574 11892
rect 3973 11883 4031 11889
rect 3973 11880 3985 11883
rect 3568 11852 3985 11880
rect 3568 11840 3574 11852
rect 3973 11849 3985 11852
rect 4019 11849 4031 11883
rect 7190 11880 7196 11892
rect 7151 11852 7196 11880
rect 3973 11843 4031 11849
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 7374 11840 7380 11892
rect 7432 11880 7438 11892
rect 7469 11883 7527 11889
rect 7469 11880 7481 11883
rect 7432 11852 7481 11880
rect 7432 11840 7438 11852
rect 7469 11849 7481 11852
rect 7515 11849 7527 11883
rect 7834 11880 7840 11892
rect 7795 11852 7840 11880
rect 7469 11843 7527 11849
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 10781 11883 10839 11889
rect 10781 11849 10793 11883
rect 10827 11880 10839 11883
rect 10962 11880 10968 11892
rect 10827 11852 10968 11880
rect 10827 11849 10839 11852
rect 10781 11843 10839 11849
rect 10962 11840 10968 11852
rect 11020 11840 11026 11892
rect 11054 11840 11060 11892
rect 11112 11880 11118 11892
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 11112 11852 11805 11880
rect 11112 11840 11118 11852
rect 11793 11849 11805 11852
rect 11839 11880 11851 11883
rect 11977 11883 12035 11889
rect 11977 11880 11989 11883
rect 11839 11852 11989 11880
rect 11839 11849 11851 11852
rect 11793 11843 11851 11849
rect 11977 11849 11989 11852
rect 12023 11849 12035 11883
rect 11977 11843 12035 11849
rect 12434 11840 12440 11892
rect 12492 11880 12498 11892
rect 12492 11852 12537 11880
rect 12492 11840 12498 11852
rect 12894 11840 12900 11892
rect 12952 11880 12958 11892
rect 14001 11883 14059 11889
rect 14001 11880 14013 11883
rect 12952 11852 14013 11880
rect 12952 11840 12958 11852
rect 14001 11849 14013 11852
rect 14047 11880 14059 11883
rect 14090 11880 14096 11892
rect 14047 11852 14096 11880
rect 14047 11849 14059 11852
rect 14001 11843 14059 11849
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 15930 11880 15936 11892
rect 15891 11852 15936 11880
rect 15930 11840 15936 11852
rect 15988 11840 15994 11892
rect 17402 11880 17408 11892
rect 17363 11852 17408 11880
rect 17402 11840 17408 11852
rect 17460 11840 17466 11892
rect 17678 11880 17684 11892
rect 17639 11852 17684 11880
rect 17678 11840 17684 11852
rect 17736 11840 17742 11892
rect 18782 11880 18788 11892
rect 18743 11852 18788 11880
rect 18782 11840 18788 11852
rect 18840 11840 18846 11892
rect 19242 11840 19248 11892
rect 19300 11880 19306 11892
rect 19429 11883 19487 11889
rect 19429 11880 19441 11883
rect 19300 11852 19441 11880
rect 19300 11840 19306 11852
rect 19429 11849 19441 11852
rect 19475 11849 19487 11883
rect 19429 11843 19487 11849
rect 21450 11840 21456 11892
rect 21508 11880 21514 11892
rect 21913 11883 21971 11889
rect 21913 11880 21925 11883
rect 21508 11852 21925 11880
rect 21508 11840 21514 11852
rect 21913 11849 21925 11852
rect 21959 11849 21971 11883
rect 21913 11843 21971 11849
rect 22373 11883 22431 11889
rect 22373 11849 22385 11883
rect 22419 11880 22431 11883
rect 22554 11880 22560 11892
rect 22419 11852 22560 11880
rect 22419 11849 22431 11852
rect 22373 11843 22431 11849
rect 22554 11840 22560 11852
rect 22612 11840 22618 11892
rect 22649 11883 22707 11889
rect 22649 11849 22661 11883
rect 22695 11880 22707 11883
rect 23382 11880 23388 11892
rect 22695 11852 23388 11880
rect 22695 11849 22707 11852
rect 22649 11843 22707 11849
rect 23382 11840 23388 11852
rect 23440 11840 23446 11892
rect 23842 11840 23848 11892
rect 23900 11880 23906 11892
rect 23937 11883 23995 11889
rect 23937 11880 23949 11883
rect 23900 11852 23949 11880
rect 23900 11840 23906 11852
rect 23937 11849 23949 11852
rect 23983 11849 23995 11883
rect 23937 11843 23995 11849
rect 24026 11840 24032 11892
rect 24084 11880 24090 11892
rect 24949 11883 25007 11889
rect 24949 11880 24961 11883
rect 24084 11852 24961 11880
rect 24084 11840 24090 11852
rect 24949 11849 24961 11852
rect 24995 11849 25007 11883
rect 25682 11880 25688 11892
rect 25643 11852 25688 11880
rect 24949 11843 25007 11849
rect 25682 11840 25688 11852
rect 25740 11840 25746 11892
rect 16758 11772 16764 11824
rect 16816 11812 16822 11824
rect 18325 11815 18383 11821
rect 18325 11812 18337 11815
rect 16816 11784 18337 11812
rect 16816 11772 16822 11784
rect 18325 11781 18337 11784
rect 18371 11812 18383 11815
rect 20162 11812 20168 11824
rect 18371 11784 20168 11812
rect 18371 11781 18383 11784
rect 18325 11775 18383 11781
rect 20162 11772 20168 11784
rect 20220 11772 20226 11824
rect 3053 11747 3111 11753
rect 3053 11713 3065 11747
rect 3099 11713 3111 11747
rect 3053 11707 3111 11713
rect 3881 11747 3939 11753
rect 3881 11713 3893 11747
rect 3927 11744 3939 11747
rect 4338 11744 4344 11756
rect 3927 11716 4344 11744
rect 3927 11713 3939 11716
rect 3881 11707 3939 11713
rect 4338 11704 4344 11716
rect 4396 11744 4402 11756
rect 4433 11747 4491 11753
rect 4433 11744 4445 11747
rect 4396 11716 4445 11744
rect 4396 11704 4402 11716
rect 4433 11713 4445 11716
rect 4479 11713 4491 11747
rect 4433 11707 4491 11713
rect 4522 11704 4528 11756
rect 4580 11744 4586 11756
rect 5537 11747 5595 11753
rect 4580 11716 4625 11744
rect 4580 11704 4586 11716
rect 5537 11713 5549 11747
rect 5583 11744 5595 11747
rect 6178 11744 6184 11756
rect 5583 11716 6184 11744
rect 5583 11713 5595 11716
rect 5537 11707 5595 11713
rect 6178 11704 6184 11716
rect 6236 11704 6242 11756
rect 8573 11747 8631 11753
rect 8573 11713 8585 11747
rect 8619 11744 8631 11747
rect 8938 11744 8944 11756
rect 8619 11716 8944 11744
rect 8619 11713 8631 11716
rect 8573 11707 8631 11713
rect 8938 11704 8944 11716
rect 8996 11704 9002 11756
rect 10686 11704 10692 11756
rect 10744 11744 10750 11756
rect 11241 11747 11299 11753
rect 11241 11744 11253 11747
rect 10744 11716 11253 11744
rect 10744 11704 10750 11716
rect 11241 11713 11253 11716
rect 11287 11713 11299 11747
rect 11241 11707 11299 11713
rect 11425 11747 11483 11753
rect 11425 11713 11437 11747
rect 11471 11744 11483 11747
rect 11698 11744 11704 11756
rect 11471 11716 11704 11744
rect 11471 11713 11483 11716
rect 11425 11707 11483 11713
rect 11698 11704 11704 11716
rect 11756 11704 11762 11756
rect 12986 11744 12992 11756
rect 12899 11716 12992 11744
rect 12986 11704 12992 11716
rect 13044 11744 13050 11756
rect 14366 11744 14372 11756
rect 13044 11716 14372 11744
rect 13044 11704 13050 11716
rect 14366 11704 14372 11716
rect 14424 11704 14430 11756
rect 15562 11744 15568 11756
rect 15475 11716 15568 11744
rect 15562 11704 15568 11716
rect 15620 11744 15626 11756
rect 15930 11744 15936 11756
rect 15620 11716 15936 11744
rect 15620 11704 15626 11716
rect 15930 11704 15936 11716
rect 15988 11704 15994 11756
rect 16298 11704 16304 11756
rect 16356 11744 16362 11756
rect 16485 11747 16543 11753
rect 16485 11744 16497 11747
rect 16356 11716 16497 11744
rect 16356 11704 16362 11716
rect 16485 11713 16497 11716
rect 16531 11713 16543 11747
rect 16485 11707 16543 11713
rect 19613 11747 19671 11753
rect 19613 11713 19625 11747
rect 19659 11744 19671 11747
rect 20438 11744 20444 11756
rect 19659 11716 20444 11744
rect 19659 11713 19671 11716
rect 19613 11707 19671 11713
rect 20438 11704 20444 11716
rect 20496 11704 20502 11756
rect 21453 11747 21511 11753
rect 21453 11713 21465 11747
rect 21499 11744 21511 11747
rect 21910 11744 21916 11756
rect 21499 11716 21916 11744
rect 21499 11713 21511 11716
rect 21453 11707 21511 11713
rect 21910 11704 21916 11716
rect 21968 11704 21974 11756
rect 23014 11744 23020 11756
rect 22975 11716 23020 11744
rect 23014 11704 23020 11716
rect 23072 11744 23078 11756
rect 23934 11744 23940 11756
rect 23072 11716 23940 11744
rect 23072 11704 23078 11716
rect 23934 11704 23940 11716
rect 23992 11744 23998 11756
rect 24489 11747 24547 11753
rect 24489 11744 24501 11747
rect 23992 11716 24501 11744
rect 23992 11704 23998 11716
rect 24489 11713 24501 11716
rect 24535 11713 24547 11747
rect 24489 11707 24547 11713
rect 10597 11679 10655 11685
rect 10597 11645 10609 11679
rect 10643 11676 10655 11679
rect 11330 11676 11336 11688
rect 10643 11648 11336 11676
rect 10643 11645 10655 11648
rect 10597 11639 10655 11645
rect 11330 11636 11336 11648
rect 11388 11636 11394 11688
rect 11977 11679 12035 11685
rect 11977 11645 11989 11679
rect 12023 11676 12035 11679
rect 12897 11679 12955 11685
rect 12023 11648 12204 11676
rect 12023 11645 12035 11648
rect 11977 11639 12035 11645
rect 2774 11568 2780 11620
rect 2832 11608 2838 11620
rect 4062 11608 4068 11620
rect 2832 11580 4068 11608
rect 2832 11568 2838 11580
rect 4062 11568 4068 11580
rect 4120 11568 4126 11620
rect 10321 11611 10379 11617
rect 10321 11577 10333 11611
rect 10367 11608 10379 11611
rect 11149 11611 11207 11617
rect 11149 11608 11161 11611
rect 10367 11580 11161 11608
rect 10367 11577 10379 11580
rect 10321 11571 10379 11577
rect 11149 11577 11161 11580
rect 11195 11608 11207 11611
rect 12066 11608 12072 11620
rect 11195 11580 12072 11608
rect 11195 11577 11207 11580
rect 11149 11571 11207 11577
rect 12066 11568 12072 11580
rect 12124 11568 12130 11620
rect 12176 11608 12204 11648
rect 12897 11645 12909 11679
rect 12943 11676 12955 11679
rect 13078 11676 13084 11688
rect 12943 11648 13084 11676
rect 12943 11645 12955 11648
rect 12897 11639 12955 11645
rect 12805 11611 12863 11617
rect 12805 11608 12817 11611
rect 12176 11580 12817 11608
rect 12805 11577 12817 11580
rect 12851 11577 12863 11611
rect 12805 11571 12863 11577
rect 3510 11540 3516 11552
rect 3471 11512 3516 11540
rect 3510 11500 3516 11512
rect 3568 11540 3574 11552
rect 4246 11540 4252 11552
rect 3568 11512 4252 11540
rect 3568 11500 3574 11512
rect 4246 11500 4252 11512
rect 4304 11540 4310 11552
rect 4341 11543 4399 11549
rect 4341 11540 4353 11543
rect 4304 11512 4353 11540
rect 4304 11500 4310 11512
rect 4341 11509 4353 11512
rect 4387 11540 4399 11543
rect 5077 11543 5135 11549
rect 5077 11540 5089 11543
rect 4387 11512 5089 11540
rect 4387 11509 4399 11512
rect 4341 11503 4399 11509
rect 5077 11509 5089 11512
rect 5123 11509 5135 11543
rect 5077 11503 5135 11509
rect 11054 11500 11060 11552
rect 11112 11540 11118 11552
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 11112 11512 12173 11540
rect 11112 11500 11118 11512
rect 12161 11509 12173 11512
rect 12207 11540 12219 11543
rect 12912 11540 12940 11639
rect 13078 11636 13084 11648
rect 13136 11636 13142 11688
rect 13633 11679 13691 11685
rect 13633 11645 13645 11679
rect 13679 11676 13691 11679
rect 13814 11676 13820 11688
rect 13679 11648 13820 11676
rect 13679 11645 13691 11648
rect 13633 11639 13691 11645
rect 13814 11636 13820 11648
rect 13872 11676 13878 11688
rect 14829 11679 14887 11685
rect 14829 11676 14841 11679
rect 13872 11648 14841 11676
rect 13872 11636 13878 11648
rect 14829 11645 14841 11648
rect 14875 11676 14887 11679
rect 15102 11676 15108 11688
rect 14875 11648 15108 11676
rect 14875 11645 14887 11648
rect 14829 11639 14887 11645
rect 15102 11636 15108 11648
rect 15160 11636 15166 11688
rect 15378 11636 15384 11688
rect 15436 11676 15442 11688
rect 15746 11676 15752 11688
rect 15436 11648 15752 11676
rect 15436 11636 15442 11648
rect 15746 11636 15752 11648
rect 15804 11676 15810 11688
rect 16393 11679 16451 11685
rect 16393 11676 16405 11679
rect 15804 11648 16405 11676
rect 15804 11636 15810 11648
rect 16393 11645 16405 11648
rect 16439 11645 16451 11679
rect 22462 11676 22468 11688
rect 22423 11648 22468 11676
rect 16393 11639 16451 11645
rect 22462 11636 22468 11648
rect 22520 11636 22526 11688
rect 23477 11679 23535 11685
rect 23477 11645 23489 11679
rect 23523 11676 23535 11679
rect 24305 11679 24363 11685
rect 24305 11676 24317 11679
rect 23523 11648 24317 11676
rect 23523 11645 23535 11648
rect 23477 11639 23535 11645
rect 24305 11645 24317 11648
rect 24351 11676 24363 11679
rect 24762 11676 24768 11688
rect 24351 11648 24768 11676
rect 24351 11645 24363 11648
rect 24305 11639 24363 11645
rect 24762 11636 24768 11648
rect 24820 11636 24826 11688
rect 25498 11676 25504 11688
rect 25459 11648 25504 11676
rect 25498 11636 25504 11648
rect 25556 11676 25562 11688
rect 26053 11679 26111 11685
rect 26053 11676 26065 11679
rect 25556 11648 26065 11676
rect 25556 11636 25562 11648
rect 26053 11645 26065 11648
rect 26099 11645 26111 11679
rect 26053 11639 26111 11645
rect 15010 11568 15016 11620
rect 15068 11608 15074 11620
rect 15289 11611 15347 11617
rect 15289 11608 15301 11611
rect 15068 11580 15301 11608
rect 15068 11568 15074 11580
rect 15289 11577 15301 11580
rect 15335 11608 15347 11611
rect 16482 11608 16488 11620
rect 15335 11580 16488 11608
rect 15335 11577 15347 11580
rect 15289 11571 15347 11577
rect 16482 11568 16488 11580
rect 16540 11568 16546 11620
rect 24118 11568 24124 11620
rect 24176 11608 24182 11620
rect 24397 11611 24455 11617
rect 24397 11608 24409 11611
rect 24176 11580 24409 11608
rect 24176 11568 24182 11580
rect 24397 11577 24409 11580
rect 24443 11577 24455 11611
rect 24397 11571 24455 11577
rect 14918 11540 14924 11552
rect 12207 11512 12940 11540
rect 14879 11512 14924 11540
rect 12207 11509 12219 11512
rect 12161 11503 12219 11509
rect 14918 11500 14924 11512
rect 14976 11500 14982 11552
rect 15102 11500 15108 11552
rect 15160 11540 15166 11552
rect 15381 11543 15439 11549
rect 15381 11540 15393 11543
rect 15160 11512 15393 11540
rect 15160 11500 15166 11512
rect 15381 11509 15393 11512
rect 15427 11540 15439 11543
rect 15562 11540 15568 11552
rect 15427 11512 15568 11540
rect 15427 11509 15439 11512
rect 15381 11503 15439 11509
rect 15562 11500 15568 11512
rect 15620 11500 15626 11552
rect 17034 11540 17040 11552
rect 16995 11512 17040 11540
rect 17034 11500 17040 11512
rect 17092 11500 17098 11552
rect 19150 11540 19156 11552
rect 19111 11512 19156 11540
rect 19150 11500 19156 11512
rect 19208 11500 19214 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1854 11336 1860 11348
rect 1815 11308 1860 11336
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 2041 11339 2099 11345
rect 2041 11305 2053 11339
rect 2087 11336 2099 11339
rect 2406 11336 2412 11348
rect 2087 11308 2412 11336
rect 2087 11305 2099 11308
rect 2041 11299 2099 11305
rect 2406 11296 2412 11308
rect 2464 11336 2470 11348
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 2464 11308 3801 11336
rect 2464 11296 2470 11308
rect 3789 11305 3801 11308
rect 3835 11305 3847 11339
rect 4062 11336 4068 11348
rect 4023 11308 4068 11336
rect 3789 11299 3847 11305
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 4154 11296 4160 11348
rect 4212 11336 4218 11348
rect 4433 11339 4491 11345
rect 4433 11336 4445 11339
rect 4212 11308 4445 11336
rect 4212 11296 4218 11308
rect 4433 11305 4445 11308
rect 4479 11336 4491 11339
rect 4798 11336 4804 11348
rect 4479 11308 4804 11336
rect 4479 11305 4491 11308
rect 4433 11299 4491 11305
rect 4798 11296 4804 11308
rect 4856 11296 4862 11348
rect 5534 11336 5540 11348
rect 5495 11308 5540 11336
rect 5534 11296 5540 11308
rect 5592 11296 5598 11348
rect 10873 11339 10931 11345
rect 10873 11305 10885 11339
rect 10919 11336 10931 11339
rect 11698 11336 11704 11348
rect 10919 11308 11704 11336
rect 10919 11305 10931 11308
rect 10873 11299 10931 11305
rect 11698 11296 11704 11308
rect 11756 11296 11762 11348
rect 12066 11336 12072 11348
rect 12027 11308 12072 11336
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 12437 11339 12495 11345
rect 12437 11305 12449 11339
rect 12483 11336 12495 11339
rect 12526 11336 12532 11348
rect 12483 11308 12532 11336
rect 12483 11305 12495 11308
rect 12437 11299 12495 11305
rect 12526 11296 12532 11308
rect 12584 11296 12590 11348
rect 12894 11296 12900 11348
rect 12952 11336 12958 11348
rect 13081 11339 13139 11345
rect 13081 11336 13093 11339
rect 12952 11308 13093 11336
rect 12952 11296 12958 11308
rect 13081 11305 13093 11308
rect 13127 11305 13139 11339
rect 13081 11299 13139 11305
rect 13998 11296 14004 11348
rect 14056 11336 14062 11348
rect 14093 11339 14151 11345
rect 14093 11336 14105 11339
rect 14056 11308 14105 11336
rect 14056 11296 14062 11308
rect 14093 11305 14105 11308
rect 14139 11305 14151 11339
rect 15010 11336 15016 11348
rect 14971 11308 15016 11336
rect 14093 11299 14151 11305
rect 15010 11296 15016 11308
rect 15068 11296 15074 11348
rect 15286 11336 15292 11348
rect 15247 11308 15292 11336
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 16390 11336 16396 11348
rect 16351 11308 16396 11336
rect 16390 11296 16396 11308
rect 16448 11296 16454 11348
rect 22370 11336 22376 11348
rect 22331 11308 22376 11336
rect 22370 11296 22376 11308
rect 22428 11296 22434 11348
rect 22462 11296 22468 11348
rect 22520 11336 22526 11348
rect 22925 11339 22983 11345
rect 22925 11336 22937 11339
rect 22520 11308 22937 11336
rect 22520 11296 22526 11308
rect 22925 11305 22937 11308
rect 22971 11336 22983 11339
rect 23382 11336 23388 11348
rect 22971 11308 23388 11336
rect 22971 11305 22983 11308
rect 22925 11299 22983 11305
rect 23382 11296 23388 11308
rect 23440 11296 23446 11348
rect 23658 11336 23664 11348
rect 23619 11308 23664 11336
rect 23658 11296 23664 11308
rect 23716 11296 23722 11348
rect 24765 11339 24823 11345
rect 24765 11305 24777 11339
rect 24811 11336 24823 11339
rect 25314 11336 25320 11348
rect 24811 11308 25320 11336
rect 24811 11305 24823 11308
rect 24765 11299 24823 11305
rect 25314 11296 25320 11308
rect 25372 11296 25378 11348
rect 2498 11228 2504 11280
rect 2556 11268 2562 11280
rect 3421 11271 3479 11277
rect 3421 11268 3433 11271
rect 2556 11240 3433 11268
rect 2556 11228 2562 11240
rect 3421 11237 3433 11240
rect 3467 11237 3479 11271
rect 3421 11231 3479 11237
rect 13541 11271 13599 11277
rect 13541 11237 13553 11271
rect 13587 11268 13599 11271
rect 13906 11268 13912 11280
rect 13587 11240 13912 11268
rect 13587 11237 13599 11240
rect 13541 11231 13599 11237
rect 13906 11228 13912 11240
rect 13964 11268 13970 11280
rect 14918 11268 14924 11280
rect 13964 11240 14924 11268
rect 13964 11228 13970 11240
rect 14918 11228 14924 11240
rect 14976 11228 14982 11280
rect 23934 11228 23940 11280
rect 23992 11268 23998 11280
rect 24121 11271 24179 11277
rect 24121 11268 24133 11271
rect 23992 11240 24133 11268
rect 23992 11228 23998 11240
rect 24121 11237 24133 11240
rect 24167 11237 24179 11271
rect 24121 11231 24179 11237
rect 1394 11160 1400 11212
rect 1452 11200 1458 11212
rect 2038 11200 2044 11212
rect 1452 11172 2044 11200
rect 1452 11160 1458 11172
rect 2038 11160 2044 11172
rect 2096 11200 2102 11212
rect 2409 11203 2467 11209
rect 2409 11200 2421 11203
rect 2096 11172 2421 11200
rect 2096 11160 2102 11172
rect 2409 11169 2421 11172
rect 2455 11169 2467 11203
rect 2409 11163 2467 11169
rect 2958 11160 2964 11212
rect 3016 11200 3022 11212
rect 3053 11203 3111 11209
rect 3053 11200 3065 11203
rect 3016 11172 3065 11200
rect 3016 11160 3022 11172
rect 3053 11169 3065 11172
rect 3099 11169 3111 11203
rect 3053 11163 3111 11169
rect 12529 11203 12587 11209
rect 12529 11169 12541 11203
rect 12575 11200 12587 11203
rect 12618 11200 12624 11212
rect 12575 11172 12624 11200
rect 12575 11169 12587 11172
rect 12529 11163 12587 11169
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 14001 11203 14059 11209
rect 14001 11169 14013 11203
rect 14047 11200 14059 11203
rect 14090 11200 14096 11212
rect 14047 11172 14096 11200
rect 14047 11169 14059 11172
rect 14001 11163 14059 11169
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 15562 11160 15568 11212
rect 15620 11200 15626 11212
rect 15657 11203 15715 11209
rect 15657 11200 15669 11203
rect 15620 11172 15669 11200
rect 15620 11160 15626 11172
rect 15657 11169 15669 11172
rect 15703 11169 15715 11203
rect 15657 11163 15715 11169
rect 15749 11203 15807 11209
rect 15749 11169 15761 11203
rect 15795 11200 15807 11203
rect 16022 11200 16028 11212
rect 15795 11172 16028 11200
rect 15795 11169 15807 11172
rect 15749 11163 15807 11169
rect 16022 11160 16028 11172
rect 16080 11160 16086 11212
rect 23477 11203 23535 11209
rect 23477 11169 23489 11203
rect 23523 11200 23535 11203
rect 24026 11200 24032 11212
rect 23523 11172 24032 11200
rect 23523 11169 23535 11172
rect 23477 11163 23535 11169
rect 24026 11160 24032 11172
rect 24084 11160 24090 11212
rect 24578 11200 24584 11212
rect 24539 11172 24584 11200
rect 24578 11160 24584 11172
rect 24636 11200 24642 11212
rect 24762 11200 24768 11212
rect 24636 11172 24768 11200
rect 24636 11160 24642 11172
rect 24762 11160 24768 11172
rect 24820 11160 24826 11212
rect 1946 11092 1952 11144
rect 2004 11132 2010 11144
rect 2314 11132 2320 11144
rect 2004 11104 2320 11132
rect 2004 11092 2010 11104
rect 2314 11092 2320 11104
rect 2372 11132 2378 11144
rect 2501 11135 2559 11141
rect 2501 11132 2513 11135
rect 2372 11104 2513 11132
rect 2372 11092 2378 11104
rect 2501 11101 2513 11104
rect 2547 11101 2559 11135
rect 2501 11095 2559 11101
rect 2593 11135 2651 11141
rect 2593 11101 2605 11135
rect 2639 11101 2651 11135
rect 4522 11132 4528 11144
rect 4483 11104 4528 11132
rect 2593 11095 2651 11101
rect 1854 11024 1860 11076
rect 1912 11064 1918 11076
rect 2608 11064 2636 11095
rect 4522 11092 4528 11104
rect 4580 11092 4586 11144
rect 4706 11132 4712 11144
rect 4667 11104 4712 11132
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 12158 11092 12164 11144
rect 12216 11132 12222 11144
rect 12713 11135 12771 11141
rect 12713 11132 12725 11135
rect 12216 11104 12725 11132
rect 12216 11092 12222 11104
rect 12713 11101 12725 11104
rect 12759 11132 12771 11135
rect 12986 11132 12992 11144
rect 12759 11104 12992 11132
rect 12759 11101 12771 11104
rect 12713 11095 12771 11101
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 14182 11132 14188 11144
rect 14143 11104 14188 11132
rect 14182 11092 14188 11104
rect 14240 11092 14246 11144
rect 15930 11132 15936 11144
rect 15891 11104 15936 11132
rect 15930 11092 15936 11104
rect 15988 11092 15994 11144
rect 16574 11092 16580 11144
rect 16632 11132 16638 11144
rect 16853 11135 16911 11141
rect 16853 11132 16865 11135
rect 16632 11104 16865 11132
rect 16632 11092 16638 11104
rect 16853 11101 16865 11104
rect 16899 11101 16911 11135
rect 16853 11095 16911 11101
rect 1912 11036 2728 11064
rect 1912 11024 1918 11036
rect 2700 10996 2728 11036
rect 3602 11024 3608 11076
rect 3660 11064 3666 11076
rect 5074 11064 5080 11076
rect 3660 11036 5080 11064
rect 3660 11024 3666 11036
rect 5074 11024 5080 11036
rect 5132 11024 5138 11076
rect 11146 11024 11152 11076
rect 11204 11064 11210 11076
rect 11241 11067 11299 11073
rect 11241 11064 11253 11067
rect 11204 11036 11253 11064
rect 11204 11024 11210 11036
rect 11241 11033 11253 11036
rect 11287 11064 11299 11067
rect 11974 11064 11980 11076
rect 11287 11036 11980 11064
rect 11287 11033 11299 11036
rect 11241 11027 11299 11033
rect 11974 11024 11980 11036
rect 12032 11024 12038 11076
rect 13633 11067 13691 11073
rect 13633 11033 13645 11067
rect 13679 11064 13691 11067
rect 13679 11036 13768 11064
rect 13679 11033 13691 11036
rect 13633 11027 13691 11033
rect 3050 10996 3056 11008
rect 2700 10968 3056 10996
rect 3050 10956 3056 10968
rect 3108 10956 3114 11008
rect 13740 10996 13768 11036
rect 24118 11024 24124 11076
rect 24176 11064 24182 11076
rect 24397 11067 24455 11073
rect 24397 11064 24409 11067
rect 24176 11036 24409 11064
rect 24176 11024 24182 11036
rect 24397 11033 24409 11036
rect 24443 11033 24455 11067
rect 24397 11027 24455 11033
rect 14642 10996 14648 11008
rect 13740 10968 14648 10996
rect 14642 10956 14648 10968
rect 14700 10956 14706 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 2409 10795 2467 10801
rect 2409 10761 2421 10795
rect 2455 10792 2467 10795
rect 2498 10792 2504 10804
rect 2455 10764 2504 10792
rect 2455 10761 2467 10764
rect 2409 10755 2467 10761
rect 2498 10752 2504 10764
rect 2556 10752 2562 10804
rect 4154 10792 4160 10804
rect 4115 10764 4160 10792
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 4522 10792 4528 10804
rect 4483 10764 4528 10792
rect 4522 10752 4528 10764
rect 4580 10752 4586 10804
rect 4706 10752 4712 10804
rect 4764 10792 4770 10804
rect 4801 10795 4859 10801
rect 4801 10792 4813 10795
rect 4764 10764 4813 10792
rect 4764 10752 4770 10764
rect 4801 10761 4813 10764
rect 4847 10761 4859 10795
rect 4801 10755 4859 10761
rect 12161 10795 12219 10801
rect 12161 10761 12173 10795
rect 12207 10792 12219 10795
rect 12342 10792 12348 10804
rect 12207 10764 12348 10792
rect 12207 10761 12219 10764
rect 12161 10755 12219 10761
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 13998 10792 14004 10804
rect 13959 10764 14004 10792
rect 13998 10752 14004 10764
rect 14056 10752 14062 10804
rect 14090 10752 14096 10804
rect 14148 10792 14154 10804
rect 14277 10795 14335 10801
rect 14277 10792 14289 10795
rect 14148 10764 14289 10792
rect 14148 10752 14154 10764
rect 14277 10761 14289 10764
rect 14323 10761 14335 10795
rect 14277 10755 14335 10761
rect 14553 10795 14611 10801
rect 14553 10761 14565 10795
rect 14599 10792 14611 10795
rect 15378 10792 15384 10804
rect 14599 10764 15384 10792
rect 14599 10761 14611 10764
rect 14553 10755 14611 10761
rect 15378 10752 15384 10764
rect 15436 10752 15442 10804
rect 23937 10795 23995 10801
rect 23937 10761 23949 10795
rect 23983 10792 23995 10795
rect 24026 10792 24032 10804
rect 23983 10764 24032 10792
rect 23983 10761 23995 10764
rect 23937 10755 23995 10761
rect 24026 10752 24032 10764
rect 24084 10752 24090 10804
rect 24489 10795 24547 10801
rect 24489 10761 24501 10795
rect 24535 10792 24547 10795
rect 24762 10792 24768 10804
rect 24535 10764 24768 10792
rect 24535 10761 24547 10764
rect 24489 10755 24547 10761
rect 24762 10752 24768 10764
rect 24820 10752 24826 10804
rect 3050 10656 3056 10668
rect 2963 10628 3056 10656
rect 3050 10616 3056 10628
rect 3108 10656 3114 10668
rect 4724 10656 4752 10752
rect 3108 10628 4752 10656
rect 11793 10659 11851 10665
rect 3108 10616 3114 10628
rect 11793 10625 11805 10659
rect 11839 10656 11851 10659
rect 12342 10656 12348 10668
rect 11839 10628 12348 10656
rect 11839 10625 11851 10628
rect 11793 10619 11851 10625
rect 12342 10616 12348 10628
rect 12400 10616 12406 10668
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10656 13231 10659
rect 13262 10656 13268 10668
rect 13219 10628 13268 10656
rect 13219 10625 13231 10628
rect 13173 10619 13231 10625
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 15102 10656 15108 10668
rect 15063 10628 15108 10656
rect 15102 10616 15108 10628
rect 15160 10656 15166 10668
rect 15930 10656 15936 10668
rect 15160 10628 15936 10656
rect 15160 10616 15166 10628
rect 15930 10616 15936 10628
rect 15988 10656 15994 10668
rect 16301 10659 16359 10665
rect 16301 10656 16313 10659
rect 15988 10628 16313 10656
rect 15988 10616 15994 10628
rect 16301 10625 16313 10628
rect 16347 10625 16359 10659
rect 16301 10619 16359 10625
rect 12894 10588 12900 10600
rect 12855 10560 12900 10588
rect 12894 10548 12900 10560
rect 12952 10548 12958 10600
rect 14826 10548 14832 10600
rect 14884 10588 14890 10600
rect 14921 10591 14979 10597
rect 14921 10588 14933 10591
rect 14884 10560 14933 10588
rect 14884 10548 14890 10560
rect 14921 10557 14933 10560
rect 14967 10557 14979 10591
rect 24578 10588 24584 10600
rect 24539 10560 24584 10588
rect 14921 10551 14979 10557
rect 24578 10548 24584 10560
rect 24636 10588 24642 10600
rect 25133 10591 25191 10597
rect 25133 10588 25145 10591
rect 24636 10560 25145 10588
rect 24636 10548 24642 10560
rect 25133 10557 25145 10560
rect 25179 10557 25191 10591
rect 25133 10551 25191 10557
rect 1765 10523 1823 10529
rect 1765 10489 1777 10523
rect 1811 10520 1823 10523
rect 2682 10520 2688 10532
rect 1811 10492 2688 10520
rect 1811 10489 1823 10492
rect 1765 10483 1823 10489
rect 2682 10480 2688 10492
rect 2740 10520 2746 10532
rect 2869 10523 2927 10529
rect 2869 10520 2881 10523
rect 2740 10492 2881 10520
rect 2740 10480 2746 10492
rect 2869 10489 2881 10492
rect 2915 10520 2927 10523
rect 2958 10520 2964 10532
rect 2915 10492 2964 10520
rect 2915 10489 2927 10492
rect 2869 10483 2927 10489
rect 2958 10480 2964 10492
rect 3016 10480 3022 10532
rect 14642 10480 14648 10532
rect 14700 10520 14706 10532
rect 15013 10523 15071 10529
rect 15013 10520 15025 10523
rect 14700 10492 15025 10520
rect 14700 10480 14706 10492
rect 15013 10489 15025 10492
rect 15059 10520 15071 10523
rect 16669 10523 16727 10529
rect 16669 10520 16681 10523
rect 15059 10492 16681 10520
rect 15059 10489 15071 10492
rect 15013 10483 15071 10489
rect 16669 10489 16681 10492
rect 16715 10489 16727 10523
rect 16669 10483 16727 10489
rect 1946 10412 1952 10464
rect 2004 10452 2010 10464
rect 2041 10455 2099 10461
rect 2041 10452 2053 10455
rect 2004 10424 2053 10452
rect 2004 10412 2010 10424
rect 2041 10421 2053 10424
rect 2087 10421 2099 10455
rect 2041 10415 2099 10421
rect 2777 10455 2835 10461
rect 2777 10421 2789 10455
rect 2823 10452 2835 10455
rect 3326 10452 3332 10464
rect 2823 10424 3332 10452
rect 2823 10421 2835 10424
rect 2777 10415 2835 10421
rect 3326 10412 3332 10424
rect 3384 10452 3390 10464
rect 3421 10455 3479 10461
rect 3421 10452 3433 10455
rect 3384 10424 3433 10452
rect 3384 10412 3390 10424
rect 3421 10421 3433 10424
rect 3467 10452 3479 10455
rect 3786 10452 3792 10464
rect 3467 10424 3792 10452
rect 3467 10421 3479 10424
rect 3421 10415 3479 10421
rect 3786 10412 3792 10424
rect 3844 10412 3850 10464
rect 12526 10452 12532 10464
rect 12487 10424 12532 10452
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 12989 10455 13047 10461
rect 12989 10421 13001 10455
rect 13035 10452 13047 10455
rect 13538 10452 13544 10464
rect 13035 10424 13544 10452
rect 13035 10421 13047 10424
rect 12989 10415 13047 10421
rect 13538 10412 13544 10424
rect 13596 10412 13602 10464
rect 15562 10452 15568 10464
rect 15523 10424 15568 10452
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 16022 10452 16028 10464
rect 15983 10424 16028 10452
rect 16022 10412 16028 10424
rect 16080 10412 16086 10464
rect 24765 10455 24823 10461
rect 24765 10421 24777 10455
rect 24811 10452 24823 10455
rect 25774 10452 25780 10464
rect 24811 10424 25780 10452
rect 24811 10421 24823 10424
rect 24765 10415 24823 10421
rect 25774 10412 25780 10424
rect 25832 10412 25838 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 2038 10248 2044 10260
rect 1999 10220 2044 10248
rect 2038 10208 2044 10220
rect 2096 10208 2102 10260
rect 3050 10248 3056 10260
rect 3011 10220 3056 10248
rect 3050 10208 3056 10220
rect 3108 10208 3114 10260
rect 12250 10248 12256 10260
rect 12211 10220 12256 10248
rect 12250 10208 12256 10220
rect 12308 10208 12314 10260
rect 12526 10208 12532 10260
rect 12584 10248 12590 10260
rect 12621 10251 12679 10257
rect 12621 10248 12633 10251
rect 12584 10220 12633 10248
rect 12584 10208 12590 10220
rect 12621 10217 12633 10220
rect 12667 10217 12679 10251
rect 12621 10211 12679 10217
rect 12710 10208 12716 10260
rect 12768 10248 12774 10260
rect 13262 10248 13268 10260
rect 12768 10220 12813 10248
rect 13223 10220 13268 10248
rect 12768 10208 12774 10220
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 14645 10251 14703 10257
rect 14645 10217 14657 10251
rect 14691 10248 14703 10251
rect 14826 10248 14832 10260
rect 14691 10220 14832 10248
rect 14691 10217 14703 10220
rect 14645 10211 14703 10217
rect 14826 10208 14832 10220
rect 14884 10208 14890 10260
rect 15013 10251 15071 10257
rect 15013 10217 15025 10251
rect 15059 10248 15071 10251
rect 15102 10248 15108 10260
rect 15059 10220 15108 10248
rect 15059 10217 15071 10220
rect 15013 10211 15071 10217
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 15289 10251 15347 10257
rect 15289 10217 15301 10251
rect 15335 10248 15347 10251
rect 15470 10248 15476 10260
rect 15335 10220 15476 10248
rect 15335 10217 15347 10220
rect 15289 10211 15347 10217
rect 15470 10208 15476 10220
rect 15528 10208 15534 10260
rect 15657 10251 15715 10257
rect 15657 10217 15669 10251
rect 15703 10248 15715 10251
rect 15746 10248 15752 10260
rect 15703 10220 15752 10248
rect 15703 10217 15715 10220
rect 15657 10211 15715 10217
rect 15746 10208 15752 10220
rect 15804 10248 15810 10260
rect 16482 10248 16488 10260
rect 15804 10220 16488 10248
rect 15804 10208 15810 10220
rect 16482 10208 16488 10220
rect 16540 10208 16546 10260
rect 24765 10251 24823 10257
rect 24765 10217 24777 10251
rect 24811 10248 24823 10251
rect 26050 10248 26056 10260
rect 24811 10220 26056 10248
rect 24811 10217 24823 10220
rect 24765 10211 24823 10217
rect 26050 10208 26056 10220
rect 26108 10208 26114 10260
rect 12158 10180 12164 10192
rect 12119 10152 12164 10180
rect 12158 10140 12164 10152
rect 12216 10140 12222 10192
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 1670 10112 1676 10124
rect 1443 10084 1676 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 2501 10115 2559 10121
rect 2501 10081 2513 10115
rect 2547 10112 2559 10115
rect 2682 10112 2688 10124
rect 2547 10084 2688 10112
rect 2547 10081 2559 10084
rect 2501 10075 2559 10081
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 15654 10072 15660 10124
rect 15712 10112 15718 10124
rect 15749 10115 15807 10121
rect 15749 10112 15761 10115
rect 15712 10084 15761 10112
rect 15712 10072 15718 10084
rect 15749 10081 15761 10084
rect 15795 10081 15807 10115
rect 15749 10075 15807 10081
rect 24581 10115 24639 10121
rect 24581 10081 24593 10115
rect 24627 10112 24639 10115
rect 24670 10112 24676 10124
rect 24627 10084 24676 10112
rect 24627 10081 24639 10084
rect 24581 10075 24639 10081
rect 24670 10072 24676 10084
rect 24728 10072 24734 10124
rect 12618 10004 12624 10056
rect 12676 10044 12682 10056
rect 12897 10047 12955 10053
rect 12897 10044 12909 10047
rect 12676 10016 12909 10044
rect 12676 10004 12682 10016
rect 12897 10013 12909 10016
rect 12943 10044 12955 10047
rect 13354 10044 13360 10056
rect 12943 10016 13360 10044
rect 12943 10013 12955 10016
rect 12897 10007 12955 10013
rect 13354 10004 13360 10016
rect 13412 10044 13418 10056
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 13412 10016 14105 10044
rect 13412 10004 13418 10016
rect 14093 10013 14105 10016
rect 14139 10044 14151 10047
rect 14642 10044 14648 10056
rect 14139 10016 14648 10044
rect 14139 10013 14151 10016
rect 14093 10007 14151 10013
rect 14642 10004 14648 10016
rect 14700 10044 14706 10056
rect 15841 10047 15899 10053
rect 15841 10044 15853 10047
rect 14700 10016 15853 10044
rect 14700 10004 14706 10016
rect 15841 10013 15853 10016
rect 15887 10044 15899 10047
rect 15930 10044 15936 10056
rect 15887 10016 15936 10044
rect 15887 10013 15899 10016
rect 15841 10007 15899 10013
rect 15930 10004 15936 10016
rect 15988 10004 15994 10056
rect 2685 9979 2743 9985
rect 2685 9945 2697 9979
rect 2731 9976 2743 9979
rect 6178 9976 6184 9988
rect 2731 9948 6184 9976
rect 2731 9945 2743 9948
rect 2685 9939 2743 9945
rect 6178 9936 6184 9948
rect 6236 9936 6242 9988
rect 13725 9911 13783 9917
rect 13725 9877 13737 9911
rect 13771 9908 13783 9911
rect 14090 9908 14096 9920
rect 13771 9880 14096 9908
rect 13771 9877 13783 9880
rect 13725 9871 13783 9877
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2590 9704 2596 9716
rect 2551 9676 2596 9704
rect 2590 9664 2596 9676
rect 2648 9664 2654 9716
rect 12618 9704 12624 9716
rect 12579 9676 12624 9704
rect 12618 9664 12624 9676
rect 12676 9664 12682 9716
rect 12710 9664 12716 9716
rect 12768 9704 12774 9716
rect 12989 9707 13047 9713
rect 12989 9704 13001 9707
rect 12768 9676 13001 9704
rect 12768 9664 12774 9676
rect 12989 9673 13001 9676
rect 13035 9673 13047 9707
rect 15746 9704 15752 9716
rect 15707 9676 15752 9704
rect 12989 9667 13047 9673
rect 15746 9664 15752 9676
rect 15804 9664 15810 9716
rect 15930 9664 15936 9716
rect 15988 9704 15994 9716
rect 16025 9707 16083 9713
rect 16025 9704 16037 9707
rect 15988 9676 16037 9704
rect 15988 9664 15994 9676
rect 16025 9673 16037 9676
rect 16071 9673 16083 9707
rect 24670 9704 24676 9716
rect 24631 9676 24676 9704
rect 16025 9667 16083 9673
rect 24670 9664 24676 9676
rect 24728 9664 24734 9716
rect 26234 9664 26240 9716
rect 26292 9704 26298 9716
rect 27065 9707 27123 9713
rect 27065 9704 27077 9707
rect 26292 9676 27077 9704
rect 26292 9664 26298 9676
rect 27065 9673 27077 9676
rect 27111 9673 27123 9707
rect 27065 9667 27123 9673
rect 14093 9639 14151 9645
rect 14093 9605 14105 9639
rect 14139 9636 14151 9639
rect 14734 9636 14740 9648
rect 14139 9608 14740 9636
rect 14139 9605 14151 9608
rect 14093 9599 14151 9605
rect 14734 9596 14740 9608
rect 14792 9596 14798 9648
rect 15381 9639 15439 9645
rect 15381 9605 15393 9639
rect 15427 9636 15439 9639
rect 15654 9636 15660 9648
rect 15427 9608 15660 9636
rect 15427 9605 15439 9608
rect 15381 9599 15439 9605
rect 15654 9596 15660 9608
rect 15712 9596 15718 9648
rect 24210 9596 24216 9648
rect 24268 9636 24274 9648
rect 25958 9636 25964 9648
rect 24268 9608 25964 9636
rect 24268 9596 24274 9608
rect 25958 9596 25964 9608
rect 26016 9596 26022 9648
rect 12253 9571 12311 9577
rect 12253 9537 12265 9571
rect 12299 9568 12311 9571
rect 12526 9568 12532 9580
rect 12299 9540 12532 9568
rect 12299 9537 12311 9540
rect 12253 9531 12311 9537
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 14642 9568 14648 9580
rect 14603 9540 14648 9568
rect 14642 9528 14648 9540
rect 14700 9528 14706 9580
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1486 9500 1492 9512
rect 1443 9472 1492 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1486 9460 1492 9472
rect 1544 9500 1550 9512
rect 1949 9503 2007 9509
rect 1949 9500 1961 9503
rect 1544 9472 1961 9500
rect 1544 9460 1550 9472
rect 1949 9469 1961 9472
rect 1995 9469 2007 9503
rect 1949 9463 2007 9469
rect 14458 9460 14464 9512
rect 14516 9460 14522 9512
rect 14182 9392 14188 9444
rect 14240 9432 14246 9444
rect 14476 9432 14504 9460
rect 14553 9435 14611 9441
rect 14553 9432 14565 9435
rect 14240 9404 14565 9432
rect 14240 9392 14246 9404
rect 14553 9401 14565 9404
rect 14599 9401 14611 9435
rect 14553 9395 14611 9401
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 13906 9324 13912 9376
rect 13964 9364 13970 9376
rect 14001 9367 14059 9373
rect 14001 9364 14013 9367
rect 13964 9336 14013 9364
rect 13964 9324 13970 9336
rect 14001 9333 14013 9336
rect 14047 9364 14059 9367
rect 14461 9367 14519 9373
rect 14461 9364 14473 9367
rect 14047 9336 14473 9364
rect 14047 9333 14059 9336
rect 14001 9327 14059 9333
rect 14461 9333 14473 9336
rect 14507 9364 14519 9367
rect 14826 9364 14832 9376
rect 14507 9336 14832 9364
rect 14507 9333 14519 9336
rect 14461 9327 14519 9333
rect 14826 9324 14832 9336
rect 14884 9324 14890 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1670 9160 1676 9172
rect 1631 9132 1676 9160
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 14182 8820 14188 8832
rect 14143 8792 14188 8820
rect 14182 8780 14188 8792
rect 14240 8780 14246 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 23845 8619 23903 8625
rect 23845 8585 23857 8619
rect 23891 8616 23903 8619
rect 25130 8616 25136 8628
rect 23891 8588 25136 8616
rect 23891 8585 23903 8588
rect 23845 8579 23903 8585
rect 25130 8576 25136 8588
rect 25188 8576 25194 8628
rect 23658 8412 23664 8424
rect 23619 8384 23664 8412
rect 23658 8372 23664 8384
rect 23716 8412 23722 8424
rect 24213 8415 24271 8421
rect 24213 8412 24225 8415
rect 23716 8384 24225 8412
rect 23716 8372 23722 8384
rect 24213 8381 24225 8384
rect 24259 8381 24271 8415
rect 24213 8375 24271 8381
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 24210 5896 24216 5908
rect 24171 5868 24216 5896
rect 24210 5856 24216 5868
rect 24268 5856 24274 5908
rect 24026 5760 24032 5772
rect 23987 5732 24032 5760
rect 24026 5720 24032 5732
rect 24084 5720 24090 5772
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 24026 5352 24032 5364
rect 23987 5324 24032 5352
rect 24026 5312 24032 5324
rect 24084 5312 24090 5364
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 24118 4808 24124 4820
rect 24079 4780 24124 4808
rect 24118 4768 24124 4780
rect 24176 4768 24182 4820
rect 24581 4743 24639 4749
rect 24581 4709 24593 4743
rect 24627 4740 24639 4743
rect 24670 4740 24676 4752
rect 24627 4712 24676 4740
rect 24627 4709 24639 4712
rect 24581 4703 24639 4709
rect 24670 4700 24676 4712
rect 24728 4700 24734 4752
rect 24118 4632 24124 4684
rect 24176 4672 24182 4684
rect 24489 4675 24547 4681
rect 24489 4672 24501 4675
rect 24176 4644 24501 4672
rect 24176 4632 24182 4644
rect 24489 4641 24501 4644
rect 24535 4641 24547 4675
rect 24489 4635 24547 4641
rect 24762 4604 24768 4616
rect 24723 4576 24768 4604
rect 24762 4564 24768 4576
rect 24820 4564 24826 4616
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 566 4224 572 4276
rect 624 4264 630 4276
rect 8202 4264 8208 4276
rect 624 4236 8208 4264
rect 624 4224 630 4236
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 17954 4156 17960 4208
rect 18012 4196 18018 4208
rect 24118 4196 24124 4208
rect 18012 4168 24124 4196
rect 18012 4156 18018 4168
rect 24118 4156 24124 4168
rect 24176 4156 24182 4208
rect 24762 4156 24768 4208
rect 24820 4156 24826 4208
rect 24780 4128 24808 4156
rect 24857 4131 24915 4137
rect 24857 4128 24869 4131
rect 24780 4100 24869 4128
rect 24857 4097 24869 4100
rect 24903 4097 24915 4131
rect 24857 4091 24915 4097
rect 24578 3924 24584 3936
rect 24539 3896 24584 3924
rect 24578 3884 24584 3896
rect 24636 3884 24642 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 934 3680 940 3732
rect 992 3720 998 3732
rect 2958 3720 2964 3732
rect 992 3692 2964 3720
rect 992 3680 998 3692
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1302 2864 1308 2916
rect 1360 2904 1366 2916
rect 3510 2904 3516 2916
rect 1360 2876 3516 2904
rect 1360 2864 1366 2876
rect 3510 2864 3516 2876
rect 3568 2864 3574 2916
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 11974 2632 11980 2644
rect 11935 2604 11980 2632
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 12434 2632 12440 2644
rect 12395 2604 12440 2632
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 14001 2635 14059 2641
rect 14001 2601 14013 2635
rect 14047 2632 14059 2635
rect 14090 2632 14096 2644
rect 14047 2604 14096 2632
rect 14047 2601 14059 2604
rect 14001 2595 14059 2601
rect 14090 2592 14096 2604
rect 14148 2592 14154 2644
rect 25317 2635 25375 2641
rect 25317 2601 25329 2635
rect 25363 2632 25375 2635
rect 26510 2632 26516 2644
rect 25363 2604 26516 2632
rect 25363 2601 25375 2604
rect 25317 2595 25375 2601
rect 26510 2592 26516 2604
rect 26568 2592 26574 2644
rect 11992 2496 12020 2592
rect 12452 2564 12480 2592
rect 12866 2567 12924 2573
rect 12866 2564 12878 2567
rect 12452 2536 12878 2564
rect 12866 2533 12878 2536
rect 12912 2533 12924 2567
rect 12866 2527 12924 2533
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 11992 2468 12633 2496
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 25130 2496 25136 2508
rect 25091 2468 25136 2496
rect 12621 2459 12679 2465
rect 25130 2456 25136 2468
rect 25188 2496 25194 2508
rect 25685 2499 25743 2505
rect 25685 2496 25697 2499
rect 25188 2468 25697 2496
rect 25188 2456 25194 2468
rect 25685 2465 25697 2468
rect 25731 2465 25743 2499
rect 25685 2459 25743 2465
rect 24213 2295 24271 2301
rect 24213 2261 24225 2295
rect 24259 2292 24271 2295
rect 25130 2292 25136 2304
rect 24259 2264 25136 2292
rect 24259 2261 24271 2264
rect 24213 2255 24271 2261
rect 25130 2252 25136 2264
rect 25188 2252 25194 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 8668 27412 8720 27464
rect 8760 27412 8812 27464
rect 27068 27455 27120 27464
rect 27068 27421 27077 27455
rect 27077 27421 27111 27455
rect 27111 27421 27120 27455
rect 27068 27412 27120 27421
rect 3516 26256 3568 26308
rect 8392 26256 8444 26308
rect 4252 25984 4304 26036
rect 17776 25984 17828 26036
rect 14372 25916 14424 25968
rect 20352 25916 20404 25968
rect 14556 25848 14608 25900
rect 24032 25848 24084 25900
rect 3608 25644 3660 25696
rect 16856 25780 16908 25832
rect 13452 25712 13504 25764
rect 25044 25712 25096 25764
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 4160 25440 4212 25492
rect 4344 25440 4396 25492
rect 14372 25440 14424 25492
rect 16120 25440 16172 25492
rect 16488 25440 16540 25492
rect 20904 25440 20956 25492
rect 24768 25483 24820 25492
rect 24768 25449 24777 25483
rect 24777 25449 24811 25483
rect 24811 25449 24820 25483
rect 24768 25440 24820 25449
rect 14004 25372 14056 25424
rect 2044 25304 2096 25356
rect 3424 25304 3476 25356
rect 4528 25304 4580 25356
rect 5172 25347 5224 25356
rect 5172 25313 5181 25347
rect 5181 25313 5215 25347
rect 5215 25313 5224 25347
rect 5172 25304 5224 25313
rect 6184 25304 6236 25356
rect 7932 25304 7984 25356
rect 10324 25347 10376 25356
rect 10324 25313 10333 25347
rect 10333 25313 10367 25347
rect 10367 25313 10376 25347
rect 10324 25304 10376 25313
rect 12072 25304 12124 25356
rect 12992 25347 13044 25356
rect 12992 25313 13001 25347
rect 13001 25313 13035 25347
rect 13035 25313 13044 25347
rect 12992 25304 13044 25313
rect 20260 25372 20312 25424
rect 19800 25304 19852 25356
rect 20076 25304 20128 25356
rect 22468 25304 22520 25356
rect 23848 25304 23900 25356
rect 25136 25304 25188 25356
rect 7748 25279 7800 25288
rect 7748 25245 7757 25279
rect 7757 25245 7791 25279
rect 7791 25245 7800 25279
rect 7748 25236 7800 25245
rect 13268 25279 13320 25288
rect 2964 25168 3016 25220
rect 7380 25168 7432 25220
rect 12256 25168 12308 25220
rect 13268 25245 13277 25279
rect 13277 25245 13311 25279
rect 13311 25245 13320 25279
rect 13268 25236 13320 25245
rect 15844 25236 15896 25288
rect 16028 25279 16080 25288
rect 16028 25245 16037 25279
rect 16037 25245 16071 25279
rect 16071 25245 16080 25279
rect 16028 25236 16080 25245
rect 16396 25236 16448 25288
rect 17684 25236 17736 25288
rect 22284 25236 22336 25288
rect 2872 25100 2924 25152
rect 4712 25143 4764 25152
rect 4712 25109 4721 25143
rect 4721 25109 4755 25143
rect 4755 25109 4764 25143
rect 4712 25100 4764 25109
rect 7104 25143 7156 25152
rect 7104 25109 7113 25143
rect 7113 25109 7147 25143
rect 7147 25109 7156 25143
rect 7104 25100 7156 25109
rect 8944 25100 8996 25152
rect 11612 25143 11664 25152
rect 11612 25109 11621 25143
rect 11621 25109 11655 25143
rect 11655 25109 11664 25143
rect 11612 25100 11664 25109
rect 13820 25100 13872 25152
rect 14372 25168 14424 25220
rect 17592 25168 17644 25220
rect 15476 25100 15528 25152
rect 16212 25100 16264 25152
rect 16580 25143 16632 25152
rect 16580 25109 16589 25143
rect 16589 25109 16623 25143
rect 16623 25109 16632 25143
rect 16580 25100 16632 25109
rect 19432 25168 19484 25220
rect 24768 25168 24820 25220
rect 18328 25143 18380 25152
rect 18328 25109 18337 25143
rect 18337 25109 18371 25143
rect 18371 25109 18380 25143
rect 18328 25100 18380 25109
rect 18696 25100 18748 25152
rect 19984 25100 20036 25152
rect 21548 25100 21600 25152
rect 21732 25143 21784 25152
rect 21732 25109 21741 25143
rect 21741 25109 21775 25143
rect 21775 25109 21784 25143
rect 21732 25100 21784 25109
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 3792 24939 3844 24948
rect 3792 24905 3801 24939
rect 3801 24905 3835 24939
rect 3835 24905 3844 24939
rect 3792 24896 3844 24905
rect 3884 24896 3936 24948
rect 10324 24896 10376 24948
rect 1860 24828 1912 24880
rect 4712 24828 4764 24880
rect 4252 24803 4304 24812
rect 4252 24769 4261 24803
rect 4261 24769 4295 24803
rect 4295 24769 4304 24803
rect 4252 24760 4304 24769
rect 2596 24692 2648 24744
rect 4160 24692 4212 24744
rect 4804 24760 4856 24812
rect 5356 24760 5408 24812
rect 7380 24803 7432 24812
rect 7380 24769 7389 24803
rect 7389 24769 7423 24803
rect 7423 24769 7432 24803
rect 7380 24760 7432 24769
rect 7840 24828 7892 24880
rect 8944 24803 8996 24812
rect 8944 24769 8953 24803
rect 8953 24769 8987 24803
rect 8987 24769 8996 24803
rect 8944 24760 8996 24769
rect 11612 24896 11664 24948
rect 13176 24828 13228 24880
rect 13636 24828 13688 24880
rect 18328 24896 18380 24948
rect 25412 24896 25464 24948
rect 19524 24828 19576 24880
rect 19800 24871 19852 24880
rect 19800 24837 19809 24871
rect 19809 24837 19843 24871
rect 19843 24837 19852 24871
rect 19800 24828 19852 24837
rect 20076 24828 20128 24880
rect 21732 24828 21784 24880
rect 25136 24871 25188 24880
rect 7104 24692 7156 24744
rect 8852 24667 8904 24676
rect 8852 24633 8861 24667
rect 8861 24633 8895 24667
rect 8895 24633 8904 24667
rect 8852 24624 8904 24633
rect 1584 24599 1636 24608
rect 1584 24565 1593 24599
rect 1593 24565 1627 24599
rect 1627 24565 1636 24599
rect 1584 24556 1636 24565
rect 2044 24599 2096 24608
rect 2044 24565 2053 24599
rect 2053 24565 2087 24599
rect 2087 24565 2096 24599
rect 2044 24556 2096 24565
rect 2412 24599 2464 24608
rect 2412 24565 2421 24599
rect 2421 24565 2455 24599
rect 2455 24565 2464 24599
rect 2412 24556 2464 24565
rect 2688 24599 2740 24608
rect 2688 24565 2697 24599
rect 2697 24565 2731 24599
rect 2731 24565 2740 24599
rect 2688 24556 2740 24565
rect 3424 24556 3476 24608
rect 4528 24599 4580 24608
rect 4528 24565 4537 24599
rect 4537 24565 4571 24599
rect 4571 24565 4580 24599
rect 4528 24556 4580 24565
rect 5172 24556 5224 24608
rect 6184 24599 6236 24608
rect 6184 24565 6193 24599
rect 6193 24565 6227 24599
rect 6227 24565 6236 24599
rect 6184 24556 6236 24565
rect 7012 24556 7064 24608
rect 7932 24599 7984 24608
rect 7932 24565 7941 24599
rect 7941 24565 7975 24599
rect 7975 24565 7984 24599
rect 7932 24556 7984 24565
rect 8484 24599 8536 24608
rect 8484 24565 8493 24599
rect 8493 24565 8527 24599
rect 8527 24565 8536 24599
rect 8484 24556 8536 24565
rect 12256 24803 12308 24812
rect 12256 24769 12265 24803
rect 12265 24769 12299 24803
rect 12299 24769 12308 24803
rect 12256 24760 12308 24769
rect 13452 24760 13504 24812
rect 14372 24760 14424 24812
rect 17776 24803 17828 24812
rect 9864 24624 9916 24676
rect 13268 24692 13320 24744
rect 13636 24692 13688 24744
rect 14004 24735 14056 24744
rect 14004 24701 14013 24735
rect 14013 24701 14047 24735
rect 14047 24701 14056 24735
rect 14004 24692 14056 24701
rect 14740 24692 14792 24744
rect 17776 24769 17785 24803
rect 17785 24769 17819 24803
rect 17819 24769 17828 24803
rect 17776 24760 17828 24769
rect 18788 24803 18840 24812
rect 18788 24769 18797 24803
rect 18797 24769 18831 24803
rect 18831 24769 18840 24803
rect 18788 24760 18840 24769
rect 25136 24837 25145 24871
rect 25145 24837 25179 24871
rect 25179 24837 25188 24871
rect 25136 24828 25188 24837
rect 12624 24624 12676 24676
rect 14096 24667 14148 24676
rect 14096 24633 14105 24667
rect 14105 24633 14139 24667
rect 14139 24633 14148 24667
rect 14096 24624 14148 24633
rect 18420 24692 18472 24744
rect 22652 24760 22704 24812
rect 23204 24760 23256 24812
rect 24032 24760 24084 24812
rect 21456 24692 21508 24744
rect 18328 24624 18380 24676
rect 21180 24667 21232 24676
rect 9956 24556 10008 24608
rect 10968 24599 11020 24608
rect 10968 24565 10977 24599
rect 10977 24565 11011 24599
rect 11011 24565 11020 24599
rect 10968 24556 11020 24565
rect 11980 24556 12032 24608
rect 12716 24599 12768 24608
rect 12716 24565 12725 24599
rect 12725 24565 12759 24599
rect 12759 24565 12768 24599
rect 12716 24556 12768 24565
rect 14004 24556 14056 24608
rect 14740 24599 14792 24608
rect 14740 24565 14749 24599
rect 14749 24565 14783 24599
rect 14783 24565 14792 24599
rect 14740 24556 14792 24565
rect 15108 24599 15160 24608
rect 15108 24565 15117 24599
rect 15117 24565 15151 24599
rect 15151 24565 15160 24599
rect 15108 24556 15160 24565
rect 15476 24556 15528 24608
rect 15844 24556 15896 24608
rect 16120 24556 16172 24608
rect 16396 24556 16448 24608
rect 17316 24556 17368 24608
rect 17684 24556 17736 24608
rect 18236 24599 18288 24608
rect 18236 24565 18245 24599
rect 18245 24565 18279 24599
rect 18279 24565 18288 24599
rect 18236 24556 18288 24565
rect 19340 24556 19392 24608
rect 19984 24556 20036 24608
rect 21180 24633 21189 24667
rect 21189 24633 21223 24667
rect 21223 24633 21232 24667
rect 21180 24624 21232 24633
rect 21548 24624 21600 24676
rect 22652 24624 22704 24676
rect 23112 24624 23164 24676
rect 20720 24556 20772 24608
rect 21364 24599 21416 24608
rect 21364 24565 21373 24599
rect 21373 24565 21407 24599
rect 21407 24565 21416 24599
rect 21364 24556 21416 24565
rect 21640 24556 21692 24608
rect 21824 24599 21876 24608
rect 21824 24565 21833 24599
rect 21833 24565 21867 24599
rect 21867 24565 21876 24599
rect 21824 24556 21876 24565
rect 22468 24599 22520 24608
rect 22468 24565 22477 24599
rect 22477 24565 22511 24599
rect 22511 24565 22520 24599
rect 22468 24556 22520 24565
rect 23388 24556 23440 24608
rect 24676 24556 24728 24608
rect 24860 24556 24912 24608
rect 25136 24556 25188 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 2044 24395 2096 24404
rect 2044 24361 2053 24395
rect 2053 24361 2087 24395
rect 2087 24361 2096 24395
rect 2044 24352 2096 24361
rect 4252 24395 4304 24404
rect 4252 24361 4261 24395
rect 4261 24361 4295 24395
rect 4295 24361 4304 24395
rect 4252 24352 4304 24361
rect 9588 24352 9640 24404
rect 9680 24352 9732 24404
rect 12440 24352 12492 24404
rect 12992 24352 13044 24404
rect 13452 24352 13504 24404
rect 14004 24352 14056 24404
rect 15292 24352 15344 24404
rect 15936 24352 15988 24404
rect 16212 24395 16264 24404
rect 16212 24361 16221 24395
rect 16221 24361 16255 24395
rect 16255 24361 16264 24395
rect 16212 24352 16264 24361
rect 18236 24352 18288 24404
rect 19984 24352 20036 24404
rect 20904 24395 20956 24404
rect 20904 24361 20913 24395
rect 20913 24361 20947 24395
rect 20947 24361 20956 24395
rect 20904 24352 20956 24361
rect 22100 24352 22152 24404
rect 23112 24352 23164 24404
rect 24124 24352 24176 24404
rect 9220 24284 9272 24336
rect 9496 24284 9548 24336
rect 10048 24327 10100 24336
rect 10048 24293 10057 24327
rect 10057 24293 10091 24327
rect 10091 24293 10100 24327
rect 10048 24284 10100 24293
rect 12072 24284 12124 24336
rect 15568 24284 15620 24336
rect 16028 24284 16080 24336
rect 16304 24284 16356 24336
rect 18420 24327 18472 24336
rect 18420 24293 18429 24327
rect 18429 24293 18463 24327
rect 18463 24293 18472 24327
rect 18420 24284 18472 24293
rect 22744 24284 22796 24336
rect 1676 24216 1728 24268
rect 2504 24259 2556 24268
rect 2504 24225 2513 24259
rect 2513 24225 2547 24259
rect 2547 24225 2556 24259
rect 2504 24216 2556 24225
rect 4068 24259 4120 24268
rect 4068 24225 4077 24259
rect 4077 24225 4111 24259
rect 4111 24225 4120 24259
rect 4068 24216 4120 24225
rect 5540 24216 5592 24268
rect 9036 24216 9088 24268
rect 10140 24216 10192 24268
rect 10876 24216 10928 24268
rect 11428 24216 11480 24268
rect 13544 24216 13596 24268
rect 14556 24216 14608 24268
rect 1400 24012 1452 24064
rect 1768 24012 1820 24064
rect 4896 24012 4948 24064
rect 9956 24080 10008 24132
rect 10692 24148 10744 24200
rect 12348 24191 12400 24200
rect 12348 24157 12357 24191
rect 12357 24157 12391 24191
rect 12391 24157 12400 24191
rect 12348 24148 12400 24157
rect 13728 24080 13780 24132
rect 6000 24012 6052 24064
rect 7104 24012 7156 24064
rect 7748 24012 7800 24064
rect 8300 24012 8352 24064
rect 8852 24012 8904 24064
rect 11336 24012 11388 24064
rect 11796 24055 11848 24064
rect 11796 24021 11805 24055
rect 11805 24021 11839 24055
rect 11839 24021 11848 24055
rect 11796 24012 11848 24021
rect 13360 24055 13412 24064
rect 13360 24021 13369 24055
rect 13369 24021 13403 24055
rect 13403 24021 13412 24055
rect 13360 24012 13412 24021
rect 14832 24012 14884 24064
rect 16580 24216 16632 24268
rect 16764 24259 16816 24268
rect 16764 24225 16798 24259
rect 16798 24225 16816 24259
rect 19340 24259 19392 24268
rect 16764 24216 16816 24225
rect 19340 24225 19349 24259
rect 19349 24225 19383 24259
rect 19383 24225 19392 24259
rect 19340 24216 19392 24225
rect 21088 24216 21140 24268
rect 22836 24259 22888 24268
rect 22836 24225 22845 24259
rect 22845 24225 22879 24259
rect 22879 24225 22888 24259
rect 22836 24216 22888 24225
rect 24676 24216 24728 24268
rect 15108 24148 15160 24200
rect 15936 24148 15988 24200
rect 19524 24191 19576 24200
rect 19524 24157 19533 24191
rect 19533 24157 19567 24191
rect 19567 24157 19576 24191
rect 19524 24148 19576 24157
rect 20444 24148 20496 24200
rect 21456 24191 21508 24200
rect 21456 24157 21465 24191
rect 21465 24157 21499 24191
rect 21499 24157 21508 24191
rect 23020 24191 23072 24200
rect 21456 24148 21508 24157
rect 23020 24157 23029 24191
rect 23029 24157 23063 24191
rect 23063 24157 23072 24191
rect 23020 24148 23072 24157
rect 17776 24080 17828 24132
rect 21272 24080 21324 24132
rect 17868 24055 17920 24064
rect 17868 24021 17877 24055
rect 17877 24021 17911 24055
rect 17911 24021 17920 24055
rect 17868 24012 17920 24021
rect 18788 24055 18840 24064
rect 18788 24021 18797 24055
rect 18797 24021 18831 24055
rect 18831 24021 18840 24055
rect 18788 24012 18840 24021
rect 20536 24055 20588 24064
rect 20536 24021 20545 24055
rect 20545 24021 20579 24055
rect 20579 24021 20588 24055
rect 20536 24012 20588 24021
rect 22192 24012 22244 24064
rect 22376 24012 22428 24064
rect 24032 24012 24084 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2504 23808 2556 23860
rect 7380 23808 7432 23860
rect 9680 23851 9732 23860
rect 9680 23817 9689 23851
rect 9689 23817 9723 23851
rect 9723 23817 9732 23851
rect 9680 23808 9732 23817
rect 10048 23851 10100 23860
rect 10048 23817 10057 23851
rect 10057 23817 10091 23851
rect 10091 23817 10100 23851
rect 10048 23808 10100 23817
rect 12348 23808 12400 23860
rect 13544 23808 13596 23860
rect 15384 23851 15436 23860
rect 15384 23817 15393 23851
rect 15393 23817 15427 23851
rect 15427 23817 15436 23851
rect 15384 23808 15436 23817
rect 16764 23851 16816 23860
rect 4068 23740 4120 23792
rect 5080 23740 5132 23792
rect 6644 23740 6696 23792
rect 10876 23740 10928 23792
rect 14372 23740 14424 23792
rect 14556 23740 14608 23792
rect 1860 23715 1912 23724
rect 1860 23681 1869 23715
rect 1869 23681 1903 23715
rect 1903 23681 1912 23715
rect 1860 23672 1912 23681
rect 3792 23715 3844 23724
rect 3792 23681 3801 23715
rect 3801 23681 3835 23715
rect 3835 23681 3844 23715
rect 3792 23672 3844 23681
rect 7288 23715 7340 23724
rect 7288 23681 7297 23715
rect 7297 23681 7331 23715
rect 7331 23681 7340 23715
rect 7288 23672 7340 23681
rect 7472 23715 7524 23724
rect 7472 23681 7481 23715
rect 7481 23681 7515 23715
rect 7515 23681 7524 23715
rect 7472 23672 7524 23681
rect 8852 23715 8904 23724
rect 8852 23681 8861 23715
rect 8861 23681 8895 23715
rect 8895 23681 8904 23715
rect 8852 23672 8904 23681
rect 2044 23604 2096 23656
rect 2872 23647 2924 23656
rect 2872 23613 2881 23647
rect 2881 23613 2915 23647
rect 2915 23613 2924 23647
rect 2872 23604 2924 23613
rect 4896 23647 4948 23656
rect 4896 23613 4905 23647
rect 4905 23613 4939 23647
rect 4939 23613 4948 23647
rect 4896 23604 4948 23613
rect 5172 23604 5224 23656
rect 6000 23604 6052 23656
rect 6736 23604 6788 23656
rect 8484 23604 8536 23656
rect 2412 23536 2464 23588
rect 3056 23511 3108 23520
rect 3056 23477 3065 23511
rect 3065 23477 3099 23511
rect 3099 23477 3108 23511
rect 3056 23468 3108 23477
rect 4436 23511 4488 23520
rect 4436 23477 4445 23511
rect 4445 23477 4479 23511
rect 4479 23477 4488 23511
rect 4436 23468 4488 23477
rect 4896 23468 4948 23520
rect 5540 23468 5592 23520
rect 6828 23511 6880 23520
rect 6828 23477 6837 23511
rect 6837 23477 6871 23511
rect 6871 23477 6880 23511
rect 6828 23468 6880 23477
rect 7288 23536 7340 23588
rect 7932 23536 7984 23588
rect 11336 23672 11388 23724
rect 16764 23817 16773 23851
rect 16773 23817 16807 23851
rect 16807 23817 16816 23851
rect 16764 23808 16816 23817
rect 19524 23808 19576 23860
rect 19984 23851 20036 23860
rect 19984 23817 19993 23851
rect 19993 23817 20027 23851
rect 20027 23817 20036 23851
rect 19984 23808 20036 23817
rect 20444 23851 20496 23860
rect 20444 23817 20453 23851
rect 20453 23817 20487 23851
rect 20487 23817 20496 23851
rect 20444 23808 20496 23817
rect 23940 23808 23992 23860
rect 16580 23740 16632 23792
rect 17224 23740 17276 23792
rect 19340 23740 19392 23792
rect 20720 23672 20772 23724
rect 22008 23672 22060 23724
rect 10784 23604 10836 23656
rect 12440 23647 12492 23656
rect 12440 23613 12449 23647
rect 12449 23613 12483 23647
rect 12483 23613 12492 23647
rect 12440 23604 12492 23613
rect 16212 23604 16264 23656
rect 18696 23604 18748 23656
rect 22192 23604 22244 23656
rect 24216 23715 24268 23724
rect 24216 23681 24225 23715
rect 24225 23681 24259 23715
rect 24259 23681 24268 23715
rect 24216 23672 24268 23681
rect 24768 23604 24820 23656
rect 7380 23468 7432 23520
rect 8300 23511 8352 23520
rect 8300 23477 8309 23511
rect 8309 23477 8343 23511
rect 8343 23477 8352 23511
rect 8300 23468 8352 23477
rect 10692 23468 10744 23520
rect 10968 23468 11020 23520
rect 11428 23511 11480 23520
rect 11428 23477 11437 23511
rect 11437 23477 11471 23511
rect 11471 23477 11480 23511
rect 11428 23468 11480 23477
rect 12348 23468 12400 23520
rect 15292 23536 15344 23588
rect 17868 23579 17920 23588
rect 17868 23545 17877 23579
rect 17877 23545 17911 23579
rect 17911 23545 17920 23579
rect 17868 23536 17920 23545
rect 18788 23536 18840 23588
rect 19156 23536 19208 23588
rect 20536 23536 20588 23588
rect 22560 23579 22612 23588
rect 22560 23545 22569 23579
rect 22569 23545 22603 23579
rect 22603 23545 22612 23579
rect 22560 23536 22612 23545
rect 23940 23536 23992 23588
rect 24676 23579 24728 23588
rect 24676 23545 24685 23579
rect 24685 23545 24719 23579
rect 24719 23545 24728 23579
rect 24676 23536 24728 23545
rect 12992 23468 13044 23520
rect 14004 23468 14056 23520
rect 15384 23468 15436 23520
rect 16948 23511 17000 23520
rect 16948 23477 16957 23511
rect 16957 23477 16991 23511
rect 16991 23477 17000 23511
rect 16948 23468 17000 23477
rect 20812 23468 20864 23520
rect 21088 23468 21140 23520
rect 22744 23468 22796 23520
rect 22928 23468 22980 23520
rect 23664 23511 23716 23520
rect 23664 23477 23673 23511
rect 23673 23477 23707 23511
rect 23707 23477 23716 23511
rect 23664 23468 23716 23477
rect 24032 23511 24084 23520
rect 24032 23477 24041 23511
rect 24041 23477 24075 23511
rect 24075 23477 24084 23511
rect 24032 23468 24084 23477
rect 25412 23511 25464 23520
rect 25412 23477 25421 23511
rect 25421 23477 25455 23511
rect 25455 23477 25464 23511
rect 25412 23468 25464 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 2872 23307 2924 23316
rect 2872 23273 2881 23307
rect 2881 23273 2915 23307
rect 2915 23273 2924 23307
rect 2872 23264 2924 23273
rect 5540 23264 5592 23316
rect 8024 23307 8076 23316
rect 8024 23273 8033 23307
rect 8033 23273 8067 23307
rect 8067 23273 8076 23307
rect 8024 23264 8076 23273
rect 8484 23264 8536 23316
rect 9680 23264 9732 23316
rect 10140 23264 10192 23316
rect 12348 23307 12400 23316
rect 12348 23273 12357 23307
rect 12357 23273 12391 23307
rect 12391 23273 12400 23307
rect 12348 23264 12400 23273
rect 13912 23307 13964 23316
rect 2596 23196 2648 23248
rect 5448 23196 5500 23248
rect 13912 23273 13921 23307
rect 13921 23273 13955 23307
rect 13955 23273 13964 23307
rect 13912 23264 13964 23273
rect 16764 23264 16816 23316
rect 17224 23307 17276 23316
rect 17224 23273 17233 23307
rect 17233 23273 17267 23307
rect 17267 23273 17276 23307
rect 17224 23264 17276 23273
rect 19524 23264 19576 23316
rect 20720 23264 20772 23316
rect 24216 23307 24268 23316
rect 24216 23273 24225 23307
rect 24225 23273 24259 23307
rect 24259 23273 24268 23307
rect 24216 23264 24268 23273
rect 25136 23264 25188 23316
rect 25320 23264 25372 23316
rect 2504 23128 2556 23180
rect 3884 23128 3936 23180
rect 5172 23128 5224 23180
rect 7932 23171 7984 23180
rect 3976 23060 4028 23112
rect 7932 23137 7941 23171
rect 7941 23137 7975 23171
rect 7975 23137 7984 23171
rect 7932 23128 7984 23137
rect 9588 23128 9640 23180
rect 11612 23128 11664 23180
rect 13268 23128 13320 23180
rect 16580 23196 16632 23248
rect 16028 23128 16080 23180
rect 16396 23128 16448 23180
rect 19248 23196 19300 23248
rect 22100 23239 22152 23248
rect 22100 23205 22134 23239
rect 22134 23205 22152 23239
rect 22100 23196 22152 23205
rect 23664 23196 23716 23248
rect 25872 23196 25924 23248
rect 19616 23171 19668 23180
rect 19616 23137 19625 23171
rect 19625 23137 19659 23171
rect 19659 23137 19668 23171
rect 19616 23128 19668 23137
rect 20076 23128 20128 23180
rect 24032 23128 24084 23180
rect 24768 23171 24820 23180
rect 24768 23137 24777 23171
rect 24777 23137 24811 23171
rect 24811 23137 24820 23171
rect 24768 23128 24820 23137
rect 7472 23060 7524 23112
rect 9036 23103 9088 23112
rect 9036 23069 9045 23103
rect 9045 23069 9079 23103
rect 9079 23069 9088 23103
rect 9036 23060 9088 23069
rect 10140 23060 10192 23112
rect 14004 23103 14056 23112
rect 14004 23069 14013 23103
rect 14013 23069 14047 23103
rect 14047 23069 14056 23103
rect 14004 23060 14056 23069
rect 18972 23060 19024 23112
rect 19708 23103 19760 23112
rect 19708 23069 19717 23103
rect 19717 23069 19751 23103
rect 19751 23069 19760 23103
rect 19708 23060 19760 23069
rect 20536 23060 20588 23112
rect 20812 23060 20864 23112
rect 21640 23060 21692 23112
rect 24860 23103 24912 23112
rect 24860 23069 24869 23103
rect 24869 23069 24903 23103
rect 24903 23069 24912 23103
rect 24860 23060 24912 23069
rect 1676 22967 1728 22976
rect 1676 22933 1685 22967
rect 1685 22933 1719 22967
rect 1719 22933 1728 22967
rect 1676 22924 1728 22933
rect 3700 22967 3752 22976
rect 3700 22933 3709 22967
rect 3709 22933 3743 22967
rect 3743 22933 3752 22967
rect 3700 22924 3752 22933
rect 4896 22924 4948 22976
rect 7472 22924 7524 22976
rect 9312 22924 9364 22976
rect 9956 22924 10008 22976
rect 10416 22967 10468 22976
rect 10416 22933 10425 22967
rect 10425 22933 10459 22967
rect 10459 22933 10468 22967
rect 10416 22924 10468 22933
rect 10784 22967 10836 22976
rect 10784 22933 10793 22967
rect 10793 22933 10827 22967
rect 10827 22933 10836 22967
rect 10784 22924 10836 22933
rect 12440 22924 12492 22976
rect 14556 22992 14608 23044
rect 14740 22992 14792 23044
rect 19156 22992 19208 23044
rect 23572 22992 23624 23044
rect 13268 22967 13320 22976
rect 13268 22933 13277 22967
rect 13277 22933 13311 22967
rect 13311 22933 13320 22967
rect 13268 22924 13320 22933
rect 15292 22924 15344 22976
rect 20352 22924 20404 22976
rect 21456 22924 21508 22976
rect 23388 22924 23440 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 5448 22720 5500 22772
rect 10968 22720 11020 22772
rect 13912 22720 13964 22772
rect 14740 22763 14792 22772
rect 14740 22729 14749 22763
rect 14749 22729 14783 22763
rect 14783 22729 14792 22763
rect 14740 22720 14792 22729
rect 2504 22695 2556 22704
rect 2504 22661 2513 22695
rect 2513 22661 2547 22695
rect 2547 22661 2556 22695
rect 2504 22652 2556 22661
rect 9956 22652 10008 22704
rect 11428 22695 11480 22704
rect 11428 22661 11437 22695
rect 11437 22661 11471 22695
rect 11471 22661 11480 22695
rect 11428 22652 11480 22661
rect 2872 22584 2924 22636
rect 4160 22627 4212 22636
rect 4160 22593 4169 22627
rect 4169 22593 4203 22627
rect 4203 22593 4212 22627
rect 16580 22720 16632 22772
rect 4160 22584 4212 22593
rect 2044 22516 2096 22568
rect 3976 22559 4028 22568
rect 3976 22525 3985 22559
rect 3985 22525 4019 22559
rect 4019 22525 4028 22559
rect 3976 22516 4028 22525
rect 3148 22423 3200 22432
rect 3148 22389 3157 22423
rect 3157 22389 3191 22423
rect 3191 22389 3200 22423
rect 3148 22380 3200 22389
rect 6000 22448 6052 22500
rect 6736 22516 6788 22568
rect 7656 22516 7708 22568
rect 9128 22516 9180 22568
rect 7104 22448 7156 22500
rect 3700 22380 3752 22432
rect 5080 22380 5132 22432
rect 6460 22380 6512 22432
rect 8208 22380 8260 22432
rect 10416 22448 10468 22500
rect 9128 22423 9180 22432
rect 9128 22389 9137 22423
rect 9137 22389 9171 22423
rect 9171 22389 9180 22423
rect 9128 22380 9180 22389
rect 9956 22380 10008 22432
rect 12440 22559 12492 22568
rect 12440 22525 12449 22559
rect 12449 22525 12483 22559
rect 12483 22525 12492 22559
rect 12440 22516 12492 22525
rect 16856 22627 16908 22636
rect 14004 22516 14056 22568
rect 14096 22516 14148 22568
rect 15292 22516 15344 22568
rect 16856 22593 16865 22627
rect 16865 22593 16899 22627
rect 16899 22593 16908 22627
rect 16856 22584 16908 22593
rect 17776 22720 17828 22772
rect 19156 22763 19208 22772
rect 19156 22729 19165 22763
rect 19165 22729 19199 22763
rect 19199 22729 19208 22763
rect 19156 22720 19208 22729
rect 19616 22720 19668 22772
rect 19984 22720 20036 22772
rect 20536 22720 20588 22772
rect 22008 22763 22060 22772
rect 22008 22729 22017 22763
rect 22017 22729 22051 22763
rect 22051 22729 22060 22763
rect 22008 22720 22060 22729
rect 22100 22720 22152 22772
rect 24768 22720 24820 22772
rect 25872 22720 25924 22772
rect 18328 22584 18380 22636
rect 19156 22584 19208 22636
rect 23020 22584 23072 22636
rect 18052 22559 18104 22568
rect 18052 22525 18061 22559
rect 18061 22525 18095 22559
rect 18095 22525 18104 22559
rect 18052 22516 18104 22525
rect 18696 22516 18748 22568
rect 19340 22559 19392 22568
rect 19340 22525 19349 22559
rect 19349 22525 19383 22559
rect 19383 22525 19392 22559
rect 19340 22516 19392 22525
rect 21456 22516 21508 22568
rect 23572 22516 23624 22568
rect 15568 22448 15620 22500
rect 15752 22448 15804 22500
rect 18328 22491 18380 22500
rect 18328 22457 18337 22491
rect 18337 22457 18371 22491
rect 18371 22457 18380 22491
rect 18328 22448 18380 22457
rect 19524 22448 19576 22500
rect 19708 22448 19760 22500
rect 11612 22380 11664 22432
rect 11888 22423 11940 22432
rect 11888 22389 11897 22423
rect 11897 22389 11931 22423
rect 11931 22389 11940 22423
rect 11888 22380 11940 22389
rect 13912 22380 13964 22432
rect 14924 22423 14976 22432
rect 14924 22389 14933 22423
rect 14933 22389 14967 22423
rect 14967 22389 14976 22423
rect 14924 22380 14976 22389
rect 15108 22380 15160 22432
rect 16028 22423 16080 22432
rect 16028 22389 16037 22423
rect 16037 22389 16071 22423
rect 16071 22389 16080 22423
rect 16028 22380 16080 22389
rect 18696 22380 18748 22432
rect 20996 22380 21048 22432
rect 24216 22516 24268 22568
rect 23756 22448 23808 22500
rect 23480 22423 23532 22432
rect 23480 22389 23489 22423
rect 23489 22389 23523 22423
rect 23523 22389 23532 22423
rect 23480 22380 23532 22389
rect 24768 22380 24820 22432
rect 26332 22423 26384 22432
rect 26332 22389 26341 22423
rect 26341 22389 26375 22423
rect 26375 22389 26384 22423
rect 26332 22380 26384 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 2780 22219 2832 22228
rect 2780 22185 2789 22219
rect 2789 22185 2823 22219
rect 2823 22185 2832 22219
rect 2780 22176 2832 22185
rect 2964 22176 3016 22228
rect 4160 22176 4212 22228
rect 5448 22219 5500 22228
rect 5448 22185 5457 22219
rect 5457 22185 5491 22219
rect 5491 22185 5500 22219
rect 5448 22176 5500 22185
rect 6000 22219 6052 22228
rect 6000 22185 6009 22219
rect 6009 22185 6043 22219
rect 6043 22185 6052 22219
rect 6000 22176 6052 22185
rect 6460 22176 6512 22228
rect 6920 22219 6972 22228
rect 6920 22185 6929 22219
rect 6929 22185 6963 22219
rect 6963 22185 6972 22219
rect 6920 22176 6972 22185
rect 7104 22176 7156 22228
rect 7472 22176 7524 22228
rect 7932 22219 7984 22228
rect 7932 22185 7941 22219
rect 7941 22185 7975 22219
rect 7975 22185 7984 22219
rect 7932 22176 7984 22185
rect 9680 22176 9732 22228
rect 13268 22176 13320 22228
rect 14004 22176 14056 22228
rect 16028 22176 16080 22228
rect 19524 22176 19576 22228
rect 20076 22176 20128 22228
rect 20536 22219 20588 22228
rect 20536 22185 20545 22219
rect 20545 22185 20579 22219
rect 20579 22185 20588 22219
rect 20536 22176 20588 22185
rect 20720 22176 20772 22228
rect 22100 22176 22152 22228
rect 23020 22176 23072 22228
rect 2228 22108 2280 22160
rect 2872 22151 2924 22160
rect 2872 22117 2881 22151
rect 2881 22117 2915 22151
rect 2915 22117 2924 22151
rect 2872 22108 2924 22117
rect 3608 22108 3660 22160
rect 3884 22108 3936 22160
rect 3976 22108 4028 22160
rect 2320 22040 2372 22092
rect 3148 22040 3200 22092
rect 5540 22108 5592 22160
rect 8024 22108 8076 22160
rect 4344 22083 4396 22092
rect 4344 22049 4378 22083
rect 4378 22049 4396 22083
rect 4344 22040 4396 22049
rect 8116 22083 8168 22092
rect 8116 22049 8125 22083
rect 8125 22049 8159 22083
rect 8159 22049 8168 22083
rect 8116 22040 8168 22049
rect 9588 22040 9640 22092
rect 9956 22040 10008 22092
rect 11244 22083 11296 22092
rect 3240 21972 3292 22024
rect 3792 21972 3844 22024
rect 6552 21972 6604 22024
rect 10048 21972 10100 22024
rect 11244 22049 11253 22083
rect 11253 22049 11287 22083
rect 11287 22049 11296 22083
rect 11244 22040 11296 22049
rect 13360 22108 13412 22160
rect 14004 22040 14056 22092
rect 14832 22040 14884 22092
rect 12808 22015 12860 22024
rect 12808 21981 12817 22015
rect 12817 21981 12851 22015
rect 12851 21981 12860 22015
rect 12808 21972 12860 21981
rect 12992 22015 13044 22024
rect 12992 21981 13001 22015
rect 13001 21981 13035 22015
rect 13035 21981 13044 22015
rect 12992 21972 13044 21981
rect 14280 21972 14332 22024
rect 15108 22040 15160 22092
rect 16580 22108 16632 22160
rect 17960 22108 18012 22160
rect 19340 22108 19392 22160
rect 16396 22040 16448 22092
rect 18420 22040 18472 22092
rect 2596 21904 2648 21956
rect 8392 21904 8444 21956
rect 10968 21904 11020 21956
rect 11428 21947 11480 21956
rect 11428 21913 11437 21947
rect 11437 21913 11471 21947
rect 11471 21913 11480 21947
rect 11428 21904 11480 21913
rect 2412 21879 2464 21888
rect 2412 21845 2421 21879
rect 2421 21845 2455 21879
rect 2455 21845 2464 21879
rect 2412 21836 2464 21845
rect 6460 21879 6512 21888
rect 6460 21845 6469 21879
rect 6469 21845 6503 21879
rect 6503 21845 6512 21879
rect 6460 21836 6512 21845
rect 7656 21836 7708 21888
rect 9036 21836 9088 21888
rect 9312 21836 9364 21888
rect 11244 21836 11296 21888
rect 12256 21836 12308 21888
rect 15292 21836 15344 21888
rect 18788 22015 18840 22024
rect 18788 21981 18797 22015
rect 18797 21981 18831 22015
rect 18831 21981 18840 22015
rect 18788 21972 18840 21981
rect 19892 21972 19944 22024
rect 20076 21972 20128 22024
rect 20260 21972 20312 22024
rect 21640 22040 21692 22092
rect 22560 22108 22612 22160
rect 23480 22108 23532 22160
rect 24768 22108 24820 22160
rect 19064 21904 19116 21956
rect 19984 21904 20036 21956
rect 23388 22040 23440 22092
rect 23756 22015 23808 22024
rect 23756 21981 23765 22015
rect 23765 21981 23799 22015
rect 23799 21981 23808 22015
rect 23756 21972 23808 21981
rect 17500 21836 17552 21888
rect 18144 21879 18196 21888
rect 18144 21845 18153 21879
rect 18153 21845 18187 21879
rect 18187 21845 18196 21879
rect 18144 21836 18196 21845
rect 20260 21836 20312 21888
rect 20536 21836 20588 21888
rect 20812 21836 20864 21888
rect 25136 21879 25188 21888
rect 25136 21845 25145 21879
rect 25145 21845 25179 21879
rect 25179 21845 25188 21879
rect 25136 21836 25188 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1860 21675 1912 21684
rect 1860 21641 1869 21675
rect 1869 21641 1903 21675
rect 1903 21641 1912 21675
rect 1860 21632 1912 21641
rect 2688 21632 2740 21684
rect 5080 21675 5132 21684
rect 5080 21641 5089 21675
rect 5089 21641 5123 21675
rect 5123 21641 5132 21675
rect 5080 21632 5132 21641
rect 6828 21632 6880 21684
rect 7104 21675 7156 21684
rect 7104 21641 7113 21675
rect 7113 21641 7147 21675
rect 7147 21641 7156 21675
rect 7104 21632 7156 21641
rect 9680 21675 9732 21684
rect 9680 21641 9689 21675
rect 9689 21641 9723 21675
rect 9723 21641 9732 21675
rect 9680 21632 9732 21641
rect 10784 21632 10836 21684
rect 11612 21632 11664 21684
rect 5540 21564 5592 21616
rect 6552 21607 6604 21616
rect 6552 21573 6561 21607
rect 6561 21573 6595 21607
rect 6595 21573 6604 21607
rect 6552 21564 6604 21573
rect 2320 21539 2372 21548
rect 2320 21505 2329 21539
rect 2329 21505 2363 21539
rect 2363 21505 2372 21539
rect 2320 21496 2372 21505
rect 5448 21496 5500 21548
rect 7564 21539 7616 21548
rect 7564 21505 7573 21539
rect 7573 21505 7607 21539
rect 7607 21505 7616 21539
rect 7564 21496 7616 21505
rect 10968 21539 11020 21548
rect 10968 21505 10977 21539
rect 10977 21505 11011 21539
rect 11011 21505 11020 21539
rect 10968 21496 11020 21505
rect 11244 21496 11296 21548
rect 12072 21632 12124 21684
rect 12992 21632 13044 21684
rect 17040 21675 17092 21684
rect 17040 21641 17049 21675
rect 17049 21641 17083 21675
rect 17083 21641 17092 21675
rect 17040 21632 17092 21641
rect 17776 21675 17828 21684
rect 17776 21641 17785 21675
rect 17785 21641 17819 21675
rect 17819 21641 17828 21675
rect 17776 21632 17828 21641
rect 20628 21632 20680 21684
rect 22008 21675 22060 21684
rect 22008 21641 22017 21675
rect 22017 21641 22051 21675
rect 22051 21641 22060 21675
rect 22008 21632 22060 21641
rect 24768 21675 24820 21684
rect 24768 21641 24777 21675
rect 24777 21641 24811 21675
rect 24811 21641 24820 21675
rect 24768 21632 24820 21641
rect 25136 21675 25188 21684
rect 25136 21641 25145 21675
rect 25145 21641 25179 21675
rect 25179 21641 25188 21675
rect 25136 21632 25188 21641
rect 12808 21564 12860 21616
rect 18788 21564 18840 21616
rect 22100 21564 22152 21616
rect 13728 21496 13780 21548
rect 14280 21496 14332 21548
rect 18144 21496 18196 21548
rect 20720 21496 20772 21548
rect 22008 21496 22060 21548
rect 24308 21539 24360 21548
rect 24308 21505 24317 21539
rect 24317 21505 24351 21539
rect 24351 21505 24360 21539
rect 25412 21539 25464 21548
rect 24308 21496 24360 21505
rect 25412 21505 25421 21539
rect 25421 21505 25455 21539
rect 25455 21505 25464 21539
rect 25412 21496 25464 21505
rect 2596 21471 2648 21480
rect 2596 21437 2630 21471
rect 2630 21437 2648 21471
rect 2596 21428 2648 21437
rect 3608 21428 3660 21480
rect 7656 21428 7708 21480
rect 8208 21428 8260 21480
rect 13084 21428 13136 21480
rect 13176 21428 13228 21480
rect 15936 21428 15988 21480
rect 18512 21471 18564 21480
rect 8116 21360 8168 21412
rect 10232 21360 10284 21412
rect 10784 21360 10836 21412
rect 14740 21360 14792 21412
rect 2688 21292 2740 21344
rect 4344 21292 4396 21344
rect 5172 21292 5224 21344
rect 8300 21292 8352 21344
rect 10048 21335 10100 21344
rect 10048 21301 10057 21335
rect 10057 21301 10091 21335
rect 10091 21301 10100 21335
rect 10048 21292 10100 21301
rect 12256 21292 12308 21344
rect 12440 21292 12492 21344
rect 15752 21335 15804 21344
rect 15752 21301 15761 21335
rect 15761 21301 15795 21335
rect 15795 21301 15804 21335
rect 15752 21292 15804 21301
rect 16396 21335 16448 21344
rect 16396 21301 16405 21335
rect 16405 21301 16439 21335
rect 16439 21301 16448 21335
rect 16396 21292 16448 21301
rect 18512 21437 18521 21471
rect 18521 21437 18555 21471
rect 18555 21437 18564 21471
rect 18512 21428 18564 21437
rect 22468 21471 22520 21480
rect 22468 21437 22477 21471
rect 22477 21437 22511 21471
rect 22511 21437 22520 21471
rect 22468 21428 22520 21437
rect 23480 21428 23532 21480
rect 25228 21471 25280 21480
rect 25228 21437 25237 21471
rect 25237 21437 25271 21471
rect 25271 21437 25280 21471
rect 25228 21428 25280 21437
rect 17500 21360 17552 21412
rect 20444 21360 20496 21412
rect 22100 21360 22152 21412
rect 16948 21292 17000 21344
rect 17868 21292 17920 21344
rect 18328 21292 18380 21344
rect 21640 21292 21692 21344
rect 22560 21292 22612 21344
rect 23480 21335 23532 21344
rect 23480 21301 23489 21335
rect 23489 21301 23523 21335
rect 23523 21301 23532 21335
rect 23480 21292 23532 21301
rect 23664 21335 23716 21344
rect 23664 21301 23673 21335
rect 23673 21301 23707 21335
rect 23707 21301 23716 21335
rect 23664 21292 23716 21301
rect 26332 21335 26384 21344
rect 26332 21301 26341 21335
rect 26341 21301 26375 21335
rect 26375 21301 26384 21335
rect 26332 21292 26384 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 2044 21131 2096 21140
rect 2044 21097 2053 21131
rect 2053 21097 2087 21131
rect 2087 21097 2096 21131
rect 2044 21088 2096 21097
rect 2964 21088 3016 21140
rect 4528 21131 4580 21140
rect 4528 21097 4537 21131
rect 4537 21097 4571 21131
rect 4571 21097 4580 21131
rect 4528 21088 4580 21097
rect 5172 21131 5224 21140
rect 5172 21097 5181 21131
rect 5181 21097 5215 21131
rect 5215 21097 5224 21131
rect 5172 21088 5224 21097
rect 5448 21131 5500 21140
rect 5448 21097 5457 21131
rect 5457 21097 5491 21131
rect 5491 21097 5500 21131
rect 5448 21088 5500 21097
rect 6460 21131 6512 21140
rect 6460 21097 6469 21131
rect 6469 21097 6503 21131
rect 6503 21097 6512 21131
rect 6460 21088 6512 21097
rect 7656 21131 7708 21140
rect 7656 21097 7665 21131
rect 7665 21097 7699 21131
rect 7699 21097 7708 21131
rect 7656 21088 7708 21097
rect 8208 21088 8260 21140
rect 8576 21088 8628 21140
rect 9036 21131 9088 21140
rect 9036 21097 9045 21131
rect 9045 21097 9079 21131
rect 9079 21097 9088 21131
rect 9036 21088 9088 21097
rect 9404 21131 9456 21140
rect 9404 21097 9413 21131
rect 9413 21097 9447 21131
rect 9447 21097 9456 21131
rect 9404 21088 9456 21097
rect 14556 21131 14608 21140
rect 14556 21097 14565 21131
rect 14565 21097 14599 21131
rect 14599 21097 14608 21131
rect 14556 21088 14608 21097
rect 16672 21131 16724 21140
rect 16672 21097 16681 21131
rect 16681 21097 16715 21131
rect 16715 21097 16724 21131
rect 16672 21088 16724 21097
rect 19156 21131 19208 21140
rect 19156 21097 19165 21131
rect 19165 21097 19199 21131
rect 19199 21097 19208 21131
rect 19156 21088 19208 21097
rect 20444 21131 20496 21140
rect 20444 21097 20453 21131
rect 20453 21097 20487 21131
rect 20487 21097 20496 21131
rect 20444 21088 20496 21097
rect 20536 21088 20588 21140
rect 22008 21088 22060 21140
rect 22192 21131 22244 21140
rect 22192 21097 22201 21131
rect 22201 21097 22235 21131
rect 22235 21097 22244 21131
rect 22192 21088 22244 21097
rect 23664 21131 23716 21140
rect 23664 21097 23673 21131
rect 23673 21097 23707 21131
rect 23707 21097 23716 21131
rect 23664 21088 23716 21097
rect 3240 21020 3292 21072
rect 4436 21063 4488 21072
rect 4436 21029 4445 21063
rect 4445 21029 4479 21063
rect 4479 21029 4488 21063
rect 4436 21020 4488 21029
rect 8116 21020 8168 21072
rect 9496 21020 9548 21072
rect 13268 21020 13320 21072
rect 15752 21020 15804 21072
rect 1860 20952 1912 21004
rect 2596 20927 2648 20936
rect 2596 20893 2605 20927
rect 2605 20893 2639 20927
rect 2639 20893 2648 20927
rect 2596 20884 2648 20893
rect 3608 20884 3660 20936
rect 6092 20884 6144 20936
rect 7012 20952 7064 21004
rect 9956 20952 10008 21004
rect 17592 20995 17644 21004
rect 17592 20961 17601 20995
rect 17601 20961 17635 20995
rect 17635 20961 17644 20995
rect 20168 21020 20220 21072
rect 17592 20952 17644 20961
rect 18052 20995 18104 21004
rect 18052 20961 18086 20995
rect 18086 20961 18104 20995
rect 21180 21020 21232 21072
rect 22376 21020 22428 21072
rect 23480 21020 23532 21072
rect 23848 21020 23900 21072
rect 24308 21020 24360 21072
rect 24676 21020 24728 21072
rect 18052 20952 18104 20961
rect 22008 20952 22060 21004
rect 23388 20952 23440 21004
rect 23756 20995 23808 21004
rect 23756 20961 23765 20995
rect 23765 20961 23799 20995
rect 23799 20961 23808 20995
rect 23756 20952 23808 20961
rect 24768 20952 24820 21004
rect 6644 20927 6696 20936
rect 6644 20893 6653 20927
rect 6653 20893 6687 20927
rect 6687 20893 6696 20927
rect 6644 20884 6696 20893
rect 9864 20884 9916 20936
rect 10048 20884 10100 20936
rect 12440 20927 12492 20936
rect 12440 20893 12449 20927
rect 12449 20893 12483 20927
rect 12483 20893 12492 20927
rect 13176 20927 13228 20936
rect 12440 20884 12492 20893
rect 13176 20893 13185 20927
rect 13185 20893 13219 20927
rect 13219 20893 13228 20927
rect 13176 20884 13228 20893
rect 13360 20927 13412 20936
rect 13360 20893 13369 20927
rect 13369 20893 13403 20927
rect 13403 20893 13412 20927
rect 13360 20884 13412 20893
rect 13912 20884 13964 20936
rect 14280 20884 14332 20936
rect 15292 20927 15344 20936
rect 15292 20893 15301 20927
rect 15301 20893 15335 20927
rect 15335 20893 15344 20927
rect 15292 20884 15344 20893
rect 19248 20884 19300 20936
rect 20720 20884 20772 20936
rect 22468 20884 22520 20936
rect 11980 20816 12032 20868
rect 12532 20816 12584 20868
rect 14096 20816 14148 20868
rect 23020 20816 23072 20868
rect 1860 20791 1912 20800
rect 1860 20757 1869 20791
rect 1869 20757 1903 20791
rect 1903 20757 1912 20791
rect 1860 20748 1912 20757
rect 3516 20791 3568 20800
rect 3516 20757 3525 20791
rect 3525 20757 3559 20791
rect 3559 20757 3568 20791
rect 3516 20748 3568 20757
rect 3976 20748 4028 20800
rect 5540 20748 5592 20800
rect 6184 20748 6236 20800
rect 8024 20791 8076 20800
rect 8024 20757 8033 20791
rect 8033 20757 8067 20791
rect 8067 20757 8076 20791
rect 8024 20748 8076 20757
rect 9956 20791 10008 20800
rect 9956 20757 9965 20791
rect 9965 20757 9999 20791
rect 9999 20757 10008 20791
rect 9956 20748 10008 20757
rect 11612 20791 11664 20800
rect 11612 20757 11621 20791
rect 11621 20757 11655 20791
rect 11655 20757 11664 20791
rect 11612 20748 11664 20757
rect 12716 20791 12768 20800
rect 12716 20757 12725 20791
rect 12725 20757 12759 20791
rect 12759 20757 12768 20791
rect 12716 20748 12768 20757
rect 13912 20748 13964 20800
rect 14004 20748 14056 20800
rect 14648 20748 14700 20800
rect 19248 20748 19300 20800
rect 20812 20748 20864 20800
rect 21824 20748 21876 20800
rect 22100 20748 22152 20800
rect 22376 20748 22428 20800
rect 22560 20748 22612 20800
rect 23480 20748 23532 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 2596 20544 2648 20596
rect 3608 20587 3660 20596
rect 3608 20553 3617 20587
rect 3617 20553 3651 20587
rect 3651 20553 3660 20587
rect 3608 20544 3660 20553
rect 6092 20544 6144 20596
rect 6460 20544 6512 20596
rect 8208 20544 8260 20596
rect 10692 20544 10744 20596
rect 4528 20408 4580 20460
rect 9956 20476 10008 20528
rect 13360 20544 13412 20596
rect 14740 20544 14792 20596
rect 15752 20587 15804 20596
rect 15752 20553 15761 20587
rect 15761 20553 15795 20587
rect 15795 20553 15804 20587
rect 15752 20544 15804 20553
rect 12348 20476 12400 20528
rect 13268 20476 13320 20528
rect 6368 20408 6420 20460
rect 7564 20408 7616 20460
rect 10968 20408 11020 20460
rect 11244 20451 11296 20460
rect 11244 20417 11253 20451
rect 11253 20417 11287 20451
rect 11287 20417 11296 20451
rect 11612 20451 11664 20460
rect 11244 20408 11296 20417
rect 11612 20417 11621 20451
rect 11621 20417 11655 20451
rect 11655 20417 11664 20451
rect 11612 20408 11664 20417
rect 12992 20408 13044 20460
rect 18052 20544 18104 20596
rect 19340 20544 19392 20596
rect 20352 20544 20404 20596
rect 21180 20587 21232 20596
rect 21180 20553 21189 20587
rect 21189 20553 21223 20587
rect 21223 20553 21232 20587
rect 21180 20544 21232 20553
rect 23020 20544 23072 20596
rect 23388 20544 23440 20596
rect 24676 20587 24728 20596
rect 24676 20553 24685 20587
rect 24685 20553 24719 20587
rect 24719 20553 24728 20587
rect 24676 20544 24728 20553
rect 25596 20544 25648 20596
rect 18236 20519 18288 20528
rect 18236 20485 18245 20519
rect 18245 20485 18279 20519
rect 18279 20485 18288 20519
rect 18236 20476 18288 20485
rect 21824 20408 21876 20460
rect 23388 20408 23440 20460
rect 24308 20451 24360 20460
rect 24308 20417 24317 20451
rect 24317 20417 24351 20451
rect 24351 20417 24360 20451
rect 24860 20476 24912 20528
rect 26332 20544 26384 20596
rect 24308 20408 24360 20417
rect 2320 20340 2372 20392
rect 3240 20340 3292 20392
rect 4712 20340 4764 20392
rect 5448 20340 5500 20392
rect 6552 20340 6604 20392
rect 6828 20383 6880 20392
rect 6828 20349 6837 20383
rect 6837 20349 6871 20383
rect 6871 20349 6880 20383
rect 6828 20340 6880 20349
rect 12440 20383 12492 20392
rect 12440 20349 12449 20383
rect 12449 20349 12483 20383
rect 12483 20349 12492 20383
rect 13268 20383 13320 20392
rect 12440 20340 12492 20349
rect 13268 20349 13277 20383
rect 13277 20349 13311 20383
rect 13311 20349 13320 20383
rect 13268 20340 13320 20349
rect 14280 20340 14332 20392
rect 16672 20383 16724 20392
rect 16672 20349 16681 20383
rect 16681 20349 16715 20383
rect 16715 20349 16724 20383
rect 16672 20340 16724 20349
rect 17868 20340 17920 20392
rect 2412 20272 2464 20324
rect 4528 20247 4580 20256
rect 4528 20213 4537 20247
rect 4537 20213 4571 20247
rect 4571 20213 4580 20247
rect 4528 20204 4580 20213
rect 5172 20247 5224 20256
rect 5172 20213 5181 20247
rect 5181 20213 5215 20247
rect 5215 20213 5224 20247
rect 5172 20204 5224 20213
rect 8208 20272 8260 20324
rect 14004 20315 14056 20324
rect 14004 20281 14038 20315
rect 14038 20281 14056 20315
rect 14004 20272 14056 20281
rect 5540 20204 5592 20256
rect 7840 20204 7892 20256
rect 9128 20204 9180 20256
rect 9772 20204 9824 20256
rect 12992 20204 13044 20256
rect 13176 20204 13228 20256
rect 16212 20247 16264 20256
rect 16212 20213 16221 20247
rect 16221 20213 16255 20247
rect 16255 20213 16264 20247
rect 16212 20204 16264 20213
rect 16396 20272 16448 20324
rect 18144 20340 18196 20392
rect 19248 20340 19300 20392
rect 19524 20272 19576 20324
rect 20536 20272 20588 20324
rect 19340 20204 19392 20256
rect 21640 20340 21692 20392
rect 21364 20272 21416 20324
rect 23572 20340 23624 20392
rect 23940 20340 23992 20392
rect 25228 20383 25280 20392
rect 25228 20349 25237 20383
rect 25237 20349 25271 20383
rect 25271 20349 25280 20383
rect 25228 20340 25280 20349
rect 22192 20272 22244 20324
rect 21640 20247 21692 20256
rect 21640 20213 21649 20247
rect 21649 20213 21683 20247
rect 21683 20213 21692 20247
rect 21640 20204 21692 20213
rect 23020 20247 23072 20256
rect 23020 20213 23029 20247
rect 23029 20213 23063 20247
rect 23063 20213 23072 20247
rect 23020 20204 23072 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 2228 20043 2280 20052
rect 2228 20009 2237 20043
rect 2237 20009 2271 20043
rect 2271 20009 2280 20043
rect 2228 20000 2280 20009
rect 2964 20043 3016 20052
rect 2964 20009 2973 20043
rect 2973 20009 3007 20043
rect 3007 20009 3016 20043
rect 2964 20000 3016 20009
rect 4436 20000 4488 20052
rect 8116 20043 8168 20052
rect 8116 20009 8125 20043
rect 8125 20009 8159 20043
rect 8159 20009 8168 20043
rect 8116 20000 8168 20009
rect 10968 20000 11020 20052
rect 12256 20000 12308 20052
rect 13452 20000 13504 20052
rect 13728 20043 13780 20052
rect 13728 20009 13737 20043
rect 13737 20009 13771 20043
rect 13771 20009 13780 20043
rect 13728 20000 13780 20009
rect 13820 20000 13872 20052
rect 14464 20043 14516 20052
rect 14464 20009 14473 20043
rect 14473 20009 14507 20043
rect 14507 20009 14516 20043
rect 14464 20000 14516 20009
rect 15384 20000 15436 20052
rect 15936 20000 15988 20052
rect 16672 20043 16724 20052
rect 16672 20009 16681 20043
rect 16681 20009 16715 20043
rect 16715 20009 16724 20043
rect 16672 20000 16724 20009
rect 17592 20043 17644 20052
rect 17592 20009 17601 20043
rect 17601 20009 17635 20043
rect 17635 20009 17644 20043
rect 17592 20000 17644 20009
rect 19524 20000 19576 20052
rect 20168 20000 20220 20052
rect 23020 20000 23072 20052
rect 24308 20043 24360 20052
rect 24308 20009 24317 20043
rect 24317 20009 24351 20043
rect 24351 20009 24360 20043
rect 24308 20000 24360 20009
rect 4528 19932 4580 19984
rect 7656 19932 7708 19984
rect 12440 19975 12492 19984
rect 12440 19941 12449 19975
rect 12449 19941 12483 19975
rect 12483 19941 12492 19975
rect 12440 19932 12492 19941
rect 1768 19864 1820 19916
rect 3516 19864 3568 19916
rect 6368 19864 6420 19916
rect 6552 19864 6604 19916
rect 9220 19864 9272 19916
rect 9680 19864 9732 19916
rect 11244 19864 11296 19916
rect 12256 19864 12308 19916
rect 14556 19932 14608 19984
rect 15476 19932 15528 19984
rect 16488 19932 16540 19984
rect 22008 19932 22060 19984
rect 22100 19932 22152 19984
rect 2412 19839 2464 19848
rect 2412 19805 2421 19839
rect 2421 19805 2455 19839
rect 2455 19805 2464 19839
rect 2412 19796 2464 19805
rect 4344 19796 4396 19848
rect 6644 19796 6696 19848
rect 7564 19839 7616 19848
rect 7012 19771 7064 19780
rect 7012 19737 7021 19771
rect 7021 19737 7055 19771
rect 7055 19737 7064 19771
rect 7012 19728 7064 19737
rect 7564 19805 7573 19839
rect 7573 19805 7607 19839
rect 7607 19805 7616 19839
rect 7564 19796 7616 19805
rect 8944 19796 8996 19848
rect 10048 19796 10100 19848
rect 12072 19796 12124 19848
rect 14096 19864 14148 19916
rect 15752 19864 15804 19916
rect 16212 19864 16264 19916
rect 17408 19864 17460 19916
rect 19156 19864 19208 19916
rect 24768 19907 24820 19916
rect 24768 19873 24777 19907
rect 24777 19873 24811 19907
rect 24811 19873 24820 19907
rect 24768 19864 24820 19873
rect 13360 19839 13412 19848
rect 13360 19805 13369 19839
rect 13369 19805 13403 19839
rect 13403 19805 13412 19839
rect 13360 19796 13412 19805
rect 14004 19796 14056 19848
rect 16672 19796 16724 19848
rect 17316 19796 17368 19848
rect 18144 19796 18196 19848
rect 21088 19796 21140 19848
rect 24860 19839 24912 19848
rect 24860 19805 24869 19839
rect 24869 19805 24903 19839
rect 24903 19805 24912 19839
rect 24860 19796 24912 19805
rect 22928 19728 22980 19780
rect 23480 19728 23532 19780
rect 24676 19728 24728 19780
rect 2228 19660 2280 19712
rect 6000 19703 6052 19712
rect 6000 19669 6009 19703
rect 6009 19669 6043 19703
rect 6043 19669 6052 19703
rect 6000 19660 6052 19669
rect 6552 19703 6604 19712
rect 6552 19669 6561 19703
rect 6561 19669 6595 19703
rect 6595 19669 6604 19703
rect 6552 19660 6604 19669
rect 7104 19703 7156 19712
rect 7104 19669 7113 19703
rect 7113 19669 7147 19703
rect 7147 19669 7156 19703
rect 7104 19660 7156 19669
rect 9036 19703 9088 19712
rect 9036 19669 9045 19703
rect 9045 19669 9079 19703
rect 9079 19669 9088 19703
rect 9036 19660 9088 19669
rect 9312 19703 9364 19712
rect 9312 19669 9321 19703
rect 9321 19669 9355 19703
rect 9355 19669 9364 19703
rect 9312 19660 9364 19669
rect 10140 19660 10192 19712
rect 11336 19660 11388 19712
rect 14096 19703 14148 19712
rect 14096 19669 14105 19703
rect 14105 19669 14139 19703
rect 14139 19669 14148 19703
rect 14096 19660 14148 19669
rect 14280 19660 14332 19712
rect 18972 19660 19024 19712
rect 20720 19660 20772 19712
rect 21364 19660 21416 19712
rect 23940 19703 23992 19712
rect 23940 19669 23949 19703
rect 23949 19669 23983 19703
rect 23983 19669 23992 19703
rect 23940 19660 23992 19669
rect 25228 19660 25280 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1860 19499 1912 19508
rect 1860 19465 1869 19499
rect 1869 19465 1903 19499
rect 1903 19465 1912 19499
rect 1860 19456 1912 19465
rect 4528 19456 4580 19508
rect 6092 19456 6144 19508
rect 9404 19456 9456 19508
rect 9680 19499 9732 19508
rect 9680 19465 9689 19499
rect 9689 19465 9723 19499
rect 9723 19465 9732 19499
rect 9680 19456 9732 19465
rect 11796 19456 11848 19508
rect 12072 19456 12124 19508
rect 15936 19456 15988 19508
rect 17408 19499 17460 19508
rect 17408 19465 17417 19499
rect 17417 19465 17451 19499
rect 17451 19465 17460 19499
rect 17408 19456 17460 19465
rect 3608 19388 3660 19440
rect 7288 19388 7340 19440
rect 9220 19388 9272 19440
rect 9496 19388 9548 19440
rect 12256 19388 12308 19440
rect 13360 19388 13412 19440
rect 7012 19320 7064 19372
rect 7472 19320 7524 19372
rect 8760 19320 8812 19372
rect 8852 19320 8904 19372
rect 9036 19320 9088 19372
rect 9588 19320 9640 19372
rect 9956 19320 10008 19372
rect 2320 19295 2372 19304
rect 2320 19261 2329 19295
rect 2329 19261 2363 19295
rect 2363 19261 2372 19295
rect 2320 19252 2372 19261
rect 2412 19252 2464 19304
rect 2596 19252 2648 19304
rect 4160 19252 4212 19304
rect 6184 19295 6236 19304
rect 6184 19261 6193 19295
rect 6193 19261 6227 19295
rect 6227 19261 6236 19295
rect 6184 19252 6236 19261
rect 7104 19252 7156 19304
rect 12072 19252 12124 19304
rect 13452 19363 13504 19372
rect 13452 19329 13461 19363
rect 13461 19329 13495 19363
rect 13495 19329 13504 19363
rect 13452 19320 13504 19329
rect 16120 19388 16172 19440
rect 19156 19431 19208 19440
rect 14556 19320 14608 19372
rect 16488 19363 16540 19372
rect 16488 19329 16497 19363
rect 16497 19329 16531 19363
rect 16531 19329 16540 19363
rect 16488 19320 16540 19329
rect 19156 19397 19165 19431
rect 19165 19397 19199 19431
rect 19199 19397 19208 19431
rect 19156 19388 19208 19397
rect 24584 19388 24636 19440
rect 24860 19388 24912 19440
rect 18972 19320 19024 19372
rect 14464 19252 14516 19304
rect 17132 19295 17184 19304
rect 17132 19261 17141 19295
rect 17141 19261 17175 19295
rect 17175 19261 17184 19295
rect 17132 19252 17184 19261
rect 19432 19252 19484 19304
rect 19616 19295 19668 19304
rect 19616 19261 19625 19295
rect 19625 19261 19659 19295
rect 19659 19261 19668 19295
rect 19616 19252 19668 19261
rect 21088 19295 21140 19304
rect 21088 19261 21097 19295
rect 21097 19261 21131 19295
rect 21131 19261 21140 19295
rect 21088 19252 21140 19261
rect 22928 19320 22980 19372
rect 23940 19320 23992 19372
rect 24676 19320 24728 19372
rect 23480 19295 23532 19304
rect 2228 19227 2280 19236
rect 2228 19193 2237 19227
rect 2237 19193 2271 19227
rect 2271 19193 2280 19227
rect 2228 19184 2280 19193
rect 4528 19227 4580 19236
rect 4528 19193 4562 19227
rect 4562 19193 4580 19227
rect 4528 19184 4580 19193
rect 12440 19184 12492 19236
rect 13544 19184 13596 19236
rect 17684 19184 17736 19236
rect 18512 19227 18564 19236
rect 18512 19193 18521 19227
rect 18521 19193 18555 19227
rect 18555 19193 18564 19227
rect 18512 19184 18564 19193
rect 23480 19261 23489 19295
rect 23489 19261 23523 19295
rect 23523 19261 23532 19295
rect 25228 19295 25280 19304
rect 23480 19252 23532 19261
rect 21732 19184 21784 19236
rect 1860 19116 1912 19168
rect 6552 19159 6604 19168
rect 6552 19125 6561 19159
rect 6561 19125 6595 19159
rect 6595 19125 6604 19159
rect 6552 19116 6604 19125
rect 6736 19116 6788 19168
rect 7748 19116 7800 19168
rect 8576 19159 8628 19168
rect 8576 19125 8585 19159
rect 8585 19125 8619 19159
rect 8619 19125 8628 19159
rect 8576 19116 8628 19125
rect 8944 19159 8996 19168
rect 8944 19125 8953 19159
rect 8953 19125 8987 19159
rect 8987 19125 8996 19159
rect 8944 19116 8996 19125
rect 9036 19159 9088 19168
rect 9036 19125 9045 19159
rect 9045 19125 9079 19159
rect 9079 19125 9088 19159
rect 9036 19116 9088 19125
rect 10048 19116 10100 19168
rect 10968 19116 11020 19168
rect 12808 19116 12860 19168
rect 13912 19159 13964 19168
rect 13912 19125 13921 19159
rect 13921 19125 13955 19159
rect 13955 19125 13964 19159
rect 13912 19116 13964 19125
rect 14464 19159 14516 19168
rect 14464 19125 14473 19159
rect 14473 19125 14507 19159
rect 14507 19125 14516 19159
rect 14464 19116 14516 19125
rect 14832 19159 14884 19168
rect 14832 19125 14841 19159
rect 14841 19125 14875 19159
rect 14875 19125 14884 19159
rect 14832 19116 14884 19125
rect 15752 19116 15804 19168
rect 16304 19116 16356 19168
rect 16856 19116 16908 19168
rect 18052 19159 18104 19168
rect 18052 19125 18061 19159
rect 18061 19125 18095 19159
rect 18095 19125 18104 19159
rect 18052 19116 18104 19125
rect 18420 19159 18472 19168
rect 18420 19125 18429 19159
rect 18429 19125 18463 19159
rect 18463 19125 18472 19159
rect 18420 19116 18472 19125
rect 20168 19116 20220 19168
rect 22468 19159 22520 19168
rect 22468 19125 22477 19159
rect 22477 19125 22511 19159
rect 22511 19125 22520 19159
rect 22468 19116 22520 19125
rect 23664 19159 23716 19168
rect 23664 19125 23673 19159
rect 23673 19125 23707 19159
rect 23707 19125 23716 19159
rect 23664 19116 23716 19125
rect 25228 19261 25237 19295
rect 25237 19261 25271 19295
rect 25271 19261 25280 19295
rect 25228 19252 25280 19261
rect 24308 19116 24360 19168
rect 24584 19116 24636 19168
rect 24768 19116 24820 19168
rect 25228 19116 25280 19168
rect 25504 19116 25556 19168
rect 26148 19159 26200 19168
rect 26148 19125 26157 19159
rect 26157 19125 26191 19159
rect 26191 19125 26200 19159
rect 26148 19116 26200 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 2320 18912 2372 18964
rect 2504 18955 2556 18964
rect 2504 18921 2513 18955
rect 2513 18921 2547 18955
rect 2547 18921 2556 18955
rect 2504 18912 2556 18921
rect 4528 18912 4580 18964
rect 5356 18912 5408 18964
rect 6828 18912 6880 18964
rect 7104 18912 7156 18964
rect 8484 18955 8536 18964
rect 8484 18921 8493 18955
rect 8493 18921 8527 18955
rect 8527 18921 8536 18955
rect 8484 18912 8536 18921
rect 8668 18912 8720 18964
rect 9588 18912 9640 18964
rect 9680 18912 9732 18964
rect 11244 18912 11296 18964
rect 11796 18912 11848 18964
rect 12072 18912 12124 18964
rect 12900 18912 12952 18964
rect 15568 18912 15620 18964
rect 16120 18912 16172 18964
rect 17868 18912 17920 18964
rect 18420 18912 18472 18964
rect 18604 18912 18656 18964
rect 19064 18912 19116 18964
rect 19340 18912 19392 18964
rect 21088 18912 21140 18964
rect 21180 18912 21232 18964
rect 22008 18955 22060 18964
rect 22008 18921 22017 18955
rect 22017 18921 22051 18955
rect 22051 18921 22060 18955
rect 22008 18912 22060 18921
rect 23296 18912 23348 18964
rect 25136 18912 25188 18964
rect 2136 18844 2188 18896
rect 3608 18844 3660 18896
rect 4160 18844 4212 18896
rect 2412 18819 2464 18828
rect 2412 18785 2421 18819
rect 2421 18785 2455 18819
rect 2455 18785 2464 18819
rect 2412 18776 2464 18785
rect 6368 18844 6420 18896
rect 5264 18776 5316 18828
rect 6552 18776 6604 18828
rect 7564 18844 7616 18896
rect 8116 18844 8168 18896
rect 9404 18844 9456 18896
rect 10140 18844 10192 18896
rect 12256 18844 12308 18896
rect 8852 18776 8904 18828
rect 9312 18776 9364 18828
rect 14740 18844 14792 18896
rect 16856 18844 16908 18896
rect 18512 18844 18564 18896
rect 2596 18751 2648 18760
rect 2596 18717 2605 18751
rect 2605 18717 2639 18751
rect 2639 18717 2648 18751
rect 2596 18708 2648 18717
rect 2780 18708 2832 18760
rect 9220 18708 9272 18760
rect 13176 18708 13228 18760
rect 13268 18708 13320 18760
rect 14832 18708 14884 18760
rect 2136 18640 2188 18692
rect 3608 18640 3660 18692
rect 16580 18776 16632 18828
rect 17868 18776 17920 18828
rect 19892 18819 19944 18828
rect 16028 18708 16080 18760
rect 17500 18751 17552 18760
rect 17500 18717 17509 18751
rect 17509 18717 17543 18751
rect 17543 18717 17552 18751
rect 17500 18708 17552 18717
rect 17776 18708 17828 18760
rect 19892 18785 19901 18819
rect 19901 18785 19935 18819
rect 19935 18785 19944 18819
rect 19892 18776 19944 18785
rect 20168 18776 20220 18828
rect 23572 18844 23624 18896
rect 21364 18819 21416 18828
rect 18972 18708 19024 18760
rect 21364 18785 21373 18819
rect 21373 18785 21407 18819
rect 21407 18785 21416 18819
rect 21364 18776 21416 18785
rect 21732 18776 21784 18828
rect 22560 18819 22612 18828
rect 22560 18785 22569 18819
rect 22569 18785 22603 18819
rect 22603 18785 22612 18819
rect 22560 18776 22612 18785
rect 23756 18776 23808 18828
rect 23940 18819 23992 18828
rect 23940 18785 23974 18819
rect 23974 18785 23992 18819
rect 23940 18776 23992 18785
rect 20904 18708 20956 18760
rect 20996 18708 21048 18760
rect 20812 18640 20864 18692
rect 23296 18708 23348 18760
rect 2688 18572 2740 18624
rect 8024 18615 8076 18624
rect 8024 18581 8033 18615
rect 8033 18581 8067 18615
rect 8067 18581 8076 18615
rect 8024 18572 8076 18581
rect 9312 18615 9364 18624
rect 9312 18581 9321 18615
rect 9321 18581 9355 18615
rect 9355 18581 9364 18615
rect 9312 18572 9364 18581
rect 9496 18572 9548 18624
rect 10968 18572 11020 18624
rect 11336 18572 11388 18624
rect 12716 18572 12768 18624
rect 14556 18615 14608 18624
rect 14556 18581 14565 18615
rect 14565 18581 14599 18615
rect 14599 18581 14608 18615
rect 14556 18572 14608 18581
rect 18420 18572 18472 18624
rect 20904 18615 20956 18624
rect 20904 18581 20913 18615
rect 20913 18581 20947 18615
rect 20947 18581 20956 18615
rect 20904 18572 20956 18581
rect 22100 18572 22152 18624
rect 23020 18572 23072 18624
rect 24768 18572 24820 18624
rect 26148 18572 26200 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 2504 18368 2556 18420
rect 4712 18411 4764 18420
rect 4712 18377 4721 18411
rect 4721 18377 4755 18411
rect 4755 18377 4764 18411
rect 4712 18368 4764 18377
rect 5540 18368 5592 18420
rect 2136 18275 2188 18284
rect 2136 18241 2145 18275
rect 2145 18241 2179 18275
rect 2179 18241 2188 18275
rect 2136 18232 2188 18241
rect 5356 18275 5408 18284
rect 5356 18241 5365 18275
rect 5365 18241 5399 18275
rect 5399 18241 5408 18275
rect 5356 18232 5408 18241
rect 5264 18164 5316 18216
rect 7196 18368 7248 18420
rect 8484 18368 8536 18420
rect 8668 18368 8720 18420
rect 9588 18368 9640 18420
rect 9680 18411 9732 18420
rect 9680 18377 9689 18411
rect 9689 18377 9723 18411
rect 9723 18377 9732 18411
rect 9680 18368 9732 18377
rect 10140 18368 10192 18420
rect 12256 18411 12308 18420
rect 12256 18377 12265 18411
rect 12265 18377 12299 18411
rect 12299 18377 12308 18411
rect 12256 18368 12308 18377
rect 13820 18411 13872 18420
rect 8116 18343 8168 18352
rect 8116 18309 8125 18343
rect 8125 18309 8159 18343
rect 8159 18309 8168 18343
rect 8116 18300 8168 18309
rect 13820 18377 13829 18411
rect 13829 18377 13863 18411
rect 13863 18377 13872 18411
rect 13820 18368 13872 18377
rect 15568 18368 15620 18420
rect 16672 18368 16724 18420
rect 17500 18368 17552 18420
rect 19064 18411 19116 18420
rect 19064 18377 19073 18411
rect 19073 18377 19107 18411
rect 19107 18377 19116 18411
rect 19064 18368 19116 18377
rect 20996 18411 21048 18420
rect 8852 18164 8904 18216
rect 9036 18164 9088 18216
rect 11060 18232 11112 18284
rect 10692 18207 10744 18216
rect 10692 18173 10701 18207
rect 10701 18173 10735 18207
rect 10735 18173 10744 18207
rect 10692 18164 10744 18173
rect 11980 18164 12032 18216
rect 12256 18164 12308 18216
rect 14740 18232 14792 18284
rect 18052 18232 18104 18284
rect 2044 18096 2096 18148
rect 5080 18139 5132 18148
rect 5080 18105 5089 18139
rect 5089 18105 5123 18139
rect 5123 18105 5132 18139
rect 5080 18096 5132 18105
rect 2596 18028 2648 18080
rect 2872 18028 2924 18080
rect 4068 18028 4120 18080
rect 4988 18028 5040 18080
rect 6828 18028 6880 18080
rect 9220 18096 9272 18148
rect 11244 18139 11296 18148
rect 8392 18028 8444 18080
rect 10784 18071 10836 18080
rect 10784 18037 10793 18071
rect 10793 18037 10827 18071
rect 10827 18037 10836 18071
rect 10784 18028 10836 18037
rect 11244 18105 11253 18139
rect 11253 18105 11287 18139
rect 11287 18105 11296 18139
rect 11244 18096 11296 18105
rect 14280 18164 14332 18216
rect 14924 18207 14976 18216
rect 14924 18173 14933 18207
rect 14933 18173 14967 18207
rect 14967 18173 14976 18207
rect 14924 18164 14976 18173
rect 17776 18207 17828 18216
rect 17776 18173 17785 18207
rect 17785 18173 17819 18207
rect 17819 18173 17828 18207
rect 17776 18164 17828 18173
rect 18420 18207 18472 18216
rect 18420 18173 18429 18207
rect 18429 18173 18463 18207
rect 18463 18173 18472 18207
rect 18420 18164 18472 18173
rect 18604 18275 18656 18284
rect 18604 18241 18613 18275
rect 18613 18241 18647 18275
rect 18647 18241 18656 18275
rect 20996 18377 21005 18411
rect 21005 18377 21039 18411
rect 21039 18377 21048 18411
rect 20996 18368 21048 18377
rect 21180 18368 21232 18420
rect 22560 18411 22612 18420
rect 22560 18377 22569 18411
rect 22569 18377 22603 18411
rect 22603 18377 22612 18411
rect 22560 18368 22612 18377
rect 23940 18368 23992 18420
rect 20720 18300 20772 18352
rect 18604 18232 18656 18241
rect 20812 18232 20864 18284
rect 20904 18232 20956 18284
rect 22100 18275 22152 18284
rect 22100 18241 22109 18275
rect 22109 18241 22143 18275
rect 22143 18241 22152 18275
rect 22100 18232 22152 18241
rect 23572 18232 23624 18284
rect 19248 18164 19300 18216
rect 19892 18164 19944 18216
rect 21456 18164 21508 18216
rect 22560 18164 22612 18216
rect 24768 18164 24820 18216
rect 12716 18139 12768 18148
rect 12716 18105 12750 18139
rect 12750 18105 12768 18139
rect 12716 18096 12768 18105
rect 14556 18096 14608 18148
rect 15384 18096 15436 18148
rect 16028 18028 16080 18080
rect 17684 18028 17736 18080
rect 17868 18028 17920 18080
rect 22100 18096 22152 18148
rect 23940 18139 23992 18148
rect 23940 18105 23974 18139
rect 23974 18105 23992 18139
rect 23940 18096 23992 18105
rect 24032 18028 24084 18080
rect 25412 18028 25464 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1676 17824 1728 17876
rect 2688 17824 2740 17876
rect 2780 17867 2832 17876
rect 2780 17833 2789 17867
rect 2789 17833 2823 17867
rect 2823 17833 2832 17867
rect 2780 17824 2832 17833
rect 6368 17867 6420 17876
rect 6368 17833 6377 17867
rect 6377 17833 6411 17867
rect 6411 17833 6420 17867
rect 6368 17824 6420 17833
rect 6736 17867 6788 17876
rect 6736 17833 6745 17867
rect 6745 17833 6779 17867
rect 6779 17833 6788 17867
rect 6736 17824 6788 17833
rect 8024 17824 8076 17876
rect 9864 17824 9916 17876
rect 12900 17867 12952 17876
rect 1308 17756 1360 17808
rect 9036 17756 9088 17808
rect 12900 17833 12909 17867
rect 12909 17833 12943 17867
rect 12943 17833 12952 17867
rect 12900 17824 12952 17833
rect 13820 17824 13872 17876
rect 14280 17824 14332 17876
rect 14740 17824 14792 17876
rect 15292 17867 15344 17876
rect 15292 17833 15301 17867
rect 15301 17833 15335 17867
rect 15335 17833 15344 17867
rect 15292 17824 15344 17833
rect 15660 17824 15712 17876
rect 16580 17867 16632 17876
rect 16580 17833 16589 17867
rect 16589 17833 16623 17867
rect 16623 17833 16632 17867
rect 16580 17824 16632 17833
rect 17868 17824 17920 17876
rect 19340 17867 19392 17876
rect 19340 17833 19349 17867
rect 19349 17833 19383 17867
rect 19383 17833 19392 17867
rect 19340 17824 19392 17833
rect 20076 17824 20128 17876
rect 20444 17824 20496 17876
rect 22100 17824 22152 17876
rect 24860 17867 24912 17876
rect 24860 17833 24869 17867
rect 24869 17833 24903 17867
rect 24903 17833 24912 17867
rect 24860 17824 24912 17833
rect 12348 17756 12400 17808
rect 14004 17756 14056 17808
rect 17408 17756 17460 17808
rect 18972 17799 19024 17808
rect 18972 17765 18981 17799
rect 18981 17765 19015 17799
rect 19015 17765 19024 17799
rect 18972 17756 19024 17765
rect 19984 17756 20036 17808
rect 20536 17756 20588 17808
rect 25044 17756 25096 17808
rect 2044 17688 2096 17740
rect 2688 17688 2740 17740
rect 3608 17688 3660 17740
rect 4160 17688 4212 17740
rect 6644 17688 6696 17740
rect 8392 17731 8444 17740
rect 8392 17697 8401 17731
rect 8401 17697 8435 17731
rect 8435 17697 8444 17731
rect 8392 17688 8444 17697
rect 9496 17688 9548 17740
rect 10692 17688 10744 17740
rect 2320 17663 2372 17672
rect 2320 17629 2329 17663
rect 2329 17629 2363 17663
rect 2363 17629 2372 17663
rect 2320 17620 2372 17629
rect 2872 17620 2924 17672
rect 8208 17620 8260 17672
rect 8668 17663 8720 17672
rect 8668 17629 8677 17663
rect 8677 17629 8711 17663
rect 8711 17629 8720 17663
rect 8668 17620 8720 17629
rect 9956 17663 10008 17672
rect 9956 17629 9965 17663
rect 9965 17629 9999 17663
rect 9999 17629 10008 17663
rect 9956 17620 10008 17629
rect 10600 17620 10652 17672
rect 11060 17688 11112 17740
rect 13728 17688 13780 17740
rect 14556 17688 14608 17740
rect 15752 17731 15804 17740
rect 15752 17697 15761 17731
rect 15761 17697 15795 17731
rect 15795 17697 15804 17731
rect 19524 17731 19576 17740
rect 15752 17688 15804 17697
rect 19524 17697 19533 17731
rect 19533 17697 19567 17731
rect 19567 17697 19576 17731
rect 19524 17688 19576 17697
rect 20812 17688 20864 17740
rect 24032 17688 24084 17740
rect 8024 17595 8076 17604
rect 8024 17561 8033 17595
rect 8033 17561 8067 17595
rect 8067 17561 8076 17595
rect 8024 17552 8076 17561
rect 8852 17552 8904 17604
rect 12440 17620 12492 17672
rect 12716 17552 12768 17604
rect 13360 17552 13412 17604
rect 14188 17620 14240 17672
rect 14740 17620 14792 17672
rect 14924 17620 14976 17672
rect 15936 17663 15988 17672
rect 15936 17629 15945 17663
rect 15945 17629 15979 17663
rect 15979 17629 15988 17663
rect 15936 17620 15988 17629
rect 19984 17620 20036 17672
rect 20536 17552 20588 17604
rect 22744 17620 22796 17672
rect 23572 17620 23624 17672
rect 23940 17663 23992 17672
rect 23940 17629 23949 17663
rect 23949 17629 23983 17663
rect 23983 17629 23992 17663
rect 23940 17620 23992 17629
rect 1768 17527 1820 17536
rect 1768 17493 1777 17527
rect 1777 17493 1811 17527
rect 1811 17493 1820 17527
rect 1768 17484 1820 17493
rect 3148 17527 3200 17536
rect 3148 17493 3157 17527
rect 3157 17493 3191 17527
rect 3191 17493 3200 17527
rect 3148 17484 3200 17493
rect 5264 17484 5316 17536
rect 9220 17484 9272 17536
rect 10968 17484 11020 17536
rect 12256 17484 12308 17536
rect 12440 17484 12492 17536
rect 13268 17527 13320 17536
rect 13268 17493 13277 17527
rect 13277 17493 13311 17527
rect 13311 17493 13320 17527
rect 13268 17484 13320 17493
rect 16120 17484 16172 17536
rect 17040 17484 17092 17536
rect 18420 17527 18472 17536
rect 18420 17493 18429 17527
rect 18429 17493 18463 17527
rect 18463 17493 18472 17527
rect 18420 17484 18472 17493
rect 20812 17484 20864 17536
rect 25688 17552 25740 17604
rect 21640 17484 21692 17536
rect 22192 17484 22244 17536
rect 23020 17484 23072 17536
rect 24676 17484 24728 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2320 17280 2372 17332
rect 4160 17323 4212 17332
rect 4160 17289 4169 17323
rect 4169 17289 4203 17323
rect 4203 17289 4212 17323
rect 4160 17280 4212 17289
rect 5080 17323 5132 17332
rect 5080 17289 5089 17323
rect 5089 17289 5123 17323
rect 5123 17289 5132 17323
rect 5080 17280 5132 17289
rect 8208 17280 8260 17332
rect 8392 17280 8444 17332
rect 5264 17144 5316 17196
rect 9588 17255 9640 17264
rect 9588 17221 9597 17255
rect 9597 17221 9631 17255
rect 9631 17221 9640 17255
rect 9588 17212 9640 17221
rect 14004 17280 14056 17332
rect 15384 17323 15436 17332
rect 15384 17289 15393 17323
rect 15393 17289 15427 17323
rect 15427 17289 15436 17323
rect 15384 17280 15436 17289
rect 15752 17280 15804 17332
rect 19432 17323 19484 17332
rect 19432 17289 19441 17323
rect 19441 17289 19475 17323
rect 19475 17289 19484 17323
rect 19432 17280 19484 17289
rect 20628 17280 20680 17332
rect 22744 17323 22796 17332
rect 22744 17289 22753 17323
rect 22753 17289 22787 17323
rect 22787 17289 22796 17323
rect 22744 17280 22796 17289
rect 23940 17280 23992 17332
rect 25688 17323 25740 17332
rect 25688 17289 25697 17323
rect 25697 17289 25731 17323
rect 25731 17289 25740 17323
rect 25688 17280 25740 17289
rect 26148 17323 26200 17332
rect 26148 17289 26157 17323
rect 26157 17289 26191 17323
rect 26191 17289 26200 17323
rect 26148 17280 26200 17289
rect 15936 17255 15988 17264
rect 2044 17076 2096 17128
rect 4436 17076 4488 17128
rect 6736 17076 6788 17128
rect 8208 17119 8260 17128
rect 8208 17085 8217 17119
rect 8217 17085 8251 17119
rect 8251 17085 8260 17119
rect 8208 17076 8260 17085
rect 9220 17144 9272 17196
rect 11336 17187 11388 17196
rect 11336 17153 11345 17187
rect 11345 17153 11379 17187
rect 11379 17153 11388 17187
rect 11336 17144 11388 17153
rect 15936 17221 15945 17255
rect 15945 17221 15979 17255
rect 15979 17221 15988 17255
rect 15936 17212 15988 17221
rect 12532 17144 12584 17196
rect 12900 17144 12952 17196
rect 13268 17144 13320 17196
rect 20536 17144 20588 17196
rect 12072 17076 12124 17128
rect 14280 17119 14332 17128
rect 14280 17085 14314 17119
rect 14314 17085 14332 17119
rect 2780 17008 2832 17060
rect 7104 17051 7156 17060
rect 7104 17017 7113 17051
rect 7113 17017 7147 17051
rect 7147 17017 7156 17051
rect 7104 17008 7156 17017
rect 14280 17076 14332 17085
rect 15200 17076 15252 17128
rect 16488 17119 16540 17128
rect 16488 17085 16497 17119
rect 16497 17085 16531 17119
rect 16531 17085 16540 17119
rect 16488 17076 16540 17085
rect 18144 17076 18196 17128
rect 20720 17076 20772 17128
rect 22192 17076 22244 17128
rect 14740 17008 14792 17060
rect 17592 17008 17644 17060
rect 3332 16983 3384 16992
rect 3332 16949 3341 16983
rect 3341 16949 3375 16983
rect 3375 16949 3384 16983
rect 3332 16940 3384 16949
rect 6184 16940 6236 16992
rect 6644 16983 6696 16992
rect 6644 16949 6653 16983
rect 6653 16949 6687 16983
rect 6687 16949 6696 16983
rect 6644 16940 6696 16949
rect 11060 16983 11112 16992
rect 11060 16949 11069 16983
rect 11069 16949 11103 16983
rect 11103 16949 11112 16983
rect 11060 16940 11112 16949
rect 12716 16940 12768 16992
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 13728 16940 13780 16992
rect 17408 16940 17460 16992
rect 17684 16940 17736 16992
rect 18420 17008 18472 17060
rect 20352 17008 20404 17060
rect 25228 17076 25280 17128
rect 24308 17008 24360 17060
rect 20812 16940 20864 16992
rect 21180 16940 21232 16992
rect 22008 16983 22060 16992
rect 22008 16949 22017 16983
rect 22017 16949 22051 16983
rect 22051 16949 22060 16983
rect 22008 16940 22060 16949
rect 24676 16940 24728 16992
rect 25228 16940 25280 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1676 16779 1728 16788
rect 1676 16745 1685 16779
rect 1685 16745 1719 16779
rect 1719 16745 1728 16779
rect 1676 16736 1728 16745
rect 3148 16736 3200 16788
rect 3516 16779 3568 16788
rect 3516 16745 3525 16779
rect 3525 16745 3559 16779
rect 3559 16745 3568 16779
rect 3516 16736 3568 16745
rect 3884 16736 3936 16788
rect 6736 16736 6788 16788
rect 7564 16779 7616 16788
rect 7564 16745 7573 16779
rect 7573 16745 7607 16779
rect 7607 16745 7616 16779
rect 7564 16736 7616 16745
rect 8668 16779 8720 16788
rect 8668 16745 8677 16779
rect 8677 16745 8711 16779
rect 8711 16745 8720 16779
rect 8668 16736 8720 16745
rect 9588 16736 9640 16788
rect 9864 16779 9916 16788
rect 9864 16745 9873 16779
rect 9873 16745 9907 16779
rect 9907 16745 9916 16779
rect 9864 16736 9916 16745
rect 10784 16736 10836 16788
rect 13636 16779 13688 16788
rect 13636 16745 13645 16779
rect 13645 16745 13679 16779
rect 13679 16745 13688 16779
rect 13636 16736 13688 16745
rect 14004 16779 14056 16788
rect 14004 16745 14013 16779
rect 14013 16745 14047 16779
rect 14047 16745 14056 16779
rect 14004 16736 14056 16745
rect 14096 16779 14148 16788
rect 14096 16745 14105 16779
rect 14105 16745 14139 16779
rect 14139 16745 14148 16779
rect 14096 16736 14148 16745
rect 14832 16736 14884 16788
rect 16488 16779 16540 16788
rect 16488 16745 16497 16779
rect 16497 16745 16531 16779
rect 16531 16745 16540 16779
rect 16488 16736 16540 16745
rect 20720 16779 20772 16788
rect 20720 16745 20729 16779
rect 20729 16745 20763 16779
rect 20763 16745 20772 16779
rect 20720 16736 20772 16745
rect 24032 16779 24084 16788
rect 24032 16745 24041 16779
rect 24041 16745 24075 16779
rect 24075 16745 24084 16779
rect 24032 16736 24084 16745
rect 9496 16711 9548 16720
rect 2044 16643 2096 16652
rect 2044 16609 2053 16643
rect 2053 16609 2087 16643
rect 2087 16609 2096 16643
rect 2044 16600 2096 16609
rect 2136 16643 2188 16652
rect 2136 16609 2145 16643
rect 2145 16609 2179 16643
rect 2179 16609 2188 16643
rect 2136 16600 2188 16609
rect 1952 16532 2004 16584
rect 2504 16600 2556 16652
rect 3332 16600 3384 16652
rect 5356 16643 5408 16652
rect 5356 16609 5390 16643
rect 5390 16609 5408 16643
rect 5356 16600 5408 16609
rect 2780 16575 2832 16584
rect 2780 16541 2789 16575
rect 2789 16541 2823 16575
rect 2823 16541 2832 16575
rect 2780 16532 2832 16541
rect 3884 16532 3936 16584
rect 4712 16396 4764 16448
rect 6092 16532 6144 16584
rect 9496 16677 9505 16711
rect 9505 16677 9539 16711
rect 9539 16677 9548 16711
rect 9496 16668 9548 16677
rect 11060 16668 11112 16720
rect 12164 16668 12216 16720
rect 14556 16668 14608 16720
rect 19432 16668 19484 16720
rect 19524 16668 19576 16720
rect 22008 16711 22060 16720
rect 22008 16677 22042 16711
rect 22042 16677 22060 16711
rect 22008 16668 22060 16677
rect 24676 16668 24728 16720
rect 7656 16600 7708 16652
rect 9404 16600 9456 16652
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 10968 16600 11020 16652
rect 11428 16643 11480 16652
rect 11428 16609 11462 16643
rect 11462 16609 11480 16643
rect 11428 16600 11480 16609
rect 7840 16532 7892 16584
rect 8116 16575 8168 16584
rect 8116 16541 8125 16575
rect 8125 16541 8159 16575
rect 8159 16541 8168 16575
rect 8116 16532 8168 16541
rect 15476 16600 15528 16652
rect 16580 16600 16632 16652
rect 6920 16464 6972 16516
rect 9036 16439 9088 16448
rect 9036 16405 9045 16439
rect 9045 16405 9079 16439
rect 9079 16405 9088 16439
rect 9036 16396 9088 16405
rect 12624 16396 12676 16448
rect 13268 16396 13320 16448
rect 13452 16439 13504 16448
rect 13452 16405 13461 16439
rect 13461 16405 13495 16439
rect 13495 16405 13504 16439
rect 13452 16396 13504 16405
rect 14188 16396 14240 16448
rect 15384 16532 15436 16584
rect 15568 16532 15620 16584
rect 15200 16464 15252 16516
rect 15936 16464 15988 16516
rect 17868 16600 17920 16652
rect 18512 16643 18564 16652
rect 18512 16609 18521 16643
rect 18521 16609 18555 16643
rect 18555 16609 18564 16643
rect 18512 16600 18564 16609
rect 23204 16600 23256 16652
rect 24860 16600 24912 16652
rect 17684 16532 17736 16584
rect 19156 16532 19208 16584
rect 20812 16532 20864 16584
rect 21088 16532 21140 16584
rect 21732 16575 21784 16584
rect 21732 16541 21741 16575
rect 21741 16541 21775 16575
rect 21775 16541 21784 16575
rect 21732 16532 21784 16541
rect 24032 16532 24084 16584
rect 20168 16464 20220 16516
rect 20536 16464 20588 16516
rect 24308 16464 24360 16516
rect 24952 16464 25004 16516
rect 14740 16396 14792 16448
rect 16856 16439 16908 16448
rect 16856 16405 16865 16439
rect 16865 16405 16899 16439
rect 16899 16405 16908 16439
rect 16856 16396 16908 16405
rect 18788 16439 18840 16448
rect 18788 16405 18797 16439
rect 18797 16405 18831 16439
rect 18831 16405 18840 16439
rect 18788 16396 18840 16405
rect 20076 16439 20128 16448
rect 20076 16405 20085 16439
rect 20085 16405 20119 16439
rect 20119 16405 20128 16439
rect 20076 16396 20128 16405
rect 21088 16439 21140 16448
rect 21088 16405 21097 16439
rect 21097 16405 21131 16439
rect 21131 16405 21140 16439
rect 21088 16396 21140 16405
rect 23112 16439 23164 16448
rect 23112 16405 23121 16439
rect 23121 16405 23155 16439
rect 23155 16405 23164 16439
rect 23112 16396 23164 16405
rect 23756 16396 23808 16448
rect 24216 16396 24268 16448
rect 24768 16396 24820 16448
rect 25228 16439 25280 16448
rect 25228 16405 25237 16439
rect 25237 16405 25271 16439
rect 25271 16405 25280 16439
rect 25228 16396 25280 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2504 16235 2556 16244
rect 2504 16201 2513 16235
rect 2513 16201 2547 16235
rect 2547 16201 2556 16235
rect 2504 16192 2556 16201
rect 2688 16235 2740 16244
rect 2688 16201 2697 16235
rect 2697 16201 2731 16235
rect 2731 16201 2740 16235
rect 2688 16192 2740 16201
rect 4620 16192 4672 16244
rect 4988 16235 5040 16244
rect 2780 16124 2832 16176
rect 3516 16124 3568 16176
rect 3332 16099 3384 16108
rect 3332 16065 3341 16099
rect 3341 16065 3375 16099
rect 3375 16065 3384 16099
rect 3332 16056 3384 16065
rect 4988 16201 4997 16235
rect 4997 16201 5031 16235
rect 5031 16201 5040 16235
rect 4988 16192 5040 16201
rect 7656 16235 7708 16244
rect 7656 16201 7665 16235
rect 7665 16201 7699 16235
rect 7699 16201 7708 16235
rect 7656 16192 7708 16201
rect 9680 16192 9732 16244
rect 14004 16192 14056 16244
rect 14648 16192 14700 16244
rect 15936 16235 15988 16244
rect 15936 16201 15945 16235
rect 15945 16201 15979 16235
rect 15979 16201 15988 16235
rect 15936 16192 15988 16201
rect 19524 16192 19576 16244
rect 7012 16167 7064 16176
rect 7012 16133 7021 16167
rect 7021 16133 7055 16167
rect 7055 16133 7064 16167
rect 7012 16124 7064 16133
rect 14740 16167 14792 16176
rect 14740 16133 14749 16167
rect 14749 16133 14783 16167
rect 14783 16133 14792 16167
rect 14740 16124 14792 16133
rect 6092 16099 6144 16108
rect 1676 15963 1728 15972
rect 1676 15929 1685 15963
rect 1685 15929 1719 15963
rect 1719 15929 1728 15963
rect 1676 15920 1728 15929
rect 3332 15920 3384 15972
rect 5264 15988 5316 16040
rect 6092 16065 6101 16099
rect 6101 16065 6135 16099
rect 6135 16065 6144 16099
rect 6092 16056 6144 16065
rect 7196 16056 7248 16108
rect 10784 16056 10836 16108
rect 11428 16099 11480 16108
rect 11428 16065 11437 16099
rect 11437 16065 11471 16099
rect 11471 16065 11480 16099
rect 11428 16056 11480 16065
rect 11888 16056 11940 16108
rect 16028 16056 16080 16108
rect 16948 16099 17000 16108
rect 16948 16065 16957 16099
rect 16957 16065 16991 16099
rect 16991 16065 17000 16099
rect 16948 16056 17000 16065
rect 17408 16056 17460 16108
rect 18788 16056 18840 16108
rect 20076 16056 20128 16108
rect 22008 16192 22060 16244
rect 23112 16235 23164 16244
rect 21732 16167 21784 16176
rect 21732 16133 21741 16167
rect 21741 16133 21775 16167
rect 21775 16133 21784 16167
rect 21732 16124 21784 16133
rect 6828 16031 6880 16040
rect 6828 15997 6837 16031
rect 6837 15997 6871 16031
rect 6871 15997 6880 16031
rect 6828 15988 6880 15997
rect 3792 15895 3844 15904
rect 3792 15861 3801 15895
rect 3801 15861 3835 15895
rect 3835 15861 3844 15895
rect 3792 15852 3844 15861
rect 4252 15852 4304 15904
rect 7932 15920 7984 15972
rect 8668 15988 8720 16040
rect 10048 15988 10100 16040
rect 12348 15988 12400 16040
rect 12532 15988 12584 16040
rect 13544 15988 13596 16040
rect 16856 15988 16908 16040
rect 18052 15988 18104 16040
rect 20628 15988 20680 16040
rect 21732 15988 21784 16040
rect 22376 16056 22428 16108
rect 23112 16201 23121 16235
rect 23121 16201 23155 16235
rect 23155 16201 23164 16235
rect 23112 16192 23164 16201
rect 24032 16192 24084 16244
rect 24952 16192 25004 16244
rect 8208 15920 8260 15972
rect 9036 15920 9088 15972
rect 12624 15920 12676 15972
rect 14648 15920 14700 15972
rect 15476 15920 15528 15972
rect 21088 15920 21140 15972
rect 21456 15920 21508 15972
rect 21824 15920 21876 15972
rect 8576 15852 8628 15904
rect 10784 15895 10836 15904
rect 10784 15861 10793 15895
rect 10793 15861 10827 15895
rect 10827 15861 10836 15895
rect 10784 15852 10836 15861
rect 11888 15895 11940 15904
rect 11888 15861 11897 15895
rect 11897 15861 11931 15895
rect 11931 15861 11940 15895
rect 11888 15852 11940 15861
rect 13268 15852 13320 15904
rect 15384 15895 15436 15904
rect 15384 15861 15393 15895
rect 15393 15861 15427 15895
rect 15427 15861 15436 15895
rect 17408 15895 17460 15904
rect 15384 15852 15436 15861
rect 17408 15861 17417 15895
rect 17417 15861 17451 15895
rect 17451 15861 17460 15895
rect 17408 15852 17460 15861
rect 17776 15895 17828 15904
rect 17776 15861 17785 15895
rect 17785 15861 17819 15895
rect 17819 15861 17828 15895
rect 17776 15852 17828 15861
rect 17960 15852 18012 15904
rect 19156 15895 19208 15904
rect 19156 15861 19165 15895
rect 19165 15861 19199 15895
rect 19199 15861 19208 15895
rect 19156 15852 19208 15861
rect 19432 15895 19484 15904
rect 19432 15861 19441 15895
rect 19441 15861 19475 15895
rect 19475 15861 19484 15895
rect 19432 15852 19484 15861
rect 22008 15895 22060 15904
rect 22008 15861 22017 15895
rect 22017 15861 22051 15895
rect 22051 15861 22060 15895
rect 22008 15852 22060 15861
rect 23756 15988 23808 16040
rect 23940 15852 23992 15904
rect 25228 15852 25280 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2044 15648 2096 15700
rect 2412 15648 2464 15700
rect 2780 15691 2832 15700
rect 2780 15657 2789 15691
rect 2789 15657 2823 15691
rect 2823 15657 2832 15691
rect 2780 15648 2832 15657
rect 3240 15648 3292 15700
rect 7840 15648 7892 15700
rect 8300 15691 8352 15700
rect 8300 15657 8309 15691
rect 8309 15657 8343 15691
rect 8343 15657 8352 15691
rect 8300 15648 8352 15657
rect 8760 15648 8812 15700
rect 10048 15691 10100 15700
rect 10048 15657 10057 15691
rect 10057 15657 10091 15691
rect 10091 15657 10100 15691
rect 10048 15648 10100 15657
rect 6092 15580 6144 15632
rect 1768 15512 1820 15564
rect 1860 15512 1912 15564
rect 5448 15555 5500 15564
rect 5448 15521 5457 15555
rect 5457 15521 5491 15555
rect 5491 15521 5500 15555
rect 5448 15512 5500 15521
rect 1952 15444 2004 15496
rect 2228 15487 2280 15496
rect 2228 15453 2237 15487
rect 2237 15453 2271 15487
rect 2271 15453 2280 15487
rect 2228 15444 2280 15453
rect 2412 15487 2464 15496
rect 2412 15453 2421 15487
rect 2421 15453 2455 15487
rect 2455 15453 2464 15487
rect 2412 15444 2464 15453
rect 5172 15444 5224 15496
rect 5632 15487 5684 15496
rect 5632 15453 5641 15487
rect 5641 15453 5675 15487
rect 5675 15453 5684 15487
rect 5632 15444 5684 15453
rect 4712 15376 4764 15428
rect 5264 15376 5316 15428
rect 3240 15351 3292 15360
rect 3240 15317 3249 15351
rect 3249 15317 3283 15351
rect 3283 15317 3292 15351
rect 3240 15308 3292 15317
rect 3332 15308 3384 15360
rect 5080 15351 5132 15360
rect 5080 15317 5089 15351
rect 5089 15317 5123 15351
rect 5123 15317 5132 15351
rect 5080 15308 5132 15317
rect 8116 15580 8168 15632
rect 6644 15555 6696 15564
rect 6644 15521 6653 15555
rect 6653 15521 6687 15555
rect 6687 15521 6696 15555
rect 6644 15512 6696 15521
rect 7656 15512 7708 15564
rect 8668 15512 8720 15564
rect 9036 15555 9088 15564
rect 9036 15521 9045 15555
rect 9045 15521 9079 15555
rect 9079 15521 9088 15555
rect 9036 15512 9088 15521
rect 9404 15512 9456 15564
rect 10968 15648 11020 15700
rect 13452 15691 13504 15700
rect 13452 15657 13461 15691
rect 13461 15657 13495 15691
rect 13495 15657 13504 15691
rect 13452 15648 13504 15657
rect 13912 15648 13964 15700
rect 14096 15691 14148 15700
rect 14096 15657 14105 15691
rect 14105 15657 14139 15691
rect 14139 15657 14148 15691
rect 14096 15648 14148 15657
rect 17408 15648 17460 15700
rect 17684 15691 17736 15700
rect 17684 15657 17693 15691
rect 17693 15657 17727 15691
rect 17727 15657 17736 15691
rect 17684 15648 17736 15657
rect 21088 15648 21140 15700
rect 22100 15648 22152 15700
rect 23480 15691 23532 15700
rect 23480 15657 23489 15691
rect 23489 15657 23523 15691
rect 23523 15657 23532 15691
rect 23480 15648 23532 15657
rect 24952 15691 25004 15700
rect 24952 15657 24961 15691
rect 24961 15657 24995 15691
rect 24995 15657 25004 15691
rect 24952 15648 25004 15657
rect 10692 15580 10744 15632
rect 13084 15580 13136 15632
rect 18604 15580 18656 15632
rect 21364 15580 21416 15632
rect 21456 15580 21508 15632
rect 21732 15580 21784 15632
rect 24584 15623 24636 15632
rect 24584 15589 24593 15623
rect 24593 15589 24627 15623
rect 24627 15589 24636 15623
rect 24584 15580 24636 15589
rect 12532 15512 12584 15564
rect 13728 15512 13780 15564
rect 16028 15555 16080 15564
rect 16028 15521 16062 15555
rect 16062 15521 16080 15555
rect 16028 15512 16080 15521
rect 20904 15512 20956 15564
rect 22100 15512 22152 15564
rect 22468 15555 22520 15564
rect 22468 15521 22477 15555
rect 22477 15521 22511 15555
rect 22511 15521 22520 15555
rect 22468 15512 22520 15521
rect 23756 15512 23808 15564
rect 25136 15555 25188 15564
rect 25136 15521 25145 15555
rect 25145 15521 25179 15555
rect 25179 15521 25188 15555
rect 25136 15512 25188 15521
rect 8576 15487 8628 15496
rect 8576 15453 8585 15487
rect 8585 15453 8619 15487
rect 8619 15453 8628 15487
rect 8576 15444 8628 15453
rect 13544 15487 13596 15496
rect 13544 15453 13553 15487
rect 13553 15453 13587 15487
rect 13587 15453 13596 15487
rect 13544 15444 13596 15453
rect 15292 15444 15344 15496
rect 18144 15444 18196 15496
rect 21364 15487 21416 15496
rect 21364 15453 21373 15487
rect 21373 15453 21407 15487
rect 21407 15453 21416 15487
rect 21364 15444 21416 15453
rect 8116 15376 8168 15428
rect 19340 15376 19392 15428
rect 20720 15376 20772 15428
rect 21456 15376 21508 15428
rect 24676 15444 24728 15496
rect 24952 15444 25004 15496
rect 23572 15419 23624 15428
rect 23572 15385 23581 15419
rect 23581 15385 23615 15419
rect 23615 15385 23624 15419
rect 23572 15376 23624 15385
rect 24860 15376 24912 15428
rect 8576 15308 8628 15360
rect 8852 15308 8904 15360
rect 11888 15351 11940 15360
rect 11888 15317 11897 15351
rect 11897 15317 11931 15351
rect 11931 15317 11940 15351
rect 11888 15308 11940 15317
rect 12164 15308 12216 15360
rect 12624 15308 12676 15360
rect 13820 15308 13872 15360
rect 14096 15308 14148 15360
rect 14648 15308 14700 15360
rect 14740 15308 14792 15360
rect 15568 15308 15620 15360
rect 18052 15351 18104 15360
rect 18052 15317 18061 15351
rect 18061 15317 18095 15351
rect 18095 15317 18104 15351
rect 18052 15308 18104 15317
rect 19984 15308 20036 15360
rect 20628 15308 20680 15360
rect 22376 15308 22428 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2136 15104 2188 15156
rect 4436 15104 4488 15156
rect 4712 15104 4764 15156
rect 7656 15147 7708 15156
rect 7656 15113 7665 15147
rect 7665 15113 7699 15147
rect 7699 15113 7708 15147
rect 7656 15104 7708 15113
rect 7840 15104 7892 15156
rect 8208 15104 8260 15156
rect 12440 15147 12492 15156
rect 12440 15113 12449 15147
rect 12449 15113 12483 15147
rect 12483 15113 12492 15147
rect 13544 15147 13596 15156
rect 12440 15104 12492 15113
rect 13544 15113 13553 15147
rect 13553 15113 13587 15147
rect 13587 15113 13596 15147
rect 13544 15104 13596 15113
rect 13912 15147 13964 15156
rect 13912 15113 13921 15147
rect 13921 15113 13955 15147
rect 13955 15113 13964 15147
rect 13912 15104 13964 15113
rect 16028 15104 16080 15156
rect 17868 15104 17920 15156
rect 18604 15104 18656 15156
rect 21456 15104 21508 15156
rect 22468 15104 22520 15156
rect 22928 15104 22980 15156
rect 1768 14968 1820 15020
rect 2412 15036 2464 15088
rect 5356 15036 5408 15088
rect 10048 15079 10100 15088
rect 10048 15045 10057 15079
rect 10057 15045 10091 15079
rect 10091 15045 10100 15079
rect 10048 15036 10100 15045
rect 13728 15036 13780 15088
rect 17224 15036 17276 15088
rect 23848 15104 23900 15156
rect 24676 15147 24728 15156
rect 24676 15113 24685 15147
rect 24685 15113 24719 15147
rect 24719 15113 24728 15147
rect 24676 15104 24728 15113
rect 25320 15104 25372 15156
rect 23112 15036 23164 15088
rect 5264 14968 5316 15020
rect 11336 14968 11388 15020
rect 13084 15011 13136 15020
rect 13084 14977 13093 15011
rect 13093 14977 13127 15011
rect 13127 14977 13136 15011
rect 13084 14968 13136 14977
rect 18604 15011 18656 15020
rect 18604 14977 18613 15011
rect 18613 14977 18647 15011
rect 18647 14977 18656 15011
rect 18604 14968 18656 14977
rect 19248 14968 19300 15020
rect 3240 14900 3292 14952
rect 5540 14900 5592 14952
rect 2320 14764 2372 14816
rect 5264 14832 5316 14884
rect 7932 14900 7984 14952
rect 8116 14943 8168 14952
rect 8116 14909 8150 14943
rect 8150 14909 8168 14943
rect 8116 14900 8168 14909
rect 10508 14943 10560 14952
rect 10508 14909 10517 14943
rect 10517 14909 10551 14943
rect 10551 14909 10560 14943
rect 10508 14900 10560 14909
rect 11520 14900 11572 14952
rect 14832 14943 14884 14952
rect 14832 14909 14841 14943
rect 14841 14909 14875 14943
rect 14875 14909 14884 14943
rect 17868 14943 17920 14952
rect 14832 14900 14884 14909
rect 17868 14909 17877 14943
rect 17877 14909 17911 14943
rect 17911 14909 17920 14943
rect 17868 14900 17920 14909
rect 18420 14943 18472 14952
rect 18420 14909 18429 14943
rect 18429 14909 18463 14943
rect 18463 14909 18472 14943
rect 18420 14900 18472 14909
rect 21088 14900 21140 14952
rect 22284 14943 22336 14952
rect 22284 14909 22293 14943
rect 22293 14909 22327 14943
rect 22327 14909 22336 14943
rect 22284 14900 22336 14909
rect 23020 14900 23072 14952
rect 23664 14968 23716 15020
rect 24032 14943 24084 14952
rect 6644 14832 6696 14884
rect 9496 14832 9548 14884
rect 12440 14832 12492 14884
rect 12624 14832 12676 14884
rect 12992 14832 13044 14884
rect 15292 14832 15344 14884
rect 18512 14875 18564 14884
rect 3148 14764 3200 14816
rect 5172 14764 5224 14816
rect 5816 14807 5868 14816
rect 5816 14773 5825 14807
rect 5825 14773 5859 14807
rect 5859 14773 5868 14807
rect 5816 14764 5868 14773
rect 6000 14764 6052 14816
rect 6828 14807 6880 14816
rect 6828 14773 6837 14807
rect 6837 14773 6871 14807
rect 6871 14773 6880 14807
rect 6828 14764 6880 14773
rect 7288 14807 7340 14816
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 10692 14764 10744 14816
rect 11336 14764 11388 14816
rect 12900 14807 12952 14816
rect 12900 14773 12909 14807
rect 12909 14773 12943 14807
rect 12943 14773 12952 14807
rect 12900 14764 12952 14773
rect 13452 14764 13504 14816
rect 14648 14807 14700 14816
rect 14648 14773 14657 14807
rect 14657 14773 14691 14807
rect 14691 14773 14700 14807
rect 14648 14764 14700 14773
rect 18512 14841 18521 14875
rect 18521 14841 18555 14875
rect 18555 14841 18564 14875
rect 18512 14832 18564 14841
rect 19248 14832 19300 14884
rect 18052 14764 18104 14816
rect 19524 14764 19576 14816
rect 20168 14832 20220 14884
rect 21180 14807 21232 14816
rect 21180 14773 21189 14807
rect 21189 14773 21223 14807
rect 21223 14773 21232 14807
rect 21180 14764 21232 14773
rect 21456 14764 21508 14816
rect 23756 14832 23808 14884
rect 24032 14909 24041 14943
rect 24041 14909 24075 14943
rect 24075 14909 24084 14943
rect 24032 14900 24084 14909
rect 25228 14943 25280 14952
rect 25228 14909 25237 14943
rect 25237 14909 25271 14943
rect 25271 14909 25280 14943
rect 25228 14900 25280 14909
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2780 14560 2832 14612
rect 3240 14560 3292 14612
rect 4528 14603 4580 14612
rect 4528 14569 4537 14603
rect 4537 14569 4571 14603
rect 4571 14569 4580 14603
rect 4528 14560 4580 14569
rect 5448 14560 5500 14612
rect 7932 14560 7984 14612
rect 8116 14560 8168 14612
rect 9404 14603 9456 14612
rect 9404 14569 9413 14603
rect 9413 14569 9447 14603
rect 9447 14569 9456 14603
rect 9404 14560 9456 14569
rect 10784 14560 10836 14612
rect 12532 14560 12584 14612
rect 16488 14560 16540 14612
rect 16856 14560 16908 14612
rect 17868 14560 17920 14612
rect 20076 14560 20128 14612
rect 20904 14603 20956 14612
rect 20904 14569 20913 14603
rect 20913 14569 20947 14603
rect 20947 14569 20956 14603
rect 20904 14560 20956 14569
rect 21088 14560 21140 14612
rect 22284 14603 22336 14612
rect 22284 14569 22293 14603
rect 22293 14569 22327 14603
rect 22327 14569 22336 14603
rect 22284 14560 22336 14569
rect 22836 14560 22888 14612
rect 24032 14560 24084 14612
rect 24124 14560 24176 14612
rect 1952 14492 2004 14544
rect 8300 14492 8352 14544
rect 8576 14492 8628 14544
rect 9680 14492 9732 14544
rect 12624 14535 12676 14544
rect 12624 14501 12633 14535
rect 12633 14501 12667 14535
rect 12667 14501 12676 14535
rect 12624 14492 12676 14501
rect 14004 14492 14056 14544
rect 20996 14492 21048 14544
rect 21364 14492 21416 14544
rect 22744 14492 22796 14544
rect 23664 14492 23716 14544
rect 24216 14492 24268 14544
rect 25136 14535 25188 14544
rect 25136 14501 25145 14535
rect 25145 14501 25179 14535
rect 25179 14501 25188 14535
rect 25136 14492 25188 14501
rect 4436 14467 4488 14476
rect 4436 14433 4445 14467
rect 4445 14433 4479 14467
rect 4479 14433 4488 14467
rect 4436 14424 4488 14433
rect 6276 14424 6328 14476
rect 7840 14424 7892 14476
rect 8208 14424 8260 14476
rect 12440 14424 12492 14476
rect 13820 14424 13872 14476
rect 17960 14424 18012 14476
rect 18604 14467 18656 14476
rect 18604 14433 18638 14467
rect 18638 14433 18656 14467
rect 18604 14424 18656 14433
rect 19064 14424 19116 14476
rect 22008 14424 22060 14476
rect 22376 14424 22428 14476
rect 24032 14467 24084 14476
rect 24032 14433 24041 14467
rect 24041 14433 24075 14467
rect 24075 14433 24084 14467
rect 24032 14424 24084 14433
rect 25504 14424 25556 14476
rect 1400 14356 1452 14408
rect 4620 14356 4672 14408
rect 5540 14356 5592 14408
rect 5264 14288 5316 14340
rect 6736 14356 6788 14408
rect 9404 14356 9456 14408
rect 12624 14356 12676 14408
rect 14188 14399 14240 14408
rect 11888 14288 11940 14340
rect 14188 14365 14197 14399
rect 14197 14365 14231 14399
rect 14231 14365 14240 14399
rect 14188 14356 14240 14365
rect 16488 14399 16540 14408
rect 16488 14365 16497 14399
rect 16497 14365 16531 14399
rect 16531 14365 16540 14399
rect 16488 14356 16540 14365
rect 17224 14399 17276 14408
rect 17224 14365 17233 14399
rect 17233 14365 17267 14399
rect 17267 14365 17276 14399
rect 17224 14356 17276 14365
rect 17408 14399 17460 14408
rect 17408 14365 17417 14399
rect 17417 14365 17451 14399
rect 17451 14365 17460 14399
rect 17408 14356 17460 14365
rect 18052 14356 18104 14408
rect 20812 14356 20864 14408
rect 21456 14399 21508 14408
rect 21456 14365 21465 14399
rect 21465 14365 21499 14399
rect 21499 14365 21508 14399
rect 21456 14356 21508 14365
rect 21824 14356 21876 14408
rect 22284 14356 22336 14408
rect 23112 14399 23164 14408
rect 23112 14365 23121 14399
rect 23121 14365 23155 14399
rect 23155 14365 23164 14399
rect 23112 14356 23164 14365
rect 24216 14399 24268 14408
rect 24216 14365 24225 14399
rect 24225 14365 24259 14399
rect 24259 14365 24268 14399
rect 24216 14356 24268 14365
rect 19708 14331 19760 14340
rect 19708 14297 19717 14331
rect 19717 14297 19751 14331
rect 19751 14297 19760 14331
rect 19708 14288 19760 14297
rect 3516 14263 3568 14272
rect 3516 14229 3525 14263
rect 3525 14229 3559 14263
rect 3559 14229 3568 14263
rect 3516 14220 3568 14229
rect 6368 14220 6420 14272
rect 6736 14220 6788 14272
rect 12164 14220 12216 14272
rect 12532 14220 12584 14272
rect 12900 14220 12952 14272
rect 14832 14220 14884 14272
rect 22008 14220 22060 14272
rect 22560 14220 22612 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1860 14059 1912 14068
rect 1860 14025 1869 14059
rect 1869 14025 1903 14059
rect 1903 14025 1912 14059
rect 1860 14016 1912 14025
rect 3976 14016 4028 14068
rect 4436 14016 4488 14068
rect 7840 14059 7892 14068
rect 4620 13948 4672 14000
rect 1860 13812 1912 13864
rect 3424 13880 3476 13932
rect 5724 13923 5776 13932
rect 5724 13889 5733 13923
rect 5733 13889 5767 13923
rect 5767 13889 5776 13923
rect 5724 13880 5776 13889
rect 7288 13923 7340 13932
rect 7288 13889 7297 13923
rect 7297 13889 7331 13923
rect 7331 13889 7340 13923
rect 7288 13880 7340 13889
rect 7840 14025 7849 14059
rect 7849 14025 7883 14059
rect 7883 14025 7892 14059
rect 7840 14016 7892 14025
rect 1400 13744 1452 13796
rect 3792 13812 3844 13864
rect 1952 13676 2004 13728
rect 2596 13676 2648 13728
rect 4436 13676 4488 13728
rect 5816 13812 5868 13864
rect 6092 13812 6144 13864
rect 9496 14016 9548 14068
rect 9680 14016 9732 14068
rect 10784 14016 10836 14068
rect 12440 14059 12492 14068
rect 12440 14025 12449 14059
rect 12449 14025 12483 14059
rect 12483 14025 12492 14059
rect 14004 14059 14056 14068
rect 12440 14016 12492 14025
rect 14004 14025 14013 14059
rect 14013 14025 14047 14059
rect 14047 14025 14056 14059
rect 14004 14016 14056 14025
rect 17224 14016 17276 14068
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 20076 14059 20128 14068
rect 20076 14025 20085 14059
rect 20085 14025 20119 14059
rect 20119 14025 20128 14059
rect 20076 14016 20128 14025
rect 20996 14059 21048 14068
rect 20996 14025 21005 14059
rect 21005 14025 21039 14059
rect 21039 14025 21048 14059
rect 20996 14016 21048 14025
rect 22744 14016 22796 14068
rect 23296 14016 23348 14068
rect 13912 13948 13964 14000
rect 16396 13991 16448 14000
rect 16396 13957 16405 13991
rect 16405 13957 16439 13991
rect 16439 13957 16448 13991
rect 16396 13948 16448 13957
rect 19064 13948 19116 14000
rect 13084 13923 13136 13932
rect 8208 13855 8260 13864
rect 8208 13821 8217 13855
rect 8217 13821 8251 13855
rect 8251 13821 8260 13855
rect 8208 13812 8260 13821
rect 13084 13889 13093 13923
rect 13093 13889 13127 13923
rect 13127 13889 13136 13923
rect 13084 13880 13136 13889
rect 18052 13923 18104 13932
rect 6368 13744 6420 13796
rect 9404 13744 9456 13796
rect 12072 13812 12124 13864
rect 12808 13812 12860 13864
rect 13912 13812 13964 13864
rect 14464 13855 14516 13864
rect 14464 13821 14473 13855
rect 14473 13821 14507 13855
rect 14507 13821 14516 13855
rect 14464 13812 14516 13821
rect 10048 13744 10100 13796
rect 11244 13744 11296 13796
rect 14924 13744 14976 13796
rect 15936 13744 15988 13796
rect 16764 13787 16816 13796
rect 16764 13753 16773 13787
rect 16773 13753 16807 13787
rect 16807 13753 16816 13787
rect 16764 13744 16816 13753
rect 18052 13889 18061 13923
rect 18061 13889 18095 13923
rect 18095 13889 18104 13923
rect 18052 13880 18104 13889
rect 22008 13991 22060 14000
rect 22008 13957 22017 13991
rect 22017 13957 22051 13991
rect 22051 13957 22060 13991
rect 22008 13948 22060 13957
rect 21456 13880 21508 13932
rect 25504 14016 25556 14068
rect 24952 13948 25004 14000
rect 19984 13744 20036 13796
rect 21824 13812 21876 13864
rect 22376 13855 22428 13864
rect 22376 13821 22385 13855
rect 22385 13821 22419 13855
rect 22419 13821 22428 13855
rect 22376 13812 22428 13821
rect 22560 13855 22612 13864
rect 22560 13821 22569 13855
rect 22569 13821 22603 13855
rect 22603 13821 22612 13855
rect 22560 13812 22612 13821
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 11060 13719 11112 13728
rect 11060 13685 11069 13719
rect 11069 13685 11103 13719
rect 11103 13685 11112 13719
rect 11060 13676 11112 13685
rect 12532 13676 12584 13728
rect 13728 13676 13780 13728
rect 17776 13676 17828 13728
rect 19340 13676 19392 13728
rect 20812 13719 20864 13728
rect 20812 13685 20821 13719
rect 20821 13685 20855 13719
rect 20855 13685 20864 13719
rect 20812 13676 20864 13685
rect 21364 13719 21416 13728
rect 21364 13685 21373 13719
rect 21373 13685 21407 13719
rect 21407 13685 21416 13719
rect 21364 13676 21416 13685
rect 22192 13676 22244 13728
rect 22744 13676 22796 13728
rect 23848 13676 23900 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1952 13515 2004 13524
rect 1952 13481 1961 13515
rect 1961 13481 1995 13515
rect 1995 13481 2004 13515
rect 1952 13472 2004 13481
rect 2504 13472 2556 13524
rect 2780 13472 2832 13524
rect 3792 13472 3844 13524
rect 3976 13472 4028 13524
rect 4528 13472 4580 13524
rect 5724 13472 5776 13524
rect 6552 13472 6604 13524
rect 8024 13515 8076 13524
rect 8024 13481 8033 13515
rect 8033 13481 8067 13515
rect 8067 13481 8076 13515
rect 8024 13472 8076 13481
rect 8392 13515 8444 13524
rect 8392 13481 8401 13515
rect 8401 13481 8435 13515
rect 8435 13481 8444 13515
rect 8392 13472 8444 13481
rect 8668 13472 8720 13524
rect 9404 13515 9456 13524
rect 9404 13481 9413 13515
rect 9413 13481 9447 13515
rect 9447 13481 9456 13515
rect 9404 13472 9456 13481
rect 12808 13472 12860 13524
rect 13544 13472 13596 13524
rect 17960 13472 18012 13524
rect 20168 13515 20220 13524
rect 20168 13481 20177 13515
rect 20177 13481 20211 13515
rect 20211 13481 20220 13515
rect 20168 13472 20220 13481
rect 21456 13472 21508 13524
rect 22652 13472 22704 13524
rect 23112 13472 23164 13524
rect 4988 13404 5040 13456
rect 5540 13404 5592 13456
rect 6828 13404 6880 13456
rect 3056 13336 3108 13388
rect 3608 13336 3660 13388
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 2964 13311 3016 13320
rect 2964 13277 2973 13311
rect 2973 13277 3007 13311
rect 3007 13277 3016 13311
rect 2964 13268 3016 13277
rect 3976 13336 4028 13388
rect 5632 13336 5684 13388
rect 6184 13336 6236 13388
rect 6736 13336 6788 13388
rect 12532 13447 12584 13456
rect 12532 13413 12541 13447
rect 12541 13413 12575 13447
rect 12575 13413 12584 13447
rect 12532 13404 12584 13413
rect 21088 13404 21140 13456
rect 10324 13336 10376 13388
rect 12164 13336 12216 13388
rect 15568 13379 15620 13388
rect 15568 13345 15602 13379
rect 15602 13345 15620 13379
rect 15568 13336 15620 13345
rect 18236 13336 18288 13388
rect 20996 13379 21048 13388
rect 20996 13345 21005 13379
rect 21005 13345 21039 13379
rect 21039 13345 21048 13379
rect 20996 13336 21048 13345
rect 22100 13379 22152 13388
rect 22100 13345 22109 13379
rect 22109 13345 22143 13379
rect 22143 13345 22152 13379
rect 22100 13336 22152 13345
rect 23940 13336 23992 13388
rect 4896 13268 4948 13320
rect 4436 13200 4488 13252
rect 5264 13200 5316 13252
rect 8576 13311 8628 13320
rect 8576 13277 8585 13311
rect 8585 13277 8619 13311
rect 8619 13277 8628 13311
rect 8576 13268 8628 13277
rect 9680 13268 9732 13320
rect 14372 13268 14424 13320
rect 14832 13268 14884 13320
rect 18512 13311 18564 13320
rect 18512 13277 18521 13311
rect 18521 13277 18555 13311
rect 18555 13277 18564 13311
rect 18512 13268 18564 13277
rect 18604 13311 18656 13320
rect 18604 13277 18613 13311
rect 18613 13277 18647 13311
rect 18647 13277 18656 13311
rect 19064 13311 19116 13320
rect 18604 13268 18656 13277
rect 19064 13277 19073 13311
rect 19073 13277 19107 13311
rect 19107 13277 19116 13311
rect 19064 13268 19116 13277
rect 19616 13311 19668 13320
rect 19616 13277 19625 13311
rect 19625 13277 19659 13311
rect 19659 13277 19668 13311
rect 19616 13268 19668 13277
rect 23480 13268 23532 13320
rect 25412 13311 25464 13320
rect 25412 13277 25421 13311
rect 25421 13277 25455 13311
rect 25455 13277 25464 13311
rect 25412 13268 25464 13277
rect 21180 13243 21232 13252
rect 2228 13175 2280 13184
rect 2228 13141 2237 13175
rect 2237 13141 2271 13175
rect 2271 13141 2280 13175
rect 2228 13132 2280 13141
rect 3700 13132 3752 13184
rect 21180 13209 21189 13243
rect 21189 13209 21223 13243
rect 21223 13209 21232 13243
rect 21180 13200 21232 13209
rect 23756 13200 23808 13252
rect 23940 13200 23992 13252
rect 6828 13132 6880 13184
rect 11612 13175 11664 13184
rect 11612 13141 11621 13175
rect 11621 13141 11655 13175
rect 11655 13141 11664 13175
rect 11612 13132 11664 13141
rect 14004 13175 14056 13184
rect 14004 13141 14013 13175
rect 14013 13141 14047 13175
rect 14047 13141 14056 13175
rect 14004 13132 14056 13141
rect 14280 13132 14332 13184
rect 16672 13175 16724 13184
rect 16672 13141 16681 13175
rect 16681 13141 16715 13175
rect 16715 13141 16724 13175
rect 16672 13132 16724 13141
rect 23848 13132 23900 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 3056 12928 3108 12980
rect 3332 12971 3384 12980
rect 3332 12937 3341 12971
rect 3341 12937 3375 12971
rect 3375 12937 3384 12971
rect 3332 12928 3384 12937
rect 4712 12928 4764 12980
rect 2228 12835 2280 12844
rect 2228 12801 2237 12835
rect 2237 12801 2271 12835
rect 2271 12801 2280 12835
rect 2228 12792 2280 12801
rect 2688 12792 2740 12844
rect 3884 12835 3936 12844
rect 3884 12801 3893 12835
rect 3893 12801 3927 12835
rect 3927 12801 3936 12835
rect 3884 12792 3936 12801
rect 5448 12928 5500 12980
rect 6184 12971 6236 12980
rect 6184 12937 6193 12971
rect 6193 12937 6227 12971
rect 6227 12937 6236 12971
rect 6184 12928 6236 12937
rect 6552 12971 6604 12980
rect 6552 12937 6561 12971
rect 6561 12937 6595 12971
rect 6595 12937 6604 12971
rect 6552 12928 6604 12937
rect 8668 12928 8720 12980
rect 9404 12928 9456 12980
rect 10048 12928 10100 12980
rect 5724 12792 5776 12844
rect 6276 12792 6328 12844
rect 10324 12903 10376 12912
rect 10324 12869 10333 12903
rect 10333 12869 10367 12903
rect 10367 12869 10376 12903
rect 10324 12860 10376 12869
rect 14096 12928 14148 12980
rect 15568 12928 15620 12980
rect 15844 12928 15896 12980
rect 18236 12971 18288 12980
rect 18236 12937 18245 12971
rect 18245 12937 18279 12971
rect 18279 12937 18288 12971
rect 18236 12928 18288 12937
rect 19248 12928 19300 12980
rect 20996 12971 21048 12980
rect 20996 12937 21005 12971
rect 21005 12937 21039 12971
rect 21039 12937 21048 12971
rect 20996 12928 21048 12937
rect 21640 12928 21692 12980
rect 22100 12971 22152 12980
rect 22100 12937 22109 12971
rect 22109 12937 22143 12971
rect 22143 12937 22152 12971
rect 22100 12928 22152 12937
rect 23204 12928 23256 12980
rect 9772 12835 9824 12844
rect 3516 12724 3568 12776
rect 5540 12767 5592 12776
rect 5540 12733 5549 12767
rect 5549 12733 5583 12767
rect 5583 12733 5592 12767
rect 5540 12724 5592 12733
rect 6828 12767 6880 12776
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 9772 12801 9781 12835
rect 9781 12801 9815 12835
rect 9815 12801 9824 12835
rect 9772 12792 9824 12801
rect 9588 12724 9640 12776
rect 11060 12792 11112 12844
rect 11244 12835 11296 12844
rect 11244 12801 11253 12835
rect 11253 12801 11287 12835
rect 11287 12801 11296 12835
rect 11244 12792 11296 12801
rect 11612 12860 11664 12912
rect 11704 12724 11756 12776
rect 12900 12835 12952 12844
rect 12900 12801 12909 12835
rect 12909 12801 12943 12835
rect 12943 12801 12952 12835
rect 12900 12792 12952 12801
rect 12992 12835 13044 12844
rect 12992 12801 13001 12835
rect 13001 12801 13035 12835
rect 13035 12801 13044 12835
rect 14096 12835 14148 12844
rect 12992 12792 13044 12801
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 14372 12835 14424 12844
rect 14372 12801 14381 12835
rect 14381 12801 14415 12835
rect 14415 12801 14424 12835
rect 14372 12792 14424 12801
rect 17776 12792 17828 12844
rect 18696 12835 18748 12844
rect 18696 12801 18705 12835
rect 18705 12801 18739 12835
rect 18739 12801 18748 12835
rect 18696 12792 18748 12801
rect 19984 12860 20036 12912
rect 19248 12792 19300 12844
rect 19708 12835 19760 12844
rect 19708 12801 19717 12835
rect 19717 12801 19751 12835
rect 19751 12801 19760 12835
rect 19708 12792 19760 12801
rect 24952 12860 25004 12912
rect 20812 12792 20864 12844
rect 12440 12724 12492 12776
rect 14280 12724 14332 12776
rect 18328 12724 18380 12776
rect 19616 12724 19668 12776
rect 19984 12724 20036 12776
rect 3976 12656 4028 12708
rect 5724 12656 5776 12708
rect 2136 12631 2188 12640
rect 2136 12597 2145 12631
rect 2145 12597 2179 12631
rect 2179 12597 2188 12631
rect 2136 12588 2188 12597
rect 2780 12631 2832 12640
rect 2780 12597 2789 12631
rect 2789 12597 2823 12631
rect 2823 12597 2832 12631
rect 3700 12631 3752 12640
rect 2780 12588 2832 12597
rect 3700 12597 3709 12631
rect 3709 12597 3743 12631
rect 3743 12597 3752 12631
rect 3700 12588 3752 12597
rect 7840 12588 7892 12640
rect 10784 12631 10836 12640
rect 10784 12597 10793 12631
rect 10793 12597 10827 12631
rect 10827 12597 10836 12631
rect 10784 12588 10836 12597
rect 11060 12588 11112 12640
rect 12164 12631 12216 12640
rect 12164 12597 12173 12631
rect 12173 12597 12207 12631
rect 12207 12597 12216 12631
rect 12164 12588 12216 12597
rect 14188 12656 14240 12708
rect 15016 12656 15068 12708
rect 15660 12656 15712 12708
rect 15936 12656 15988 12708
rect 16580 12656 16632 12708
rect 19524 12656 19576 12708
rect 20260 12724 20312 12776
rect 21088 12724 21140 12776
rect 23848 12767 23900 12776
rect 23848 12733 23857 12767
rect 23857 12733 23891 12767
rect 23891 12733 23900 12767
rect 23848 12724 23900 12733
rect 24032 12656 24084 12708
rect 25412 12656 25464 12708
rect 13912 12631 13964 12640
rect 13912 12597 13921 12631
rect 13921 12597 13955 12631
rect 13955 12597 13964 12631
rect 13912 12588 13964 12597
rect 15108 12588 15160 12640
rect 16488 12588 16540 12640
rect 19984 12588 20036 12640
rect 20628 12588 20680 12640
rect 24768 12588 24820 12640
rect 24860 12588 24912 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2136 12384 2188 12436
rect 3884 12384 3936 12436
rect 3976 12384 4028 12436
rect 5172 12384 5224 12436
rect 6092 12427 6144 12436
rect 6092 12393 6101 12427
rect 6101 12393 6135 12427
rect 6135 12393 6144 12427
rect 6092 12384 6144 12393
rect 6828 12427 6880 12436
rect 6828 12393 6837 12427
rect 6837 12393 6871 12427
rect 6871 12393 6880 12427
rect 6828 12384 6880 12393
rect 7380 12384 7432 12436
rect 8392 12384 8444 12436
rect 8576 12427 8628 12436
rect 8576 12393 8585 12427
rect 8585 12393 8619 12427
rect 8619 12393 8628 12427
rect 8576 12384 8628 12393
rect 10876 12384 10928 12436
rect 12992 12384 13044 12436
rect 14096 12384 14148 12436
rect 14648 12384 14700 12436
rect 2964 12316 3016 12368
rect 4528 12316 4580 12368
rect 5264 12316 5316 12368
rect 10692 12316 10744 12368
rect 2412 12291 2464 12300
rect 2412 12257 2421 12291
rect 2421 12257 2455 12291
rect 2455 12257 2464 12291
rect 2412 12248 2464 12257
rect 2596 12248 2648 12300
rect 2136 12180 2188 12232
rect 2504 12223 2556 12232
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 5080 12248 5132 12300
rect 7196 12248 7248 12300
rect 7472 12291 7524 12300
rect 7472 12257 7481 12291
rect 7481 12257 7515 12291
rect 7515 12257 7524 12291
rect 7472 12248 7524 12257
rect 9404 12248 9456 12300
rect 11152 12248 11204 12300
rect 11336 12291 11388 12300
rect 11336 12257 11370 12291
rect 11370 12257 11388 12291
rect 11336 12248 11388 12257
rect 12992 12248 13044 12300
rect 13084 12248 13136 12300
rect 13544 12248 13596 12300
rect 13820 12248 13872 12300
rect 2504 12180 2556 12189
rect 4252 12180 4304 12232
rect 5724 12223 5776 12232
rect 5724 12189 5733 12223
rect 5733 12189 5767 12223
rect 5767 12189 5776 12223
rect 5724 12180 5776 12189
rect 7840 12180 7892 12232
rect 14096 12180 14148 12232
rect 14372 12180 14424 12232
rect 11060 12112 11112 12164
rect 12900 12112 12952 12164
rect 15384 12384 15436 12436
rect 15568 12384 15620 12436
rect 16120 12384 16172 12436
rect 16764 12384 16816 12436
rect 17408 12384 17460 12436
rect 18328 12427 18380 12436
rect 18328 12393 18337 12427
rect 18337 12393 18371 12427
rect 18371 12393 18380 12427
rect 18328 12384 18380 12393
rect 18512 12384 18564 12436
rect 19524 12384 19576 12436
rect 20168 12427 20220 12436
rect 20168 12393 20177 12427
rect 20177 12393 20211 12427
rect 20211 12393 20220 12427
rect 20168 12384 20220 12393
rect 21732 12384 21784 12436
rect 22744 12427 22796 12436
rect 22744 12393 22753 12427
rect 22753 12393 22787 12427
rect 22787 12393 22796 12427
rect 22744 12384 22796 12393
rect 15844 12316 15896 12368
rect 16396 12248 16448 12300
rect 15752 12223 15804 12232
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15752 12180 15804 12189
rect 15936 12112 15988 12164
rect 16672 12112 16724 12164
rect 18604 12316 18656 12368
rect 19156 12316 19208 12368
rect 23020 12316 23072 12368
rect 24860 12384 24912 12436
rect 24584 12316 24636 12368
rect 17040 12248 17092 12300
rect 21456 12291 21508 12300
rect 21456 12257 21465 12291
rect 21465 12257 21499 12291
rect 21499 12257 21508 12291
rect 21456 12248 21508 12257
rect 22560 12291 22612 12300
rect 22560 12257 22569 12291
rect 22569 12257 22603 12291
rect 22603 12257 22612 12291
rect 22560 12248 22612 12257
rect 23296 12248 23348 12300
rect 23572 12248 23624 12300
rect 24860 12248 24912 12300
rect 17684 12180 17736 12232
rect 18788 12180 18840 12232
rect 19248 12223 19300 12232
rect 19248 12189 19257 12223
rect 19257 12189 19291 12223
rect 19291 12189 19300 12223
rect 19248 12180 19300 12189
rect 2780 12044 2832 12096
rect 2964 12044 3016 12096
rect 12992 12087 13044 12096
rect 12992 12053 13001 12087
rect 13001 12053 13035 12087
rect 13035 12053 13044 12087
rect 12992 12044 13044 12053
rect 14188 12044 14240 12096
rect 15568 12044 15620 12096
rect 16488 12044 16540 12096
rect 16764 12087 16816 12096
rect 16764 12053 16773 12087
rect 16773 12053 16807 12087
rect 16807 12053 16816 12087
rect 16764 12044 16816 12053
rect 24032 12044 24084 12096
rect 25044 12087 25096 12096
rect 25044 12053 25053 12087
rect 25053 12053 25087 12087
rect 25087 12053 25096 12087
rect 25044 12044 25096 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2228 11840 2280 11892
rect 2596 11840 2648 11892
rect 2596 11704 2648 11756
rect 2964 11704 3016 11756
rect 3516 11840 3568 11892
rect 7196 11883 7248 11892
rect 7196 11849 7205 11883
rect 7205 11849 7239 11883
rect 7239 11849 7248 11883
rect 7196 11840 7248 11849
rect 7380 11840 7432 11892
rect 7840 11883 7892 11892
rect 7840 11849 7849 11883
rect 7849 11849 7883 11883
rect 7883 11849 7892 11883
rect 7840 11840 7892 11849
rect 10968 11840 11020 11892
rect 11060 11840 11112 11892
rect 12440 11883 12492 11892
rect 12440 11849 12449 11883
rect 12449 11849 12483 11883
rect 12483 11849 12492 11883
rect 12440 11840 12492 11849
rect 12900 11840 12952 11892
rect 14096 11840 14148 11892
rect 15936 11883 15988 11892
rect 15936 11849 15945 11883
rect 15945 11849 15979 11883
rect 15979 11849 15988 11883
rect 15936 11840 15988 11849
rect 17408 11883 17460 11892
rect 17408 11849 17417 11883
rect 17417 11849 17451 11883
rect 17451 11849 17460 11883
rect 17408 11840 17460 11849
rect 17684 11883 17736 11892
rect 17684 11849 17693 11883
rect 17693 11849 17727 11883
rect 17727 11849 17736 11883
rect 17684 11840 17736 11849
rect 18788 11883 18840 11892
rect 18788 11849 18797 11883
rect 18797 11849 18831 11883
rect 18831 11849 18840 11883
rect 18788 11840 18840 11849
rect 19248 11840 19300 11892
rect 21456 11840 21508 11892
rect 22560 11840 22612 11892
rect 23388 11840 23440 11892
rect 23848 11840 23900 11892
rect 24032 11840 24084 11892
rect 25688 11883 25740 11892
rect 25688 11849 25697 11883
rect 25697 11849 25731 11883
rect 25731 11849 25740 11883
rect 25688 11840 25740 11849
rect 16764 11772 16816 11824
rect 20168 11772 20220 11824
rect 4344 11704 4396 11756
rect 4528 11747 4580 11756
rect 4528 11713 4537 11747
rect 4537 11713 4571 11747
rect 4571 11713 4580 11747
rect 4528 11704 4580 11713
rect 6184 11704 6236 11756
rect 8944 11704 8996 11756
rect 10692 11704 10744 11756
rect 11704 11704 11756 11756
rect 12992 11747 13044 11756
rect 12992 11713 13001 11747
rect 13001 11713 13035 11747
rect 13035 11713 13044 11747
rect 14372 11747 14424 11756
rect 12992 11704 13044 11713
rect 14372 11713 14381 11747
rect 14381 11713 14415 11747
rect 14415 11713 14424 11747
rect 14372 11704 14424 11713
rect 15568 11747 15620 11756
rect 15568 11713 15577 11747
rect 15577 11713 15611 11747
rect 15611 11713 15620 11747
rect 15568 11704 15620 11713
rect 15936 11704 15988 11756
rect 16304 11704 16356 11756
rect 20444 11704 20496 11756
rect 21916 11704 21968 11756
rect 23020 11747 23072 11756
rect 23020 11713 23029 11747
rect 23029 11713 23063 11747
rect 23063 11713 23072 11747
rect 23020 11704 23072 11713
rect 23940 11704 23992 11756
rect 11336 11636 11388 11688
rect 2780 11611 2832 11620
rect 2780 11577 2789 11611
rect 2789 11577 2823 11611
rect 2823 11577 2832 11611
rect 2780 11568 2832 11577
rect 4068 11568 4120 11620
rect 12072 11568 12124 11620
rect 3516 11543 3568 11552
rect 3516 11509 3525 11543
rect 3525 11509 3559 11543
rect 3559 11509 3568 11543
rect 3516 11500 3568 11509
rect 4252 11500 4304 11552
rect 11060 11500 11112 11552
rect 13084 11636 13136 11688
rect 13820 11636 13872 11688
rect 15108 11636 15160 11688
rect 15384 11636 15436 11688
rect 15752 11636 15804 11688
rect 22468 11679 22520 11688
rect 22468 11645 22477 11679
rect 22477 11645 22511 11679
rect 22511 11645 22520 11679
rect 22468 11636 22520 11645
rect 24768 11636 24820 11688
rect 25504 11679 25556 11688
rect 25504 11645 25513 11679
rect 25513 11645 25547 11679
rect 25547 11645 25556 11679
rect 25504 11636 25556 11645
rect 15016 11568 15068 11620
rect 16488 11568 16540 11620
rect 24124 11568 24176 11620
rect 14924 11543 14976 11552
rect 14924 11509 14933 11543
rect 14933 11509 14967 11543
rect 14967 11509 14976 11543
rect 14924 11500 14976 11509
rect 15108 11500 15160 11552
rect 15568 11500 15620 11552
rect 17040 11543 17092 11552
rect 17040 11509 17049 11543
rect 17049 11509 17083 11543
rect 17083 11509 17092 11543
rect 17040 11500 17092 11509
rect 19156 11543 19208 11552
rect 19156 11509 19165 11543
rect 19165 11509 19199 11543
rect 19199 11509 19208 11543
rect 19156 11500 19208 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 1860 11296 1912 11305
rect 2412 11296 2464 11348
rect 4068 11339 4120 11348
rect 4068 11305 4077 11339
rect 4077 11305 4111 11339
rect 4111 11305 4120 11339
rect 4068 11296 4120 11305
rect 4160 11296 4212 11348
rect 4804 11296 4856 11348
rect 5540 11339 5592 11348
rect 5540 11305 5549 11339
rect 5549 11305 5583 11339
rect 5583 11305 5592 11339
rect 5540 11296 5592 11305
rect 11704 11296 11756 11348
rect 12072 11339 12124 11348
rect 12072 11305 12081 11339
rect 12081 11305 12115 11339
rect 12115 11305 12124 11339
rect 12072 11296 12124 11305
rect 12532 11296 12584 11348
rect 12900 11296 12952 11348
rect 14004 11296 14056 11348
rect 15016 11339 15068 11348
rect 15016 11305 15025 11339
rect 15025 11305 15059 11339
rect 15059 11305 15068 11339
rect 15016 11296 15068 11305
rect 15292 11339 15344 11348
rect 15292 11305 15301 11339
rect 15301 11305 15335 11339
rect 15335 11305 15344 11339
rect 15292 11296 15344 11305
rect 16396 11339 16448 11348
rect 16396 11305 16405 11339
rect 16405 11305 16439 11339
rect 16439 11305 16448 11339
rect 16396 11296 16448 11305
rect 22376 11339 22428 11348
rect 22376 11305 22385 11339
rect 22385 11305 22419 11339
rect 22419 11305 22428 11339
rect 22376 11296 22428 11305
rect 22468 11296 22520 11348
rect 23388 11296 23440 11348
rect 23664 11339 23716 11348
rect 23664 11305 23673 11339
rect 23673 11305 23707 11339
rect 23707 11305 23716 11339
rect 23664 11296 23716 11305
rect 25320 11296 25372 11348
rect 2504 11228 2556 11280
rect 13912 11228 13964 11280
rect 14924 11228 14976 11280
rect 23940 11228 23992 11280
rect 1400 11160 1452 11212
rect 2044 11160 2096 11212
rect 2964 11160 3016 11212
rect 12624 11160 12676 11212
rect 14096 11160 14148 11212
rect 15568 11160 15620 11212
rect 16028 11160 16080 11212
rect 24032 11160 24084 11212
rect 24584 11203 24636 11212
rect 24584 11169 24593 11203
rect 24593 11169 24627 11203
rect 24627 11169 24636 11203
rect 24584 11160 24636 11169
rect 24768 11160 24820 11212
rect 1952 11092 2004 11144
rect 2320 11092 2372 11144
rect 4528 11135 4580 11144
rect 1860 11024 1912 11076
rect 4528 11101 4537 11135
rect 4537 11101 4571 11135
rect 4571 11101 4580 11135
rect 4528 11092 4580 11101
rect 4712 11135 4764 11144
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4712 11092 4764 11101
rect 12164 11092 12216 11144
rect 12992 11092 13044 11144
rect 14188 11135 14240 11144
rect 14188 11101 14197 11135
rect 14197 11101 14231 11135
rect 14231 11101 14240 11135
rect 14188 11092 14240 11101
rect 15936 11135 15988 11144
rect 15936 11101 15945 11135
rect 15945 11101 15979 11135
rect 15979 11101 15988 11135
rect 15936 11092 15988 11101
rect 16580 11092 16632 11144
rect 3608 11024 3660 11076
rect 5080 11067 5132 11076
rect 5080 11033 5089 11067
rect 5089 11033 5123 11067
rect 5123 11033 5132 11067
rect 5080 11024 5132 11033
rect 11152 11024 11204 11076
rect 11980 11024 12032 11076
rect 3056 10956 3108 11008
rect 24124 11024 24176 11076
rect 14648 10956 14700 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2504 10752 2556 10804
rect 4160 10795 4212 10804
rect 4160 10761 4169 10795
rect 4169 10761 4203 10795
rect 4203 10761 4212 10795
rect 4160 10752 4212 10761
rect 4528 10795 4580 10804
rect 4528 10761 4537 10795
rect 4537 10761 4571 10795
rect 4571 10761 4580 10795
rect 4528 10752 4580 10761
rect 4712 10752 4764 10804
rect 12348 10752 12400 10804
rect 14004 10795 14056 10804
rect 14004 10761 14013 10795
rect 14013 10761 14047 10795
rect 14047 10761 14056 10795
rect 14004 10752 14056 10761
rect 14096 10752 14148 10804
rect 15384 10752 15436 10804
rect 24032 10752 24084 10804
rect 24768 10752 24820 10804
rect 3056 10659 3108 10668
rect 3056 10625 3065 10659
rect 3065 10625 3099 10659
rect 3099 10625 3108 10659
rect 3056 10616 3108 10625
rect 12348 10616 12400 10668
rect 13268 10616 13320 10668
rect 15108 10659 15160 10668
rect 15108 10625 15117 10659
rect 15117 10625 15151 10659
rect 15151 10625 15160 10659
rect 15108 10616 15160 10625
rect 15936 10616 15988 10668
rect 12900 10591 12952 10600
rect 12900 10557 12909 10591
rect 12909 10557 12943 10591
rect 12943 10557 12952 10591
rect 12900 10548 12952 10557
rect 14832 10548 14884 10600
rect 24584 10591 24636 10600
rect 24584 10557 24593 10591
rect 24593 10557 24627 10591
rect 24627 10557 24636 10591
rect 24584 10548 24636 10557
rect 2688 10480 2740 10532
rect 2964 10480 3016 10532
rect 14648 10480 14700 10532
rect 1952 10412 2004 10464
rect 3332 10412 3384 10464
rect 3792 10412 3844 10464
rect 12532 10455 12584 10464
rect 12532 10421 12541 10455
rect 12541 10421 12575 10455
rect 12575 10421 12584 10455
rect 12532 10412 12584 10421
rect 13544 10455 13596 10464
rect 13544 10421 13553 10455
rect 13553 10421 13587 10455
rect 13587 10421 13596 10455
rect 13544 10412 13596 10421
rect 15568 10455 15620 10464
rect 15568 10421 15577 10455
rect 15577 10421 15611 10455
rect 15611 10421 15620 10455
rect 15568 10412 15620 10421
rect 16028 10455 16080 10464
rect 16028 10421 16037 10455
rect 16037 10421 16071 10455
rect 16071 10421 16080 10455
rect 16028 10412 16080 10421
rect 25780 10412 25832 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 2044 10251 2096 10260
rect 2044 10217 2053 10251
rect 2053 10217 2087 10251
rect 2087 10217 2096 10251
rect 2044 10208 2096 10217
rect 3056 10251 3108 10260
rect 3056 10217 3065 10251
rect 3065 10217 3099 10251
rect 3099 10217 3108 10251
rect 3056 10208 3108 10217
rect 12256 10251 12308 10260
rect 12256 10217 12265 10251
rect 12265 10217 12299 10251
rect 12299 10217 12308 10251
rect 12256 10208 12308 10217
rect 12532 10208 12584 10260
rect 12716 10251 12768 10260
rect 12716 10217 12725 10251
rect 12725 10217 12759 10251
rect 12759 10217 12768 10251
rect 13268 10251 13320 10260
rect 12716 10208 12768 10217
rect 13268 10217 13277 10251
rect 13277 10217 13311 10251
rect 13311 10217 13320 10251
rect 13268 10208 13320 10217
rect 14832 10208 14884 10260
rect 15108 10208 15160 10260
rect 15476 10208 15528 10260
rect 15752 10208 15804 10260
rect 16488 10208 16540 10260
rect 26056 10208 26108 10260
rect 12164 10183 12216 10192
rect 12164 10149 12173 10183
rect 12173 10149 12207 10183
rect 12207 10149 12216 10183
rect 12164 10140 12216 10149
rect 1676 10072 1728 10124
rect 2688 10072 2740 10124
rect 15660 10072 15712 10124
rect 24676 10072 24728 10124
rect 12624 10004 12676 10056
rect 13360 10004 13412 10056
rect 14648 10004 14700 10056
rect 15936 10004 15988 10056
rect 6184 9936 6236 9988
rect 14096 9868 14148 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2596 9707 2648 9716
rect 2596 9673 2605 9707
rect 2605 9673 2639 9707
rect 2639 9673 2648 9707
rect 2596 9664 2648 9673
rect 12624 9707 12676 9716
rect 12624 9673 12633 9707
rect 12633 9673 12667 9707
rect 12667 9673 12676 9707
rect 12624 9664 12676 9673
rect 12716 9664 12768 9716
rect 15752 9707 15804 9716
rect 15752 9673 15761 9707
rect 15761 9673 15795 9707
rect 15795 9673 15804 9707
rect 15752 9664 15804 9673
rect 15936 9664 15988 9716
rect 24676 9707 24728 9716
rect 24676 9673 24685 9707
rect 24685 9673 24719 9707
rect 24719 9673 24728 9707
rect 24676 9664 24728 9673
rect 26240 9664 26292 9716
rect 14740 9596 14792 9648
rect 15660 9596 15712 9648
rect 24216 9596 24268 9648
rect 25964 9596 26016 9648
rect 12532 9528 12584 9580
rect 14648 9571 14700 9580
rect 14648 9537 14657 9571
rect 14657 9537 14691 9571
rect 14691 9537 14700 9571
rect 14648 9528 14700 9537
rect 1492 9460 1544 9512
rect 14464 9460 14516 9512
rect 14188 9392 14240 9444
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 13912 9324 13964 9376
rect 14832 9324 14884 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1676 9163 1728 9172
rect 1676 9129 1685 9163
rect 1685 9129 1719 9163
rect 1719 9129 1728 9163
rect 1676 9120 1728 9129
rect 14188 8823 14240 8832
rect 14188 8789 14197 8823
rect 14197 8789 14231 8823
rect 14231 8789 14240 8823
rect 14188 8780 14240 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 25136 8576 25188 8628
rect 23664 8415 23716 8424
rect 23664 8381 23673 8415
rect 23673 8381 23707 8415
rect 23707 8381 23716 8415
rect 23664 8372 23716 8381
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 24216 5899 24268 5908
rect 24216 5865 24225 5899
rect 24225 5865 24259 5899
rect 24259 5865 24268 5899
rect 24216 5856 24268 5865
rect 24032 5763 24084 5772
rect 24032 5729 24041 5763
rect 24041 5729 24075 5763
rect 24075 5729 24084 5763
rect 24032 5720 24084 5729
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 24032 5355 24084 5364
rect 24032 5321 24041 5355
rect 24041 5321 24075 5355
rect 24075 5321 24084 5355
rect 24032 5312 24084 5321
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 24124 4811 24176 4820
rect 24124 4777 24133 4811
rect 24133 4777 24167 4811
rect 24167 4777 24176 4811
rect 24124 4768 24176 4777
rect 24676 4700 24728 4752
rect 24124 4632 24176 4684
rect 24768 4607 24820 4616
rect 24768 4573 24777 4607
rect 24777 4573 24811 4607
rect 24811 4573 24820 4607
rect 24768 4564 24820 4573
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 572 4224 624 4276
rect 8208 4224 8260 4276
rect 17960 4156 18012 4208
rect 24124 4199 24176 4208
rect 24124 4165 24133 4199
rect 24133 4165 24167 4199
rect 24167 4165 24176 4199
rect 24124 4156 24176 4165
rect 24768 4156 24820 4208
rect 24584 3927 24636 3936
rect 24584 3893 24593 3927
rect 24593 3893 24627 3927
rect 24627 3893 24636 3927
rect 24584 3884 24636 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 940 3680 992 3732
rect 2964 3680 3016 3732
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1308 2864 1360 2916
rect 3516 2864 3568 2916
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 11980 2635 12032 2644
rect 11980 2601 11989 2635
rect 11989 2601 12023 2635
rect 12023 2601 12032 2635
rect 11980 2592 12032 2601
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12440 2592 12492 2601
rect 14096 2592 14148 2644
rect 26516 2592 26568 2644
rect 25136 2499 25188 2508
rect 25136 2465 25145 2499
rect 25145 2465 25179 2499
rect 25179 2465 25188 2499
rect 25136 2456 25188 2465
rect 25136 2252 25188 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 1950 27520 2006 28000
rect 2502 27520 2558 28000
rect 3054 27520 3110 28000
rect 3514 27704 3570 27713
rect 3514 27639 3570 27648
rect 308 27418 336 27520
rect 216 27390 336 27418
rect 216 15881 244 27390
rect 860 22681 888 27520
rect 1412 24154 1440 27520
rect 1964 25809 1992 27520
rect 1950 25800 2006 25809
rect 1950 25735 2006 25744
rect 2044 25356 2096 25362
rect 2044 25298 2096 25304
rect 1860 24880 1912 24886
rect 1860 24822 1912 24828
rect 1584 24608 1636 24614
rect 1584 24550 1636 24556
rect 1412 24126 1532 24154
rect 1400 24064 1452 24070
rect 1400 24006 1452 24012
rect 846 22672 902 22681
rect 846 22607 902 22616
rect 1412 20369 1440 24006
rect 1504 23769 1532 24126
rect 1490 23760 1546 23769
rect 1490 23695 1546 23704
rect 1596 21593 1624 24550
rect 1676 24268 1728 24274
rect 1676 24210 1728 24216
rect 1688 22982 1716 24210
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1582 21584 1638 21593
rect 1582 21519 1638 21528
rect 1398 20360 1454 20369
rect 1398 20295 1454 20304
rect 1688 20097 1716 22918
rect 1780 22273 1808 24006
rect 1872 23730 1900 24822
rect 2056 24614 2084 25298
rect 2516 24834 2544 27520
rect 3068 25945 3096 27520
rect 3528 26314 3556 27639
rect 3606 27520 3662 28000
rect 4158 27520 4214 28000
rect 4710 27520 4766 28000
rect 5262 27520 5318 28000
rect 5814 27520 5870 28000
rect 6366 27520 6422 28000
rect 6918 27520 6974 28000
rect 7562 27520 7618 28000
rect 8114 27520 8170 28000
rect 8666 27520 8722 28000
rect 9218 27520 9274 28000
rect 9770 27520 9826 28000
rect 10322 27520 10378 28000
rect 10874 27520 10930 28000
rect 11426 27520 11482 28000
rect 11978 27520 12034 28000
rect 12530 27520 12586 28000
rect 13082 27520 13138 28000
rect 13634 27520 13690 28000
rect 14278 27520 14334 28000
rect 14830 27520 14886 28000
rect 15382 27520 15438 28000
rect 15934 27520 15990 28000
rect 16486 27520 16542 28000
rect 17038 27520 17094 28000
rect 17590 27520 17646 28000
rect 18142 27520 18198 28000
rect 18694 27520 18750 28000
rect 19246 27520 19302 28000
rect 19798 27520 19854 28000
rect 20350 27520 20406 28000
rect 20902 27520 20958 28000
rect 21546 27520 21602 28000
rect 22098 27520 22154 28000
rect 22650 27520 22706 28000
rect 23202 27520 23258 28000
rect 23754 27520 23810 28000
rect 24122 27704 24178 27713
rect 24122 27639 24178 27648
rect 3516 26308 3568 26314
rect 3516 26250 3568 26256
rect 3054 25936 3110 25945
rect 3054 25871 3110 25880
rect 3620 25702 3648 27520
rect 4066 27160 4122 27169
rect 4172 27146 4200 27520
rect 4172 27118 4660 27146
rect 4066 27095 4122 27104
rect 4080 27010 4108 27095
rect 4080 26982 4384 27010
rect 4066 26480 4122 26489
rect 4122 26438 4200 26466
rect 4066 26415 4122 26424
rect 3608 25696 3660 25702
rect 3608 25638 3660 25644
rect 3882 25664 3938 25673
rect 3882 25599 3938 25608
rect 3424 25356 3476 25362
rect 3424 25298 3476 25304
rect 2964 25220 3016 25226
rect 2964 25162 3016 25168
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 2332 24806 2544 24834
rect 2044 24608 2096 24614
rect 2042 24576 2044 24585
rect 2096 24576 2098 24585
rect 2042 24511 2098 24520
rect 2042 24440 2098 24449
rect 2042 24375 2044 24384
rect 2096 24375 2098 24384
rect 2044 24346 2096 24352
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 2056 23662 2084 24346
rect 2332 24177 2360 24806
rect 2596 24744 2648 24750
rect 2596 24686 2648 24692
rect 2412 24608 2464 24614
rect 2412 24550 2464 24556
rect 2318 24168 2374 24177
rect 2318 24103 2374 24112
rect 2044 23656 2096 23662
rect 2044 23598 2096 23604
rect 2424 23594 2452 24550
rect 2504 24268 2556 24274
rect 2504 24210 2556 24216
rect 2516 23866 2544 24210
rect 2504 23860 2556 23866
rect 2504 23802 2556 23808
rect 2412 23588 2464 23594
rect 2412 23530 2464 23536
rect 2608 23254 2636 24686
rect 2688 24608 2740 24614
rect 2688 24550 2740 24556
rect 2700 23497 2728 24550
rect 2884 24041 2912 25094
rect 2870 24032 2926 24041
rect 2870 23967 2926 23976
rect 2872 23656 2924 23662
rect 2872 23598 2924 23604
rect 2686 23488 2742 23497
rect 2686 23423 2742 23432
rect 2884 23322 2912 23598
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 2596 23248 2648 23254
rect 2596 23190 2648 23196
rect 2504 23180 2556 23186
rect 2504 23122 2556 23128
rect 2516 22710 2544 23122
rect 2504 22704 2556 22710
rect 2504 22646 2556 22652
rect 2884 22642 2912 23258
rect 2976 22817 3004 25162
rect 3436 24614 3464 25298
rect 3790 25256 3846 25265
rect 3790 25191 3846 25200
rect 3804 24954 3832 25191
rect 3896 24954 3924 25599
rect 4172 25498 4200 26438
rect 4252 26036 4304 26042
rect 4252 25978 4304 25984
rect 4160 25492 4212 25498
rect 4160 25434 4212 25440
rect 3792 24948 3844 24954
rect 3792 24890 3844 24896
rect 3884 24948 3936 24954
rect 3884 24890 3936 24896
rect 4264 24818 4292 25978
rect 4356 25498 4384 26982
rect 4344 25492 4396 25498
rect 4344 25434 4396 25440
rect 4528 25356 4580 25362
rect 4528 25298 4580 25304
rect 4252 24812 4304 24818
rect 4252 24754 4304 24760
rect 4160 24744 4212 24750
rect 4160 24686 4212 24692
rect 4250 24712 4306 24721
rect 3424 24608 3476 24614
rect 3424 24550 3476 24556
rect 3056 23520 3108 23526
rect 3056 23462 3108 23468
rect 2962 22808 3018 22817
rect 2962 22743 3018 22752
rect 2872 22636 2924 22642
rect 2872 22578 2924 22584
rect 2044 22568 2096 22574
rect 2044 22510 2096 22516
rect 1766 22264 1822 22273
rect 1766 22199 1822 22208
rect 1858 22128 1914 22137
rect 1858 22063 1914 22072
rect 1872 21690 1900 22063
rect 1860 21684 1912 21690
rect 1860 21626 1912 21632
rect 2056 21146 2084 22510
rect 2962 22264 3018 22273
rect 2780 22228 2832 22234
rect 2700 22188 2780 22216
rect 2228 22160 2280 22166
rect 2228 22102 2280 22108
rect 2044 21140 2096 21146
rect 2044 21082 2096 21088
rect 1860 21004 1912 21010
rect 1860 20946 1912 20952
rect 1872 20806 1900 20946
rect 1860 20800 1912 20806
rect 1860 20742 1912 20748
rect 1674 20088 1730 20097
rect 1674 20023 1730 20032
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1780 19394 1808 19858
rect 1872 19514 1900 20742
rect 2240 20058 2268 22102
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 2332 21554 2360 22034
rect 2596 21956 2648 21962
rect 2596 21898 2648 21904
rect 2412 21888 2464 21894
rect 2412 21830 2464 21836
rect 2320 21548 2372 21554
rect 2320 21490 2372 21496
rect 2332 20398 2360 21490
rect 2424 21185 2452 21830
rect 2608 21486 2636 21898
rect 2700 21690 2728 22188
rect 2962 22199 2964 22208
rect 2780 22170 2832 22176
rect 3016 22199 3018 22208
rect 2964 22170 3016 22176
rect 2872 22160 2924 22166
rect 2870 22128 2872 22137
rect 2924 22128 2926 22137
rect 2870 22063 2926 22072
rect 2688 21684 2740 21690
rect 2688 21626 2740 21632
rect 2596 21480 2648 21486
rect 2596 21422 2648 21428
rect 2688 21344 2740 21350
rect 2608 21292 2688 21298
rect 2608 21286 2740 21292
rect 2608 21270 2728 21286
rect 2410 21176 2466 21185
rect 2410 21111 2466 21120
rect 2608 20942 2636 21270
rect 2964 21140 3016 21146
rect 2964 21082 3016 21088
rect 2596 20936 2648 20942
rect 2596 20878 2648 20884
rect 2608 20602 2636 20878
rect 2596 20596 2648 20602
rect 2596 20538 2648 20544
rect 2320 20392 2372 20398
rect 2320 20334 2372 20340
rect 2412 20324 2464 20330
rect 2412 20266 2464 20272
rect 2228 20052 2280 20058
rect 2148 20012 2228 20040
rect 1860 19508 1912 19514
rect 1860 19450 1912 19456
rect 1780 19366 1900 19394
rect 1872 19174 1900 19366
rect 1860 19168 1912 19174
rect 1860 19110 1912 19116
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1308 17808 1360 17814
rect 1308 17750 1360 17756
rect 202 15872 258 15881
rect 202 15807 258 15816
rect 1320 10033 1348 17750
rect 1688 16794 1716 17818
rect 1768 17536 1820 17542
rect 1768 17478 1820 17484
rect 1780 17241 1808 17478
rect 1766 17232 1822 17241
rect 1766 17167 1822 17176
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1872 16436 1900 19110
rect 2148 18902 2176 20012
rect 2228 19994 2280 20000
rect 2424 19854 2452 20266
rect 2976 20058 3004 21082
rect 3068 21049 3096 23462
rect 3148 22432 3200 22438
rect 3148 22374 3200 22380
rect 3160 22098 3188 22374
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 3240 22024 3292 22030
rect 3240 21966 3292 21972
rect 3252 21078 3280 21966
rect 3240 21072 3292 21078
rect 3054 21040 3110 21049
rect 3240 21014 3292 21020
rect 3054 20975 3110 20984
rect 3252 20398 3280 21014
rect 3240 20392 3292 20398
rect 3240 20334 3292 20340
rect 2964 20052 3016 20058
rect 2964 19994 3016 20000
rect 2412 19848 2464 19854
rect 2412 19790 2464 19796
rect 2228 19712 2280 19718
rect 2228 19654 2280 19660
rect 2240 19242 2268 19654
rect 2424 19310 2452 19790
rect 2320 19304 2372 19310
rect 2320 19246 2372 19252
rect 2412 19304 2464 19310
rect 2596 19304 2648 19310
rect 2412 19246 2464 19252
rect 2594 19272 2596 19281
rect 2648 19272 2650 19281
rect 2228 19236 2280 19242
rect 2228 19178 2280 19184
rect 2332 18970 2360 19246
rect 2594 19207 2650 19216
rect 2502 19000 2558 19009
rect 2320 18964 2372 18970
rect 2502 18935 2504 18944
rect 2320 18906 2372 18912
rect 2556 18935 2558 18944
rect 2504 18906 2556 18912
rect 2136 18896 2188 18902
rect 2136 18838 2188 18844
rect 2412 18828 2464 18834
rect 2412 18770 2464 18776
rect 2136 18692 2188 18698
rect 2136 18634 2188 18640
rect 2148 18290 2176 18634
rect 2136 18284 2188 18290
rect 2136 18226 2188 18232
rect 2044 18148 2096 18154
rect 2044 18090 2096 18096
rect 2056 17746 2084 18090
rect 2044 17740 2096 17746
rect 2044 17682 2096 17688
rect 2056 17354 2084 17682
rect 1964 17326 2084 17354
rect 1964 16590 1992 17326
rect 2148 17218 2176 18226
rect 2424 18068 2452 18770
rect 2516 18426 2544 18906
rect 2608 18766 2636 19207
rect 2596 18760 2648 18766
rect 2596 18702 2648 18708
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 2688 18624 2740 18630
rect 2688 18566 2740 18572
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 2596 18080 2648 18086
rect 2424 18040 2596 18068
rect 2596 18022 2648 18028
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 2332 17338 2360 17614
rect 2320 17332 2372 17338
rect 2320 17274 2372 17280
rect 2056 17190 2176 17218
rect 2056 17134 2084 17190
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 2136 16652 2188 16658
rect 2136 16594 2188 16600
rect 2504 16652 2556 16658
rect 2504 16594 2556 16600
rect 1952 16584 2004 16590
rect 1952 16526 2004 16532
rect 1872 16408 1992 16436
rect 1582 16144 1638 16153
rect 1582 16079 1638 16088
rect 1490 15464 1546 15473
rect 1490 15399 1546 15408
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1412 13802 1440 14350
rect 1400 13796 1452 13802
rect 1400 13738 1452 13744
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 11218 1440 13262
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1306 10024 1362 10033
rect 1306 9959 1362 9968
rect 1504 9518 1532 15399
rect 1596 10266 1624 16079
rect 1676 15972 1728 15978
rect 1676 15914 1728 15920
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1688 10130 1716 15914
rect 1766 15600 1822 15609
rect 1766 15535 1768 15544
rect 1820 15535 1822 15544
rect 1860 15564 1912 15570
rect 1768 15506 1820 15512
rect 1860 15506 1912 15512
rect 1780 15026 1808 15506
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1872 14074 1900 15506
rect 1964 15502 1992 16408
rect 2056 15706 2084 16594
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 1952 15496 2004 15502
rect 1952 15438 2004 15444
rect 2148 15162 2176 16594
rect 2516 16250 2544 16594
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 2608 16130 2636 18022
rect 2700 17882 2728 18566
rect 2792 17882 2820 18702
rect 2872 18080 2924 18086
rect 2872 18022 2924 18028
rect 2688 17876 2740 17882
rect 2688 17818 2740 17824
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2688 17740 2740 17746
rect 2688 17682 2740 17688
rect 2700 16250 2728 17682
rect 2884 17678 2912 18022
rect 3238 17912 3294 17921
rect 3238 17847 3294 17856
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 2780 17060 2832 17066
rect 2780 17002 2832 17008
rect 2792 16590 2820 17002
rect 3160 16794 3188 17478
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 2792 16182 2820 16526
rect 2516 16102 2636 16130
rect 2780 16176 2832 16182
rect 2780 16118 2832 16124
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2424 15502 2452 15642
rect 2228 15496 2280 15502
rect 2228 15438 2280 15444
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2136 15156 2188 15162
rect 2136 15098 2188 15104
rect 2240 14804 2268 15438
rect 2424 15094 2452 15438
rect 2412 15088 2464 15094
rect 2412 15030 2464 15036
rect 2320 14816 2372 14822
rect 2240 14776 2320 14804
rect 2320 14758 2372 14764
rect 1952 14544 2004 14550
rect 1952 14486 2004 14492
rect 1860 14068 1912 14074
rect 1860 14010 1912 14016
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 1872 11354 1900 13806
rect 1964 13734 1992 14486
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1964 13530 1992 13670
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2240 12850 2268 13126
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 2148 12442 2176 12582
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2148 12238 2176 12378
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2240 11898 2268 12786
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1872 11082 1900 11290
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1964 10470 1992 11086
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1582 9480 1638 9489
rect 1582 9415 1638 9424
rect 1596 9382 1624 9415
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1688 9178 1716 10066
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 570 4584 626 4593
rect 570 4519 626 4528
rect 584 4282 612 4519
rect 572 4276 624 4282
rect 572 4218 624 4224
rect 940 3732 992 3738
rect 940 3674 992 3680
rect 952 921 980 3674
rect 1964 3233 1992 10406
rect 2056 10266 2084 11154
rect 2332 11150 2360 14758
rect 2516 13530 2544 16102
rect 2792 15706 2820 16118
rect 3252 15706 3280 17847
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 3344 16658 3372 16934
rect 3332 16652 3384 16658
rect 3332 16594 3384 16600
rect 3344 16114 3372 16594
rect 3332 16108 3384 16114
rect 3332 16050 3384 16056
rect 3332 15972 3384 15978
rect 3332 15914 3384 15920
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 3344 15366 3372 15914
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 3252 14958 3280 15302
rect 3240 14952 3292 14958
rect 3240 14894 3292 14900
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2792 14226 2820 14554
rect 2700 14198 2820 14226
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2608 12306 2636 13670
rect 2700 12850 2728 14198
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2792 12646 2820 13466
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 2870 13152 2926 13161
rect 2870 13087 2926 13096
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2792 12458 2820 12582
rect 2700 12430 2820 12458
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 2424 11354 2452 12242
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2516 11286 2544 12174
rect 2608 11898 2636 12242
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2608 11762 2636 11834
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2516 10810 2544 11222
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2700 10538 2728 12430
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2792 11626 2820 12038
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2688 10532 2740 10538
rect 2688 10474 2740 10480
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 2884 10146 2912 13087
rect 2976 12374 3004 13262
rect 3068 12986 3096 13330
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 2964 12368 3016 12374
rect 2964 12310 3016 12316
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 2976 11762 3004 12038
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2976 11218 3004 11698
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 3056 11008 3108 11014
rect 3056 10950 3108 10956
rect 3068 10674 3096 10950
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2608 10124 2912 10146
rect 2608 10118 2688 10124
rect 2608 9722 2636 10118
rect 2740 10118 2912 10124
rect 2688 10066 2740 10072
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2778 4040 2834 4049
rect 2778 3975 2834 3984
rect 1950 3224 2006 3233
rect 1950 3159 2006 3168
rect 1308 2916 1360 2922
rect 1308 2858 1360 2864
rect 938 912 994 921
rect 938 847 994 856
rect 1320 377 1348 2858
rect 2792 480 2820 3975
rect 2976 3738 3004 10474
rect 3068 10266 3096 10610
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3160 2825 3188 14758
rect 3252 14618 3280 14894
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3344 12986 3372 15302
rect 3436 13938 3464 24550
rect 4172 24290 4200 24686
rect 4250 24647 4306 24656
rect 4264 24410 4292 24647
rect 4540 24614 4568 25298
rect 4632 24698 4660 27118
rect 4724 25242 4752 27520
rect 5172 25356 5224 25362
rect 5172 25298 5224 25304
rect 4724 25214 4844 25242
rect 4712 25152 4764 25158
rect 4712 25094 4764 25100
rect 4724 24886 4752 25094
rect 4712 24880 4764 24886
rect 4712 24822 4764 24828
rect 4816 24818 4844 25214
rect 4804 24812 4856 24818
rect 4804 24754 4856 24760
rect 4632 24670 4844 24698
rect 4528 24608 4580 24614
rect 4528 24550 4580 24556
rect 4252 24404 4304 24410
rect 4252 24346 4304 24352
rect 4068 24268 4120 24274
rect 4172 24262 4292 24290
rect 4068 24210 4120 24216
rect 4080 23798 4108 24210
rect 4068 23792 4120 23798
rect 4068 23734 4120 23740
rect 3792 23724 3844 23730
rect 3792 23666 3844 23672
rect 3606 23488 3662 23497
rect 3606 23423 3662 23432
rect 3620 22166 3648 23423
rect 3700 22976 3752 22982
rect 3700 22918 3752 22924
rect 3712 22438 3740 22918
rect 3700 22432 3752 22438
rect 3700 22374 3752 22380
rect 3608 22160 3660 22166
rect 3608 22102 3660 22108
rect 3804 22030 3832 23666
rect 3884 23180 3936 23186
rect 3884 23122 3936 23128
rect 3896 22386 3924 23122
rect 3976 23112 4028 23118
rect 3976 23054 4028 23060
rect 3988 22574 4016 23054
rect 4160 22636 4212 22642
rect 4160 22578 4212 22584
rect 3976 22568 4028 22574
rect 3976 22510 4028 22516
rect 3896 22358 4016 22386
rect 3988 22166 4016 22358
rect 4172 22234 4200 22578
rect 4160 22228 4212 22234
rect 4160 22170 4212 22176
rect 3884 22160 3936 22166
rect 3884 22102 3936 22108
rect 3976 22160 4028 22166
rect 3976 22102 4028 22108
rect 3792 22024 3844 22030
rect 3792 21966 3844 21972
rect 3608 21480 3660 21486
rect 3608 21422 3660 21428
rect 3620 20942 3648 21422
rect 3608 20936 3660 20942
rect 3608 20878 3660 20884
rect 3516 20800 3568 20806
rect 3516 20742 3568 20748
rect 3528 19922 3556 20742
rect 3620 20602 3648 20878
rect 3608 20596 3660 20602
rect 3608 20538 3660 20544
rect 3516 19916 3568 19922
rect 3516 19858 3568 19864
rect 3620 19446 3648 20538
rect 3608 19440 3660 19446
rect 3608 19382 3660 19388
rect 3698 19136 3754 19145
rect 3698 19071 3754 19080
rect 3608 18896 3660 18902
rect 3608 18838 3660 18844
rect 3620 18698 3648 18838
rect 3608 18692 3660 18698
rect 3608 18634 3660 18640
rect 3514 18048 3570 18057
rect 3514 17983 3570 17992
rect 3528 16794 3556 17983
rect 3620 17746 3648 18634
rect 3608 17740 3660 17746
rect 3608 17682 3660 17688
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3528 16182 3556 16730
rect 3516 16176 3568 16182
rect 3516 16118 3568 16124
rect 3606 15600 3662 15609
rect 3606 15535 3662 15544
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3528 12782 3556 14214
rect 3620 13512 3648 15535
rect 3712 14929 3740 19071
rect 3790 18592 3846 18601
rect 3790 18527 3846 18536
rect 3804 16153 3832 18527
rect 3896 16794 3924 22102
rect 3976 20800 4028 20806
rect 3976 20742 4028 20748
rect 3988 20505 4016 20742
rect 3974 20496 4030 20505
rect 3974 20431 4030 20440
rect 3974 19816 4030 19825
rect 3974 19751 4030 19760
rect 3988 17921 4016 19751
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 4172 18902 4200 19246
rect 4160 18896 4212 18902
rect 4160 18838 4212 18844
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 3974 17912 4030 17921
rect 3974 17847 4030 17856
rect 4080 17728 4108 18022
rect 4160 17740 4212 17746
rect 4080 17700 4160 17728
rect 4160 17682 4212 17688
rect 4172 17338 4200 17682
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 4264 17218 4292 24262
rect 4436 23520 4488 23526
rect 4436 23462 4488 23468
rect 4344 22092 4396 22098
rect 4344 22034 4396 22040
rect 4356 21350 4384 22034
rect 4344 21344 4396 21350
rect 4344 21286 4396 21292
rect 4448 21078 4476 23462
rect 4540 22817 4568 24550
rect 4526 22808 4582 22817
rect 4526 22743 4582 22752
rect 4540 21298 4568 22743
rect 4540 21270 4752 21298
rect 4526 21176 4582 21185
rect 4526 21111 4528 21120
rect 4580 21111 4582 21120
rect 4528 21082 4580 21088
rect 4436 21072 4488 21078
rect 4356 21032 4436 21060
rect 4356 19854 4384 21032
rect 4436 21014 4488 21020
rect 4540 20584 4568 21082
rect 4448 20556 4568 20584
rect 4448 20058 4476 20556
rect 4724 20482 4752 21270
rect 4528 20460 4580 20466
rect 4528 20402 4580 20408
rect 4632 20454 4752 20482
rect 4540 20262 4568 20402
rect 4528 20256 4580 20262
rect 4528 20198 4580 20204
rect 4436 20052 4488 20058
rect 4436 19994 4488 20000
rect 4540 19990 4568 20198
rect 4528 19984 4580 19990
rect 4528 19926 4580 19932
rect 4344 19848 4396 19854
rect 4344 19790 4396 19796
rect 4540 19514 4568 19926
rect 4528 19508 4580 19514
rect 4528 19450 4580 19456
rect 4528 19236 4580 19242
rect 4528 19178 4580 19184
rect 4540 18970 4568 19178
rect 4528 18964 4580 18970
rect 4528 18906 4580 18912
rect 4264 17190 4384 17218
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3790 16144 3846 16153
rect 3790 16079 3846 16088
rect 3792 15904 3844 15910
rect 3792 15846 3844 15852
rect 3698 14920 3754 14929
rect 3698 14855 3754 14864
rect 3804 13870 3832 15846
rect 3792 13864 3844 13870
rect 3792 13806 3844 13812
rect 3790 13696 3846 13705
rect 3790 13631 3846 13640
rect 3804 13530 3832 13631
rect 3792 13524 3844 13530
rect 3620 13484 3740 13512
rect 3712 13410 3740 13484
rect 3792 13466 3844 13472
rect 3608 13388 3660 13394
rect 3712 13382 3832 13410
rect 3608 13330 3660 13336
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3528 11898 3556 12718
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3146 2816 3202 2825
rect 3146 2751 3202 2760
rect 3344 2145 3372 10406
rect 3528 2922 3556 11494
rect 3620 11082 3648 13330
rect 3700 13184 3752 13190
rect 3700 13126 3752 13132
rect 3712 12646 3740 13126
rect 3700 12640 3752 12646
rect 3698 12608 3700 12617
rect 3752 12608 3754 12617
rect 3698 12543 3754 12552
rect 3608 11076 3660 11082
rect 3608 11018 3660 11024
rect 3620 6202 3648 11018
rect 3804 10470 3832 13382
rect 3896 12850 3924 16526
rect 4252 15904 4304 15910
rect 4252 15846 4304 15852
rect 4066 15056 4122 15065
rect 4066 14991 4122 15000
rect 4080 14385 4108 14991
rect 4066 14376 4122 14385
rect 4066 14311 4122 14320
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 3988 13530 4016 14010
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 3976 13388 4028 13394
rect 3976 13330 4028 13336
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3896 12442 3924 12786
rect 3988 12714 4016 13330
rect 3976 12708 4028 12714
rect 3976 12650 4028 12656
rect 3988 12442 4016 12650
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 4264 12238 4292 15846
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 3974 11656 4030 11665
rect 3974 11591 4030 11600
rect 4068 11620 4120 11626
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3698 10160 3754 10169
rect 3698 10095 3754 10104
rect 3712 6361 3740 10095
rect 3882 9072 3938 9081
rect 3882 9007 3938 9016
rect 3896 7041 3924 9007
rect 3882 7032 3938 7041
rect 3882 6967 3938 6976
rect 3698 6352 3754 6361
rect 3698 6287 3754 6296
rect 3620 6174 3740 6202
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3330 2136 3386 2145
rect 3330 2071 3386 2080
rect 3712 1465 3740 6174
rect 3988 5137 4016 11591
rect 4068 11562 4120 11568
rect 4080 11354 4108 11562
rect 4264 11558 4292 12174
rect 4356 11762 4384 17190
rect 4436 17128 4488 17134
rect 4436 17070 4488 17076
rect 4448 15162 4476 17070
rect 4526 16824 4582 16833
rect 4526 16759 4582 16768
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 4540 14618 4568 16759
rect 4632 16250 4660 20454
rect 4712 20392 4764 20398
rect 4712 20334 4764 20340
rect 4724 18426 4752 20334
rect 4816 19145 4844 24670
rect 5184 24614 5212 25298
rect 5172 24608 5224 24614
rect 5172 24550 5224 24556
rect 5184 24154 5212 24550
rect 5276 24313 5304 27520
rect 5828 25242 5856 27520
rect 6184 25356 6236 25362
rect 6184 25298 6236 25304
rect 5828 25214 6132 25242
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5356 24812 5408 24818
rect 5356 24754 5408 24760
rect 5262 24304 5318 24313
rect 5262 24239 5318 24248
rect 5184 24126 5304 24154
rect 4896 24064 4948 24070
rect 4896 24006 4948 24012
rect 4908 23662 4936 24006
rect 5080 23792 5132 23798
rect 5080 23734 5132 23740
rect 4896 23656 4948 23662
rect 4894 23624 4896 23633
rect 4948 23624 4950 23633
rect 4894 23559 4950 23568
rect 4896 23520 4948 23526
rect 4896 23462 4948 23468
rect 4908 22982 4936 23462
rect 5092 23338 5120 23734
rect 5172 23656 5224 23662
rect 5172 23598 5224 23604
rect 5000 23310 5120 23338
rect 4896 22976 4948 22982
rect 4896 22918 4948 22924
rect 4908 21593 4936 22918
rect 4894 21584 4950 21593
rect 4894 21519 4950 21528
rect 4802 19136 4858 19145
rect 4802 19071 4858 19080
rect 4712 18420 4764 18426
rect 4712 18362 4764 18368
rect 5000 18170 5028 23310
rect 5184 23186 5212 23598
rect 5172 23180 5224 23186
rect 5172 23122 5224 23128
rect 5276 22545 5304 24126
rect 5262 22536 5318 22545
rect 5262 22471 5318 22480
rect 5080 22432 5132 22438
rect 5080 22374 5132 22380
rect 5092 21690 5120 22374
rect 5080 21684 5132 21690
rect 5080 21626 5132 21632
rect 5172 21344 5224 21350
rect 5172 21286 5224 21292
rect 5184 21146 5212 21286
rect 5172 21140 5224 21146
rect 5172 21082 5224 21088
rect 5184 20584 5212 21082
rect 5092 20556 5212 20584
rect 5092 18306 5120 20556
rect 5170 20496 5226 20505
rect 5170 20431 5226 20440
rect 5184 20262 5212 20431
rect 5172 20256 5224 20262
rect 5172 20198 5224 20204
rect 5276 19009 5304 22471
rect 5368 19122 5396 24754
rect 5540 24268 5592 24274
rect 5540 24210 5592 24216
rect 5552 23526 5580 24210
rect 6000 24064 6052 24070
rect 6000 24006 6052 24012
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 6012 23662 6040 24006
rect 6000 23656 6052 23662
rect 6000 23598 6052 23604
rect 5540 23520 5592 23526
rect 5540 23462 5592 23468
rect 5552 23322 5580 23462
rect 6104 23361 6132 25214
rect 6196 24614 6224 25298
rect 6184 24608 6236 24614
rect 6184 24550 6236 24556
rect 6196 23497 6224 24550
rect 6182 23488 6238 23497
rect 6182 23423 6238 23432
rect 6090 23352 6146 23361
rect 5540 23316 5592 23322
rect 6090 23287 6146 23296
rect 5540 23258 5592 23264
rect 5448 23248 5500 23254
rect 5448 23190 5500 23196
rect 5460 22778 5488 23190
rect 5448 22772 5500 22778
rect 5448 22714 5500 22720
rect 5460 22234 5488 22714
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 5460 21554 5488 22170
rect 5552 22166 5580 23258
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 6274 22672 6330 22681
rect 6274 22607 6330 22616
rect 6000 22500 6052 22506
rect 6000 22442 6052 22448
rect 6012 22234 6040 22442
rect 6000 22228 6052 22234
rect 6000 22170 6052 22176
rect 5540 22160 5592 22166
rect 5540 22102 5592 22108
rect 5552 21622 5580 22102
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5540 21616 5592 21622
rect 5540 21558 5592 21564
rect 5448 21548 5500 21554
rect 5448 21490 5500 21496
rect 5460 21146 5488 21490
rect 5448 21140 5500 21146
rect 5448 21082 5500 21088
rect 6092 20936 6144 20942
rect 6092 20878 6144 20884
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5448 20392 5500 20398
rect 5552 20380 5580 20742
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6104 20602 6132 20878
rect 6184 20800 6236 20806
rect 6184 20742 6236 20748
rect 6092 20596 6144 20602
rect 6092 20538 6144 20544
rect 5500 20352 5580 20380
rect 5448 20334 5500 20340
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 5368 19094 5488 19122
rect 5262 19000 5318 19009
rect 5262 18935 5318 18944
rect 5356 18964 5408 18970
rect 5356 18906 5408 18912
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 5092 18278 5212 18306
rect 4816 18142 5028 18170
rect 5080 18148 5132 18154
rect 4712 16448 4764 16454
rect 4712 16390 4764 16396
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4724 15434 4752 16390
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4436 14476 4488 14482
rect 4436 14418 4488 14424
rect 4448 14074 4476 14418
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4448 13258 4476 13670
rect 4540 13530 4568 14554
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4632 14006 4660 14350
rect 4620 14000 4672 14006
rect 4620 13942 4672 13948
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4436 13252 4488 13258
rect 4436 13194 4488 13200
rect 4724 12986 4752 15098
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4528 12368 4580 12374
rect 4528 12310 4580 12316
rect 4540 11762 4568 12310
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4710 11384 4766 11393
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4160 11348 4212 11354
rect 4816 11354 4844 18142
rect 5080 18090 5132 18096
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 5000 16250 5028 18022
rect 5092 17338 5120 18090
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 5184 15586 5212 18278
rect 5276 18222 5304 18770
rect 5368 18290 5396 18906
rect 5356 18284 5408 18290
rect 5356 18226 5408 18232
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 5276 17542 5304 18158
rect 5264 17536 5316 17542
rect 5264 17478 5316 17484
rect 5276 17202 5304 17478
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 5276 16046 5304 17138
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 4908 15558 5212 15586
rect 4908 13326 4936 15558
rect 5172 15496 5224 15502
rect 5172 15438 5224 15444
rect 5080 15360 5132 15366
rect 5080 15302 5132 15308
rect 4986 13832 5042 13841
rect 4986 13767 5042 13776
rect 5000 13462 5028 13767
rect 5092 13705 5120 15302
rect 5184 14822 5212 15438
rect 5264 15428 5316 15434
rect 5264 15370 5316 15376
rect 5276 15026 5304 15370
rect 5368 15094 5396 16594
rect 5460 15745 5488 19094
rect 5552 18426 5580 20198
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6012 19281 6040 19654
rect 6092 19508 6144 19514
rect 6092 19450 6144 19456
rect 5998 19272 6054 19281
rect 5998 19207 6054 19216
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 6104 16674 6132 19450
rect 6196 19310 6224 20742
rect 6184 19304 6236 19310
rect 6288 19281 6316 22607
rect 6380 22137 6408 27520
rect 6642 24032 6698 24041
rect 6642 23967 6698 23976
rect 6656 23798 6684 23967
rect 6644 23792 6696 23798
rect 6644 23734 6696 23740
rect 6736 23656 6788 23662
rect 6736 23598 6788 23604
rect 6748 22574 6776 23598
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 6736 22568 6788 22574
rect 6736 22510 6788 22516
rect 6460 22432 6512 22438
rect 6460 22374 6512 22380
rect 6472 22234 6500 22374
rect 6460 22228 6512 22234
rect 6460 22170 6512 22176
rect 6840 22216 6868 23462
rect 6932 23338 6960 27520
rect 7576 25378 7604 27520
rect 7208 25350 7604 25378
rect 7932 25356 7984 25362
rect 7104 25152 7156 25158
rect 7104 25094 7156 25100
rect 7116 24750 7144 25094
rect 7104 24744 7156 24750
rect 7104 24686 7156 24692
rect 7012 24608 7064 24614
rect 7012 24550 7064 24556
rect 7024 24449 7052 24550
rect 7010 24440 7066 24449
rect 7010 24375 7066 24384
rect 7104 24064 7156 24070
rect 7104 24006 7156 24012
rect 6932 23310 7052 23338
rect 6920 22228 6972 22234
rect 6840 22188 6920 22216
rect 6366 22128 6422 22137
rect 6366 22063 6422 22072
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6460 21888 6512 21894
rect 6460 21830 6512 21836
rect 6472 21298 6500 21830
rect 6564 21622 6592 21966
rect 6840 21690 6868 22188
rect 6920 22170 6972 22176
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 6552 21616 6604 21622
rect 6552 21558 6604 21564
rect 7024 21321 7052 23310
rect 7116 22506 7144 24006
rect 7104 22500 7156 22506
rect 7104 22442 7156 22448
rect 7104 22228 7156 22234
rect 7104 22170 7156 22176
rect 7116 21690 7144 22170
rect 7104 21684 7156 21690
rect 7104 21626 7156 21632
rect 7010 21312 7066 21321
rect 6472 21270 6592 21298
rect 6458 21176 6514 21185
rect 6458 21111 6460 21120
rect 6512 21111 6514 21120
rect 6460 21082 6512 21088
rect 6472 20602 6500 21082
rect 6460 20596 6512 20602
rect 6460 20538 6512 20544
rect 6368 20460 6420 20466
rect 6368 20402 6420 20408
rect 6380 19922 6408 20402
rect 6564 20398 6592 21270
rect 7010 21247 7066 21256
rect 7024 21010 7052 21247
rect 7012 21004 7064 21010
rect 7012 20946 7064 20952
rect 6644 20936 6696 20942
rect 6644 20878 6696 20884
rect 6552 20392 6604 20398
rect 6552 20334 6604 20340
rect 6564 19922 6592 20334
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6552 19916 6604 19922
rect 6552 19858 6604 19864
rect 6184 19246 6236 19252
rect 6274 19272 6330 19281
rect 6274 19207 6330 19216
rect 6380 18902 6408 19858
rect 6656 19854 6684 20878
rect 6734 20496 6790 20505
rect 6734 20431 6790 20440
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 6552 19712 6604 19718
rect 6552 19654 6604 19660
rect 6564 19174 6592 19654
rect 6748 19174 6776 20431
rect 6828 20392 6880 20398
rect 6826 20360 6828 20369
rect 6880 20360 6882 20369
rect 6826 20295 6882 20304
rect 7012 19780 7064 19786
rect 7012 19722 7064 19728
rect 7024 19378 7052 19722
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 6552 19168 6604 19174
rect 6552 19110 6604 19116
rect 6736 19168 6788 19174
rect 6736 19110 6788 19116
rect 6368 18896 6420 18902
rect 6368 18838 6420 18844
rect 6380 17882 6408 18838
rect 6564 18834 6592 19110
rect 7024 18986 7052 19314
rect 7116 19310 7144 19654
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 6840 18970 7052 18986
rect 7116 18970 7144 19246
rect 6828 18964 7052 18970
rect 6880 18958 7052 18964
rect 7104 18964 7156 18970
rect 6828 18906 6880 18912
rect 7104 18906 7156 18912
rect 6552 18828 6604 18834
rect 6552 18770 6604 18776
rect 7208 18426 7236 25350
rect 7932 25298 7984 25304
rect 7748 25288 7800 25294
rect 7748 25230 7800 25236
rect 7380 25220 7432 25226
rect 7380 25162 7432 25168
rect 7392 24818 7420 25162
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 7286 23896 7342 23905
rect 7392 23866 7420 24754
rect 7760 24070 7788 25230
rect 7840 24880 7892 24886
rect 7840 24822 7892 24828
rect 7748 24064 7800 24070
rect 7748 24006 7800 24012
rect 7286 23831 7342 23840
rect 7380 23860 7432 23866
rect 7300 23730 7328 23831
rect 7380 23802 7432 23808
rect 7288 23724 7340 23730
rect 7288 23666 7340 23672
rect 7472 23724 7524 23730
rect 7472 23666 7524 23672
rect 7288 23588 7340 23594
rect 7288 23530 7340 23536
rect 7300 19446 7328 23530
rect 7380 23520 7432 23526
rect 7378 23488 7380 23497
rect 7432 23488 7434 23497
rect 7378 23423 7434 23432
rect 7484 23118 7512 23666
rect 7472 23112 7524 23118
rect 7472 23054 7524 23060
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7484 22234 7512 22918
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7668 21894 7696 22510
rect 7656 21888 7708 21894
rect 7576 21848 7656 21876
rect 7576 21554 7604 21848
rect 7656 21830 7708 21836
rect 7564 21548 7616 21554
rect 7564 21490 7616 21496
rect 7576 20466 7604 21490
rect 7656 21480 7708 21486
rect 7656 21422 7708 21428
rect 7668 21146 7696 21422
rect 7656 21140 7708 21146
rect 7656 21082 7708 21088
rect 7564 20460 7616 20466
rect 7564 20402 7616 20408
rect 7852 20262 7880 24822
rect 7944 24614 7972 25298
rect 7932 24608 7984 24614
rect 7932 24550 7984 24556
rect 7944 23594 7972 24550
rect 7932 23588 7984 23594
rect 7932 23530 7984 23536
rect 8022 23352 8078 23361
rect 8022 23287 8024 23296
rect 8076 23287 8078 23296
rect 8024 23258 8076 23264
rect 7932 23180 7984 23186
rect 7932 23122 7984 23128
rect 7944 22817 7972 23122
rect 8036 22953 8064 23258
rect 8022 22944 8078 22953
rect 8022 22879 8078 22888
rect 7930 22808 7986 22817
rect 7930 22743 7986 22752
rect 7944 22234 7972 22743
rect 7932 22228 7984 22234
rect 7932 22170 7984 22176
rect 8036 22166 8064 22879
rect 8128 22409 8156 27520
rect 8680 27470 8708 27520
rect 8668 27464 8720 27470
rect 8668 27406 8720 27412
rect 8760 27464 8812 27470
rect 8760 27406 8812 27412
rect 8392 26308 8444 26314
rect 8392 26250 8444 26256
rect 8300 24064 8352 24070
rect 8300 24006 8352 24012
rect 8312 23526 8340 24006
rect 8300 23520 8352 23526
rect 8300 23462 8352 23468
rect 8208 22432 8260 22438
rect 8114 22400 8170 22409
rect 8208 22374 8260 22380
rect 8114 22335 8170 22344
rect 8024 22160 8076 22166
rect 8024 22102 8076 22108
rect 8116 22092 8168 22098
rect 8116 22034 8168 22040
rect 8128 21457 8156 22034
rect 8220 21486 8248 22374
rect 8208 21480 8260 21486
rect 8114 21448 8170 21457
rect 8208 21422 8260 21428
rect 8114 21383 8116 21392
rect 8168 21383 8170 21392
rect 8116 21354 8168 21360
rect 8128 21323 8156 21354
rect 8312 21350 8340 23462
rect 8404 21962 8432 26250
rect 8484 24608 8536 24614
rect 8484 24550 8536 24556
rect 8496 23662 8524 24550
rect 8574 24304 8630 24313
rect 8574 24239 8630 24248
rect 8484 23656 8536 23662
rect 8484 23598 8536 23604
rect 8496 23322 8524 23598
rect 8484 23316 8536 23322
rect 8484 23258 8536 23264
rect 8392 21956 8444 21962
rect 8392 21898 8444 21904
rect 8300 21344 8352 21350
rect 8300 21286 8352 21292
rect 8208 21140 8260 21146
rect 8208 21082 8260 21088
rect 8116 21072 8168 21078
rect 8116 21014 8168 21020
rect 8024 20800 8076 20806
rect 8024 20742 8076 20748
rect 7840 20256 7892 20262
rect 7840 20198 7892 20204
rect 7654 20088 7710 20097
rect 7654 20023 7710 20032
rect 7668 19990 7696 20023
rect 7656 19984 7708 19990
rect 7656 19926 7708 19932
rect 7564 19848 7616 19854
rect 7564 19790 7616 19796
rect 7288 19440 7340 19446
rect 7576 19417 7604 19790
rect 7288 19382 7340 19388
rect 7378 19408 7434 19417
rect 7562 19408 7618 19417
rect 7378 19343 7434 19352
rect 7472 19372 7524 19378
rect 7196 18420 7248 18426
rect 7196 18362 7248 18368
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 6734 17912 6790 17921
rect 6368 17876 6420 17882
rect 6734 17847 6736 17856
rect 6368 17818 6420 17824
rect 6788 17847 6790 17856
rect 6736 17818 6788 17824
rect 6644 17740 6696 17746
rect 6644 17682 6696 17688
rect 6656 16998 6684 17682
rect 6734 17232 6790 17241
rect 6734 17167 6790 17176
rect 6748 17134 6776 17167
rect 6736 17128 6788 17134
rect 6736 17070 6788 17076
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6012 16646 6132 16674
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5446 15736 5502 15745
rect 5446 15671 5502 15680
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5356 15088 5408 15094
rect 5356 15030 5408 15036
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5276 14890 5304 14962
rect 5264 14884 5316 14890
rect 5264 14826 5316 14832
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5078 13696 5134 13705
rect 5078 13631 5134 13640
rect 4988 13456 5040 13462
rect 4988 13398 5040 13404
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 5184 12442 5212 14758
rect 5276 14346 5304 14826
rect 5264 14340 5316 14346
rect 5264 14282 5316 14288
rect 5276 13258 5304 14282
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 5368 12594 5396 15030
rect 5460 14618 5488 15506
rect 5632 15496 5684 15502
rect 5552 15456 5632 15484
rect 5552 14958 5580 15456
rect 5632 15438 5684 15444
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5814 14920 5870 14929
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 5460 12986 5488 14554
rect 5552 14414 5580 14894
rect 6012 14906 6040 16646
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6104 16114 6132 16526
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6092 15632 6144 15638
rect 6092 15574 6144 15580
rect 5814 14855 5870 14864
rect 5920 14878 6040 14906
rect 5828 14822 5856 14855
rect 5816 14816 5868 14822
rect 5920 14793 5948 14878
rect 6000 14816 6052 14822
rect 5816 14758 5868 14764
rect 5906 14784 5962 14793
rect 6000 14758 6052 14764
rect 5906 14719 5962 14728
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5552 14056 5580 14350
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5552 14028 5672 14056
rect 5540 13728 5592 13734
rect 5538 13696 5540 13705
rect 5592 13696 5594 13705
rect 5538 13631 5594 13640
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 5552 12782 5580 13398
rect 5644 13394 5672 14028
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5736 13530 5764 13874
rect 5816 13864 5868 13870
rect 5816 13806 5868 13812
rect 5828 13705 5856 13806
rect 5814 13696 5870 13705
rect 5814 13631 5870 13640
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5736 12714 5764 12786
rect 5724 12708 5776 12714
rect 5724 12650 5776 12656
rect 5276 12566 5396 12594
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5276 12374 5304 12566
rect 5264 12368 5316 12374
rect 5264 12310 5316 12316
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 4710 11319 4766 11328
rect 4804 11348 4856 11354
rect 4160 11290 4212 11296
rect 4172 10810 4200 11290
rect 4724 11150 4752 11319
rect 4804 11290 4856 11296
rect 4528 11144 4580 11150
rect 4526 11112 4528 11121
rect 4712 11144 4764 11150
rect 4580 11112 4582 11121
rect 4712 11086 4764 11092
rect 4526 11047 4582 11056
rect 4540 10810 4568 11047
rect 4724 10810 4752 11086
rect 5092 11082 5120 12242
rect 5736 12238 5764 12650
rect 5724 12232 5776 12238
rect 5552 12192 5724 12220
rect 5552 11354 5580 12192
rect 5724 12174 5776 12180
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 6012 11121 6040 14758
rect 6104 13870 6132 15574
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6196 13716 6224 16934
rect 6656 16561 6684 16934
rect 6748 16794 6776 17070
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6734 16688 6790 16697
rect 6734 16623 6790 16632
rect 6642 16552 6698 16561
rect 6642 16487 6698 16496
rect 6458 15872 6514 15881
rect 6458 15807 6514 15816
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 6104 13688 6224 13716
rect 6104 12866 6132 13688
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 6196 12986 6224 13330
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6104 12838 6224 12866
rect 6288 12850 6316 14418
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6380 13802 6408 14214
rect 6368 13796 6420 13802
rect 6368 13738 6420 13744
rect 6472 12889 6500 15807
rect 6644 15564 6696 15570
rect 6644 15506 6696 15512
rect 6656 14890 6684 15506
rect 6644 14884 6696 14890
rect 6644 14826 6696 14832
rect 6748 14414 6776 16623
rect 6840 16046 6868 18022
rect 6918 17912 6974 17921
rect 6918 17847 6974 17856
rect 6932 16522 6960 17847
rect 7104 17060 7156 17066
rect 7104 17002 7156 17008
rect 7116 16697 7144 17002
rect 7102 16688 7158 16697
rect 7102 16623 7158 16632
rect 6920 16516 6972 16522
rect 6920 16458 6972 16464
rect 6918 16416 6974 16425
rect 6918 16351 6974 16360
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 6564 12986 6592 13466
rect 6748 13394 6776 14214
rect 6840 13462 6868 14758
rect 6932 13569 6960 16351
rect 7012 16176 7064 16182
rect 7010 16144 7012 16153
rect 7064 16144 7066 16153
rect 7010 16079 7066 16088
rect 7194 16144 7250 16153
rect 7194 16079 7196 16088
rect 7248 16079 7250 16088
rect 7196 16050 7248 16056
rect 7392 15065 7420 19343
rect 7562 19343 7618 19352
rect 7472 19314 7524 19320
rect 7484 15609 7512 19314
rect 7576 18902 7604 19343
rect 7668 19156 7696 19926
rect 7748 19168 7800 19174
rect 7668 19128 7748 19156
rect 7748 19110 7800 19116
rect 7564 18896 7616 18902
rect 7564 18838 7616 18844
rect 7562 16824 7618 16833
rect 7562 16759 7564 16768
rect 7616 16759 7618 16768
rect 7564 16730 7616 16736
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7668 16250 7696 16594
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7654 15736 7710 15745
rect 7654 15671 7710 15680
rect 7470 15600 7526 15609
rect 7668 15570 7696 15671
rect 7470 15535 7526 15544
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7668 15162 7696 15506
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7378 15056 7434 15065
rect 7378 14991 7434 15000
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7300 13977 7328 14758
rect 7286 13968 7342 13977
rect 7286 13903 7288 13912
rect 7340 13903 7342 13912
rect 7288 13874 7340 13880
rect 6918 13560 6974 13569
rect 6918 13495 6974 13504
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6458 12880 6514 12889
rect 6090 12608 6146 12617
rect 6090 12543 6146 12552
rect 6104 12442 6132 12543
rect 6092 12436 6144 12442
rect 6092 12378 6144 12384
rect 6196 11762 6224 12838
rect 6276 12844 6328 12850
rect 6458 12815 6514 12824
rect 6276 12786 6328 12792
rect 6840 12782 6868 13126
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6840 12442 6868 12718
rect 7392 12442 7420 14991
rect 7470 14920 7526 14929
rect 7470 14855 7526 14864
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7208 11898 7236 12242
rect 7392 11898 7420 12378
rect 7484 12306 7512 14855
rect 7760 14385 7788 19110
rect 8036 18737 8064 20742
rect 8128 20058 8156 21014
rect 8220 20602 8248 21082
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 8312 20482 8340 21286
rect 8588 21146 8616 24239
rect 8772 22114 8800 27406
rect 8944 25152 8996 25158
rect 8944 25094 8996 25100
rect 8956 24857 8984 25094
rect 8942 24848 8998 24857
rect 8942 24783 8944 24792
rect 8996 24783 8998 24792
rect 8944 24754 8996 24760
rect 8850 24712 8906 24721
rect 8850 24647 8852 24656
rect 8904 24647 8906 24656
rect 8852 24618 8904 24624
rect 9232 24342 9260 27520
rect 9678 24440 9734 24449
rect 9588 24404 9640 24410
rect 9678 24375 9680 24384
rect 9588 24346 9640 24352
rect 9732 24375 9734 24384
rect 9680 24346 9732 24352
rect 9220 24336 9272 24342
rect 9220 24278 9272 24284
rect 9496 24336 9548 24342
rect 9600 24313 9628 24346
rect 9496 24278 9548 24284
rect 9586 24304 9642 24313
rect 9036 24268 9088 24274
rect 9036 24210 9088 24216
rect 8852 24064 8904 24070
rect 8852 24006 8904 24012
rect 8864 23730 8892 24006
rect 8852 23724 8904 23730
rect 8852 23666 8904 23672
rect 9048 23118 9076 24210
rect 9036 23112 9088 23118
rect 9034 23080 9036 23089
rect 9088 23080 9090 23089
rect 9034 23015 9090 23024
rect 9312 22976 9364 22982
rect 9312 22918 9364 22924
rect 9128 22568 9180 22574
rect 9128 22510 9180 22516
rect 9140 22438 9168 22510
rect 9128 22432 9180 22438
rect 9128 22374 9180 22380
rect 9140 22137 9168 22374
rect 9126 22128 9182 22137
rect 8772 22086 8892 22114
rect 8576 21140 8628 21146
rect 8576 21082 8628 21088
rect 8220 20454 8340 20482
rect 8220 20330 8248 20454
rect 8208 20324 8260 20330
rect 8208 20266 8260 20272
rect 8116 20052 8168 20058
rect 8116 19994 8168 20000
rect 8864 19378 8892 22086
rect 9126 22063 9182 22072
rect 9324 21894 9352 22918
rect 9402 21992 9458 22001
rect 9402 21927 9458 21936
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9048 21146 9076 21830
rect 9036 21140 9088 21146
rect 9036 21082 9088 21088
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 8760 19372 8812 19378
rect 8760 19314 8812 19320
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8482 19000 8538 19009
rect 8482 18935 8484 18944
rect 8536 18935 8538 18944
rect 8484 18906 8536 18912
rect 8116 18896 8168 18902
rect 8116 18838 8168 18844
rect 8022 18728 8078 18737
rect 8022 18663 8078 18672
rect 8024 18624 8076 18630
rect 8024 18566 8076 18572
rect 8036 17882 8064 18566
rect 8128 18358 8156 18838
rect 8390 18728 8446 18737
rect 8390 18663 8446 18672
rect 8116 18352 8168 18358
rect 8116 18294 8168 18300
rect 8114 18184 8170 18193
rect 8114 18119 8170 18128
rect 8024 17876 8076 17882
rect 8024 17818 8076 17824
rect 8022 17776 8078 17785
rect 8022 17711 8078 17720
rect 8036 17610 8064 17711
rect 8024 17604 8076 17610
rect 8024 17546 8076 17552
rect 8128 17490 8156 18119
rect 8404 18086 8432 18663
rect 8496 18426 8524 18906
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8036 17462 8156 17490
rect 7840 16584 7892 16590
rect 7840 16526 7892 16532
rect 7852 15706 7880 16526
rect 7932 15972 7984 15978
rect 7932 15914 7984 15920
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7852 14482 7880 15098
rect 7944 14958 7972 15914
rect 7932 14952 7984 14958
rect 7932 14894 7984 14900
rect 7944 14618 7972 14894
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 7746 14376 7802 14385
rect 7746 14311 7802 14320
rect 7852 14074 7880 14418
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 8036 13530 8064 17462
rect 8220 17338 8248 17614
rect 8404 17338 8432 17682
rect 8588 17513 8616 19110
rect 8668 18964 8720 18970
rect 8668 18906 8720 18912
rect 8680 18426 8708 18906
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 8680 17678 8708 18362
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8574 17504 8630 17513
rect 8574 17439 8630 17448
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 8128 15638 8156 16526
rect 8220 15978 8248 17070
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8680 16046 8708 16730
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 8576 15904 8628 15910
rect 8576 15846 8628 15852
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8116 15632 8168 15638
rect 8168 15592 8248 15620
rect 8116 15574 8168 15580
rect 8116 15428 8168 15434
rect 8116 15370 8168 15376
rect 8128 14958 8156 15370
rect 8220 15162 8248 15592
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 8128 14618 8156 14894
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 8312 14550 8340 15642
rect 8588 15502 8616 15846
rect 8772 15706 8800 19314
rect 8956 19174 8984 19790
rect 9036 19712 9088 19718
rect 9036 19654 9088 19660
rect 9048 19378 9076 19654
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 8864 18222 8892 18770
rect 8852 18216 8904 18222
rect 8852 18158 8904 18164
rect 8864 17610 8892 18158
rect 8852 17604 8904 17610
rect 8852 17546 8904 17552
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8668 15564 8720 15570
rect 8668 15506 8720 15512
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8588 14550 8616 15302
rect 8300 14544 8352 14550
rect 8300 14486 8352 14492
rect 8576 14544 8628 14550
rect 8576 14486 8628 14492
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8220 13870 8248 14418
rect 8312 14226 8340 14486
rect 8312 14198 8432 14226
rect 8208 13864 8260 13870
rect 8206 13832 8208 13841
rect 8260 13832 8262 13841
rect 8206 13767 8262 13776
rect 8404 13530 8432 14198
rect 8680 13530 8708 15506
rect 8864 15366 8892 17546
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7852 12238 7880 12582
rect 8404 12442 8432 13466
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8588 12442 8616 13262
rect 8680 12986 8708 13466
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7852 11898 7880 12174
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 7852 11393 7880 11834
rect 8956 11762 8984 19110
rect 9048 18222 9076 19110
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 9048 17814 9076 18158
rect 9036 17808 9088 17814
rect 9036 17750 9088 17756
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 9048 15978 9076 16390
rect 9036 15972 9088 15978
rect 9036 15914 9088 15920
rect 9048 15570 9076 15914
rect 9036 15564 9088 15570
rect 9036 15506 9088 15512
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 7838 11384 7894 11393
rect 7838 11319 7894 11328
rect 5998 11112 6054 11121
rect 5080 11076 5132 11082
rect 5998 11047 6054 11056
rect 5080 11018 5132 11024
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 6182 10024 6238 10033
rect 6182 9959 6184 9968
rect 6236 9959 6238 9968
rect 6184 9930 6236 9936
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 4066 8256 4122 8265
rect 4066 8191 4122 8200
rect 4080 7449 4108 8191
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 4066 7440 4122 7449
rect 4066 7375 4122 7384
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 3974 5128 4030 5137
rect 3974 5063 4030 5072
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8220 4185 8248 4218
rect 8206 4176 8262 4185
rect 8206 4111 8262 4120
rect 9140 3641 9168 20198
rect 9220 19916 9272 19922
rect 9220 19858 9272 19864
rect 9232 19689 9260 19858
rect 9324 19718 9352 21830
rect 9416 21146 9444 21927
rect 9404 21140 9456 21146
rect 9404 21082 9456 21088
rect 9508 21078 9536 24278
rect 9586 24239 9642 24248
rect 9692 23866 9720 24346
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 9680 23316 9732 23322
rect 9680 23258 9732 23264
rect 9588 23180 9640 23186
rect 9588 23122 9640 23128
rect 9600 22098 9628 23122
rect 9692 22234 9720 23258
rect 9784 22817 9812 27520
rect 10336 26081 10364 27520
rect 10322 26072 10378 26081
rect 10322 26007 10378 26016
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10324 25356 10376 25362
rect 10324 25298 10376 25304
rect 10336 24954 10364 25298
rect 10324 24948 10376 24954
rect 10324 24890 10376 24896
rect 9864 24676 9916 24682
rect 9864 24618 9916 24624
rect 9770 22808 9826 22817
rect 9770 22743 9826 22752
rect 9680 22228 9732 22234
rect 9680 22170 9732 22176
rect 9588 22092 9640 22098
rect 9588 22034 9640 22040
rect 9692 21690 9720 22170
rect 9876 22137 9904 24618
rect 9956 24608 10008 24614
rect 9956 24550 10008 24556
rect 9968 24138 9996 24550
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10782 24440 10838 24449
rect 10782 24375 10838 24384
rect 10048 24336 10100 24342
rect 10048 24278 10100 24284
rect 9956 24132 10008 24138
rect 9956 24074 10008 24080
rect 9968 22982 9996 24074
rect 10060 23866 10088 24278
rect 10140 24268 10192 24274
rect 10140 24210 10192 24216
rect 10048 23860 10100 23866
rect 10048 23802 10100 23808
rect 10152 23322 10180 24210
rect 10692 24200 10744 24206
rect 10796 24177 10824 24375
rect 10888 24274 10916 27520
rect 11440 24834 11468 27520
rect 11612 25152 11664 25158
rect 11612 25094 11664 25100
rect 11624 24954 11652 25094
rect 11612 24948 11664 24954
rect 11612 24890 11664 24896
rect 11992 24834 12020 27520
rect 12072 25356 12124 25362
rect 12072 25298 12124 25304
rect 11072 24806 11468 24834
rect 11532 24806 12020 24834
rect 10968 24608 11020 24614
rect 10966 24576 10968 24585
rect 11020 24576 11022 24585
rect 10966 24511 11022 24520
rect 10876 24268 10928 24274
rect 10876 24210 10928 24216
rect 10692 24142 10744 24148
rect 10782 24168 10838 24177
rect 10704 23526 10732 24142
rect 10782 24103 10838 24112
rect 10966 24032 11022 24041
rect 10966 23967 11022 23976
rect 10876 23792 10928 23798
rect 10876 23734 10928 23740
rect 10784 23656 10836 23662
rect 10784 23598 10836 23604
rect 10692 23520 10744 23526
rect 10692 23462 10744 23468
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10140 23316 10192 23322
rect 10140 23258 10192 23264
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 9956 22976 10008 22982
rect 9956 22918 10008 22924
rect 9968 22710 9996 22741
rect 9956 22704 10008 22710
rect 9954 22672 9956 22681
rect 10008 22672 10010 22681
rect 9954 22607 10010 22616
rect 9968 22438 9996 22607
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 9968 22273 9996 22374
rect 9954 22264 10010 22273
rect 9954 22199 10010 22208
rect 10152 22216 10180 23054
rect 10416 22976 10468 22982
rect 10416 22918 10468 22924
rect 10428 22506 10456 22918
rect 10416 22500 10468 22506
rect 10416 22442 10468 22448
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10152 22188 10272 22216
rect 9862 22128 9918 22137
rect 9862 22063 9918 22072
rect 9956 22092 10008 22098
rect 9956 22034 10008 22040
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9692 21185 9720 21626
rect 9678 21176 9734 21185
rect 9678 21111 9734 21120
rect 9496 21072 9548 21078
rect 9496 21014 9548 21020
rect 9968 21010 9996 22034
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 10060 21350 10088 21966
rect 10244 21418 10272 22188
rect 10704 21536 10732 23462
rect 10796 22982 10824 23598
rect 10784 22976 10836 22982
rect 10784 22918 10836 22924
rect 10796 21690 10824 22918
rect 10784 21684 10836 21690
rect 10784 21626 10836 21632
rect 10612 21508 10732 21536
rect 10232 21412 10284 21418
rect 10232 21354 10284 21360
rect 10048 21344 10100 21350
rect 10046 21312 10048 21321
rect 10612 21332 10640 21508
rect 10784 21412 10836 21418
rect 10784 21354 10836 21360
rect 10100 21312 10102 21321
rect 10612 21304 10732 21332
rect 10046 21247 10102 21256
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 9864 20936 9916 20942
rect 9864 20878 9916 20884
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9494 19816 9550 19825
rect 9416 19774 9494 19802
rect 9312 19712 9364 19718
rect 9218 19680 9274 19689
rect 9312 19654 9364 19660
rect 9218 19615 9274 19624
rect 9232 19446 9260 19615
rect 9220 19440 9272 19446
rect 9220 19382 9272 19388
rect 9324 18834 9352 19654
rect 9416 19514 9444 19774
rect 9494 19751 9550 19760
rect 9692 19514 9720 19858
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9496 19440 9548 19446
rect 9496 19382 9548 19388
rect 9404 18896 9456 18902
rect 9404 18838 9456 18844
rect 9312 18828 9364 18834
rect 9312 18770 9364 18776
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 9232 18154 9260 18702
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9220 18148 9272 18154
rect 9220 18090 9272 18096
rect 9232 17542 9260 18090
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 9232 17202 9260 17478
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9324 13705 9352 18566
rect 9416 18442 9444 18838
rect 9508 18630 9536 19382
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9600 18970 9628 19314
rect 9678 19136 9734 19145
rect 9678 19071 9734 19080
rect 9692 18970 9720 19071
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 9680 18964 9732 18970
rect 9680 18906 9732 18912
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 9494 18456 9550 18465
rect 9416 18414 9494 18442
rect 9494 18391 9550 18400
rect 9588 18420 9640 18426
rect 9680 18420 9732 18426
rect 9640 18380 9680 18408
rect 9588 18362 9640 18368
rect 9680 18362 9732 18368
rect 9402 18320 9458 18329
rect 9402 18255 9458 18264
rect 9416 16658 9444 18255
rect 9496 17740 9548 17746
rect 9496 17682 9548 17688
rect 9508 16726 9536 17682
rect 9588 17264 9640 17270
rect 9586 17232 9588 17241
rect 9640 17232 9642 17241
rect 9586 17167 9642 17176
rect 9600 16794 9628 17167
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 9678 16688 9734 16697
rect 9404 16652 9456 16658
rect 9678 16623 9680 16632
rect 9404 16594 9456 16600
rect 9732 16623 9734 16632
rect 9680 16594 9732 16600
rect 9692 16250 9720 16594
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 9416 14618 9444 15506
rect 9496 14884 9548 14890
rect 9496 14826 9548 14832
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9416 14414 9444 14554
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9416 13802 9444 14350
rect 9508 14074 9536 14826
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 9692 14074 9720 14486
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9404 13796 9456 13802
rect 9404 13738 9456 13744
rect 9310 13696 9366 13705
rect 9310 13631 9366 13640
rect 9416 13530 9444 13738
rect 9586 13696 9642 13705
rect 9586 13631 9642 13640
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9416 12986 9444 13466
rect 9600 13025 9628 13631
rect 9692 13326 9720 14010
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9586 13016 9642 13025
rect 9404 12980 9456 12986
rect 9586 12951 9642 12960
rect 9404 12922 9456 12928
rect 9416 12306 9444 12922
rect 9600 12782 9628 12951
rect 9784 12850 9812 20198
rect 9876 17882 9904 20878
rect 9968 20806 9996 20946
rect 10048 20936 10100 20942
rect 10048 20878 10100 20884
rect 9956 20800 10008 20806
rect 9956 20742 10008 20748
rect 9968 20534 9996 20742
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 10060 19854 10088 20878
rect 10704 20602 10732 21304
rect 10692 20596 10744 20602
rect 10692 20538 10744 20544
rect 10796 20482 10824 21354
rect 10888 20641 10916 23734
rect 10980 23633 11008 23967
rect 10966 23624 11022 23633
rect 10966 23559 11022 23568
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 10980 22778 11008 23462
rect 10968 22772 11020 22778
rect 10968 22714 11020 22720
rect 10968 21956 11020 21962
rect 10968 21898 11020 21904
rect 10980 21554 11008 21898
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 10874 20632 10930 20641
rect 10874 20567 10930 20576
rect 10966 20496 11022 20505
rect 10796 20454 10916 20482
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10048 19848 10100 19854
rect 10048 19790 10100 19796
rect 10140 19712 10192 19718
rect 10140 19654 10192 19660
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 9968 17921 9996 19314
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 10060 18057 10088 19110
rect 10152 18902 10180 19654
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10140 18896 10192 18902
rect 10140 18838 10192 18844
rect 10152 18426 10180 18838
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10690 18320 10746 18329
rect 10690 18255 10746 18264
rect 10704 18222 10732 18255
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10784 18080 10836 18086
rect 10046 18048 10102 18057
rect 10784 18022 10836 18028
rect 10046 17983 10102 17992
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 9954 17912 10010 17921
rect 9864 17876 9916 17882
rect 10289 17904 10585 17924
rect 10690 17912 10746 17921
rect 9954 17847 10010 17856
rect 10690 17847 10746 17856
rect 9864 17818 9916 17824
rect 10704 17746 10732 17847
rect 10692 17740 10744 17746
rect 10692 17682 10744 17688
rect 9956 17672 10008 17678
rect 9862 17640 9918 17649
rect 9956 17614 10008 17620
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 9862 17575 9918 17584
rect 9876 16794 9904 17575
rect 9968 17377 9996 17614
rect 9954 17368 10010 17377
rect 9954 17303 10010 17312
rect 10612 16980 10640 17614
rect 10612 16952 10732 16980
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 10060 15706 10088 15982
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10704 15638 10732 16952
rect 10796 16794 10824 18022
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10796 16114 10824 16730
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10796 15745 10824 15846
rect 10782 15736 10838 15745
rect 10782 15671 10838 15680
rect 10692 15632 10744 15638
rect 10744 15592 10824 15620
rect 10692 15574 10744 15580
rect 10048 15088 10100 15094
rect 10046 15056 10048 15065
rect 10100 15056 10102 15065
rect 10046 14991 10102 15000
rect 10508 14952 10560 14958
rect 10506 14920 10508 14929
rect 10560 14920 10562 14929
rect 10506 14855 10562 14864
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 10060 12986 10088 13738
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10336 12918 10364 13330
rect 10324 12912 10376 12918
rect 10324 12854 10376 12860
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10704 12374 10732 14758
rect 10796 14618 10824 15592
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10796 14074 10824 14554
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10888 13977 10916 20454
rect 10966 20431 10968 20440
rect 11020 20431 11022 20440
rect 10968 20402 11020 20408
rect 10980 20058 11008 20402
rect 10968 20052 11020 20058
rect 10968 19994 11020 20000
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 10980 18630 11008 19110
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 10980 17649 11008 18566
rect 11072 18465 11100 24806
rect 11428 24268 11480 24274
rect 11428 24210 11480 24216
rect 11150 24168 11206 24177
rect 11150 24103 11206 24112
rect 11058 18456 11114 18465
rect 11058 18391 11114 18400
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 11072 17746 11100 18226
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 10966 17640 11022 17649
rect 10966 17575 11022 17584
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10980 16658 11008 17478
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 11072 16726 11100 16934
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10966 16280 11022 16289
rect 10966 16215 11022 16224
rect 10980 15706 11008 16215
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 10874 13968 10930 13977
rect 10874 13903 10930 13912
rect 11164 13818 11192 24103
rect 11336 24064 11388 24070
rect 11336 24006 11388 24012
rect 11348 23730 11376 24006
rect 11336 23724 11388 23730
rect 11336 23666 11388 23672
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 11256 22001 11284 22034
rect 11242 21992 11298 22001
rect 11242 21927 11298 21936
rect 11244 21888 11296 21894
rect 11244 21830 11296 21836
rect 11256 21554 11284 21830
rect 11244 21548 11296 21554
rect 11244 21490 11296 21496
rect 11256 20466 11284 21490
rect 11244 20460 11296 20466
rect 11244 20402 11296 20408
rect 11256 19922 11284 20402
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11348 19718 11376 23666
rect 11440 23526 11468 24210
rect 11428 23520 11480 23526
rect 11428 23462 11480 23468
rect 11428 22704 11480 22710
rect 11426 22672 11428 22681
rect 11480 22672 11482 22681
rect 11426 22607 11482 22616
rect 11426 21992 11482 22001
rect 11426 21927 11428 21936
rect 11480 21927 11482 21936
rect 11428 21898 11480 21904
rect 11336 19712 11388 19718
rect 11336 19654 11388 19660
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11256 18329 11284 18906
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11242 18320 11298 18329
rect 11242 18255 11298 18264
rect 11242 18184 11298 18193
rect 11242 18119 11244 18128
rect 11296 18119 11298 18128
rect 11244 18090 11296 18096
rect 11348 17202 11376 18566
rect 11426 18456 11482 18465
rect 11426 18391 11482 18400
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11440 16833 11468 18391
rect 11426 16824 11482 16833
rect 11426 16759 11482 16768
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11440 16114 11468 16594
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 11336 15020 11388 15026
rect 11336 14962 11388 14968
rect 11348 14822 11376 14962
rect 11532 14958 11560 24806
rect 11980 24608 12032 24614
rect 12084 24596 12112 25298
rect 12256 25220 12308 25226
rect 12256 25162 12308 25168
rect 12268 24818 12296 25162
rect 12256 24812 12308 24818
rect 12256 24754 12308 24760
rect 12032 24568 12112 24596
rect 11980 24550 12032 24556
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11808 23361 11836 24006
rect 11794 23352 11850 23361
rect 11794 23287 11850 23296
rect 11612 23180 11664 23186
rect 11612 23122 11664 23128
rect 11624 22438 11652 23122
rect 11612 22432 11664 22438
rect 11612 22374 11664 22380
rect 11888 22432 11940 22438
rect 11888 22374 11940 22380
rect 11624 21690 11652 22374
rect 11612 21684 11664 21690
rect 11612 21626 11664 21632
rect 11702 21584 11758 21593
rect 11702 21519 11758 21528
rect 11612 20800 11664 20806
rect 11612 20742 11664 20748
rect 11624 20466 11652 20742
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 11716 16017 11744 21519
rect 11900 21049 11928 22374
rect 11992 21321 12020 24550
rect 12176 24410 12480 24426
rect 12176 24404 12492 24410
rect 12176 24398 12440 24404
rect 12072 24336 12124 24342
rect 12072 24278 12124 24284
rect 12084 21690 12112 24278
rect 12072 21684 12124 21690
rect 12072 21626 12124 21632
rect 11978 21312 12034 21321
rect 11978 21247 12034 21256
rect 11886 21040 11942 21049
rect 11886 20975 11942 20984
rect 11980 20868 12032 20874
rect 11980 20810 12032 20816
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 11808 18970 11836 19450
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 11992 18222 12020 20810
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 12084 19514 12112 19790
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 12070 19408 12126 19417
rect 12070 19343 12126 19352
rect 12084 19310 12112 19343
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 12072 18964 12124 18970
rect 12072 18906 12124 18912
rect 11980 18216 12032 18222
rect 11980 18158 12032 18164
rect 12084 17134 12112 18906
rect 12176 17218 12204 24398
rect 12440 24346 12492 24352
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12360 23866 12388 24142
rect 12348 23860 12400 23866
rect 12348 23802 12400 23808
rect 12360 23526 12388 23802
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 12348 23520 12400 23526
rect 12348 23462 12400 23468
rect 12360 23322 12388 23462
rect 12348 23316 12400 23322
rect 12348 23258 12400 23264
rect 12452 22982 12480 23598
rect 12440 22976 12492 22982
rect 12440 22918 12492 22924
rect 12452 22574 12480 22918
rect 12440 22568 12492 22574
rect 12440 22510 12492 22516
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 12268 21350 12296 21830
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12268 20058 12296 21286
rect 12452 20942 12480 21286
rect 12440 20936 12492 20942
rect 12440 20878 12492 20884
rect 12452 20754 12480 20878
rect 12544 20874 12572 27520
rect 12992 25356 13044 25362
rect 12992 25298 13044 25304
rect 12714 24712 12770 24721
rect 12624 24676 12676 24682
rect 12714 24647 12770 24656
rect 12624 24618 12676 24624
rect 12532 20868 12584 20874
rect 12532 20810 12584 20816
rect 12452 20726 12572 20754
rect 12438 20632 12494 20641
rect 12438 20567 12494 20576
rect 12348 20528 12400 20534
rect 12348 20470 12400 20476
rect 12256 20052 12308 20058
rect 12256 19994 12308 20000
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 12268 19446 12296 19858
rect 12360 19825 12388 20470
rect 12452 20398 12480 20567
rect 12440 20392 12492 20398
rect 12440 20334 12492 20340
rect 12452 19990 12480 20334
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 12346 19816 12402 19825
rect 12346 19751 12402 19760
rect 12256 19440 12308 19446
rect 12256 19382 12308 19388
rect 12440 19236 12492 19242
rect 12440 19178 12492 19184
rect 12256 18896 12308 18902
rect 12256 18838 12308 18844
rect 12268 18426 12296 18838
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12268 17542 12296 18158
rect 12348 17808 12400 17814
rect 12348 17750 12400 17756
rect 12256 17536 12308 17542
rect 12360 17524 12388 17750
rect 12452 17678 12480 19178
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12440 17536 12492 17542
rect 12360 17496 12440 17524
rect 12256 17478 12308 17484
rect 12440 17478 12492 17484
rect 12176 17190 12296 17218
rect 12544 17202 12572 20726
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11702 16008 11758 16017
rect 11702 15943 11758 15952
rect 11900 15910 11928 16050
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11900 15366 11928 15846
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11520 14952 11572 14958
rect 11520 14894 11572 14900
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11164 13802 11284 13818
rect 11164 13796 11296 13802
rect 11164 13790 11244 13796
rect 11244 13738 11296 13744
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 11072 12850 11100 13670
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 10782 12744 10838 12753
rect 10782 12679 10838 12688
rect 10796 12646 10824 12679
rect 10784 12640 10836 12646
rect 11060 12640 11112 12646
rect 10784 12582 10836 12588
rect 10888 12588 11060 12594
rect 10888 12582 11112 12588
rect 10888 12566 11100 12582
rect 10888 12442 10916 12566
rect 10876 12436 10928 12442
rect 11256 12424 11284 12786
rect 10876 12378 10928 12384
rect 11072 12396 11284 12424
rect 10692 12368 10744 12374
rect 10692 12310 10744 12316
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 10704 11762 10732 12310
rect 11072 12288 11100 12396
rect 11348 12306 11376 14758
rect 11900 14346 11928 15302
rect 11888 14340 11940 14346
rect 11888 14282 11940 14288
rect 12084 14260 12112 17070
rect 12164 16720 12216 16726
rect 12164 16662 12216 16668
rect 12176 15366 12204 16662
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 12164 14272 12216 14278
rect 12084 14232 12164 14260
rect 12164 14214 12216 14220
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11624 12918 11652 13126
rect 11612 12912 11664 12918
rect 11612 12854 11664 12860
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 10980 12260 11100 12288
rect 11152 12300 11204 12306
rect 10980 11898 11008 12260
rect 11152 12242 11204 12248
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 11072 11898 11100 12106
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 11072 11257 11100 11494
rect 11058 11248 11114 11257
rect 11058 11183 11114 11192
rect 11164 11082 11192 12242
rect 11348 11694 11376 12242
rect 11716 11762 11744 12718
rect 12084 12209 12112 13806
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12176 12646 12204 13330
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12070 12200 12126 12209
rect 12070 12135 12126 12144
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11716 11354 11744 11698
rect 12072 11620 12124 11626
rect 12072 11562 12124 11568
rect 12084 11354 12112 11562
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 12176 11234 12204 12582
rect 12084 11206 12204 11234
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 9678 9752 9734 9761
rect 9678 9687 9734 9696
rect 9692 4049 9720 9687
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 9678 4040 9734 4049
rect 9678 3975 9734 3984
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 9126 3632 9182 3641
rect 9126 3567 9182 3576
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 8298 2952 8354 2961
rect 8298 2887 8354 2896
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 3698 1456 3754 1465
rect 3698 1391 3754 1400
rect 8312 480 8340 2887
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 11992 2650 12020 11018
rect 12084 9761 12112 11206
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12176 10198 12204 11086
rect 12268 10266 12296 17190
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12636 17082 12664 24618
rect 12728 24614 12756 24647
rect 12716 24608 12768 24614
rect 12716 24550 12768 24556
rect 13004 24410 13032 25298
rect 13096 24857 13124 27520
rect 13452 25764 13504 25770
rect 13452 25706 13504 25712
rect 13268 25288 13320 25294
rect 13268 25230 13320 25236
rect 13176 24880 13228 24886
rect 13082 24848 13138 24857
rect 13176 24822 13228 24828
rect 13082 24783 13138 24792
rect 12992 24404 13044 24410
rect 12992 24346 13044 24352
rect 13096 24290 13124 24783
rect 12912 24262 13124 24290
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 12820 21622 12848 21966
rect 12808 21616 12860 21622
rect 12808 21558 12860 21564
rect 12716 20800 12768 20806
rect 12716 20742 12768 20748
rect 12728 20505 12756 20742
rect 12714 20496 12770 20505
rect 12714 20431 12770 20440
rect 12820 19174 12848 21558
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12912 18970 12940 24262
rect 13188 23905 13216 24822
rect 13280 24750 13308 25230
rect 13464 24818 13492 25706
rect 13648 24886 13676 27520
rect 14004 25424 14056 25430
rect 14004 25366 14056 25372
rect 13820 25152 13872 25158
rect 13820 25094 13872 25100
rect 13636 24880 13688 24886
rect 13636 24822 13688 24828
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13268 24744 13320 24750
rect 13268 24686 13320 24692
rect 13464 24410 13492 24754
rect 13636 24744 13688 24750
rect 13636 24686 13688 24692
rect 13452 24404 13504 24410
rect 13452 24346 13504 24352
rect 13544 24268 13596 24274
rect 13544 24210 13596 24216
rect 13556 24177 13584 24210
rect 13542 24168 13598 24177
rect 13542 24103 13598 24112
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 13174 23896 13230 23905
rect 13174 23831 13230 23840
rect 12992 23520 13044 23526
rect 12992 23462 13044 23468
rect 13082 23488 13138 23497
rect 13004 22030 13032 23462
rect 13082 23423 13138 23432
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 13004 21690 13032 21966
rect 12992 21684 13044 21690
rect 12992 21626 13044 21632
rect 13096 21486 13124 23423
rect 13188 21486 13216 23831
rect 13268 23180 13320 23186
rect 13268 23122 13320 23128
rect 13280 22982 13308 23122
rect 13268 22976 13320 22982
rect 13268 22918 13320 22924
rect 13280 22234 13308 22918
rect 13268 22228 13320 22234
rect 13268 22170 13320 22176
rect 13372 22166 13400 24006
rect 13556 23866 13584 24103
rect 13544 23860 13596 23866
rect 13544 23802 13596 23808
rect 13360 22160 13412 22166
rect 13360 22102 13412 22108
rect 13084 21480 13136 21486
rect 13084 21422 13136 21428
rect 13176 21480 13228 21486
rect 13176 21422 13228 21428
rect 13268 21072 13320 21078
rect 13268 21014 13320 21020
rect 13176 20936 13228 20942
rect 13176 20878 13228 20884
rect 12990 20496 13046 20505
rect 12990 20431 12992 20440
rect 13044 20431 13046 20440
rect 12992 20402 13044 20408
rect 13188 20262 13216 20878
rect 13280 20534 13308 21014
rect 13360 20936 13412 20942
rect 13360 20878 13412 20884
rect 13372 20602 13400 20878
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 13268 20528 13320 20534
rect 13268 20470 13320 20476
rect 13280 20398 13308 20470
rect 13268 20392 13320 20398
rect 13266 20360 13268 20369
rect 13320 20360 13322 20369
rect 13266 20295 13322 20304
rect 12992 20256 13044 20262
rect 12992 20198 13044 20204
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 12900 18964 12952 18970
rect 12900 18906 12952 18912
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12728 18154 12756 18566
rect 12716 18148 12768 18154
rect 12716 18090 12768 18096
rect 12728 17610 12756 18090
rect 12912 17882 12940 18906
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 12636 17054 12848 17082
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12530 16280 12586 16289
rect 12530 16215 12586 16224
rect 12544 16046 12572 16215
rect 12348 16040 12400 16046
rect 12532 16040 12584 16046
rect 12400 16000 12480 16028
rect 12348 15982 12400 15988
rect 12452 15162 12480 16000
rect 12532 15982 12584 15988
rect 12636 15978 12664 16390
rect 12624 15972 12676 15978
rect 12624 15914 12676 15920
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12438 15056 12494 15065
rect 12438 14991 12494 15000
rect 12452 14890 12480 14991
rect 12440 14884 12492 14890
rect 12440 14826 12492 14832
rect 12544 14618 12572 15506
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12636 14890 12664 15302
rect 12624 14884 12676 14890
rect 12624 14826 12676 14832
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12452 14074 12480 14418
rect 12636 14414 12664 14486
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12544 13954 12572 14214
rect 12452 13926 12572 13954
rect 12452 13274 12480 13926
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12544 13462 12572 13670
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12452 13246 12572 13274
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12452 11898 12480 12718
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12544 11354 12572 13246
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12438 10840 12494 10849
rect 12360 10810 12438 10826
rect 12348 10804 12438 10810
rect 12400 10798 12438 10804
rect 12438 10775 12494 10784
rect 12348 10746 12400 10752
rect 12544 10690 12572 11290
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12636 10849 12664 11154
rect 12622 10840 12678 10849
rect 12622 10775 12678 10784
rect 12360 10674 12572 10690
rect 12348 10668 12572 10674
rect 12400 10662 12572 10668
rect 12348 10610 12400 10616
rect 12452 10577 12480 10662
rect 12438 10568 12494 10577
rect 12438 10503 12494 10512
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12544 10266 12572 10406
rect 12728 10266 12756 16934
rect 12820 13870 12848 17054
rect 12912 16998 12940 17138
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12912 14822 12940 16934
rect 13004 15609 13032 20198
rect 13372 19854 13400 20538
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13372 19446 13400 19790
rect 13360 19440 13412 19446
rect 13360 19382 13412 19388
rect 13464 19378 13492 19994
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 13544 19236 13596 19242
rect 13544 19178 13596 19184
rect 13174 19136 13230 19145
rect 13174 19071 13230 19080
rect 13188 18766 13216 19071
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 13084 15632 13136 15638
rect 12990 15600 13046 15609
rect 13084 15574 13136 15580
rect 12990 15535 13046 15544
rect 13096 15026 13124 15574
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 12992 14884 13044 14890
rect 12992 14826 13044 14832
rect 12900 14816 12952 14822
rect 12900 14758 12952 14764
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12164 10192 12216 10198
rect 12164 10134 12216 10140
rect 12070 9752 12126 9761
rect 12070 9687 12126 9696
rect 12544 9586 12572 10202
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12636 9722 12664 9998
rect 12728 9722 12756 10202
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12820 9625 12848 13466
rect 12912 12850 12940 14214
rect 13004 13818 13032 14826
rect 13096 13938 13124 14962
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 13004 13790 13124 13818
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 12912 12170 12940 12786
rect 13004 12442 13032 12786
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 13096 12306 13124 13790
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 12900 12164 12952 12170
rect 12900 12106 12952 12112
rect 13004 12102 13032 12242
rect 13082 12200 13138 12209
rect 13082 12135 13138 12144
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12912 11354 12940 11834
rect 13004 11762 13032 12038
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12912 10606 12940 11290
rect 13004 11150 13032 11698
rect 13096 11694 13124 12135
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 13188 10849 13216 18702
rect 13280 17542 13308 18702
rect 13360 17604 13412 17610
rect 13360 17546 13412 17552
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13280 17202 13308 17478
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 13280 16454 13308 17138
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 13280 15910 13308 16390
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 13174 10840 13230 10849
rect 13174 10775 13230 10784
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12806 9616 12862 9625
rect 12532 9580 12584 9586
rect 12806 9551 12862 9560
rect 12532 9522 12584 9528
rect 12438 2952 12494 2961
rect 12438 2887 12494 2896
rect 12452 2650 12480 2887
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 1306 368 1362 377
rect 1306 303 1362 312
rect 2778 0 2834 480
rect 8298 0 8354 480
rect 13188 241 13216 10775
rect 13280 10674 13308 15846
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13280 10266 13308 10610
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13372 10062 13400 17546
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13464 16153 13492 16390
rect 13450 16144 13506 16153
rect 13556 16130 13584 19178
rect 13648 18408 13676 24686
rect 13728 24132 13780 24138
rect 13728 24074 13780 24080
rect 13740 21593 13768 24074
rect 13726 21584 13782 21593
rect 13726 21519 13728 21528
rect 13780 21519 13782 21528
rect 13728 21490 13780 21496
rect 13740 20058 13768 21490
rect 13832 20058 13860 25094
rect 14016 24750 14044 25366
rect 14004 24744 14056 24750
rect 14004 24686 14056 24692
rect 14096 24676 14148 24682
rect 14096 24618 14148 24624
rect 14004 24608 14056 24614
rect 14004 24550 14056 24556
rect 14016 24410 14044 24550
rect 14004 24404 14056 24410
rect 14004 24346 14056 24352
rect 14108 24177 14136 24618
rect 14094 24168 14150 24177
rect 14094 24103 14150 24112
rect 14004 23520 14056 23526
rect 14292 23497 14320 27520
rect 14372 25968 14424 25974
rect 14372 25910 14424 25916
rect 14384 25498 14412 25910
rect 14556 25900 14608 25906
rect 14556 25842 14608 25848
rect 14372 25492 14424 25498
rect 14372 25434 14424 25440
rect 14372 25220 14424 25226
rect 14372 25162 14424 25168
rect 14384 24857 14412 25162
rect 14370 24848 14426 24857
rect 14370 24783 14372 24792
rect 14424 24783 14426 24792
rect 14372 24754 14424 24760
rect 14568 24274 14596 25842
rect 14844 24834 14872 27520
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14660 24806 14872 24834
rect 15396 24834 15424 27520
rect 15844 25288 15896 25294
rect 15844 25230 15896 25236
rect 15476 25152 15528 25158
rect 15528 25100 15792 25106
rect 15476 25094 15792 25100
rect 15488 25078 15792 25094
rect 15396 24806 15700 24834
rect 14556 24268 14608 24274
rect 14556 24210 14608 24216
rect 14568 23798 14596 24210
rect 14372 23792 14424 23798
rect 14372 23734 14424 23740
rect 14556 23792 14608 23798
rect 14556 23734 14608 23740
rect 14004 23462 14056 23468
rect 14278 23488 14334 23497
rect 13910 23352 13966 23361
rect 13910 23287 13912 23296
rect 13964 23287 13966 23296
rect 13912 23258 13964 23264
rect 13924 22778 13952 23258
rect 14016 23118 14044 23462
rect 14278 23423 14334 23432
rect 14004 23112 14056 23118
rect 14004 23054 14056 23060
rect 13912 22772 13964 22778
rect 13912 22714 13964 22720
rect 14016 22574 14044 23054
rect 14278 22808 14334 22817
rect 14278 22743 14334 22752
rect 14004 22568 14056 22574
rect 14004 22510 14056 22516
rect 14096 22568 14148 22574
rect 14096 22510 14148 22516
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 13924 20942 13952 22374
rect 14016 22234 14044 22510
rect 14004 22228 14056 22234
rect 14004 22170 14056 22176
rect 14004 22092 14056 22098
rect 14004 22034 14056 22040
rect 13912 20936 13964 20942
rect 13912 20878 13964 20884
rect 14016 20806 14044 22034
rect 14108 20874 14136 22510
rect 14292 22030 14320 22743
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 14280 21548 14332 21554
rect 14280 21490 14332 21496
rect 14292 20942 14320 21490
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14096 20868 14148 20874
rect 14096 20810 14148 20816
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 14004 20800 14056 20806
rect 14004 20742 14056 20748
rect 13924 20312 13952 20742
rect 14292 20398 14320 20878
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 14004 20324 14056 20330
rect 13924 20284 14004 20312
rect 14004 20266 14056 20272
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 14016 19854 14044 20266
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 14108 19718 14136 19858
rect 14292 19718 14320 20334
rect 14096 19712 14148 19718
rect 14094 19680 14096 19689
rect 14280 19712 14332 19718
rect 14148 19680 14150 19689
rect 14280 19654 14332 19660
rect 14094 19615 14150 19624
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 13820 18420 13872 18426
rect 13648 18380 13820 18408
rect 13820 18362 13872 18368
rect 13832 17882 13860 18362
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13634 17640 13690 17649
rect 13634 17575 13690 17584
rect 13648 16794 13676 17575
rect 13740 16998 13768 17682
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 13740 16561 13768 16934
rect 13726 16552 13782 16561
rect 13726 16487 13782 16496
rect 13634 16144 13690 16153
rect 13556 16102 13634 16130
rect 13450 16079 13506 16088
rect 13634 16079 13690 16088
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13450 15736 13506 15745
rect 13450 15671 13452 15680
rect 13504 15671 13506 15680
rect 13452 15642 13504 15648
rect 13450 15600 13506 15609
rect 13450 15535 13506 15544
rect 13464 15042 13492 15535
rect 13556 15502 13584 15982
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 13556 15162 13584 15438
rect 13544 15156 13596 15162
rect 13544 15098 13596 15104
rect 13464 15014 13584 15042
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 13174 232 13230 241
rect 13174 167 13230 176
rect 13464 105 13492 14758
rect 13556 13530 13584 15014
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13544 12300 13596 12306
rect 13544 12242 13596 12248
rect 13556 10470 13584 12242
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13556 5137 13584 10406
rect 13648 8945 13676 16079
rect 13740 15881 13768 16487
rect 13726 15872 13782 15881
rect 13924 15858 13952 19110
rect 14094 18864 14150 18873
rect 14094 18799 14150 18808
rect 14004 17808 14056 17814
rect 14004 17750 14056 17756
rect 14016 17338 14044 17750
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 14002 16824 14058 16833
rect 14108 16794 14136 18799
rect 14292 18222 14320 19654
rect 14280 18216 14332 18222
rect 14280 18158 14332 18164
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14002 16759 14004 16768
rect 14056 16759 14058 16768
rect 14096 16788 14148 16794
rect 14004 16730 14056 16736
rect 14096 16730 14148 16736
rect 14016 16250 14044 16730
rect 14004 16244 14056 16250
rect 14004 16186 14056 16192
rect 13924 15830 14044 15858
rect 13726 15807 13782 15816
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13740 15094 13768 15506
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 13832 14482 13860 15302
rect 13924 15162 13952 15642
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 14016 14634 14044 15830
rect 14108 15706 14136 16730
rect 14200 16454 14228 17614
rect 14292 17134 14320 17818
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 14188 16448 14240 16454
rect 14188 16390 14240 16396
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14384 15586 14412 23734
rect 14556 23044 14608 23050
rect 14556 22986 14608 22992
rect 14568 21146 14596 22986
rect 14556 21140 14608 21146
rect 14556 21082 14608 21088
rect 14660 20992 14688 24806
rect 14740 24744 14792 24750
rect 14740 24686 14792 24692
rect 14752 24614 14780 24686
rect 14740 24608 14792 24614
rect 14740 24550 14792 24556
rect 15108 24608 15160 24614
rect 15476 24608 15528 24614
rect 15108 24550 15160 24556
rect 15382 24576 15438 24585
rect 14752 23050 14780 24550
rect 15120 24206 15148 24550
rect 15476 24550 15528 24556
rect 15382 24511 15438 24520
rect 15292 24404 15344 24410
rect 15292 24346 15344 24352
rect 15108 24200 15160 24206
rect 15108 24142 15160 24148
rect 14832 24064 14884 24070
rect 14832 24006 14884 24012
rect 14740 23044 14792 23050
rect 14740 22986 14792 22992
rect 14738 22944 14794 22953
rect 14738 22879 14794 22888
rect 14752 22778 14780 22879
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 14844 22098 14872 24006
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15304 23594 15332 24346
rect 15396 23866 15424 24511
rect 15384 23860 15436 23866
rect 15384 23802 15436 23808
rect 15292 23588 15344 23594
rect 15292 23530 15344 23536
rect 15384 23520 15436 23526
rect 15384 23462 15436 23468
rect 15292 22976 15344 22982
rect 15292 22918 15344 22924
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15304 22574 15332 22918
rect 15292 22568 15344 22574
rect 15292 22510 15344 22516
rect 14924 22432 14976 22438
rect 14924 22374 14976 22380
rect 15108 22432 15160 22438
rect 15108 22374 15160 22380
rect 14936 22273 14964 22374
rect 14922 22264 14978 22273
rect 14922 22199 14978 22208
rect 15120 22098 15148 22374
rect 14832 22092 14884 22098
rect 14832 22034 14884 22040
rect 15108 22092 15160 22098
rect 15108 22034 15160 22040
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14740 21412 14792 21418
rect 14740 21354 14792 21360
rect 14568 20964 14688 20992
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 14476 19310 14504 19994
rect 14568 19990 14596 20964
rect 14752 20913 14780 21354
rect 15304 20942 15332 21830
rect 15396 21593 15424 23462
rect 15382 21584 15438 21593
rect 15382 21519 15438 21528
rect 15292 20936 15344 20942
rect 14738 20904 14794 20913
rect 15292 20878 15344 20884
rect 14738 20839 14794 20848
rect 14648 20800 14700 20806
rect 14648 20742 14700 20748
rect 14556 19984 14608 19990
rect 14556 19926 14608 19932
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14476 17649 14504 19110
rect 14568 18630 14596 19314
rect 14556 18624 14608 18630
rect 14556 18566 14608 18572
rect 14568 18154 14596 18566
rect 14556 18148 14608 18154
rect 14556 18090 14608 18096
rect 14556 17740 14608 17746
rect 14556 17682 14608 17688
rect 14462 17640 14518 17649
rect 14462 17575 14518 17584
rect 14568 17513 14596 17682
rect 14554 17504 14610 17513
rect 14554 17439 14610 17448
rect 14568 16726 14596 17439
rect 14556 16720 14608 16726
rect 14556 16662 14608 16668
rect 14660 16250 14688 20742
rect 14752 20602 14780 20839
rect 15382 20768 15438 20777
rect 14956 20700 15252 20720
rect 15382 20703 15438 20712
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 15396 20058 15424 20703
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15488 19990 15516 24550
rect 15566 24440 15622 24449
rect 15566 24375 15622 24384
rect 15580 24342 15608 24375
rect 15568 24336 15620 24342
rect 15568 24278 15620 24284
rect 15568 22500 15620 22506
rect 15568 22442 15620 22448
rect 15476 19984 15528 19990
rect 15476 19926 15528 19932
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14740 18896 14792 18902
rect 14740 18838 14792 18844
rect 14752 18290 14780 18838
rect 14844 18766 14872 19110
rect 15580 18970 15608 22442
rect 15568 18964 15620 18970
rect 15568 18906 15620 18912
rect 14832 18760 14884 18766
rect 14832 18702 14884 18708
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14752 17882 14780 18226
rect 14740 17876 14792 17882
rect 14740 17818 14792 17824
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14752 17066 14780 17614
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 14844 16794 14872 18702
rect 15566 18592 15622 18601
rect 14956 18524 15252 18544
rect 15566 18527 15622 18536
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15580 18426 15608 18527
rect 15568 18420 15620 18426
rect 15568 18362 15620 18368
rect 14924 18216 14976 18222
rect 14924 18158 14976 18164
rect 14936 17678 14964 18158
rect 15384 18148 15436 18154
rect 15384 18090 15436 18096
rect 15290 17912 15346 17921
rect 15290 17847 15292 17856
rect 15344 17847 15346 17856
rect 15292 17818 15344 17824
rect 14924 17672 14976 17678
rect 14924 17614 14976 17620
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15396 17338 15424 18090
rect 15672 17882 15700 24806
rect 15764 22506 15792 25078
rect 15856 24614 15884 25230
rect 15844 24608 15896 24614
rect 15844 24550 15896 24556
rect 15752 22500 15804 22506
rect 15752 22442 15804 22448
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 15764 21078 15792 21286
rect 15752 21072 15804 21078
rect 15752 21014 15804 21020
rect 15764 20602 15792 21014
rect 15752 20596 15804 20602
rect 15752 20538 15804 20544
rect 15752 19916 15804 19922
rect 15752 19858 15804 19864
rect 15764 19174 15792 19858
rect 15752 19168 15804 19174
rect 15750 19136 15752 19145
rect 15804 19136 15806 19145
rect 15750 19071 15806 19080
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 15750 17776 15806 17785
rect 15750 17711 15752 17720
rect 15804 17711 15806 17720
rect 15752 17682 15804 17688
rect 15764 17338 15792 17682
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15752 17332 15804 17338
rect 15752 17274 15804 17280
rect 15856 17218 15884 24550
rect 15948 24410 15976 27520
rect 16500 25498 16528 27520
rect 16856 25832 16908 25838
rect 16856 25774 16908 25780
rect 16120 25492 16172 25498
rect 16120 25434 16172 25440
rect 16488 25492 16540 25498
rect 16488 25434 16540 25440
rect 16028 25288 16080 25294
rect 16028 25230 16080 25236
rect 15936 24404 15988 24410
rect 15936 24346 15988 24352
rect 16040 24342 16068 25230
rect 16132 24614 16160 25434
rect 16396 25288 16448 25294
rect 16396 25230 16448 25236
rect 16212 25152 16264 25158
rect 16212 25094 16264 25100
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 16028 24336 16080 24342
rect 16028 24278 16080 24284
rect 15936 24200 15988 24206
rect 15936 24142 15988 24148
rect 15948 22114 15976 24142
rect 16132 23633 16160 24550
rect 16224 24410 16252 25094
rect 16408 24857 16436 25230
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 16394 24848 16450 24857
rect 16394 24783 16450 24792
rect 16408 24614 16436 24783
rect 16396 24608 16448 24614
rect 16396 24550 16448 24556
rect 16212 24404 16264 24410
rect 16212 24346 16264 24352
rect 16224 23662 16252 24346
rect 16304 24336 16356 24342
rect 16304 24278 16356 24284
rect 16212 23656 16264 23662
rect 16118 23624 16174 23633
rect 16212 23598 16264 23604
rect 16118 23559 16174 23568
rect 16028 23180 16080 23186
rect 16028 23122 16080 23128
rect 16040 22438 16068 23122
rect 16028 22432 16080 22438
rect 16028 22374 16080 22380
rect 16040 22234 16068 22374
rect 16028 22228 16080 22234
rect 16028 22170 16080 22176
rect 15948 22086 16068 22114
rect 15936 21480 15988 21486
rect 15936 21422 15988 21428
rect 15948 20058 15976 21422
rect 15936 20052 15988 20058
rect 15936 19994 15988 20000
rect 15948 19514 15976 19994
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 16040 18850 16068 22086
rect 16118 20904 16174 20913
rect 16118 20839 16174 20848
rect 16132 19446 16160 20839
rect 16212 20256 16264 20262
rect 16212 20198 16264 20204
rect 16224 19922 16252 20198
rect 16212 19916 16264 19922
rect 16212 19858 16264 19864
rect 16316 19666 16344 24278
rect 16408 23186 16436 24550
rect 16592 24274 16620 25094
rect 16580 24268 16632 24274
rect 16580 24210 16632 24216
rect 16764 24268 16816 24274
rect 16764 24210 16816 24216
rect 16592 23798 16620 24210
rect 16776 23866 16804 24210
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 16580 23792 16632 23798
rect 16580 23734 16632 23740
rect 16486 23624 16542 23633
rect 16486 23559 16542 23568
rect 16396 23180 16448 23186
rect 16396 23122 16448 23128
rect 16396 22092 16448 22098
rect 16396 22034 16448 22040
rect 16408 21350 16436 22034
rect 16396 21344 16448 21350
rect 16396 21286 16448 21292
rect 16408 21185 16436 21286
rect 16394 21176 16450 21185
rect 16394 21111 16450 21120
rect 16396 20324 16448 20330
rect 16396 20266 16448 20272
rect 16224 19638 16344 19666
rect 16120 19440 16172 19446
rect 16120 19382 16172 19388
rect 16132 18970 16160 19382
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 16040 18822 16160 18850
rect 16028 18760 16080 18766
rect 16028 18702 16080 18708
rect 16040 18086 16068 18702
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 15948 17270 15976 17614
rect 16132 17542 16160 18822
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 15936 17264 15988 17270
rect 15764 17190 15884 17218
rect 15934 17232 15936 17241
rect 15988 17232 15990 17241
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 15212 16522 15240 17070
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15200 16516 15252 16522
rect 15200 16458 15252 16464
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 14752 16182 14780 16390
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14740 16176 14792 16182
rect 14740 16118 14792 16124
rect 14648 15972 14700 15978
rect 14648 15914 14700 15920
rect 14292 15558 14412 15586
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 13924 14606 14044 14634
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13924 14006 13952 14606
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 14016 14074 14044 14486
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 13924 13870 13952 13942
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 14002 13696 14058 13705
rect 13740 10169 13768 13670
rect 14002 13631 14058 13640
rect 14016 13190 14044 13631
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 14016 13025 14044 13126
rect 14002 13016 14058 13025
rect 14108 12986 14136 15302
rect 14292 15201 14320 15558
rect 14660 15366 14688 15914
rect 15396 15910 15424 16526
rect 15488 15978 15516 16594
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15476 15972 15528 15978
rect 15476 15914 15528 15920
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14278 15192 14334 15201
rect 14278 15127 14334 15136
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 14200 13297 14228 14350
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14372 13320 14424 13326
rect 14186 13288 14242 13297
rect 14372 13262 14424 13268
rect 14186 13223 14242 13232
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14002 12951 14058 12960
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14002 12880 14058 12889
rect 14002 12815 14058 12824
rect 14096 12844 14148 12850
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13832 11694 13860 12242
rect 13820 11688 13872 11694
rect 13818 11656 13820 11665
rect 13872 11656 13874 11665
rect 13818 11591 13874 11600
rect 13924 11286 13952 12582
rect 14016 11354 14044 12815
rect 14096 12786 14148 12792
rect 14108 12442 14136 12786
rect 14292 12782 14320 13126
rect 14384 12850 14412 13262
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 14094 12336 14150 12345
rect 14094 12271 14150 12280
rect 14108 12238 14136 12271
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 14108 11898 14136 12174
rect 14200 12102 14228 12650
rect 14384 12481 14412 12786
rect 14370 12472 14426 12481
rect 14370 12407 14426 12416
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14094 11384 14150 11393
rect 14004 11348 14056 11354
rect 14094 11319 14150 11328
rect 14004 11290 14056 11296
rect 13912 11280 13964 11286
rect 13912 11222 13964 11228
rect 14016 10810 14044 11290
rect 14108 11218 14136 11319
rect 14096 11212 14148 11218
rect 14096 11154 14148 11160
rect 14108 10810 14136 11154
rect 14200 11150 14228 12038
rect 14384 11801 14412 12174
rect 14370 11792 14426 11801
rect 14370 11727 14372 11736
rect 14424 11727 14426 11736
rect 14372 11698 14424 11704
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14004 10804 14056 10810
rect 14004 10746 14056 10752
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 13726 10160 13782 10169
rect 13726 10095 13782 10104
rect 14200 10010 14228 11086
rect 14108 9982 14228 10010
rect 14108 9926 14136 9982
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13924 9081 13952 9318
rect 13910 9072 13966 9081
rect 13910 9007 13966 9016
rect 13634 8936 13690 8945
rect 13634 8871 13690 8880
rect 13542 5128 13598 5137
rect 13542 5063 13598 5072
rect 13910 3632 13966 3641
rect 13910 3567 13966 3576
rect 13924 480 13952 3567
rect 14108 2650 14136 9862
rect 14476 9518 14504 13806
rect 14554 13560 14610 13569
rect 14554 13495 14610 13504
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14188 9444 14240 9450
rect 14188 9386 14240 9392
rect 14200 8838 14228 9386
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14200 3777 14228 8774
rect 14568 7857 14596 13495
rect 14660 12442 14688 14758
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14660 10538 14688 10950
rect 14648 10532 14700 10538
rect 14648 10474 14700 10480
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14660 9586 14688 9998
rect 14752 9654 14780 15302
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14844 14278 14872 14894
rect 15304 14890 15332 15438
rect 15292 14884 15344 14890
rect 15292 14826 15344 14832
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14844 13326 14872 14214
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14924 13796 14976 13802
rect 14924 13738 14976 13744
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 14936 13172 14964 13738
rect 14844 13144 14964 13172
rect 14844 10606 14872 13144
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15016 12708 15068 12714
rect 15016 12650 15068 12656
rect 15028 12617 15056 12650
rect 15108 12640 15160 12646
rect 15014 12608 15070 12617
rect 15160 12617 15332 12628
rect 15160 12608 15346 12617
rect 15160 12600 15290 12608
rect 15108 12582 15160 12588
rect 15014 12543 15070 12552
rect 15290 12543 15346 12552
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 14924 11552 14976 11558
rect 14924 11494 14976 11500
rect 14936 11286 14964 11494
rect 15028 11354 15056 11562
rect 15120 11558 15148 11630
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15304 11354 15332 12543
rect 15396 12442 15424 15846
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 14924 11280 14976 11286
rect 14924 11222 14976 11228
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15396 10810 15424 11630
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14844 10266 14872 10542
rect 15120 10266 15148 10610
rect 15488 10266 15516 15914
rect 15580 15366 15608 16526
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15658 13832 15714 13841
rect 15658 13767 15714 13776
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15580 12986 15608 13330
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15672 12866 15700 13767
rect 15580 12838 15700 12866
rect 15580 12442 15608 12838
rect 15660 12708 15712 12714
rect 15660 12650 15712 12656
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15580 11762 15608 12038
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15566 11656 15622 11665
rect 15566 11591 15622 11600
rect 15580 11558 15608 11591
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15580 10470 15608 11154
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15476 10260 15528 10266
rect 15476 10202 15528 10208
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14830 9616 14886 9625
rect 14648 9580 14700 9586
rect 14830 9551 14886 9560
rect 14648 9522 14700 9528
rect 14844 9382 14872 9551
rect 14832 9376 14884 9382
rect 14832 9318 14884 9324
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14554 7848 14610 7857
rect 14554 7783 14610 7792
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14186 3768 14242 3777
rect 14186 3703 14242 3712
rect 15580 3505 15608 10406
rect 15672 10130 15700 12650
rect 15764 12345 15792 17190
rect 15934 17167 15990 17176
rect 15936 16516 15988 16522
rect 16224 16504 16252 19638
rect 16408 19530 16436 20266
rect 16500 20074 16528 23559
rect 16592 23254 16620 23734
rect 16776 23322 16804 23802
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 16580 23248 16632 23254
rect 16868 23202 16896 25774
rect 16948 23520 17000 23526
rect 16948 23462 17000 23468
rect 16580 23190 16632 23196
rect 16592 22778 16620 23190
rect 16776 23174 16896 23202
rect 16580 22772 16632 22778
rect 16580 22714 16632 22720
rect 16592 22166 16620 22714
rect 16776 22409 16804 23174
rect 16854 23080 16910 23089
rect 16854 23015 16910 23024
rect 16868 22642 16896 23015
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 16762 22400 16818 22409
rect 16762 22335 16818 22344
rect 16580 22160 16632 22166
rect 16580 22102 16632 22108
rect 16670 21584 16726 21593
rect 16670 21519 16726 21528
rect 16684 21146 16712 21519
rect 16672 21140 16724 21146
rect 16672 21082 16724 21088
rect 16672 20392 16724 20398
rect 16672 20334 16724 20340
rect 16500 20046 16620 20074
rect 16684 20058 16712 20334
rect 16488 19984 16540 19990
rect 16488 19926 16540 19932
rect 16316 19502 16436 19530
rect 16316 19174 16344 19502
rect 16394 19408 16450 19417
rect 16500 19378 16528 19926
rect 16394 19343 16450 19352
rect 16488 19372 16540 19378
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16408 18329 16436 19343
rect 16488 19314 16540 19320
rect 16592 19258 16620 20046
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16684 19553 16712 19790
rect 16670 19544 16726 19553
rect 16670 19479 16726 19488
rect 16500 19230 16620 19258
rect 16394 18320 16450 18329
rect 16394 18255 16450 18264
rect 16500 17785 16528 19230
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16592 17882 16620 18770
rect 16684 18426 16712 19479
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16486 17776 16542 17785
rect 16486 17711 16542 17720
rect 16486 17640 16542 17649
rect 16486 17575 16542 17584
rect 16302 17504 16358 17513
rect 16302 17439 16358 17448
rect 15936 16458 15988 16464
rect 16132 16476 16252 16504
rect 15948 16250 15976 16458
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 16040 15570 16068 16050
rect 16028 15564 16080 15570
rect 16028 15506 16080 15512
rect 16040 15162 16068 15506
rect 16028 15156 16080 15162
rect 16028 15098 16080 15104
rect 16132 14090 16160 16476
rect 16210 16416 16266 16425
rect 16210 16351 16266 16360
rect 15948 14062 16160 14090
rect 15948 13802 15976 14062
rect 16026 13968 16082 13977
rect 16026 13903 16082 13912
rect 15936 13796 15988 13802
rect 15936 13738 15988 13744
rect 15934 13152 15990 13161
rect 15934 13087 15990 13096
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15856 12374 15884 12922
rect 15948 12714 15976 13087
rect 15936 12708 15988 12714
rect 15936 12650 15988 12656
rect 15844 12368 15896 12374
rect 15750 12336 15806 12345
rect 15844 12310 15896 12316
rect 15750 12271 15806 12280
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15764 11694 15792 12174
rect 15856 11778 15884 12310
rect 15936 12164 15988 12170
rect 15936 12106 15988 12112
rect 15948 11898 15976 12106
rect 15936 11892 15988 11898
rect 15936 11834 15988 11840
rect 16040 11801 16068 13903
rect 16120 12436 16172 12442
rect 16120 12378 16172 12384
rect 16026 11792 16082 11801
rect 15856 11762 15976 11778
rect 15856 11756 15988 11762
rect 15856 11750 15936 11756
rect 16026 11727 16082 11736
rect 15936 11698 15988 11704
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15948 11150 15976 11698
rect 16132 11642 16160 12378
rect 16224 12209 16252 16351
rect 16210 12200 16266 12209
rect 16210 12135 16266 12144
rect 16210 12064 16266 12073
rect 16210 11999 16266 12008
rect 16040 11614 16160 11642
rect 16040 11218 16068 11614
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 15948 10674 15976 11086
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 16040 10470 16068 11154
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15672 9654 15700 10066
rect 15764 9722 15792 10202
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15948 9722 15976 9998
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15936 9716 15988 9722
rect 15936 9658 15988 9664
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 16040 8945 16068 10406
rect 16026 8936 16082 8945
rect 16026 8871 16082 8880
rect 16224 7857 16252 11999
rect 16316 11762 16344 17439
rect 16500 17134 16528 17575
rect 16488 17128 16540 17134
rect 16488 17070 16540 17076
rect 16500 16794 16528 17070
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16592 16658 16620 17818
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16486 15328 16542 15337
rect 16486 15263 16542 15272
rect 16500 14618 16528 15263
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 16776 14498 16804 22335
rect 16960 21865 16988 23462
rect 16946 21856 17002 21865
rect 16946 21791 17002 21800
rect 17052 21690 17080 27520
rect 17604 25226 17632 27520
rect 17776 26036 17828 26042
rect 17776 25978 17828 25984
rect 17684 25288 17736 25294
rect 17684 25230 17736 25236
rect 17592 25220 17644 25226
rect 17592 25162 17644 25168
rect 17314 24848 17370 24857
rect 17314 24783 17370 24792
rect 17328 24614 17356 24783
rect 17696 24614 17724 25230
rect 17788 24818 17816 25978
rect 17776 24812 17828 24818
rect 17776 24754 17828 24760
rect 18156 24721 18184 27520
rect 18418 25936 18474 25945
rect 18418 25871 18474 25880
rect 18328 25152 18380 25158
rect 18328 25094 18380 25100
rect 18340 24954 18368 25094
rect 18328 24948 18380 24954
rect 18328 24890 18380 24896
rect 18432 24750 18460 25871
rect 18708 25344 18736 27520
rect 18524 25316 18736 25344
rect 18420 24744 18472 24750
rect 18142 24712 18198 24721
rect 18420 24686 18472 24692
rect 18142 24647 18198 24656
rect 18328 24676 18380 24682
rect 18328 24618 18380 24624
rect 17316 24608 17368 24614
rect 17316 24550 17368 24556
rect 17684 24608 17736 24614
rect 17684 24550 17736 24556
rect 18236 24608 18288 24614
rect 18236 24550 18288 24556
rect 17224 23792 17276 23798
rect 17224 23734 17276 23740
rect 17236 23322 17264 23734
rect 17224 23316 17276 23322
rect 17224 23258 17276 23264
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 17040 21684 17092 21690
rect 17040 21626 17092 21632
rect 17512 21418 17540 21830
rect 17500 21412 17552 21418
rect 17500 21354 17552 21360
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 16868 18902 16896 19110
rect 16856 18896 16908 18902
rect 16854 18864 16856 18873
rect 16908 18864 16910 18873
rect 16854 18799 16910 18808
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 16868 16046 16896 16390
rect 16960 16114 16988 21286
rect 17512 20777 17540 21354
rect 17696 21185 17724 24550
rect 18248 24410 18276 24550
rect 18236 24404 18288 24410
rect 18236 24346 18288 24352
rect 17776 24132 17828 24138
rect 17776 24074 17828 24080
rect 17788 22778 17816 24074
rect 17868 24064 17920 24070
rect 17868 24006 17920 24012
rect 17880 23594 17908 24006
rect 17868 23588 17920 23594
rect 17868 23530 17920 23536
rect 17776 22772 17828 22778
rect 17776 22714 17828 22720
rect 18340 22642 18368 24618
rect 18432 24342 18460 24686
rect 18420 24336 18472 24342
rect 18420 24278 18472 24284
rect 18432 22658 18460 24278
rect 18524 22817 18552 25316
rect 19260 25242 19288 27520
rect 19812 26194 19840 27520
rect 18616 25214 19288 25242
rect 19536 26166 19840 26194
rect 19432 25220 19484 25226
rect 18616 23361 18644 25214
rect 19432 25162 19484 25168
rect 18696 25152 18748 25158
rect 18696 25094 18748 25100
rect 18708 23662 18736 25094
rect 18788 24812 18840 24818
rect 18788 24754 18840 24760
rect 18800 24070 18828 24754
rect 19340 24608 19392 24614
rect 18892 24568 19340 24596
rect 18788 24064 18840 24070
rect 18788 24006 18840 24012
rect 18696 23656 18748 23662
rect 18696 23598 18748 23604
rect 18602 23352 18658 23361
rect 18602 23287 18658 23296
rect 18510 22808 18566 22817
rect 18510 22743 18566 22752
rect 18328 22636 18380 22642
rect 18432 22630 18644 22658
rect 18328 22578 18380 22584
rect 18052 22568 18104 22574
rect 18050 22536 18052 22545
rect 18104 22536 18106 22545
rect 18050 22471 18106 22480
rect 18328 22500 18380 22506
rect 18328 22442 18380 22448
rect 17960 22160 18012 22166
rect 17774 22128 17830 22137
rect 17830 22108 17960 22114
rect 17830 22102 18012 22108
rect 17830 22086 18000 22102
rect 17774 22063 17830 22072
rect 17788 21690 17816 22063
rect 18340 22001 18368 22442
rect 18510 22264 18566 22273
rect 18510 22199 18566 22208
rect 18420 22092 18472 22098
rect 18420 22034 18472 22040
rect 18326 21992 18382 22001
rect 18326 21927 18382 21936
rect 18144 21888 18196 21894
rect 18432 21842 18460 22034
rect 18144 21830 18196 21836
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 18156 21554 18184 21830
rect 18340 21814 18460 21842
rect 18144 21548 18196 21554
rect 18144 21490 18196 21496
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17682 21176 17738 21185
rect 17682 21111 17738 21120
rect 17592 21004 17644 21010
rect 17592 20946 17644 20952
rect 17498 20768 17554 20777
rect 17498 20703 17554 20712
rect 17604 20058 17632 20946
rect 17880 20398 17908 21286
rect 18052 21004 18104 21010
rect 18052 20946 18104 20952
rect 18064 20602 18092 20946
rect 18156 20913 18184 21490
rect 18340 21350 18368 21814
rect 18524 21486 18552 22199
rect 18512 21480 18564 21486
rect 18512 21422 18564 21428
rect 18328 21344 18380 21350
rect 18328 21286 18380 21292
rect 18142 20904 18198 20913
rect 18142 20839 18198 20848
rect 18052 20596 18104 20602
rect 18052 20538 18104 20544
rect 18236 20528 18288 20534
rect 18234 20496 18236 20505
rect 18288 20496 18290 20505
rect 18234 20431 18290 20440
rect 17868 20392 17920 20398
rect 17868 20334 17920 20340
rect 18144 20392 18196 20398
rect 18144 20334 18196 20340
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 17408 19916 17460 19922
rect 17408 19858 17460 19864
rect 17316 19848 17368 19854
rect 17316 19790 17368 19796
rect 17130 19544 17186 19553
rect 17130 19479 17186 19488
rect 17144 19310 17172 19479
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 17040 17536 17092 17542
rect 17040 17478 17092 17484
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16856 16040 16908 16046
rect 16856 15982 16908 15988
rect 16868 14618 16896 15982
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 16500 14470 16804 14498
rect 16500 14414 16528 14470
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16394 14104 16450 14113
rect 16394 14039 16450 14048
rect 16408 14006 16436 14039
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 16776 13802 16804 14470
rect 16764 13796 16816 13802
rect 16764 13738 16816 13744
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 16580 12708 16632 12714
rect 16580 12650 16632 12656
rect 16488 12640 16540 12646
rect 16486 12608 16488 12617
rect 16540 12608 16542 12617
rect 16486 12543 16542 12552
rect 16486 12472 16542 12481
rect 16486 12407 16542 12416
rect 16396 12300 16448 12306
rect 16396 12242 16448 12248
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16408 11354 16436 12242
rect 16500 12102 16528 12407
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16488 11620 16540 11626
rect 16592 11608 16620 12650
rect 16684 12170 16712 13126
rect 16776 12442 16804 13738
rect 17052 13569 17080 17478
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17236 14414 17264 15030
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17236 14074 17264 14350
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 17038 13560 17094 13569
rect 17038 13495 17094 13504
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 17328 12345 17356 19790
rect 17420 19514 17448 19858
rect 18156 19854 18184 20334
rect 18340 19961 18368 21286
rect 18326 19952 18382 19961
rect 18326 19887 18382 19896
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 17408 19508 17460 19514
rect 17408 19450 17460 19456
rect 17682 19272 17738 19281
rect 17682 19207 17684 19216
rect 17736 19207 17738 19216
rect 17866 19272 17922 19281
rect 17866 19207 17922 19216
rect 17684 19178 17736 19184
rect 17880 18970 17908 19207
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 17868 18964 17920 18970
rect 17868 18906 17920 18912
rect 17868 18828 17920 18834
rect 17868 18770 17920 18776
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17512 18426 17540 18702
rect 17500 18420 17552 18426
rect 17500 18362 17552 18368
rect 17408 17808 17460 17814
rect 17408 17750 17460 17756
rect 17420 16998 17448 17750
rect 17512 17377 17540 18362
rect 17788 18222 17816 18702
rect 17776 18216 17828 18222
rect 17774 18184 17776 18193
rect 17828 18184 17830 18193
rect 17774 18119 17830 18128
rect 17880 18086 17908 18770
rect 18064 18290 18092 19110
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 17684 18080 17736 18086
rect 17684 18022 17736 18028
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17498 17368 17554 17377
rect 17498 17303 17554 17312
rect 17592 17060 17644 17066
rect 17592 17002 17644 17008
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17420 16114 17448 16934
rect 17408 16108 17460 16114
rect 17408 16050 17460 16056
rect 17420 15910 17448 16050
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17420 15706 17448 15846
rect 17408 15700 17460 15706
rect 17408 15642 17460 15648
rect 17408 14408 17460 14414
rect 17406 14376 17408 14385
rect 17460 14376 17462 14385
rect 17406 14311 17462 14320
rect 17420 14074 17448 14311
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17604 13433 17632 17002
rect 17696 16998 17724 18022
rect 17880 17882 17908 18022
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 18156 17134 18184 19790
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17696 16590 17724 16934
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17696 15706 17724 16526
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17880 15858 17908 16594
rect 18052 16040 18104 16046
rect 18052 15982 18104 15988
rect 17960 15904 18012 15910
rect 17880 15852 17960 15858
rect 17880 15846 18012 15852
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17788 13734 17816 15846
rect 17880 15830 18000 15846
rect 17880 15162 17908 15830
rect 18064 15366 18092 15982
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 18052 15360 18104 15366
rect 18050 15328 18052 15337
rect 18104 15328 18106 15337
rect 18050 15263 18106 15272
rect 18156 15178 18184 15438
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 18064 15150 18184 15178
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17880 14618 17908 14894
rect 18064 14822 18092 15150
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17776 13728 17828 13734
rect 17880 13705 17908 14554
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17776 13670 17828 13676
rect 17866 13696 17922 13705
rect 17866 13631 17922 13640
rect 17972 13530 18000 14418
rect 18064 14414 18092 14758
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 18064 13938 18092 14350
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 17590 13424 17646 13433
rect 17590 13359 17646 13368
rect 18236 13388 18288 13394
rect 18236 13330 18288 13336
rect 18248 12986 18276 13330
rect 18340 13161 18368 19887
rect 18512 19236 18564 19242
rect 18512 19178 18564 19184
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 18432 18970 18460 19110
rect 18420 18964 18472 18970
rect 18420 18906 18472 18912
rect 18432 18737 18460 18906
rect 18524 18902 18552 19178
rect 18616 18970 18644 22630
rect 18708 22574 18736 23598
rect 18800 23594 18828 24006
rect 18788 23588 18840 23594
rect 18788 23530 18840 23536
rect 18696 22568 18748 22574
rect 18696 22510 18748 22516
rect 18696 22432 18748 22438
rect 18694 22400 18696 22409
rect 18748 22400 18750 22409
rect 18694 22335 18750 22344
rect 18800 22030 18828 23530
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18800 21622 18828 21966
rect 18788 21616 18840 21622
rect 18788 21558 18840 21564
rect 18892 20233 18920 24568
rect 19340 24550 19392 24556
rect 19340 24268 19392 24274
rect 19340 24210 19392 24216
rect 19352 23882 19380 24210
rect 19076 23854 19380 23882
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 18878 20224 18934 20233
rect 18878 20159 18934 20168
rect 18984 19802 19012 23054
rect 19076 21962 19104 23854
rect 19340 23792 19392 23798
rect 19340 23734 19392 23740
rect 19156 23588 19208 23594
rect 19156 23530 19208 23536
rect 19168 23050 19196 23530
rect 19248 23248 19300 23254
rect 19352 23236 19380 23734
rect 19300 23208 19380 23236
rect 19248 23190 19300 23196
rect 19156 23044 19208 23050
rect 19156 22986 19208 22992
rect 19154 22808 19210 22817
rect 19154 22743 19156 22752
rect 19208 22743 19210 22752
rect 19156 22714 19208 22720
rect 19156 22636 19208 22642
rect 19156 22578 19208 22584
rect 19064 21956 19116 21962
rect 19064 21898 19116 21904
rect 19168 21298 19196 22578
rect 19340 22568 19392 22574
rect 19340 22510 19392 22516
rect 19352 22166 19380 22510
rect 19340 22160 19392 22166
rect 19340 22102 19392 22108
rect 18892 19774 19012 19802
rect 19076 21270 19196 21298
rect 18604 18964 18656 18970
rect 18604 18906 18656 18912
rect 18512 18896 18564 18902
rect 18512 18838 18564 18844
rect 18418 18728 18474 18737
rect 18418 18663 18474 18672
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18432 18222 18460 18566
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 18420 17536 18472 17542
rect 18616 17524 18644 18226
rect 18472 17496 18644 17524
rect 18420 17478 18472 17484
rect 18432 17066 18460 17478
rect 18602 17368 18658 17377
rect 18602 17303 18658 17312
rect 18420 17060 18472 17066
rect 18420 17002 18472 17008
rect 18512 16652 18564 16658
rect 18512 16594 18564 16600
rect 18420 14952 18472 14958
rect 18420 14894 18472 14900
rect 18432 14113 18460 14894
rect 18524 14890 18552 16594
rect 18616 15638 18644 17303
rect 18892 16697 18920 19774
rect 18972 19712 19024 19718
rect 18972 19654 19024 19660
rect 18984 19378 19012 19654
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 18984 18766 19012 19314
rect 19076 19258 19104 21270
rect 19154 21176 19210 21185
rect 19154 21111 19156 21120
rect 19208 21111 19210 21120
rect 19156 21082 19208 21088
rect 19248 20936 19300 20942
rect 19300 20896 19380 20924
rect 19248 20878 19300 20884
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 19260 20398 19288 20742
rect 19352 20602 19380 20896
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19444 20516 19472 25162
rect 19536 24886 19564 26166
rect 20364 25974 20392 27520
rect 20352 25968 20404 25974
rect 20352 25910 20404 25916
rect 20442 25800 20498 25809
rect 20442 25735 20498 25744
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 20260 25424 20312 25430
rect 20260 25366 20312 25372
rect 19800 25356 19852 25362
rect 19800 25298 19852 25304
rect 20076 25356 20128 25362
rect 20076 25298 20128 25304
rect 19812 24886 19840 25298
rect 19984 25152 20036 25158
rect 19984 25094 20036 25100
rect 19524 24880 19576 24886
rect 19524 24822 19576 24828
rect 19800 24880 19852 24886
rect 19800 24822 19852 24828
rect 19996 24614 20024 25094
rect 20088 24886 20116 25298
rect 20076 24880 20128 24886
rect 20076 24822 20128 24828
rect 19984 24608 20036 24614
rect 19984 24550 20036 24556
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19984 24404 20036 24410
rect 19984 24346 20036 24352
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19536 23866 19564 24142
rect 19996 23866 20024 24346
rect 20088 24177 20116 24822
rect 20074 24168 20130 24177
rect 20074 24103 20130 24112
rect 19524 23860 19576 23866
rect 19524 23802 19576 23808
rect 19984 23860 20036 23866
rect 19984 23802 20036 23808
rect 19536 23322 19564 23802
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19524 23316 19576 23322
rect 19524 23258 19576 23264
rect 19536 22506 19564 23258
rect 19616 23180 19668 23186
rect 19616 23122 19668 23128
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 19628 22778 19656 23122
rect 19708 23112 19760 23118
rect 19708 23054 19760 23060
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19720 22506 19748 23054
rect 19984 22772 20036 22778
rect 19984 22714 20036 22720
rect 19524 22500 19576 22506
rect 19524 22442 19576 22448
rect 19708 22500 19760 22506
rect 19708 22442 19760 22448
rect 19536 22234 19564 22442
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19524 22228 19576 22234
rect 19996 22216 20024 22714
rect 20088 22234 20116 23122
rect 19524 22170 19576 22176
rect 19904 22188 20024 22216
rect 20076 22228 20128 22234
rect 19904 22030 19932 22188
rect 20076 22170 20128 22176
rect 20272 22030 20300 25366
rect 20456 24206 20484 25735
rect 20916 25650 20944 27520
rect 20824 25622 20944 25650
rect 20720 24608 20772 24614
rect 20720 24550 20772 24556
rect 20444 24200 20496 24206
rect 20444 24142 20496 24148
rect 20456 23866 20484 24142
rect 20536 24064 20588 24070
rect 20536 24006 20588 24012
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 20442 23760 20498 23769
rect 20442 23695 20498 23704
rect 20352 22976 20404 22982
rect 20352 22918 20404 22924
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 20076 22024 20128 22030
rect 20076 21966 20128 21972
rect 20260 22024 20312 22030
rect 20260 21966 20312 21972
rect 19984 21956 20036 21962
rect 19984 21898 20036 21904
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19435 20488 19472 20516
rect 19435 20448 19463 20488
rect 19435 20420 19472 20448
rect 19248 20392 19300 20398
rect 19248 20334 19300 20340
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19168 19446 19196 19858
rect 19156 19440 19208 19446
rect 19154 19408 19156 19417
rect 19208 19408 19210 19417
rect 19154 19343 19210 19352
rect 19076 19230 19196 19258
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 18984 17814 19012 18702
rect 19076 18426 19104 18906
rect 19064 18420 19116 18426
rect 19064 18362 19116 18368
rect 18972 17808 19024 17814
rect 18972 17750 19024 17756
rect 19168 17320 19196 19230
rect 19260 18952 19288 20334
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19352 19156 19380 20198
rect 19444 19310 19472 20420
rect 19524 20324 19576 20330
rect 19524 20266 19576 20272
rect 19536 20058 19564 20266
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 19432 19304 19484 19310
rect 19616 19304 19668 19310
rect 19432 19246 19484 19252
rect 19614 19272 19616 19281
rect 19668 19272 19670 19281
rect 19614 19207 19670 19216
rect 19352 19128 19472 19156
rect 19340 18964 19392 18970
rect 19260 18924 19340 18952
rect 19340 18906 19392 18912
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 19260 17864 19288 18158
rect 19340 17876 19392 17882
rect 19260 17836 19340 17864
rect 19340 17818 19392 17824
rect 19444 17762 19472 19128
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19892 18828 19944 18834
rect 19892 18770 19944 18776
rect 19904 18222 19932 18770
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19996 17814 20024 21898
rect 20088 17882 20116 21966
rect 20260 21888 20312 21894
rect 20260 21830 20312 21836
rect 20168 21072 20220 21078
rect 20168 21014 20220 21020
rect 20180 20058 20208 21014
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 20180 18834 20208 19110
rect 20168 18828 20220 18834
rect 20168 18770 20220 18776
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 19352 17734 19472 17762
rect 19984 17808 20036 17814
rect 20180 17762 20208 18770
rect 19984 17750 20036 17756
rect 19524 17740 19576 17746
rect 19168 17292 19288 17320
rect 18878 16688 18934 16697
rect 18878 16623 18934 16632
rect 19156 16584 19208 16590
rect 19156 16526 19208 16532
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18800 16114 18828 16390
rect 18788 16108 18840 16114
rect 18788 16050 18840 16056
rect 19168 15910 19196 16526
rect 19156 15904 19208 15910
rect 18786 15872 18842 15881
rect 19156 15846 19208 15852
rect 18786 15807 18842 15816
rect 18604 15632 18656 15638
rect 18604 15574 18656 15580
rect 18616 15162 18644 15574
rect 18604 15156 18656 15162
rect 18604 15098 18656 15104
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18512 14884 18564 14890
rect 18512 14826 18564 14832
rect 18616 14482 18644 14962
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18418 14104 18474 14113
rect 18418 14039 18474 14048
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 18326 13152 18382 13161
rect 18326 13087 18382 13096
rect 18236 12980 18288 12986
rect 18236 12922 18288 12928
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17314 12336 17370 12345
rect 17040 12300 17092 12306
rect 17314 12271 17370 12280
rect 17040 12242 17092 12248
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 16776 11830 16804 12038
rect 16764 11824 16816 11830
rect 16764 11766 16816 11772
rect 16540 11580 16620 11608
rect 16488 11562 16540 11568
rect 17052 11558 17080 12242
rect 17420 11898 17448 12378
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17696 11898 17724 12174
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17684 11892 17736 11898
rect 17684 11834 17736 11840
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16488 10260 16540 10266
rect 16592 10248 16620 11086
rect 16540 10220 16620 10248
rect 16488 10202 16540 10208
rect 16210 7848 16266 7857
rect 16210 7783 16266 7792
rect 17052 4593 17080 11494
rect 17788 9625 17816 12786
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18340 12442 18368 12718
rect 18524 12442 18552 13262
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18616 12374 18644 13262
rect 18694 12880 18750 12889
rect 18694 12815 18696 12824
rect 18748 12815 18750 12824
rect 18696 12786 18748 12792
rect 18604 12368 18656 12374
rect 18604 12310 18656 12316
rect 18800 12238 18828 15807
rect 19168 15337 19196 15846
rect 19154 15328 19210 15337
rect 19154 15263 19210 15272
rect 19260 15178 19288 17292
rect 19352 16561 19380 17734
rect 19524 17682 19576 17688
rect 20088 17734 20208 17762
rect 19430 17368 19486 17377
rect 19430 17303 19432 17312
rect 19484 17303 19486 17312
rect 19432 17274 19484 17280
rect 19536 16726 19564 17682
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19432 16720 19484 16726
rect 19432 16662 19484 16668
rect 19524 16720 19576 16726
rect 19524 16662 19576 16668
rect 19338 16552 19394 16561
rect 19338 16487 19394 16496
rect 19444 15910 19472 16662
rect 19536 16250 19564 16662
rect 19996 16425 20024 17614
rect 20088 16561 20116 17734
rect 20166 17640 20222 17649
rect 20166 17575 20222 17584
rect 20074 16552 20130 16561
rect 20180 16522 20208 17575
rect 20074 16487 20130 16496
rect 20168 16516 20220 16522
rect 20168 16458 20220 16464
rect 20076 16448 20128 16454
rect 19982 16416 20038 16425
rect 20076 16390 20128 16396
rect 20166 16416 20222 16425
rect 19982 16351 20038 16360
rect 19524 16244 19576 16250
rect 19524 16186 19576 16192
rect 20088 16114 20116 16390
rect 20166 16351 20222 16360
rect 20076 16108 20128 16114
rect 20076 16050 20128 16056
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19168 15150 19288 15178
rect 19064 14476 19116 14482
rect 19064 14418 19116 14424
rect 19076 14006 19104 14418
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 19076 13326 19104 13942
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 19168 13025 19196 15150
rect 19352 15042 19380 15370
rect 19260 15026 19380 15042
rect 19248 15020 19380 15026
rect 19300 15014 19380 15020
rect 19248 14962 19300 14968
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19154 13016 19210 13025
rect 19260 12986 19288 14826
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 19352 13569 19380 13670
rect 19338 13560 19394 13569
rect 19338 13495 19394 13504
rect 19444 13410 19472 15846
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 20074 15600 20130 15609
rect 20180 15586 20208 16351
rect 20130 15558 20208 15586
rect 20074 15535 20130 15544
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19536 14385 19564 14758
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19522 14376 19578 14385
rect 19522 14311 19578 14320
rect 19706 14376 19762 14385
rect 19706 14311 19708 14320
rect 19760 14311 19762 14320
rect 19708 14282 19760 14288
rect 19996 13802 20024 15302
rect 20088 14618 20116 15535
rect 20168 14884 20220 14890
rect 20168 14826 20220 14832
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 20074 14240 20130 14249
rect 20074 14175 20130 14184
rect 20088 14074 20116 14175
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 19984 13796 20036 13802
rect 19984 13738 20036 13744
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19352 13382 19472 13410
rect 19154 12951 19210 12960
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19248 12844 19300 12850
rect 19248 12786 19300 12792
rect 19156 12368 19208 12374
rect 19156 12310 19208 12316
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 18800 11937 18828 12174
rect 18786 11928 18842 11937
rect 18786 11863 18788 11872
rect 18840 11863 18842 11872
rect 18788 11834 18840 11840
rect 18800 11803 18828 11834
rect 19168 11558 19196 12310
rect 19260 12238 19288 12786
rect 19248 12232 19300 12238
rect 19248 12174 19300 12180
rect 19260 11898 19288 12174
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 17774 9616 17830 9625
rect 17774 9551 17830 9560
rect 19168 8537 19196 11494
rect 19352 11121 19380 13382
rect 19616 13320 19668 13326
rect 19616 13262 19668 13268
rect 19628 12782 19656 13262
rect 19706 13152 19762 13161
rect 19706 13087 19762 13096
rect 19720 12850 19748 13087
rect 19996 12918 20024 13738
rect 20180 13530 20208 14826
rect 20168 13524 20220 13530
rect 20168 13466 20220 13472
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 19708 12844 19760 12850
rect 19708 12786 19760 12792
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 19524 12708 19576 12714
rect 19524 12650 19576 12656
rect 19536 12442 19564 12650
rect 19996 12646 20024 12718
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 20180 12442 20208 13466
rect 20272 12782 20300 21830
rect 20364 20602 20392 22918
rect 20456 22114 20484 23695
rect 20548 23594 20576 24006
rect 20732 23848 20760 24550
rect 20824 24313 20852 25622
rect 20904 25492 20956 25498
rect 20904 25434 20956 25440
rect 20916 24410 20944 25434
rect 21560 25242 21588 27520
rect 21560 25214 21956 25242
rect 21548 25152 21600 25158
rect 21732 25152 21784 25158
rect 21600 25100 21680 25106
rect 21548 25094 21680 25100
rect 21732 25094 21784 25100
rect 21560 25078 21680 25094
rect 21456 24744 21508 24750
rect 21178 24712 21234 24721
rect 21456 24686 21508 24692
rect 21178 24647 21180 24656
rect 21232 24647 21234 24656
rect 21180 24618 21232 24624
rect 21364 24608 21416 24614
rect 21364 24550 21416 24556
rect 20904 24404 20956 24410
rect 20904 24346 20956 24352
rect 20810 24304 20866 24313
rect 20810 24239 20866 24248
rect 21088 24268 21140 24274
rect 21088 24210 21140 24216
rect 20732 23820 20944 23848
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20536 23588 20588 23594
rect 20536 23530 20588 23536
rect 20732 23322 20760 23666
rect 20812 23520 20864 23526
rect 20812 23462 20864 23468
rect 20720 23316 20772 23322
rect 20720 23258 20772 23264
rect 20824 23118 20852 23462
rect 20536 23112 20588 23118
rect 20812 23112 20864 23118
rect 20536 23054 20588 23060
rect 20640 23060 20812 23066
rect 20640 23054 20864 23060
rect 20548 22778 20576 23054
rect 20640 23038 20852 23054
rect 20536 22772 20588 22778
rect 20536 22714 20588 22720
rect 20548 22234 20576 22714
rect 20536 22228 20588 22234
rect 20536 22170 20588 22176
rect 20456 22086 20576 22114
rect 20548 21894 20576 22086
rect 20536 21888 20588 21894
rect 20442 21856 20498 21865
rect 20536 21830 20588 21836
rect 20442 21791 20498 21800
rect 20456 21418 20484 21791
rect 20640 21690 20668 23038
rect 20824 22989 20852 23038
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 20628 21684 20680 21690
rect 20628 21626 20680 21632
rect 20732 21554 20760 22170
rect 20812 21888 20864 21894
rect 20812 21830 20864 21836
rect 20720 21548 20772 21554
rect 20720 21490 20772 21496
rect 20444 21412 20496 21418
rect 20444 21354 20496 21360
rect 20456 21146 20484 21354
rect 20444 21140 20496 21146
rect 20444 21082 20496 21088
rect 20536 21140 20588 21146
rect 20536 21082 20588 21088
rect 20352 20596 20404 20602
rect 20352 20538 20404 20544
rect 20548 20330 20576 21082
rect 20718 21040 20774 21049
rect 20718 20975 20774 20984
rect 20732 20942 20760 20975
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20824 20806 20852 21830
rect 20812 20800 20864 20806
rect 20812 20742 20864 20748
rect 20916 20618 20944 23820
rect 21100 23526 21128 24210
rect 21272 24132 21324 24138
rect 21272 24074 21324 24080
rect 21088 23520 21140 23526
rect 21088 23462 21140 23468
rect 20996 22432 21048 22438
rect 20996 22374 21048 22380
rect 20824 20590 20944 20618
rect 20536 20324 20588 20330
rect 20536 20266 20588 20272
rect 20824 20210 20852 20590
rect 21008 20516 21036 22374
rect 20548 20182 20852 20210
rect 20916 20488 21036 20516
rect 20548 19145 20576 20182
rect 20720 19712 20772 19718
rect 20640 19660 20720 19666
rect 20640 19654 20772 19660
rect 20640 19638 20760 19654
rect 20534 19136 20590 19145
rect 20534 19071 20590 19080
rect 20444 17876 20496 17882
rect 20444 17818 20496 17824
rect 20352 17060 20404 17066
rect 20352 17002 20404 17008
rect 20364 13444 20392 17002
rect 20456 13705 20484 17818
rect 20548 17814 20576 19071
rect 20536 17808 20588 17814
rect 20536 17750 20588 17756
rect 20536 17604 20588 17610
rect 20536 17546 20588 17552
rect 20548 17202 20576 17546
rect 20640 17513 20668 19638
rect 20916 18766 20944 20488
rect 21100 20346 21128 23462
rect 21180 21072 21232 21078
rect 21180 21014 21232 21020
rect 21192 20602 21220 21014
rect 21180 20596 21232 20602
rect 21180 20538 21232 20544
rect 21008 20318 21128 20346
rect 21008 18850 21036 20318
rect 21284 19938 21312 24074
rect 21376 22137 21404 24550
rect 21468 24206 21496 24686
rect 21548 24676 21600 24682
rect 21548 24618 21600 24624
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21468 22982 21496 24142
rect 21456 22976 21508 22982
rect 21456 22918 21508 22924
rect 21454 22672 21510 22681
rect 21454 22607 21510 22616
rect 21468 22574 21496 22607
rect 21456 22568 21508 22574
rect 21456 22510 21508 22516
rect 21362 22128 21418 22137
rect 21362 22063 21418 22072
rect 21364 20324 21416 20330
rect 21364 20266 21416 20272
rect 21192 19910 21312 19938
rect 21088 19848 21140 19854
rect 21088 19790 21140 19796
rect 21100 19310 21128 19790
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 21100 18970 21128 19246
rect 21192 18970 21220 19910
rect 21270 19816 21326 19825
rect 21270 19751 21326 19760
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 21180 18964 21232 18970
rect 21180 18906 21232 18912
rect 21008 18822 21128 18850
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 20812 18692 20864 18698
rect 20812 18634 20864 18640
rect 20720 18352 20772 18358
rect 20720 18294 20772 18300
rect 20626 17504 20682 17513
rect 20626 17439 20682 17448
rect 20628 17332 20680 17338
rect 20732 17320 20760 18294
rect 20824 18290 20852 18634
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 20916 18290 20944 18566
rect 21008 18426 21036 18702
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20824 17746 20852 18226
rect 20812 17740 20864 17746
rect 20812 17682 20864 17688
rect 20824 17542 20852 17682
rect 20812 17536 20864 17542
rect 20812 17478 20864 17484
rect 20680 17292 20760 17320
rect 20628 17274 20680 17280
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20536 16516 20588 16522
rect 20536 16458 20588 16464
rect 20442 13696 20498 13705
rect 20442 13631 20498 13640
rect 20364 13416 20484 13444
rect 20350 13016 20406 13025
rect 20350 12951 20406 12960
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20364 12481 20392 12951
rect 20350 12472 20406 12481
rect 19524 12436 19576 12442
rect 19524 12378 19576 12384
rect 20168 12436 20220 12442
rect 20350 12407 20406 12416
rect 20168 12378 20220 12384
rect 19536 11540 19564 12378
rect 20180 11830 20208 12378
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 20456 11762 20484 13416
rect 20548 12209 20576 16458
rect 20640 16046 20668 17274
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20732 16794 20760 17070
rect 20824 16998 20852 17478
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20628 16040 20680 16046
rect 20628 15982 20680 15988
rect 20732 15434 20760 16730
rect 21100 16590 21128 18822
rect 21192 18737 21220 18906
rect 21178 18728 21234 18737
rect 21178 18663 21234 18672
rect 21192 18426 21220 18663
rect 21180 18420 21232 18426
rect 21180 18362 21232 18368
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20628 15360 20680 15366
rect 20628 15302 20680 15308
rect 20640 12646 20668 15302
rect 20824 14793 20852 16526
rect 21088 16448 21140 16454
rect 21088 16390 21140 16396
rect 21100 15978 21128 16390
rect 21088 15972 21140 15978
rect 21088 15914 21140 15920
rect 21100 15706 21128 15914
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 20810 14784 20866 14793
rect 20810 14719 20866 14728
rect 20916 14618 20944 15506
rect 21088 14952 21140 14958
rect 21088 14894 21140 14900
rect 21100 14618 21128 14894
rect 21192 14822 21220 16934
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 21284 14634 21312 19751
rect 21376 19718 21404 20266
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 21364 18828 21416 18834
rect 21364 18770 21416 18776
rect 21376 15638 21404 18770
rect 21468 18222 21496 22510
rect 21456 18216 21508 18222
rect 21456 18158 21508 18164
rect 21454 16008 21510 16017
rect 21454 15943 21456 15952
rect 21508 15943 21510 15952
rect 21456 15914 21508 15920
rect 21364 15632 21416 15638
rect 21456 15632 21508 15638
rect 21364 15574 21416 15580
rect 21454 15600 21456 15609
rect 21508 15600 21510 15609
rect 21454 15535 21510 15544
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 20904 14612 20956 14618
rect 20904 14554 20956 14560
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 21192 14606 21312 14634
rect 20996 14544 21048 14550
rect 20996 14486 21048 14492
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20824 13734 20852 14350
rect 21008 14074 21036 14486
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 20812 13728 20864 13734
rect 20812 13670 20864 13676
rect 20824 12850 20852 13670
rect 21088 13456 21140 13462
rect 21086 13424 21088 13433
rect 21140 13424 21142 13433
rect 20996 13388 21048 13394
rect 21086 13359 21142 13368
rect 20996 13330 21048 13336
rect 21008 12986 21036 13330
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 21008 12889 21036 12922
rect 20994 12880 21050 12889
rect 20812 12844 20864 12850
rect 20994 12815 21050 12824
rect 20812 12786 20864 12792
rect 21100 12782 21128 13359
rect 21192 13258 21220 14606
rect 21376 14550 21404 15438
rect 21456 15428 21508 15434
rect 21456 15370 21508 15376
rect 21468 15162 21496 15370
rect 21456 15156 21508 15162
rect 21456 15098 21508 15104
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21364 14544 21416 14550
rect 21364 14486 21416 14492
rect 21468 14414 21496 14758
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 21468 13938 21496 14350
rect 21456 13932 21508 13938
rect 21456 13874 21508 13880
rect 21364 13728 21416 13734
rect 21364 13670 21416 13676
rect 21376 13433 21404 13670
rect 21468 13530 21496 13874
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 21362 13424 21418 13433
rect 21362 13359 21418 13368
rect 21180 13252 21232 13258
rect 21180 13194 21232 13200
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 21456 12300 21508 12306
rect 21456 12242 21508 12248
rect 20534 12200 20590 12209
rect 20534 12135 20590 12144
rect 21468 11898 21496 12242
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 21468 11665 21496 11834
rect 21454 11656 21510 11665
rect 21454 11591 21510 11600
rect 19444 11512 19564 11540
rect 19444 11393 19472 11512
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19430 11384 19486 11393
rect 19622 11376 19918 11396
rect 19430 11319 19486 11328
rect 19338 11112 19394 11121
rect 19338 11047 19394 11056
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 21560 10033 21588 24618
rect 21652 24614 21680 25078
rect 21744 24886 21772 25094
rect 21732 24880 21784 24886
rect 21732 24822 21784 24828
rect 21640 24608 21692 24614
rect 21640 24550 21692 24556
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21652 22098 21680 23054
rect 21640 22092 21692 22098
rect 21640 22034 21692 22040
rect 21640 21344 21692 21350
rect 21640 21286 21692 21292
rect 21652 20398 21680 21286
rect 21640 20392 21692 20398
rect 21640 20334 21692 20340
rect 21640 20256 21692 20262
rect 21640 20198 21692 20204
rect 21652 18873 21680 20198
rect 21744 19417 21772 24822
rect 21824 24608 21876 24614
rect 21824 24550 21876 24556
rect 21836 23769 21864 24550
rect 21822 23760 21878 23769
rect 21822 23695 21878 23704
rect 21824 20800 21876 20806
rect 21824 20742 21876 20748
rect 21836 20466 21864 20742
rect 21824 20460 21876 20466
rect 21824 20402 21876 20408
rect 21836 19553 21864 20402
rect 21822 19544 21878 19553
rect 21822 19479 21878 19488
rect 21730 19408 21786 19417
rect 21730 19343 21786 19352
rect 21732 19236 21784 19242
rect 21732 19178 21784 19184
rect 21638 18864 21694 18873
rect 21744 18834 21772 19178
rect 21638 18799 21694 18808
rect 21732 18828 21784 18834
rect 21732 18770 21784 18776
rect 21640 17536 21692 17542
rect 21692 17496 21772 17524
rect 21640 17478 21692 17484
rect 21744 16590 21772 17496
rect 21732 16584 21784 16590
rect 21638 16552 21694 16561
rect 21732 16526 21784 16532
rect 21638 16487 21694 16496
rect 21652 12986 21680 16487
rect 21744 16182 21772 16526
rect 21732 16176 21784 16182
rect 21732 16118 21784 16124
rect 21732 16040 21784 16046
rect 21732 15982 21784 15988
rect 21928 15994 21956 25214
rect 22112 24410 22140 27520
rect 22468 25356 22520 25362
rect 22468 25298 22520 25304
rect 22284 25288 22336 25294
rect 22284 25230 22336 25236
rect 22100 24404 22152 24410
rect 22100 24346 22152 24352
rect 22192 24064 22244 24070
rect 22192 24006 22244 24012
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 22020 23338 22048 23666
rect 22204 23662 22232 24006
rect 22192 23656 22244 23662
rect 22192 23598 22244 23604
rect 22020 23310 22140 23338
rect 22112 23254 22140 23310
rect 22100 23248 22152 23254
rect 22100 23190 22152 23196
rect 22006 23080 22062 23089
rect 22006 23015 22062 23024
rect 22020 22778 22048 23015
rect 22112 22778 22140 23190
rect 22008 22772 22060 22778
rect 22008 22714 22060 22720
rect 22100 22772 22152 22778
rect 22100 22714 22152 22720
rect 22006 22536 22062 22545
rect 22006 22471 22062 22480
rect 22020 21690 22048 22471
rect 22112 22234 22140 22714
rect 22100 22228 22152 22234
rect 22100 22170 22152 22176
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 22100 21616 22152 21622
rect 22020 21564 22100 21570
rect 22020 21558 22152 21564
rect 22020 21554 22140 21558
rect 22008 21548 22140 21554
rect 22060 21542 22140 21548
rect 22008 21490 22060 21496
rect 22020 21146 22048 21490
rect 22100 21412 22152 21418
rect 22100 21354 22152 21360
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 22008 21004 22060 21010
rect 22008 20946 22060 20952
rect 22020 19990 22048 20946
rect 22112 20806 22140 21354
rect 22204 21146 22232 23598
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 22190 21040 22246 21049
rect 22190 20975 22246 20984
rect 22100 20800 22152 20806
rect 22100 20742 22152 20748
rect 22204 20330 22232 20975
rect 22192 20324 22244 20330
rect 22192 20266 22244 20272
rect 22008 19984 22060 19990
rect 22008 19926 22060 19932
rect 22100 19984 22152 19990
rect 22100 19926 22152 19932
rect 22006 19000 22062 19009
rect 22112 18986 22140 19926
rect 22062 18958 22140 18986
rect 22006 18935 22008 18944
rect 22060 18935 22062 18944
rect 22008 18906 22060 18912
rect 22020 18875 22048 18906
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 22112 18290 22140 18566
rect 22100 18284 22152 18290
rect 22152 18244 22232 18272
rect 22100 18226 22152 18232
rect 22100 18148 22152 18154
rect 22100 18090 22152 18096
rect 22112 17882 22140 18090
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 22204 17542 22232 18244
rect 22192 17536 22244 17542
rect 22192 17478 22244 17484
rect 22204 17134 22232 17478
rect 22192 17128 22244 17134
rect 22192 17070 22244 17076
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 22020 16726 22048 16934
rect 22190 16824 22246 16833
rect 22190 16759 22246 16768
rect 22008 16720 22060 16726
rect 22008 16662 22060 16668
rect 22020 16250 22048 16662
rect 22008 16244 22060 16250
rect 22008 16186 22060 16192
rect 21744 15638 21772 15982
rect 21824 15972 21876 15978
rect 21928 15966 22140 15994
rect 21824 15914 21876 15920
rect 21732 15632 21784 15638
rect 21732 15574 21784 15580
rect 21730 15192 21786 15201
rect 21730 15127 21786 15136
rect 21640 12980 21692 12986
rect 21640 12922 21692 12928
rect 21744 12442 21772 15127
rect 21836 14414 21864 15914
rect 22008 15904 22060 15910
rect 22008 15846 22060 15852
rect 22020 15745 22048 15846
rect 22006 15736 22062 15745
rect 22112 15706 22140 15966
rect 22006 15671 22062 15680
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 21914 15600 21970 15609
rect 21914 15535 21970 15544
rect 22100 15564 22152 15570
rect 21824 14408 21876 14414
rect 21824 14350 21876 14356
rect 21824 13864 21876 13870
rect 21822 13832 21824 13841
rect 21876 13832 21878 13841
rect 21822 13767 21878 13776
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21638 12064 21694 12073
rect 21638 11999 21694 12008
rect 21652 11665 21680 11999
rect 21928 11762 21956 15535
rect 22100 15506 22152 15512
rect 22008 14476 22060 14482
rect 22008 14418 22060 14424
rect 22020 14278 22048 14418
rect 22008 14272 22060 14278
rect 22008 14214 22060 14220
rect 22020 14006 22048 14214
rect 22008 14000 22060 14006
rect 22008 13942 22060 13948
rect 22112 13394 22140 15506
rect 22204 13734 22232 16759
rect 22296 14958 22324 25230
rect 22480 24614 22508 25298
rect 22664 24818 22692 27520
rect 23216 24970 23244 27520
rect 23124 24942 23244 24970
rect 22652 24812 22704 24818
rect 22652 24754 22704 24760
rect 23124 24682 23152 24942
rect 23768 24857 23796 27520
rect 24032 25900 24084 25906
rect 24032 25842 24084 25848
rect 23848 25356 23900 25362
rect 23848 25298 23900 25304
rect 23754 24848 23810 24857
rect 23204 24812 23256 24818
rect 23754 24783 23810 24792
rect 23204 24754 23256 24760
rect 22652 24676 22704 24682
rect 22652 24618 22704 24624
rect 23112 24676 23164 24682
rect 23112 24618 23164 24624
rect 22468 24608 22520 24614
rect 22468 24550 22520 24556
rect 22376 24064 22428 24070
rect 22376 24006 22428 24012
rect 22388 21078 22416 24006
rect 22560 23588 22612 23594
rect 22560 23530 22612 23536
rect 22572 22166 22600 23530
rect 22560 22160 22612 22166
rect 22466 22128 22522 22137
rect 22560 22102 22612 22108
rect 22466 22063 22522 22072
rect 22480 21486 22508 22063
rect 22468 21480 22520 21486
rect 22468 21422 22520 21428
rect 22376 21072 22428 21078
rect 22376 21014 22428 21020
rect 22480 20942 22508 21422
rect 22560 21344 22612 21350
rect 22560 21286 22612 21292
rect 22468 20936 22520 20942
rect 22468 20878 22520 20884
rect 22572 20806 22600 21286
rect 22376 20800 22428 20806
rect 22376 20742 22428 20748
rect 22560 20800 22612 20806
rect 22560 20742 22612 20748
rect 22388 16114 22416 20742
rect 22466 19408 22522 19417
rect 22466 19343 22522 19352
rect 22480 19174 22508 19343
rect 22468 19168 22520 19174
rect 22468 19110 22520 19116
rect 22558 19136 22614 19145
rect 22558 19071 22614 19080
rect 22572 18834 22600 19071
rect 22560 18828 22612 18834
rect 22560 18770 22612 18776
rect 22572 18426 22600 18770
rect 22560 18420 22612 18426
rect 22560 18362 22612 18368
rect 22560 18216 22612 18222
rect 22560 18158 22612 18164
rect 22466 16688 22522 16697
rect 22466 16623 22522 16632
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22388 15366 22416 16050
rect 22480 15570 22508 16623
rect 22468 15564 22520 15570
rect 22468 15506 22520 15512
rect 22376 15360 22428 15366
rect 22376 15302 22428 15308
rect 22480 15162 22508 15506
rect 22468 15156 22520 15162
rect 22468 15098 22520 15104
rect 22284 14952 22336 14958
rect 22284 14894 22336 14900
rect 22296 14618 22324 14894
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22376 14476 22428 14482
rect 22376 14418 22428 14424
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22192 13728 22244 13734
rect 22192 13670 22244 13676
rect 22100 13388 22152 13394
rect 22100 13330 22152 13336
rect 22112 12986 22140 13330
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 21916 11756 21968 11762
rect 21916 11698 21968 11704
rect 21638 11656 21694 11665
rect 21638 11591 21694 11600
rect 21546 10024 21602 10033
rect 21546 9959 21602 9968
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 22296 9081 22324 14350
rect 22388 13870 22416 14418
rect 22572 14385 22600 18158
rect 22558 14376 22614 14385
rect 22558 14311 22614 14320
rect 22560 14272 22612 14278
rect 22560 14214 22612 14220
rect 22572 13870 22600 14214
rect 22376 13864 22428 13870
rect 22376 13806 22428 13812
rect 22560 13864 22612 13870
rect 22560 13806 22612 13812
rect 22388 11354 22416 13806
rect 22664 13530 22692 24618
rect 23112 24404 23164 24410
rect 23112 24346 23164 24352
rect 22744 24336 22796 24342
rect 22744 24278 22796 24284
rect 22756 23526 22784 24278
rect 22836 24268 22888 24274
rect 22836 24210 22888 24216
rect 22744 23520 22796 23526
rect 22744 23462 22796 23468
rect 22756 18193 22784 23462
rect 22742 18184 22798 18193
rect 22742 18119 22798 18128
rect 22744 17672 22796 17678
rect 22744 17614 22796 17620
rect 22756 17338 22784 17614
rect 22744 17332 22796 17338
rect 22744 17274 22796 17280
rect 22742 16008 22798 16017
rect 22742 15943 22798 15952
rect 22756 14550 22784 15943
rect 22848 14618 22876 24210
rect 23020 24200 23072 24206
rect 23020 24142 23072 24148
rect 23032 23610 23060 24142
rect 22940 23582 23060 23610
rect 22940 23526 22968 23582
rect 22928 23520 22980 23526
rect 22928 23462 22980 23468
rect 22940 19786 22968 23462
rect 23020 22636 23072 22642
rect 23020 22578 23072 22584
rect 23032 22234 23060 22578
rect 23020 22228 23072 22234
rect 23020 22170 23072 22176
rect 23020 20868 23072 20874
rect 23020 20810 23072 20816
rect 23032 20602 23060 20810
rect 23020 20596 23072 20602
rect 23020 20538 23072 20544
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 23032 20058 23060 20198
rect 23020 20052 23072 20058
rect 23020 19994 23072 20000
rect 22928 19780 22980 19786
rect 22928 19722 22980 19728
rect 22940 19378 22968 19722
rect 22928 19372 22980 19378
rect 22928 19314 22980 19320
rect 22926 19000 22982 19009
rect 22926 18935 22982 18944
rect 22940 15162 22968 18935
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 23032 17542 23060 18566
rect 23020 17536 23072 17542
rect 23020 17478 23072 17484
rect 23124 16708 23152 24346
rect 23032 16680 23152 16708
rect 22928 15156 22980 15162
rect 22928 15098 22980 15104
rect 23032 14958 23060 16680
rect 23216 16658 23244 24754
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23294 23760 23350 23769
rect 23294 23695 23350 23704
rect 23308 18970 23336 23695
rect 23400 22982 23428 24550
rect 23664 23520 23716 23526
rect 23664 23462 23716 23468
rect 23676 23254 23704 23462
rect 23664 23248 23716 23254
rect 23664 23190 23716 23196
rect 23572 23044 23624 23050
rect 23572 22986 23624 22992
rect 23388 22976 23440 22982
rect 23388 22918 23440 22924
rect 23584 22574 23612 22986
rect 23572 22568 23624 22574
rect 23572 22510 23624 22516
rect 23756 22500 23808 22506
rect 23756 22442 23808 22448
rect 23480 22432 23532 22438
rect 23480 22374 23532 22380
rect 23492 22166 23520 22374
rect 23570 22264 23626 22273
rect 23570 22199 23626 22208
rect 23480 22160 23532 22166
rect 23480 22102 23532 22108
rect 23388 22092 23440 22098
rect 23388 22034 23440 22040
rect 23400 21162 23428 22034
rect 23478 21720 23534 21729
rect 23478 21655 23534 21664
rect 23492 21486 23520 21655
rect 23480 21480 23532 21486
rect 23480 21422 23532 21428
rect 23492 21350 23520 21422
rect 23480 21344 23532 21350
rect 23478 21312 23480 21321
rect 23532 21312 23534 21321
rect 23478 21247 23534 21256
rect 23400 21134 23520 21162
rect 23492 21078 23520 21134
rect 23480 21072 23532 21078
rect 23480 21014 23532 21020
rect 23388 21004 23440 21010
rect 23388 20946 23440 20952
rect 23400 20602 23428 20946
rect 23480 20800 23532 20806
rect 23480 20742 23532 20748
rect 23388 20596 23440 20602
rect 23388 20538 23440 20544
rect 23388 20460 23440 20466
rect 23388 20402 23440 20408
rect 23296 18964 23348 18970
rect 23296 18906 23348 18912
rect 23296 18760 23348 18766
rect 23296 18702 23348 18708
rect 23204 16652 23256 16658
rect 23204 16594 23256 16600
rect 23112 16448 23164 16454
rect 23112 16390 23164 16396
rect 23124 16250 23152 16390
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 23308 16028 23336 18702
rect 23216 16000 23336 16028
rect 23112 15088 23164 15094
rect 23112 15030 23164 15036
rect 23020 14952 23072 14958
rect 23020 14894 23072 14900
rect 22836 14612 22888 14618
rect 22836 14554 22888 14560
rect 22744 14544 22796 14550
rect 22744 14486 22796 14492
rect 22756 14074 22784 14486
rect 23124 14414 23152 15030
rect 23112 14408 23164 14414
rect 23112 14350 23164 14356
rect 22744 14068 22796 14074
rect 22744 14010 22796 14016
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22652 13524 22704 13530
rect 22652 13466 22704 13472
rect 22756 12442 22784 13670
rect 23124 13530 23152 14350
rect 23112 13524 23164 13530
rect 23112 13466 23164 13472
rect 23216 12986 23244 16000
rect 23400 15960 23428 20402
rect 23492 19786 23520 20742
rect 23584 20505 23612 22199
rect 23768 22030 23796 22442
rect 23756 22024 23808 22030
rect 23756 21966 23808 21972
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23676 21146 23704 21286
rect 23664 21140 23716 21146
rect 23664 21082 23716 21088
rect 23768 21010 23796 21966
rect 23860 21185 23888 25298
rect 24044 24818 24072 25842
rect 24032 24812 24084 24818
rect 24032 24754 24084 24760
rect 24044 24154 24072 24754
rect 24136 24410 24164 27639
rect 24306 27520 24362 28000
rect 24858 27520 24914 28000
rect 25410 27520 25466 28000
rect 25962 27520 26018 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 24320 25140 24348 27520
rect 24674 27160 24730 27169
rect 24674 27095 24730 27104
rect 24228 25112 24348 25140
rect 24228 24721 24256 25112
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24214 24712 24270 24721
rect 24214 24647 24270 24656
rect 24688 24614 24716 27095
rect 24766 26480 24822 26489
rect 24766 26415 24822 26424
rect 24780 25498 24808 26415
rect 24768 25492 24820 25498
rect 24768 25434 24820 25440
rect 24768 25220 24820 25226
rect 24768 25162 24820 25168
rect 24780 24721 24808 25162
rect 24766 24712 24822 24721
rect 24766 24647 24822 24656
rect 24872 24614 24900 27520
rect 25424 25922 25452 27520
rect 24964 25894 25452 25922
rect 25502 25936 25558 25945
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 24860 24608 24912 24614
rect 24860 24550 24912 24556
rect 24124 24404 24176 24410
rect 24124 24346 24176 24352
rect 24676 24268 24728 24274
rect 24676 24210 24728 24216
rect 23952 24126 24072 24154
rect 23952 23866 23980 24126
rect 24032 24064 24084 24070
rect 24032 24006 24084 24012
rect 23940 23860 23992 23866
rect 23940 23802 23992 23808
rect 23940 23588 23992 23594
rect 23940 23530 23992 23536
rect 23846 21176 23902 21185
rect 23846 21111 23902 21120
rect 23848 21072 23900 21078
rect 23848 21014 23900 21020
rect 23756 21004 23808 21010
rect 23756 20946 23808 20952
rect 23570 20496 23626 20505
rect 23570 20431 23626 20440
rect 23572 20392 23624 20398
rect 23570 20360 23572 20369
rect 23624 20360 23626 20369
rect 23570 20295 23626 20304
rect 23754 20360 23810 20369
rect 23754 20295 23810 20304
rect 23480 19780 23532 19786
rect 23480 19722 23532 19728
rect 23480 19304 23532 19310
rect 23480 19246 23532 19252
rect 23492 18329 23520 19246
rect 23664 19168 23716 19174
rect 23664 19110 23716 19116
rect 23572 18896 23624 18902
rect 23572 18838 23624 18844
rect 23478 18320 23534 18329
rect 23584 18290 23612 18838
rect 23478 18255 23534 18264
rect 23572 18284 23624 18290
rect 23572 18226 23624 18232
rect 23478 17912 23534 17921
rect 23478 17847 23534 17856
rect 23308 15932 23428 15960
rect 23308 14074 23336 15932
rect 23492 15858 23520 17847
rect 23572 17672 23624 17678
rect 23572 17614 23624 17620
rect 23400 15830 23520 15858
rect 23400 15201 23428 15830
rect 23478 15736 23534 15745
rect 23478 15671 23480 15680
rect 23532 15671 23534 15680
rect 23480 15642 23532 15648
rect 23584 15434 23612 17614
rect 23572 15428 23624 15434
rect 23572 15370 23624 15376
rect 23386 15192 23442 15201
rect 23386 15127 23442 15136
rect 23386 15056 23442 15065
rect 23676 15026 23704 19110
rect 23768 18834 23796 20295
rect 23860 18873 23888 21014
rect 23952 20398 23980 23530
rect 24044 23526 24072 24006
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24216 23724 24268 23730
rect 24216 23666 24268 23672
rect 24032 23520 24084 23526
rect 24032 23462 24084 23468
rect 24044 23186 24072 23462
rect 24228 23322 24256 23666
rect 24688 23594 24716 24210
rect 24768 23656 24820 23662
rect 24768 23598 24820 23604
rect 24676 23588 24728 23594
rect 24676 23530 24728 23536
rect 24780 23474 24808 23598
rect 24688 23446 24808 23474
rect 24216 23316 24268 23322
rect 24216 23258 24268 23264
rect 24032 23180 24084 23186
rect 24032 23122 24084 23128
rect 24122 22672 24178 22681
rect 24122 22607 24178 22616
rect 24030 21584 24086 21593
rect 24030 21519 24086 21528
rect 23940 20392 23992 20398
rect 23940 20334 23992 20340
rect 23940 19712 23992 19718
rect 23940 19654 23992 19660
rect 23952 19378 23980 19654
rect 23940 19372 23992 19378
rect 23940 19314 23992 19320
rect 23846 18864 23902 18873
rect 23756 18828 23808 18834
rect 23952 18834 23980 19314
rect 23846 18799 23902 18808
rect 23940 18828 23992 18834
rect 23756 18770 23808 18776
rect 23940 18770 23992 18776
rect 23952 18426 23980 18770
rect 23940 18420 23992 18426
rect 23940 18362 23992 18368
rect 23754 18320 23810 18329
rect 23754 18255 23810 18264
rect 23768 16833 23796 18255
rect 23846 18184 23902 18193
rect 23846 18119 23902 18128
rect 23940 18148 23992 18154
rect 23754 16824 23810 16833
rect 23754 16759 23810 16768
rect 23756 16448 23808 16454
rect 23756 16390 23808 16396
rect 23768 16046 23796 16390
rect 23756 16040 23808 16046
rect 23756 15982 23808 15988
rect 23756 15564 23808 15570
rect 23756 15506 23808 15512
rect 23386 14991 23442 15000
rect 23664 15020 23716 15026
rect 23296 14068 23348 14074
rect 23296 14010 23348 14016
rect 23294 13016 23350 13025
rect 23204 12980 23256 12986
rect 23294 12951 23350 12960
rect 23204 12922 23256 12928
rect 22744 12436 22796 12442
rect 23308 12424 23336 12951
rect 22744 12378 22796 12384
rect 23216 12396 23336 12424
rect 23020 12368 23072 12374
rect 22558 12336 22614 12345
rect 23216 12322 23244 12396
rect 23020 12310 23072 12316
rect 22558 12271 22560 12280
rect 22612 12271 22614 12280
rect 22560 12242 22612 12248
rect 22572 11898 22600 12242
rect 22560 11892 22612 11898
rect 22560 11834 22612 11840
rect 23032 11762 23060 12310
rect 23124 12294 23244 12322
rect 23296 12300 23348 12306
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 22468 11688 22520 11694
rect 22468 11630 22520 11636
rect 22480 11354 22508 11630
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 23124 11234 23152 12294
rect 23296 12242 23348 12248
rect 23202 11928 23258 11937
rect 23202 11863 23258 11872
rect 23216 11529 23244 11863
rect 23202 11520 23258 11529
rect 23202 11455 23258 11464
rect 23308 11234 23336 12242
rect 23400 11898 23428 14991
rect 23664 14962 23716 14968
rect 23768 14890 23796 15506
rect 23860 15162 23888 18119
rect 23940 18090 23992 18096
rect 23952 17678 23980 18090
rect 24044 18086 24072 21519
rect 24032 18080 24084 18086
rect 24032 18022 24084 18028
rect 24032 17740 24084 17746
rect 24032 17682 24084 17688
rect 23940 17672 23992 17678
rect 23940 17614 23992 17620
rect 23952 17338 23980 17614
rect 23940 17332 23992 17338
rect 23940 17274 23992 17280
rect 24044 16794 24072 17682
rect 24032 16788 24084 16794
rect 24032 16730 24084 16736
rect 24032 16584 24084 16590
rect 24032 16526 24084 16532
rect 24044 16250 24072 16526
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 24044 16017 24072 16186
rect 24030 16008 24086 16017
rect 24030 15943 24086 15952
rect 23940 15904 23992 15910
rect 23940 15846 23992 15852
rect 23848 15156 23900 15162
rect 23848 15098 23900 15104
rect 23756 14884 23808 14890
rect 23756 14826 23808 14832
rect 23664 14544 23716 14550
rect 23664 14486 23716 14492
rect 23570 13424 23626 13433
rect 23570 13359 23626 13368
rect 23480 13320 23532 13326
rect 23480 13262 23532 13268
rect 23388 11892 23440 11898
rect 23388 11834 23440 11840
rect 23492 11370 23520 13262
rect 23584 12306 23612 13359
rect 23572 12300 23624 12306
rect 23572 12242 23624 12248
rect 23570 11520 23626 11529
rect 23570 11455 23626 11464
rect 23400 11354 23520 11370
rect 23388 11348 23520 11354
rect 23440 11342 23520 11348
rect 23388 11290 23440 11296
rect 23124 11206 23244 11234
rect 23308 11206 23520 11234
rect 23216 10418 23244 11206
rect 23492 10577 23520 11206
rect 23478 10568 23534 10577
rect 23478 10503 23534 10512
rect 23216 10390 23520 10418
rect 22282 9072 22338 9081
rect 22282 9007 22338 9016
rect 19154 8528 19210 8537
rect 19154 8463 19210 8472
rect 17958 8392 18014 8401
rect 17958 8327 18014 8336
rect 17972 7449 18000 8327
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 17958 7440 18014 7449
rect 17958 7375 18014 7384
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 23492 6089 23520 10390
rect 23584 7041 23612 11455
rect 23676 11354 23704 14486
rect 23768 13433 23796 14826
rect 23848 13728 23900 13734
rect 23952 13716 23980 15846
rect 24030 15464 24086 15473
rect 24030 15399 24086 15408
rect 24044 14958 24072 15399
rect 24032 14952 24084 14958
rect 24032 14894 24084 14900
rect 24044 14618 24072 14894
rect 24136 14618 24164 22607
rect 24228 22574 24256 23258
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24216 22568 24268 22574
rect 24216 22510 24268 22516
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24688 21672 24716 23446
rect 24768 23180 24820 23186
rect 24768 23122 24820 23128
rect 24780 23089 24808 23122
rect 24860 23112 24912 23118
rect 24766 23080 24822 23089
rect 24860 23054 24912 23060
rect 24766 23015 24822 23024
rect 24780 22778 24808 23015
rect 24768 22772 24820 22778
rect 24768 22714 24820 22720
rect 24872 22522 24900 23054
rect 24780 22494 24900 22522
rect 24780 22438 24808 22494
rect 24768 22432 24820 22438
rect 24768 22374 24820 22380
rect 24780 22166 24808 22374
rect 24768 22160 24820 22166
rect 24768 22102 24820 22108
rect 24780 21690 24808 22102
rect 24596 21644 24716 21672
rect 24768 21684 24820 21690
rect 24308 21548 24360 21554
rect 24308 21490 24360 21496
rect 24320 21078 24348 21490
rect 24308 21072 24360 21078
rect 24214 21040 24270 21049
rect 24308 21014 24360 21020
rect 24214 20975 24270 20984
rect 24228 16454 24256 20975
rect 24596 20913 24624 21644
rect 24768 21626 24820 21632
rect 24676 21072 24728 21078
rect 24676 21014 24728 21020
rect 24582 20904 24638 20913
rect 24582 20839 24638 20848
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24688 20602 24716 21014
rect 24768 21004 24820 21010
rect 24768 20946 24820 20952
rect 24780 20618 24808 20946
rect 24676 20596 24728 20602
rect 24780 20590 24900 20618
rect 24676 20538 24728 20544
rect 24872 20534 24900 20590
rect 24860 20528 24912 20534
rect 24860 20470 24912 20476
rect 24308 20460 24360 20466
rect 24308 20402 24360 20408
rect 24320 20058 24348 20402
rect 24308 20052 24360 20058
rect 24308 19994 24360 20000
rect 24768 19916 24820 19922
rect 24768 19858 24820 19864
rect 24676 19780 24728 19786
rect 24676 19722 24728 19728
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24584 19440 24636 19446
rect 24688 19417 24716 19722
rect 24584 19382 24636 19388
rect 24674 19408 24730 19417
rect 24596 19174 24624 19382
rect 24674 19343 24676 19352
rect 24728 19343 24730 19352
rect 24676 19314 24728 19320
rect 24688 19283 24716 19314
rect 24780 19174 24808 19858
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 24872 19446 24900 19790
rect 24860 19440 24912 19446
rect 24860 19382 24912 19388
rect 24308 19168 24360 19174
rect 24306 19136 24308 19145
rect 24584 19168 24636 19174
rect 24360 19136 24362 19145
rect 24584 19110 24636 19116
rect 24768 19168 24820 19174
rect 24768 19110 24820 19116
rect 24306 19071 24362 19080
rect 24596 18737 24624 19110
rect 24582 18728 24638 18737
rect 24582 18663 24638 18672
rect 24768 18624 24820 18630
rect 24768 18566 24820 18572
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24780 18222 24808 18566
rect 24768 18216 24820 18222
rect 24768 18158 24820 18164
rect 24780 17898 24808 18158
rect 24780 17882 24900 17898
rect 24780 17876 24912 17882
rect 24780 17870 24860 17876
rect 24860 17818 24912 17824
rect 24676 17536 24728 17542
rect 24676 17478 24728 17484
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24308 17060 24360 17066
rect 24308 17002 24360 17008
rect 24320 16522 24348 17002
rect 24688 16998 24716 17478
rect 24766 17368 24822 17377
rect 24766 17303 24822 17312
rect 24676 16992 24728 16998
rect 24676 16934 24728 16940
rect 24676 16720 24728 16726
rect 24676 16662 24728 16668
rect 24308 16516 24360 16522
rect 24308 16458 24360 16464
rect 24216 16448 24268 16454
rect 24216 16390 24268 16396
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24214 16144 24270 16153
rect 24214 16079 24270 16088
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 24124 14612 24176 14618
rect 24124 14554 24176 14560
rect 24228 14550 24256 16079
rect 24584 15632 24636 15638
rect 24582 15600 24584 15609
rect 24688 15620 24716 16662
rect 24780 16561 24808 17303
rect 24964 17218 24992 25894
rect 25502 25871 25558 25880
rect 25044 25764 25096 25770
rect 25044 25706 25096 25712
rect 25056 17814 25084 25706
rect 25136 25356 25188 25362
rect 25136 25298 25188 25304
rect 25148 24886 25176 25298
rect 25412 24948 25464 24954
rect 25412 24890 25464 24896
rect 25136 24880 25188 24886
rect 25136 24822 25188 24828
rect 25136 24608 25188 24614
rect 25136 24550 25188 24556
rect 25148 23322 25176 24550
rect 25424 23610 25452 24890
rect 25240 23582 25452 23610
rect 25136 23316 25188 23322
rect 25136 23258 25188 23264
rect 25136 21888 25188 21894
rect 25136 21830 25188 21836
rect 25148 21690 25176 21830
rect 25136 21684 25188 21690
rect 25136 21626 25188 21632
rect 25240 21486 25268 23582
rect 25412 23520 25464 23526
rect 25410 23488 25412 23497
rect 25464 23488 25466 23497
rect 25410 23423 25466 23432
rect 25320 23316 25372 23322
rect 25320 23258 25372 23264
rect 25228 21480 25280 21486
rect 25228 21422 25280 21428
rect 25228 20392 25280 20398
rect 25228 20334 25280 20340
rect 25240 19961 25268 20334
rect 25226 19952 25282 19961
rect 25226 19887 25282 19896
rect 25228 19712 25280 19718
rect 25228 19654 25280 19660
rect 25240 19310 25268 19654
rect 25228 19304 25280 19310
rect 25226 19272 25228 19281
rect 25280 19272 25282 19281
rect 25226 19207 25282 19216
rect 25228 19168 25280 19174
rect 25228 19110 25280 19116
rect 25134 19000 25190 19009
rect 25134 18935 25136 18944
rect 25188 18935 25190 18944
rect 25136 18906 25188 18912
rect 25134 18864 25190 18873
rect 25134 18799 25190 18808
rect 25044 17808 25096 17814
rect 25044 17750 25096 17756
rect 24964 17190 25084 17218
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 24766 16552 24822 16561
rect 24766 16487 24822 16496
rect 24768 16448 24820 16454
rect 24768 16390 24820 16396
rect 24636 15600 24716 15620
rect 24638 15592 24716 15600
rect 24582 15535 24638 15544
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24688 15162 24716 15438
rect 24676 15156 24728 15162
rect 24676 15098 24728 15104
rect 24216 14544 24268 14550
rect 24216 14486 24268 14492
rect 24032 14476 24084 14482
rect 24032 14418 24084 14424
rect 23900 13688 23980 13716
rect 23848 13670 23900 13676
rect 23754 13424 23810 13433
rect 23754 13359 23810 13368
rect 23756 13252 23808 13258
rect 23756 13194 23808 13200
rect 23768 12628 23796 13194
rect 23860 13190 23888 13670
rect 23940 13388 23992 13394
rect 23940 13330 23992 13336
rect 23952 13258 23980 13330
rect 23940 13252 23992 13258
rect 23940 13194 23992 13200
rect 23848 13184 23900 13190
rect 23848 13126 23900 13132
rect 23860 12782 23888 13126
rect 24044 13025 24072 14418
rect 24216 14408 24268 14414
rect 24216 14350 24268 14356
rect 24122 13832 24178 13841
rect 24122 13767 24178 13776
rect 24030 13016 24086 13025
rect 24030 12951 24086 12960
rect 24136 12889 24164 13767
rect 24122 12880 24178 12889
rect 24122 12815 24178 12824
rect 23848 12776 23900 12782
rect 23848 12718 23900 12724
rect 24032 12708 24084 12714
rect 24032 12650 24084 12656
rect 23768 12600 23888 12628
rect 23860 11898 23888 12600
rect 24044 12102 24072 12650
rect 24228 12322 24256 14350
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24780 13410 24808 16390
rect 24872 15434 24900 16594
rect 24952 16516 25004 16522
rect 24952 16458 25004 16464
rect 24964 16250 24992 16458
rect 24952 16244 25004 16250
rect 24952 16186 25004 16192
rect 24964 15706 24992 16186
rect 24952 15700 25004 15706
rect 24952 15642 25004 15648
rect 24964 15502 24992 15642
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 24860 15428 24912 15434
rect 24860 15370 24912 15376
rect 24952 14000 25004 14006
rect 24952 13942 25004 13948
rect 24780 13382 24900 13410
rect 24674 13288 24730 13297
rect 24674 13223 24730 13232
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24688 12866 24716 13223
rect 24136 12294 24256 12322
rect 24504 12838 24716 12866
rect 24032 12096 24084 12102
rect 24032 12038 24084 12044
rect 24044 11898 24072 12038
rect 23848 11892 23900 11898
rect 23848 11834 23900 11840
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 23940 11756 23992 11762
rect 24136 11744 24164 12294
rect 24504 12186 24532 12838
rect 24582 12744 24638 12753
rect 24872 12730 24900 13382
rect 24964 12918 24992 13942
rect 24952 12912 25004 12918
rect 24952 12854 25004 12860
rect 24582 12679 24638 12688
rect 24688 12702 24900 12730
rect 24596 12374 24624 12679
rect 24584 12368 24636 12374
rect 24688 12345 24716 12702
rect 24768 12640 24820 12646
rect 24768 12582 24820 12588
rect 24860 12640 24912 12646
rect 24860 12582 24912 12588
rect 24584 12310 24636 12316
rect 24674 12336 24730 12345
rect 24674 12271 24730 12280
rect 24504 12158 24716 12186
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 23940 11698 23992 11704
rect 24044 11716 24164 11744
rect 23664 11348 23716 11354
rect 23664 11290 23716 11296
rect 23952 11286 23980 11698
rect 23940 11280 23992 11286
rect 23940 11222 23992 11228
rect 24044 11218 24072 11716
rect 24124 11620 24176 11626
rect 24124 11562 24176 11568
rect 24032 11212 24084 11218
rect 24032 11154 24084 11160
rect 23754 11112 23810 11121
rect 23754 11047 23810 11056
rect 23664 8424 23716 8430
rect 23662 8392 23664 8401
rect 23716 8392 23718 8401
rect 23662 8327 23718 8336
rect 23662 7848 23718 7857
rect 23662 7783 23718 7792
rect 23570 7032 23626 7041
rect 23570 6967 23626 6976
rect 23478 6080 23534 6089
rect 19622 6012 19918 6032
rect 23478 6015 23534 6024
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 23478 5128 23534 5137
rect 23478 5063 23534 5072
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 17038 4584 17094 4593
rect 17038 4519 17094 4528
rect 17958 4210 18014 4219
rect 17958 4145 18014 4154
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 15566 3496 15622 3505
rect 15566 3431 15622 3440
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 19522 2952 19578 2961
rect 19522 2887 19578 2896
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 19536 480 19564 2887
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 23492 2417 23520 5063
rect 23676 2689 23704 7783
rect 23768 6361 23796 11047
rect 23938 10840 23994 10849
rect 24044 10810 24072 11154
rect 24136 11082 24164 11562
rect 24582 11248 24638 11257
rect 24582 11183 24584 11192
rect 24636 11183 24638 11192
rect 24584 11154 24636 11160
rect 24124 11076 24176 11082
rect 24124 11018 24176 11024
rect 23938 10775 23994 10784
rect 24032 10804 24084 10810
rect 23754 6352 23810 6361
rect 23754 6287 23810 6296
rect 23662 2680 23718 2689
rect 23662 2615 23718 2624
rect 23478 2408 23534 2417
rect 23478 2343 23534 2352
rect 23952 1465 23980 10775
rect 24032 10746 24084 10752
rect 24030 5808 24086 5817
rect 24030 5743 24032 5752
rect 24084 5743 24086 5752
rect 24032 5714 24084 5720
rect 24044 5370 24072 5714
rect 24032 5364 24084 5370
rect 24032 5306 24084 5312
rect 24136 4826 24164 11018
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24582 10704 24638 10713
rect 24582 10639 24638 10648
rect 24596 10606 24624 10639
rect 24584 10600 24636 10606
rect 24584 10542 24636 10548
rect 24688 10130 24716 12158
rect 24780 11694 24808 12582
rect 24872 12442 24900 12582
rect 24860 12436 24912 12442
rect 24860 12378 24912 12384
rect 24860 12300 24912 12306
rect 24860 12242 24912 12248
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24768 11212 24820 11218
rect 24768 11154 24820 11160
rect 24780 10810 24808 11154
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24872 10690 24900 12242
rect 24780 10662 24900 10690
rect 24676 10124 24728 10130
rect 24676 10066 24728 10072
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24688 9722 24716 10066
rect 24676 9716 24728 9722
rect 24676 9658 24728 9664
rect 24216 9648 24268 9654
rect 24216 9590 24268 9596
rect 24228 5914 24256 9590
rect 24674 8936 24730 8945
rect 24674 8871 24730 8880
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24216 5908 24268 5914
rect 24216 5850 24268 5856
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5137 24716 8871
rect 24780 7585 24808 10662
rect 24766 7576 24822 7585
rect 24766 7511 24822 7520
rect 24964 5250 24992 12854
rect 25056 12186 25084 17190
rect 25148 15570 25176 18799
rect 25240 17134 25268 19110
rect 25228 17128 25280 17134
rect 25228 17070 25280 17076
rect 25228 16992 25280 16998
rect 25228 16934 25280 16940
rect 25240 16454 25268 16934
rect 25228 16448 25280 16454
rect 25228 16390 25280 16396
rect 25240 15910 25268 16390
rect 25228 15904 25280 15910
rect 25228 15846 25280 15852
rect 25136 15564 25188 15570
rect 25136 15506 25188 15512
rect 25148 14550 25176 15506
rect 25332 15162 25360 23258
rect 25412 21548 25464 21554
rect 25412 21490 25464 21496
rect 25424 21457 25452 21490
rect 25410 21448 25466 21457
rect 25410 21383 25466 21392
rect 25516 19174 25544 25871
rect 25594 25256 25650 25265
rect 25594 25191 25650 25200
rect 25608 20602 25636 25191
rect 25872 23248 25924 23254
rect 25872 23190 25924 23196
rect 25884 22778 25912 23190
rect 25872 22772 25924 22778
rect 25872 22714 25924 22720
rect 25596 20596 25648 20602
rect 25596 20538 25648 20544
rect 25504 19168 25556 19174
rect 25504 19110 25556 19116
rect 25778 19136 25834 19145
rect 25778 19071 25834 19080
rect 25502 18728 25558 18737
rect 25502 18663 25558 18672
rect 25412 18080 25464 18086
rect 25412 18022 25464 18028
rect 25320 15156 25372 15162
rect 25320 15098 25372 15104
rect 25228 14952 25280 14958
rect 25228 14894 25280 14900
rect 25136 14544 25188 14550
rect 25136 14486 25188 14492
rect 25056 12158 25176 12186
rect 25044 12096 25096 12102
rect 25044 12038 25096 12044
rect 25056 11665 25084 12038
rect 25042 11656 25098 11665
rect 25042 11591 25098 11600
rect 25148 8634 25176 12158
rect 25240 10985 25268 14894
rect 25424 13410 25452 18022
rect 25516 14482 25544 18663
rect 25688 17604 25740 17610
rect 25688 17546 25740 17552
rect 25700 17338 25728 17546
rect 25688 17332 25740 17338
rect 25688 17274 25740 17280
rect 25594 14784 25650 14793
rect 25594 14719 25650 14728
rect 25504 14476 25556 14482
rect 25504 14418 25556 14424
rect 25516 14074 25544 14418
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25332 13382 25452 13410
rect 25332 11354 25360 13382
rect 25412 13320 25464 13326
rect 25412 13262 25464 13268
rect 25424 12714 25452 13262
rect 25412 12708 25464 12714
rect 25412 12650 25464 12656
rect 25502 11792 25558 11801
rect 25502 11727 25558 11736
rect 25516 11694 25544 11727
rect 25504 11688 25556 11694
rect 25504 11630 25556 11636
rect 25320 11348 25372 11354
rect 25320 11290 25372 11296
rect 25608 11257 25636 14719
rect 25686 12336 25742 12345
rect 25686 12271 25742 12280
rect 25700 11898 25728 12271
rect 25688 11892 25740 11898
rect 25688 11834 25740 11840
rect 25594 11248 25650 11257
rect 25594 11183 25650 11192
rect 25226 10976 25282 10985
rect 25226 10911 25282 10920
rect 25792 10470 25820 19071
rect 25780 10464 25832 10470
rect 25780 10406 25832 10412
rect 25976 9654 26004 27520
rect 26332 22432 26384 22438
rect 26332 22374 26384 22380
rect 26344 21350 26372 22374
rect 26332 21344 26384 21350
rect 26332 21286 26384 21292
rect 26344 20602 26372 21286
rect 26332 20596 26384 20602
rect 26332 20538 26384 20544
rect 26148 19168 26200 19174
rect 26148 19110 26200 19116
rect 26160 18630 26188 19110
rect 26148 18624 26200 18630
rect 26148 18566 26200 18572
rect 26160 17338 26188 18566
rect 26148 17332 26200 17338
rect 26148 17274 26200 17280
rect 26054 16688 26110 16697
rect 26054 16623 26110 16632
rect 26068 10266 26096 16623
rect 26528 15337 26556 27520
rect 27080 27470 27108 27520
rect 27068 27464 27120 27470
rect 27068 27406 27120 27412
rect 27342 24576 27398 24585
rect 27632 24562 27660 27520
rect 27398 24534 27660 24562
rect 27342 24511 27398 24520
rect 26514 15328 26570 15337
rect 26514 15263 26570 15272
rect 26056 10260 26108 10266
rect 26056 10202 26108 10208
rect 26240 9716 26292 9722
rect 26240 9658 26292 9664
rect 25964 9648 26016 9654
rect 26252 9625 26280 9658
rect 25964 9590 26016 9596
rect 26238 9616 26294 9625
rect 26238 9551 26294 9560
rect 26514 9616 26570 9625
rect 26514 9551 26570 9560
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 24780 5222 24992 5250
rect 24674 5128 24730 5137
rect 24674 5063 24730 5072
rect 24124 4820 24176 4826
rect 24124 4762 24176 4768
rect 24676 4752 24728 4758
rect 24676 4694 24728 4700
rect 24124 4684 24176 4690
rect 24124 4626 24176 4632
rect 24136 4214 24164 4626
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24124 4208 24176 4214
rect 24688 4162 24716 4694
rect 24780 4622 24808 5222
rect 24768 4616 24820 4622
rect 24768 4558 24820 4564
rect 24780 4214 24808 4558
rect 24124 4150 24176 4156
rect 24596 4134 24716 4162
rect 24768 4208 24820 4214
rect 24768 4150 24820 4156
rect 24596 3942 24624 4134
rect 24584 3936 24636 3942
rect 24582 3904 24584 3913
rect 24636 3904 24638 3913
rect 24582 3839 24638 3848
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 25134 2952 25190 2961
rect 25134 2887 25190 2896
rect 25148 2514 25176 2887
rect 26528 2650 26556 9551
rect 26516 2644 26568 2650
rect 26516 2586 26568 2592
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 23938 1456 23994 1465
rect 23938 1391 23994 1400
rect 20350 912 20406 921
rect 20350 847 20406 856
rect 13450 96 13506 105
rect 13450 31 13506 40
rect 13910 0 13966 480
rect 19522 0 19578 480
rect 20364 105 20392 847
rect 25148 480 25176 2246
rect 20350 96 20406 105
rect 20350 31 20406 40
rect 25134 0 25190 480
<< via2 >>
rect 3514 27648 3570 27704
rect 1950 25744 2006 25800
rect 846 22616 902 22672
rect 1490 23704 1546 23760
rect 1582 21528 1638 21584
rect 1398 20304 1454 20360
rect 24122 27648 24178 27704
rect 3054 25880 3110 25936
rect 4066 27104 4122 27160
rect 4066 26424 4122 26480
rect 3882 25608 3938 25664
rect 2042 24556 2044 24576
rect 2044 24556 2096 24576
rect 2096 24556 2098 24576
rect 2042 24520 2098 24556
rect 2042 24404 2098 24440
rect 2042 24384 2044 24404
rect 2044 24384 2096 24404
rect 2096 24384 2098 24404
rect 2318 24112 2374 24168
rect 2870 23976 2926 24032
rect 2686 23432 2742 23488
rect 3790 25200 3846 25256
rect 2962 22752 3018 22808
rect 1766 22208 1822 22264
rect 1858 22072 1914 22128
rect 1674 20032 1730 20088
rect 2962 22228 3018 22264
rect 2962 22208 2964 22228
rect 2964 22208 3016 22228
rect 3016 22208 3018 22228
rect 2870 22108 2872 22128
rect 2872 22108 2924 22128
rect 2924 22108 2926 22128
rect 2870 22072 2926 22108
rect 2410 21120 2466 21176
rect 202 15816 258 15872
rect 1766 17176 1822 17232
rect 3054 20984 3110 21040
rect 2594 19252 2596 19272
rect 2596 19252 2648 19272
rect 2648 19252 2650 19272
rect 2594 19216 2650 19252
rect 2502 18964 2558 19000
rect 2502 18944 2504 18964
rect 2504 18944 2556 18964
rect 2556 18944 2558 18964
rect 1582 16088 1638 16144
rect 1490 15408 1546 15464
rect 1306 9968 1362 10024
rect 1766 15564 1822 15600
rect 1766 15544 1768 15564
rect 1768 15544 1820 15564
rect 1820 15544 1822 15564
rect 3238 17856 3294 17912
rect 1582 9424 1638 9480
rect 570 4528 626 4584
rect 2870 13096 2926 13152
rect 2778 3984 2834 4040
rect 1950 3168 2006 3224
rect 938 856 994 912
rect 4250 24656 4306 24712
rect 3606 23432 3662 23488
rect 3698 19080 3754 19136
rect 3514 17992 3570 18048
rect 3606 15544 3662 15600
rect 3790 18536 3846 18592
rect 3974 20440 4030 20496
rect 3974 19760 4030 19816
rect 3974 17856 4030 17912
rect 4526 22752 4582 22808
rect 4526 21140 4582 21176
rect 4526 21120 4528 21140
rect 4528 21120 4580 21140
rect 4580 21120 4582 21140
rect 3790 16088 3846 16144
rect 3698 14864 3754 14920
rect 3790 13640 3846 13696
rect 3146 2760 3202 2816
rect 3698 12588 3700 12608
rect 3700 12588 3752 12608
rect 3752 12588 3754 12608
rect 3698 12552 3754 12588
rect 4066 15000 4122 15056
rect 4066 14320 4122 14376
rect 3974 11600 4030 11656
rect 3698 10104 3754 10160
rect 3882 9016 3938 9072
rect 3882 6976 3938 7032
rect 3698 6296 3754 6352
rect 3330 2080 3386 2136
rect 4526 16768 4582 16824
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5262 24248 5318 24304
rect 4894 23604 4896 23624
rect 4896 23604 4948 23624
rect 4948 23604 4950 23624
rect 4894 23568 4950 23604
rect 4894 21528 4950 21584
rect 4802 19080 4858 19136
rect 5262 22480 5318 22536
rect 5170 20440 5226 20496
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 6182 23432 6238 23488
rect 6090 23296 6146 23352
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 6274 22616 6330 22672
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5262 18944 5318 19000
rect 4710 11328 4766 11384
rect 4986 13776 5042 13832
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5998 19216 6054 19272
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 6642 23976 6698 24032
rect 7010 24384 7066 24440
rect 6366 22072 6422 22128
rect 6458 21140 6514 21176
rect 6458 21120 6460 21140
rect 6460 21120 6512 21140
rect 6512 21120 6514 21140
rect 7010 21256 7066 21312
rect 6274 19216 6330 19272
rect 6734 20440 6790 20496
rect 6826 20340 6828 20360
rect 6828 20340 6880 20360
rect 6880 20340 6882 20360
rect 6826 20304 6882 20340
rect 7286 23840 7342 23896
rect 7378 23468 7380 23488
rect 7380 23468 7432 23488
rect 7432 23468 7434 23488
rect 7378 23432 7434 23468
rect 8022 23316 8078 23352
rect 8022 23296 8024 23316
rect 8024 23296 8076 23316
rect 8076 23296 8078 23316
rect 8022 22888 8078 22944
rect 7930 22752 7986 22808
rect 8114 22344 8170 22400
rect 8114 21412 8170 21448
rect 8114 21392 8116 21412
rect 8116 21392 8168 21412
rect 8168 21392 8170 21412
rect 8574 24248 8630 24304
rect 7654 20032 7710 20088
rect 7378 19352 7434 19408
rect 6734 17876 6790 17912
rect 6734 17856 6736 17876
rect 6736 17856 6788 17876
rect 6788 17856 6790 17876
rect 6734 17176 6790 17232
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5446 15680 5502 15736
rect 5078 13640 5134 13696
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5814 14864 5870 14920
rect 5906 14728 5962 14784
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5538 13676 5540 13696
rect 5540 13676 5592 13696
rect 5592 13676 5594 13696
rect 5538 13640 5594 13676
rect 5814 13640 5870 13696
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 4526 11092 4528 11112
rect 4528 11092 4580 11112
rect 4580 11092 4582 11112
rect 4526 11056 4582 11092
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 6734 16632 6790 16688
rect 6642 16496 6698 16552
rect 6458 15816 6514 15872
rect 6918 17856 6974 17912
rect 7102 16632 7158 16688
rect 6918 16360 6974 16416
rect 7010 16124 7012 16144
rect 7012 16124 7064 16144
rect 7064 16124 7066 16144
rect 7010 16088 7066 16124
rect 7194 16108 7250 16144
rect 7194 16088 7196 16108
rect 7196 16088 7248 16108
rect 7248 16088 7250 16108
rect 7562 19352 7618 19408
rect 7562 16788 7618 16824
rect 7562 16768 7564 16788
rect 7564 16768 7616 16788
rect 7616 16768 7618 16788
rect 7654 15680 7710 15736
rect 7470 15544 7526 15600
rect 7378 15000 7434 15056
rect 7286 13932 7342 13968
rect 7286 13912 7288 13932
rect 7288 13912 7340 13932
rect 7340 13912 7342 13932
rect 6918 13504 6974 13560
rect 6090 12552 6146 12608
rect 6458 12824 6514 12880
rect 7470 14864 7526 14920
rect 8942 24812 8998 24848
rect 8942 24792 8944 24812
rect 8944 24792 8996 24812
rect 8996 24792 8998 24812
rect 8850 24676 8906 24712
rect 8850 24656 8852 24676
rect 8852 24656 8904 24676
rect 8904 24656 8906 24676
rect 9678 24404 9734 24440
rect 9678 24384 9680 24404
rect 9680 24384 9732 24404
rect 9732 24384 9734 24404
rect 9034 23060 9036 23080
rect 9036 23060 9088 23080
rect 9088 23060 9090 23080
rect 9034 23024 9090 23060
rect 9126 22072 9182 22128
rect 9402 21936 9458 21992
rect 8482 18964 8538 19000
rect 8482 18944 8484 18964
rect 8484 18944 8536 18964
rect 8536 18944 8538 18964
rect 8022 18672 8078 18728
rect 8390 18672 8446 18728
rect 8114 18128 8170 18184
rect 8022 17720 8078 17776
rect 7746 14320 7802 14376
rect 8574 17448 8630 17504
rect 8206 13812 8208 13832
rect 8208 13812 8260 13832
rect 8260 13812 8262 13832
rect 8206 13776 8262 13812
rect 7838 11328 7894 11384
rect 5998 11056 6054 11112
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 6182 9988 6238 10024
rect 6182 9968 6184 9988
rect 6184 9968 6236 9988
rect 6236 9968 6238 9988
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 4066 8200 4122 8256
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 4066 7384 4122 7440
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 3974 5072 4030 5128
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 8206 4120 8262 4176
rect 9586 24248 9642 24304
rect 10322 26016 10378 26072
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 9770 22752 9826 22808
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10782 24384 10838 24440
rect 10966 24556 10968 24576
rect 10968 24556 11020 24576
rect 11020 24556 11022 24576
rect 10966 24520 11022 24556
rect 10782 24112 10838 24168
rect 10966 23976 11022 24032
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 9954 22652 9956 22672
rect 9956 22652 10008 22672
rect 10008 22652 10010 22672
rect 9954 22616 10010 22652
rect 9954 22208 10010 22264
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 9862 22072 9918 22128
rect 9678 21120 9734 21176
rect 10046 21292 10048 21312
rect 10048 21292 10100 21312
rect 10100 21292 10102 21312
rect 10046 21256 10102 21292
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 9218 19624 9274 19680
rect 9494 19760 9550 19816
rect 9678 19080 9734 19136
rect 9494 18400 9550 18456
rect 9402 18264 9458 18320
rect 9586 17212 9588 17232
rect 9588 17212 9640 17232
rect 9640 17212 9642 17232
rect 9586 17176 9642 17212
rect 9678 16652 9734 16688
rect 9678 16632 9680 16652
rect 9680 16632 9732 16652
rect 9732 16632 9734 16652
rect 9310 13640 9366 13696
rect 9586 13640 9642 13696
rect 9586 12960 9642 13016
rect 10966 23568 11022 23624
rect 10874 20576 10930 20632
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10690 18264 10746 18320
rect 10046 17992 10102 18048
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 9954 17856 10010 17912
rect 10690 17856 10746 17912
rect 9862 17584 9918 17640
rect 9954 17312 10010 17368
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10782 15680 10838 15736
rect 10046 15036 10048 15056
rect 10048 15036 10100 15056
rect 10100 15036 10102 15056
rect 10046 15000 10102 15036
rect 10506 14900 10508 14920
rect 10508 14900 10560 14920
rect 10560 14900 10562 14920
rect 10506 14864 10562 14900
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10966 20460 11022 20496
rect 10966 20440 10968 20460
rect 10968 20440 11020 20460
rect 11020 20440 11022 20460
rect 11150 24112 11206 24168
rect 11058 18400 11114 18456
rect 10966 17584 11022 17640
rect 10966 16224 11022 16280
rect 10874 13912 10930 13968
rect 11242 21936 11298 21992
rect 11426 22652 11428 22672
rect 11428 22652 11480 22672
rect 11480 22652 11482 22672
rect 11426 22616 11482 22652
rect 11426 21956 11482 21992
rect 11426 21936 11428 21956
rect 11428 21936 11480 21956
rect 11480 21936 11482 21956
rect 11242 18264 11298 18320
rect 11242 18148 11298 18184
rect 11242 18128 11244 18148
rect 11244 18128 11296 18148
rect 11296 18128 11298 18148
rect 11426 18400 11482 18456
rect 11426 16768 11482 16824
rect 11794 23296 11850 23352
rect 11702 21528 11758 21584
rect 11978 21256 12034 21312
rect 11886 20984 11942 21040
rect 12070 19352 12126 19408
rect 12714 24656 12770 24712
rect 12438 20576 12494 20632
rect 12346 19760 12402 19816
rect 11702 15952 11758 16008
rect 10782 12688 10838 12744
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 11058 11192 11114 11248
rect 12070 12144 12126 12200
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 9678 9696 9734 9752
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 9678 3984 9734 4040
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 9126 3576 9182 3632
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 8298 2896 8354 2952
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 3698 1400 3754 1456
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 13082 24792 13138 24848
rect 12714 20440 12770 20496
rect 13542 24112 13598 24168
rect 13174 23840 13230 23896
rect 13082 23432 13138 23488
rect 12990 20460 13046 20496
rect 12990 20440 12992 20460
rect 12992 20440 13044 20460
rect 13044 20440 13046 20460
rect 13266 20340 13268 20360
rect 13268 20340 13320 20360
rect 13320 20340 13322 20360
rect 13266 20304 13322 20340
rect 12530 16224 12586 16280
rect 12438 15000 12494 15056
rect 12438 10784 12494 10840
rect 12622 10784 12678 10840
rect 12438 10512 12494 10568
rect 13174 19080 13230 19136
rect 12990 15544 13046 15600
rect 12070 9696 12126 9752
rect 13082 12144 13138 12200
rect 13174 10784 13230 10840
rect 12806 9560 12862 9616
rect 12438 2896 12494 2952
rect 1306 312 1362 368
rect 13450 16088 13506 16144
rect 13726 21548 13782 21584
rect 13726 21528 13728 21548
rect 13728 21528 13780 21548
rect 13780 21528 13782 21548
rect 14094 24112 14150 24168
rect 14370 24812 14426 24848
rect 14370 24792 14372 24812
rect 14372 24792 14424 24812
rect 14424 24792 14426 24812
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 13910 23316 13966 23352
rect 13910 23296 13912 23316
rect 13912 23296 13964 23316
rect 13964 23296 13966 23316
rect 14278 23432 14334 23488
rect 14278 22752 14334 22808
rect 14094 19660 14096 19680
rect 14096 19660 14148 19680
rect 14148 19660 14150 19680
rect 14094 19624 14150 19660
rect 13634 17584 13690 17640
rect 13726 16496 13782 16552
rect 13634 16088 13690 16144
rect 13450 15700 13506 15736
rect 13450 15680 13452 15700
rect 13452 15680 13504 15700
rect 13504 15680 13506 15700
rect 13450 15544 13506 15600
rect 13174 176 13230 232
rect 13726 15816 13782 15872
rect 14094 18808 14150 18864
rect 14002 16788 14058 16824
rect 14002 16768 14004 16788
rect 14004 16768 14056 16788
rect 14056 16768 14058 16788
rect 15382 24520 15438 24576
rect 14738 22888 14794 22944
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14922 22208 14978 22264
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15382 21528 15438 21584
rect 14738 20848 14794 20904
rect 14462 17584 14518 17640
rect 14554 17448 14610 17504
rect 15382 20712 15438 20768
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 15566 24384 15622 24440
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 15566 18536 15622 18592
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 15290 17876 15346 17912
rect 15290 17856 15292 17876
rect 15292 17856 15344 17876
rect 15344 17856 15346 17876
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 15750 19116 15752 19136
rect 15752 19116 15804 19136
rect 15804 19116 15806 19136
rect 15750 19080 15806 19116
rect 15750 17740 15806 17776
rect 15750 17720 15752 17740
rect 15752 17720 15804 17740
rect 15804 17720 15806 17740
rect 16394 24792 16450 24848
rect 16118 23568 16174 23624
rect 16118 20848 16174 20904
rect 16486 23568 16542 23624
rect 16394 21120 16450 21176
rect 15934 17212 15936 17232
rect 15936 17212 15988 17232
rect 15988 17212 15990 17232
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14002 13640 14058 13696
rect 14002 12960 14058 13016
rect 14278 15136 14334 15192
rect 14186 13232 14242 13288
rect 14002 12824 14058 12880
rect 13818 11636 13820 11656
rect 13820 11636 13872 11656
rect 13872 11636 13874 11656
rect 13818 11600 13874 11636
rect 14094 12280 14150 12336
rect 14370 12416 14426 12472
rect 14094 11328 14150 11384
rect 14370 11756 14426 11792
rect 14370 11736 14372 11756
rect 14372 11736 14424 11756
rect 14424 11736 14426 11756
rect 13726 10104 13782 10160
rect 13910 9016 13966 9072
rect 13634 8880 13690 8936
rect 13542 5072 13598 5128
rect 13910 3576 13966 3632
rect 14554 13504 14610 13560
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15014 12552 15070 12608
rect 15290 12552 15346 12608
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15658 13776 15714 13832
rect 15566 11600 15622 11656
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14830 9560 14886 9616
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14554 7792 14610 7848
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14186 3712 14242 3768
rect 15934 17176 15990 17212
rect 16854 23024 16910 23080
rect 16762 22344 16818 22400
rect 16670 21528 16726 21584
rect 16394 19352 16450 19408
rect 16670 19488 16726 19544
rect 16394 18264 16450 18320
rect 16486 17720 16542 17776
rect 16486 17584 16542 17640
rect 16302 17448 16358 17504
rect 16210 16360 16266 16416
rect 16026 13912 16082 13968
rect 15934 13096 15990 13152
rect 15750 12280 15806 12336
rect 16026 11736 16082 11792
rect 16210 12144 16266 12200
rect 16210 12008 16266 12064
rect 16026 8880 16082 8936
rect 16486 15272 16542 15328
rect 16946 21800 17002 21856
rect 17314 24792 17370 24848
rect 18418 25880 18474 25936
rect 18142 24656 18198 24712
rect 16854 18844 16856 18864
rect 16856 18844 16908 18864
rect 16908 18844 16910 18864
rect 16854 18808 16910 18844
rect 18602 23296 18658 23352
rect 18510 22752 18566 22808
rect 18050 22516 18052 22536
rect 18052 22516 18104 22536
rect 18104 22516 18106 22536
rect 18050 22480 18106 22516
rect 17774 22072 17830 22128
rect 18510 22208 18566 22264
rect 18326 21936 18382 21992
rect 17682 21120 17738 21176
rect 17498 20712 17554 20768
rect 18142 20848 18198 20904
rect 18234 20476 18236 20496
rect 18236 20476 18288 20496
rect 18288 20476 18290 20496
rect 18234 20440 18290 20476
rect 17130 19488 17186 19544
rect 16394 14048 16450 14104
rect 16486 12588 16488 12608
rect 16488 12588 16540 12608
rect 16540 12588 16542 12608
rect 16486 12552 16542 12588
rect 16486 12416 16542 12472
rect 17038 13504 17094 13560
rect 18326 19896 18382 19952
rect 17682 19236 17738 19272
rect 17682 19216 17684 19236
rect 17684 19216 17736 19236
rect 17736 19216 17738 19236
rect 17866 19216 17922 19272
rect 17774 18164 17776 18184
rect 17776 18164 17828 18184
rect 17828 18164 17830 18184
rect 17774 18128 17830 18164
rect 17498 17312 17554 17368
rect 17406 14356 17408 14376
rect 17408 14356 17460 14376
rect 17460 14356 17462 14376
rect 17406 14320 17462 14356
rect 18050 15308 18052 15328
rect 18052 15308 18104 15328
rect 18104 15308 18106 15328
rect 18050 15272 18106 15308
rect 17866 13640 17922 13696
rect 17590 13368 17646 13424
rect 18694 22380 18696 22400
rect 18696 22380 18748 22400
rect 18748 22380 18750 22400
rect 18694 22344 18750 22380
rect 18878 20168 18934 20224
rect 19154 22772 19210 22808
rect 19154 22752 19156 22772
rect 19156 22752 19208 22772
rect 19208 22752 19210 22772
rect 18418 18672 18474 18728
rect 18602 17312 18658 17368
rect 19154 21140 19210 21176
rect 19154 21120 19156 21140
rect 19156 21120 19208 21140
rect 19208 21120 19210 21140
rect 20442 25744 20498 25800
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 20074 24112 20130 24168
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 20442 23704 20498 23760
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19154 19388 19156 19408
rect 19156 19388 19208 19408
rect 19208 19388 19210 19408
rect 19154 19352 19210 19388
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19614 19252 19616 19272
rect 19616 19252 19668 19272
rect 19668 19252 19670 19272
rect 19614 19216 19670 19252
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 18878 16632 18934 16688
rect 18786 15816 18842 15872
rect 18418 14048 18474 14104
rect 18326 13096 18382 13152
rect 17314 12280 17370 12336
rect 16210 7792 16266 7848
rect 18694 12844 18750 12880
rect 18694 12824 18696 12844
rect 18696 12824 18748 12844
rect 18748 12824 18750 12844
rect 19154 15272 19210 15328
rect 19430 17332 19486 17368
rect 19430 17312 19432 17332
rect 19432 17312 19484 17332
rect 19484 17312 19486 17332
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19338 16496 19394 16552
rect 20166 17584 20222 17640
rect 20074 16496 20130 16552
rect 19982 16360 20038 16416
rect 20166 16360 20222 16416
rect 19154 12960 19210 13016
rect 19338 13504 19394 13560
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 20074 15544 20130 15600
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19522 14320 19578 14376
rect 19706 14340 19762 14376
rect 19706 14320 19708 14340
rect 19708 14320 19760 14340
rect 19760 14320 19762 14340
rect 20074 14184 20130 14240
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 18786 11892 18842 11928
rect 18786 11872 18788 11892
rect 18788 11872 18840 11892
rect 18840 11872 18842 11892
rect 17774 9560 17830 9616
rect 19706 13096 19762 13152
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 21178 24676 21234 24712
rect 21178 24656 21180 24676
rect 21180 24656 21232 24676
rect 21232 24656 21234 24676
rect 20810 24248 20866 24304
rect 20442 21800 20498 21856
rect 20718 20984 20774 21040
rect 20534 19080 20590 19136
rect 21454 22616 21510 22672
rect 21362 22072 21418 22128
rect 21270 19760 21326 19816
rect 20626 17448 20682 17504
rect 20442 13640 20498 13696
rect 20350 12960 20406 13016
rect 20350 12416 20406 12472
rect 21178 18672 21234 18728
rect 20810 14728 20866 14784
rect 21454 15972 21510 16008
rect 21454 15952 21456 15972
rect 21456 15952 21508 15972
rect 21508 15952 21510 15972
rect 21454 15580 21456 15600
rect 21456 15580 21508 15600
rect 21508 15580 21510 15600
rect 21454 15544 21510 15580
rect 21086 13404 21088 13424
rect 21088 13404 21140 13424
rect 21140 13404 21142 13424
rect 21086 13368 21142 13404
rect 20994 12824 21050 12880
rect 21362 13368 21418 13424
rect 20534 12144 20590 12200
rect 21454 11600 21510 11656
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19430 11328 19486 11384
rect 19338 11056 19394 11112
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 21822 23704 21878 23760
rect 21822 19488 21878 19544
rect 21730 19352 21786 19408
rect 21638 18808 21694 18864
rect 21638 16496 21694 16552
rect 22006 23024 22062 23080
rect 22006 22480 22062 22536
rect 22190 20984 22246 21040
rect 22006 18964 22062 19000
rect 22006 18944 22008 18964
rect 22008 18944 22060 18964
rect 22060 18944 22062 18964
rect 22190 16768 22246 16824
rect 21730 15136 21786 15192
rect 22006 15680 22062 15736
rect 21914 15544 21970 15600
rect 21822 13812 21824 13832
rect 21824 13812 21876 13832
rect 21876 13812 21878 13832
rect 21822 13776 21878 13812
rect 21638 12008 21694 12064
rect 23754 24792 23810 24848
rect 22466 22072 22522 22128
rect 22466 19352 22522 19408
rect 22558 19080 22614 19136
rect 22466 16632 22522 16688
rect 21638 11600 21694 11656
rect 21546 9968 21602 10024
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 22558 14320 22614 14376
rect 22742 18128 22798 18184
rect 22742 15952 22798 16008
rect 22926 18944 22982 19000
rect 23294 23704 23350 23760
rect 23570 22208 23626 22264
rect 23478 21664 23534 21720
rect 23478 21292 23480 21312
rect 23480 21292 23532 21312
rect 23532 21292 23534 21312
rect 23478 21256 23534 21292
rect 24674 27104 24730 27160
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24214 24656 24270 24712
rect 24766 26424 24822 26480
rect 24766 24656 24822 24712
rect 23846 21120 23902 21176
rect 23570 20440 23626 20496
rect 23570 20340 23572 20360
rect 23572 20340 23624 20360
rect 23624 20340 23626 20360
rect 23570 20304 23626 20340
rect 23754 20304 23810 20360
rect 23478 18264 23534 18320
rect 23478 17856 23534 17912
rect 23478 15700 23534 15736
rect 23478 15680 23480 15700
rect 23480 15680 23532 15700
rect 23532 15680 23534 15700
rect 23386 15136 23442 15192
rect 23386 15000 23442 15056
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24122 22616 24178 22672
rect 24030 21528 24086 21584
rect 23846 18808 23902 18864
rect 23754 18264 23810 18320
rect 23846 18128 23902 18184
rect 23754 16768 23810 16824
rect 23294 12960 23350 13016
rect 22558 12300 22614 12336
rect 22558 12280 22560 12300
rect 22560 12280 22612 12300
rect 22612 12280 22614 12300
rect 23202 11872 23258 11928
rect 23202 11464 23258 11520
rect 24030 15952 24086 16008
rect 23570 13368 23626 13424
rect 23570 11464 23626 11520
rect 23478 10512 23534 10568
rect 22282 9016 22338 9072
rect 19154 8472 19210 8528
rect 17958 8336 18014 8392
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 17958 7384 18014 7440
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 24030 15408 24086 15464
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24766 23024 24822 23080
rect 24214 20984 24270 21040
rect 24582 20848 24638 20904
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24674 19372 24730 19408
rect 24674 19352 24676 19372
rect 24676 19352 24728 19372
rect 24728 19352 24730 19372
rect 24306 19116 24308 19136
rect 24308 19116 24360 19136
rect 24360 19116 24362 19136
rect 24306 19080 24362 19116
rect 24582 18672 24638 18728
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24766 17312 24822 17368
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24214 16088 24270 16144
rect 25502 25880 25558 25936
rect 25410 23468 25412 23488
rect 25412 23468 25464 23488
rect 25464 23468 25466 23488
rect 25410 23432 25466 23468
rect 25226 19896 25282 19952
rect 25226 19252 25228 19272
rect 25228 19252 25280 19272
rect 25280 19252 25282 19272
rect 25226 19216 25282 19252
rect 25134 18964 25190 19000
rect 25134 18944 25136 18964
rect 25136 18944 25188 18964
rect 25188 18944 25190 18964
rect 25134 18808 25190 18864
rect 24766 16496 24822 16552
rect 24582 15580 24584 15600
rect 24584 15580 24636 15600
rect 24636 15580 24638 15600
rect 24582 15544 24638 15580
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 23754 13368 23810 13424
rect 24122 13776 24178 13832
rect 24030 12960 24086 13016
rect 24122 12824 24178 12880
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24674 13232 24730 13288
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24582 12688 24638 12744
rect 24674 12280 24730 12336
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 23754 11056 23810 11112
rect 23662 8372 23664 8392
rect 23664 8372 23716 8392
rect 23716 8372 23718 8392
rect 23662 8336 23718 8372
rect 23662 7792 23718 7848
rect 23570 6976 23626 7032
rect 23478 6024 23534 6080
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 23478 5072 23534 5128
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 17038 4528 17094 4584
rect 17958 4208 18014 4210
rect 17958 4156 17960 4208
rect 17960 4156 18012 4208
rect 18012 4156 18014 4208
rect 17958 4154 18014 4156
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 15566 3440 15622 3496
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 19522 2896 19578 2952
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 23938 10784 23994 10840
rect 24582 11212 24638 11248
rect 24582 11192 24584 11212
rect 24584 11192 24636 11212
rect 24636 11192 24638 11212
rect 23754 6296 23810 6352
rect 23662 2624 23718 2680
rect 23478 2352 23534 2408
rect 24030 5772 24086 5808
rect 24030 5752 24032 5772
rect 24032 5752 24084 5772
rect 24084 5752 24086 5772
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24582 10648 24638 10704
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24674 8880 24730 8936
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24766 7520 24822 7576
rect 25410 21392 25466 21448
rect 25594 25200 25650 25256
rect 25778 19080 25834 19136
rect 25502 18672 25558 18728
rect 25042 11600 25098 11656
rect 25594 14728 25650 14784
rect 25502 11736 25558 11792
rect 25686 12280 25742 12336
rect 25594 11192 25650 11248
rect 25226 10920 25282 10976
rect 26054 16632 26110 16688
rect 27342 24520 27398 24576
rect 26514 15272 26570 15328
rect 26238 9560 26294 9616
rect 26514 9560 26570 9616
rect 24674 5072 24730 5128
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24582 3884 24584 3904
rect 24584 3884 24636 3904
rect 24636 3884 24638 3904
rect 24582 3848 24638 3884
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 25134 2896 25190 2952
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 23938 1400 23994 1456
rect 20350 856 20406 912
rect 13450 40 13506 96
rect 20350 40 20406 96
<< metal3 >>
rect 0 27706 480 27736
rect 3509 27706 3575 27709
rect 0 27704 3575 27706
rect 0 27648 3514 27704
rect 3570 27648 3575 27704
rect 0 27646 3575 27648
rect 0 27616 480 27646
rect 3509 27643 3575 27646
rect 24117 27706 24183 27709
rect 27520 27706 28000 27736
rect 24117 27704 28000 27706
rect 24117 27648 24122 27704
rect 24178 27648 28000 27704
rect 24117 27646 28000 27648
rect 24117 27643 24183 27646
rect 27520 27616 28000 27646
rect 0 27162 480 27192
rect 4061 27162 4127 27165
rect 0 27160 4127 27162
rect 0 27104 4066 27160
rect 4122 27104 4127 27160
rect 0 27102 4127 27104
rect 0 27072 480 27102
rect 4061 27099 4127 27102
rect 24669 27162 24735 27165
rect 27520 27162 28000 27192
rect 24669 27160 28000 27162
rect 24669 27104 24674 27160
rect 24730 27104 28000 27160
rect 24669 27102 28000 27104
rect 24669 27099 24735 27102
rect 27520 27072 28000 27102
rect 0 26482 480 26512
rect 4061 26482 4127 26485
rect 0 26480 4127 26482
rect 0 26424 4066 26480
rect 4122 26424 4127 26480
rect 0 26422 4127 26424
rect 0 26392 480 26422
rect 4061 26419 4127 26422
rect 24761 26482 24827 26485
rect 27520 26482 28000 26512
rect 24761 26480 28000 26482
rect 24761 26424 24766 26480
rect 24822 26424 28000 26480
rect 24761 26422 28000 26424
rect 24761 26419 24827 26422
rect 27520 26392 28000 26422
rect 9990 26012 9996 26076
rect 10060 26074 10066 26076
rect 10317 26074 10383 26077
rect 10060 26072 10383 26074
rect 10060 26016 10322 26072
rect 10378 26016 10383 26072
rect 10060 26014 10383 26016
rect 10060 26012 10066 26014
rect 10317 26011 10383 26014
rect 0 25938 480 25968
rect 3049 25938 3115 25941
rect 18413 25938 18479 25941
rect 0 25878 1410 25938
rect 0 25848 480 25878
rect 1350 25666 1410 25878
rect 3049 25936 18479 25938
rect 3049 25880 3054 25936
rect 3110 25880 18418 25936
rect 18474 25880 18479 25936
rect 3049 25878 18479 25880
rect 3049 25875 3115 25878
rect 18413 25875 18479 25878
rect 25497 25938 25563 25941
rect 27520 25938 28000 25968
rect 25497 25936 28000 25938
rect 25497 25880 25502 25936
rect 25558 25880 28000 25936
rect 25497 25878 28000 25880
rect 25497 25875 25563 25878
rect 27520 25848 28000 25878
rect 1945 25802 2011 25805
rect 20437 25802 20503 25805
rect 1945 25800 20503 25802
rect 1945 25744 1950 25800
rect 2006 25744 20442 25800
rect 20498 25744 20503 25800
rect 1945 25742 20503 25744
rect 1945 25739 2011 25742
rect 20437 25739 20503 25742
rect 3877 25666 3943 25669
rect 1350 25664 3943 25666
rect 1350 25608 3882 25664
rect 3938 25608 3943 25664
rect 1350 25606 3943 25608
rect 3877 25603 3943 25606
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25258 480 25288
rect 3785 25258 3851 25261
rect 0 25256 3851 25258
rect 0 25200 3790 25256
rect 3846 25200 3851 25256
rect 0 25198 3851 25200
rect 0 25168 480 25198
rect 3785 25195 3851 25198
rect 25589 25258 25655 25261
rect 27520 25258 28000 25288
rect 25589 25256 28000 25258
rect 25589 25200 25594 25256
rect 25650 25200 28000 25256
rect 25589 25198 28000 25200
rect 25589 25195 25655 25198
rect 27520 25168 28000 25198
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 8937 24850 9003 24853
rect 13077 24850 13143 24853
rect 8937 24848 13143 24850
rect 8937 24792 8942 24848
rect 8998 24792 13082 24848
rect 13138 24792 13143 24848
rect 8937 24790 13143 24792
rect 8937 24787 9003 24790
rect 13077 24787 13143 24790
rect 14365 24850 14431 24853
rect 16389 24850 16455 24853
rect 14365 24848 16455 24850
rect 14365 24792 14370 24848
rect 14426 24792 16394 24848
rect 16450 24792 16455 24848
rect 14365 24790 16455 24792
rect 14365 24787 14431 24790
rect 16389 24787 16455 24790
rect 17309 24850 17375 24853
rect 17309 24848 23536 24850
rect 17309 24792 17314 24848
rect 17370 24792 23536 24848
rect 17309 24790 23536 24792
rect 17309 24787 17375 24790
rect 0 24714 480 24744
rect 4245 24714 4311 24717
rect 8845 24716 8911 24717
rect 8845 24714 8892 24716
rect 0 24712 4311 24714
rect 0 24656 4250 24712
rect 4306 24656 4311 24712
rect 0 24654 4311 24656
rect 0 24624 480 24654
rect 4245 24651 4311 24654
rect 7974 24712 8892 24714
rect 7974 24656 8850 24712
rect 7974 24654 8892 24656
rect 2037 24578 2103 24581
rect 7974 24578 8034 24654
rect 8845 24652 8892 24654
rect 8956 24652 8962 24716
rect 12709 24714 12775 24717
rect 18137 24714 18203 24717
rect 12709 24712 18203 24714
rect 12709 24656 12714 24712
rect 12770 24656 18142 24712
rect 18198 24656 18203 24712
rect 12709 24654 18203 24656
rect 8845 24651 8911 24652
rect 12709 24651 12775 24654
rect 18137 24651 18203 24654
rect 21030 24652 21036 24716
rect 21100 24714 21106 24716
rect 21173 24714 21239 24717
rect 21100 24712 21239 24714
rect 21100 24656 21178 24712
rect 21234 24656 21239 24712
rect 21100 24654 21239 24656
rect 21100 24652 21106 24654
rect 21173 24651 21239 24654
rect 2037 24576 8034 24578
rect 2037 24520 2042 24576
rect 2098 24520 8034 24576
rect 2037 24518 8034 24520
rect 10961 24578 11027 24581
rect 15377 24578 15443 24581
rect 10961 24576 15443 24578
rect 10961 24520 10966 24576
rect 11022 24520 15382 24576
rect 15438 24520 15443 24576
rect 10961 24518 15443 24520
rect 23476 24578 23536 24790
rect 23606 24788 23612 24852
rect 23676 24850 23682 24852
rect 23749 24850 23815 24853
rect 23676 24848 23815 24850
rect 23676 24792 23754 24848
rect 23810 24792 23815 24848
rect 23676 24790 23815 24792
rect 23676 24788 23682 24790
rect 23749 24787 23815 24790
rect 23790 24652 23796 24716
rect 23860 24714 23866 24716
rect 24209 24714 24275 24717
rect 23860 24712 24275 24714
rect 23860 24656 24214 24712
rect 24270 24656 24275 24712
rect 23860 24654 24275 24656
rect 23860 24652 23866 24654
rect 24209 24651 24275 24654
rect 24761 24714 24827 24717
rect 27520 24714 28000 24744
rect 24761 24712 28000 24714
rect 24761 24656 24766 24712
rect 24822 24656 28000 24712
rect 24761 24654 28000 24656
rect 24761 24651 24827 24654
rect 27520 24624 28000 24654
rect 27337 24578 27403 24581
rect 23476 24576 27403 24578
rect 23476 24520 27342 24576
rect 27398 24520 27403 24576
rect 23476 24518 27403 24520
rect 2037 24515 2103 24518
rect 10961 24515 11027 24518
rect 15377 24515 15443 24518
rect 27337 24515 27403 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 2037 24442 2103 24445
rect 7005 24442 7071 24445
rect 9673 24442 9739 24445
rect 2037 24440 7071 24442
rect 2037 24384 2042 24440
rect 2098 24384 7010 24440
rect 7066 24384 7071 24440
rect 2037 24382 7071 24384
rect 2037 24379 2103 24382
rect 7005 24379 7071 24382
rect 9446 24440 9739 24442
rect 9446 24384 9678 24440
rect 9734 24384 9739 24440
rect 9446 24382 9739 24384
rect 5257 24306 5323 24309
rect 8569 24306 8635 24309
rect 9446 24306 9506 24382
rect 9673 24379 9739 24382
rect 10777 24442 10843 24445
rect 15561 24442 15627 24445
rect 10777 24440 15627 24442
rect 10777 24384 10782 24440
rect 10838 24384 15566 24440
rect 15622 24384 15627 24440
rect 10777 24382 15627 24384
rect 10777 24379 10843 24382
rect 15561 24379 15627 24382
rect 5257 24304 9506 24306
rect 5257 24248 5262 24304
rect 5318 24248 8574 24304
rect 8630 24248 9506 24304
rect 5257 24246 9506 24248
rect 9581 24306 9647 24309
rect 20805 24306 20871 24309
rect 9581 24304 20871 24306
rect 9581 24248 9586 24304
rect 9642 24248 20810 24304
rect 20866 24248 20871 24304
rect 9581 24246 20871 24248
rect 5257 24243 5323 24246
rect 8569 24243 8635 24246
rect 9581 24243 9647 24246
rect 20805 24243 20871 24246
rect 2313 24170 2379 24173
rect 10777 24170 10843 24173
rect 2313 24168 10843 24170
rect 2313 24112 2318 24168
rect 2374 24112 10782 24168
rect 10838 24112 10843 24168
rect 2313 24110 10843 24112
rect 2313 24107 2379 24110
rect 10777 24107 10843 24110
rect 11145 24170 11211 24173
rect 13537 24170 13603 24173
rect 11145 24168 13603 24170
rect 11145 24112 11150 24168
rect 11206 24112 13542 24168
rect 13598 24112 13603 24168
rect 11145 24110 13603 24112
rect 11145 24107 11211 24110
rect 13537 24107 13603 24110
rect 14089 24170 14155 24173
rect 20069 24170 20135 24173
rect 14089 24168 20135 24170
rect 14089 24112 14094 24168
rect 14150 24112 20074 24168
rect 20130 24112 20135 24168
rect 14089 24110 20135 24112
rect 14089 24107 14155 24110
rect 20069 24107 20135 24110
rect 0 24034 480 24064
rect 2865 24034 2931 24037
rect 0 24032 2931 24034
rect 0 23976 2870 24032
rect 2926 23976 2931 24032
rect 0 23974 2931 23976
rect 0 23944 480 23974
rect 2865 23971 2931 23974
rect 6637 24034 6703 24037
rect 10961 24034 11027 24037
rect 27520 24034 28000 24064
rect 6637 24032 11027 24034
rect 6637 23976 6642 24032
rect 6698 23976 10966 24032
rect 11022 23976 11027 24032
rect 6637 23974 11027 23976
rect 6637 23971 6703 23974
rect 10961 23971 11027 23974
rect 24718 23974 28000 24034
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 7281 23898 7347 23901
rect 13169 23898 13235 23901
rect 7281 23896 13235 23898
rect 7281 23840 7286 23896
rect 7342 23840 13174 23896
rect 13230 23840 13235 23896
rect 7281 23838 13235 23840
rect 7281 23835 7347 23838
rect 13169 23835 13235 23838
rect 1485 23762 1551 23765
rect 20437 23762 20503 23765
rect 21817 23762 21883 23765
rect 1485 23760 21883 23762
rect 1485 23704 1490 23760
rect 1546 23704 20442 23760
rect 20498 23704 21822 23760
rect 21878 23704 21883 23760
rect 1485 23702 21883 23704
rect 1485 23699 1551 23702
rect 20437 23699 20503 23702
rect 21817 23699 21883 23702
rect 23289 23762 23355 23765
rect 24718 23762 24778 23974
rect 27520 23944 28000 23974
rect 23289 23760 24778 23762
rect 23289 23704 23294 23760
rect 23350 23704 24778 23760
rect 23289 23702 24778 23704
rect 23289 23699 23355 23702
rect 4889 23626 4955 23629
rect 10961 23626 11027 23629
rect 16113 23626 16179 23629
rect 16481 23626 16547 23629
rect 4889 23624 10794 23626
rect 4889 23568 4894 23624
rect 4950 23568 10794 23624
rect 4889 23566 10794 23568
rect 4889 23563 4955 23566
rect 0 23490 480 23520
rect 2681 23490 2747 23493
rect 0 23488 2747 23490
rect 0 23432 2686 23488
rect 2742 23432 2747 23488
rect 0 23430 2747 23432
rect 0 23400 480 23430
rect 2681 23427 2747 23430
rect 3601 23490 3667 23493
rect 6177 23490 6243 23493
rect 3601 23488 6243 23490
rect 3601 23432 3606 23488
rect 3662 23432 6182 23488
rect 6238 23432 6243 23488
rect 3601 23430 6243 23432
rect 3601 23427 3667 23430
rect 6177 23427 6243 23430
rect 7373 23490 7439 23493
rect 9438 23490 9444 23492
rect 7373 23488 9444 23490
rect 7373 23432 7378 23488
rect 7434 23432 9444 23488
rect 7373 23430 9444 23432
rect 7373 23427 7439 23430
rect 9438 23428 9444 23430
rect 9508 23428 9514 23492
rect 10734 23490 10794 23566
rect 10961 23624 16547 23626
rect 10961 23568 10966 23624
rect 11022 23568 16118 23624
rect 16174 23568 16486 23624
rect 16542 23568 16547 23624
rect 10961 23566 16547 23568
rect 10961 23563 11027 23566
rect 16113 23563 16179 23566
rect 16481 23563 16547 23566
rect 13077 23490 13143 23493
rect 14273 23490 14339 23493
rect 10734 23488 14339 23490
rect 10734 23432 13082 23488
rect 13138 23432 14278 23488
rect 14334 23432 14339 23488
rect 10734 23430 14339 23432
rect 13077 23427 13143 23430
rect 14273 23427 14339 23430
rect 25405 23490 25471 23493
rect 27520 23490 28000 23520
rect 25405 23488 28000 23490
rect 25405 23432 25410 23488
rect 25466 23432 28000 23488
rect 25405 23430 28000 23432
rect 25405 23427 25471 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 27520 23400 28000 23430
rect 19610 23359 19930 23360
rect 6085 23354 6151 23357
rect 8017 23354 8083 23357
rect 6085 23352 8083 23354
rect 6085 23296 6090 23352
rect 6146 23296 8022 23352
rect 8078 23296 8083 23352
rect 6085 23294 8083 23296
rect 6085 23291 6151 23294
rect 8017 23291 8083 23294
rect 11789 23354 11855 23357
rect 13905 23354 13971 23357
rect 11789 23352 13971 23354
rect 11789 23296 11794 23352
rect 11850 23296 13910 23352
rect 13966 23296 13971 23352
rect 11789 23294 13971 23296
rect 11789 23291 11855 23294
rect 13905 23291 13971 23294
rect 14038 23292 14044 23356
rect 14108 23354 14114 23356
rect 18597 23354 18663 23357
rect 14108 23352 18663 23354
rect 14108 23296 18602 23352
rect 18658 23296 18663 23352
rect 14108 23294 18663 23296
rect 14108 23292 14114 23294
rect 18597 23291 18663 23294
rect 9029 23082 9095 23085
rect 16849 23082 16915 23085
rect 9029 23080 16915 23082
rect 9029 23024 9034 23080
rect 9090 23024 16854 23080
rect 16910 23024 16915 23080
rect 9029 23022 16915 23024
rect 9029 23019 9095 23022
rect 16849 23019 16915 23022
rect 22001 23082 22067 23085
rect 24761 23082 24827 23085
rect 22001 23080 24827 23082
rect 22001 23024 22006 23080
rect 22062 23024 24766 23080
rect 24822 23024 24827 23080
rect 22001 23022 24827 23024
rect 22001 23019 22067 23022
rect 24761 23019 24827 23022
rect 8017 22946 8083 22949
rect 14733 22946 14799 22949
rect 8017 22944 14799 22946
rect 8017 22888 8022 22944
rect 8078 22888 14738 22944
rect 14794 22888 14799 22944
rect 8017 22886 14799 22888
rect 8017 22883 8083 22886
rect 14733 22883 14799 22886
rect 5610 22880 5930 22881
rect 0 22810 480 22840
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 2957 22810 3023 22813
rect 0 22808 3023 22810
rect 0 22752 2962 22808
rect 3018 22752 3023 22808
rect 0 22750 3023 22752
rect 0 22720 480 22750
rect 2957 22747 3023 22750
rect 4521 22810 4587 22813
rect 5022 22810 5028 22812
rect 4521 22808 5028 22810
rect 4521 22752 4526 22808
rect 4582 22752 5028 22808
rect 4521 22750 5028 22752
rect 4521 22747 4587 22750
rect 5022 22748 5028 22750
rect 5092 22748 5098 22812
rect 7925 22810 7991 22813
rect 9765 22810 9831 22813
rect 14273 22810 14339 22813
rect 18505 22810 18571 22813
rect 7925 22808 14339 22810
rect 7925 22752 7930 22808
rect 7986 22752 9770 22808
rect 9826 22752 14278 22808
rect 14334 22752 14339 22808
rect 7925 22750 14339 22752
rect 7925 22747 7991 22750
rect 9765 22747 9831 22750
rect 14273 22747 14339 22750
rect 15518 22808 18571 22810
rect 15518 22752 18510 22808
rect 18566 22752 18571 22808
rect 15518 22750 18571 22752
rect 841 22674 907 22677
rect 6269 22674 6335 22677
rect 9949 22676 10015 22677
rect 9949 22674 9996 22676
rect 841 22672 6335 22674
rect 841 22616 846 22672
rect 902 22616 6274 22672
rect 6330 22616 6335 22672
rect 841 22614 6335 22616
rect 9904 22672 9996 22674
rect 9904 22616 9954 22672
rect 9904 22614 9996 22616
rect 841 22611 907 22614
rect 6269 22611 6335 22614
rect 9949 22612 9996 22614
rect 10060 22612 10066 22676
rect 11421 22674 11487 22677
rect 15518 22674 15578 22750
rect 18505 22747 18571 22750
rect 19006 22748 19012 22812
rect 19076 22810 19082 22812
rect 19149 22810 19215 22813
rect 27520 22810 28000 22840
rect 19076 22808 19215 22810
rect 19076 22752 19154 22808
rect 19210 22752 19215 22808
rect 19076 22750 19215 22752
rect 19076 22748 19082 22750
rect 19149 22747 19215 22750
rect 24718 22750 28000 22810
rect 21449 22674 21515 22677
rect 11421 22672 15578 22674
rect 11421 22616 11426 22672
rect 11482 22616 15578 22672
rect 11421 22614 15578 22616
rect 17910 22672 21515 22674
rect 17910 22616 21454 22672
rect 21510 22616 21515 22672
rect 17910 22614 21515 22616
rect 9949 22611 10015 22612
rect 11421 22611 11487 22614
rect 5257 22538 5323 22541
rect 17910 22538 17970 22614
rect 21449 22611 21515 22614
rect 24117 22674 24183 22677
rect 24718 22674 24778 22750
rect 27520 22720 28000 22750
rect 24117 22672 24778 22674
rect 24117 22616 24122 22672
rect 24178 22616 24778 22672
rect 24117 22614 24778 22616
rect 24117 22611 24183 22614
rect 5257 22536 17970 22538
rect 5257 22480 5262 22536
rect 5318 22480 17970 22536
rect 5257 22478 17970 22480
rect 18045 22538 18111 22541
rect 22001 22538 22067 22541
rect 18045 22536 22067 22538
rect 18045 22480 18050 22536
rect 18106 22480 22006 22536
rect 22062 22480 22067 22536
rect 18045 22478 22067 22480
rect 5257 22475 5323 22478
rect 18045 22475 18111 22478
rect 22001 22475 22067 22478
rect 7414 22340 7420 22404
rect 7484 22402 7490 22404
rect 8109 22402 8175 22405
rect 7484 22400 8175 22402
rect 7484 22344 8114 22400
rect 8170 22344 8175 22400
rect 7484 22342 8175 22344
rect 7484 22340 7490 22342
rect 8109 22339 8175 22342
rect 16757 22402 16823 22405
rect 18689 22402 18755 22405
rect 16757 22400 18755 22402
rect 16757 22344 16762 22400
rect 16818 22344 18694 22400
rect 18750 22344 18755 22400
rect 16757 22342 18755 22344
rect 16757 22339 16823 22342
rect 18689 22339 18755 22342
rect 10277 22336 10597 22337
rect 0 22266 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 1761 22266 1827 22269
rect 0 22264 1827 22266
rect 0 22208 1766 22264
rect 1822 22208 1827 22264
rect 0 22206 1827 22208
rect 0 22176 480 22206
rect 1761 22203 1827 22206
rect 2957 22266 3023 22269
rect 9949 22266 10015 22269
rect 2957 22264 10015 22266
rect 2957 22208 2962 22264
rect 3018 22208 9954 22264
rect 10010 22208 10015 22264
rect 2957 22206 10015 22208
rect 2957 22203 3023 22206
rect 9949 22203 10015 22206
rect 14917 22266 14983 22269
rect 18505 22266 18571 22269
rect 14917 22264 18571 22266
rect 14917 22208 14922 22264
rect 14978 22208 18510 22264
rect 18566 22208 18571 22264
rect 14917 22206 18571 22208
rect 14917 22203 14983 22206
rect 18505 22203 18571 22206
rect 23565 22266 23631 22269
rect 27520 22266 28000 22296
rect 23565 22264 28000 22266
rect 23565 22208 23570 22264
rect 23626 22208 28000 22264
rect 23565 22206 28000 22208
rect 23565 22203 23631 22206
rect 27520 22176 28000 22206
rect 1853 22130 1919 22133
rect 2865 22130 2931 22133
rect 6361 22130 6427 22133
rect 9121 22130 9187 22133
rect 1853 22128 9187 22130
rect 1853 22072 1858 22128
rect 1914 22072 2870 22128
rect 2926 22072 6366 22128
rect 6422 22072 9126 22128
rect 9182 22072 9187 22128
rect 1853 22070 9187 22072
rect 1853 22067 1919 22070
rect 2865 22067 2931 22070
rect 6361 22067 6427 22070
rect 9121 22067 9187 22070
rect 9857 22130 9923 22133
rect 17769 22130 17835 22133
rect 9857 22128 17835 22130
rect 9857 22072 9862 22128
rect 9918 22072 17774 22128
rect 17830 22072 17835 22128
rect 9857 22070 17835 22072
rect 9857 22067 9923 22070
rect 17769 22067 17835 22070
rect 21357 22130 21423 22133
rect 22461 22130 22527 22133
rect 21357 22128 22527 22130
rect 21357 22072 21362 22128
rect 21418 22072 22466 22128
rect 22522 22072 22527 22128
rect 21357 22070 22527 22072
rect 21357 22067 21423 22070
rect 22461 22067 22527 22070
rect 9397 21994 9463 21997
rect 11237 21994 11303 21997
rect 11421 21994 11487 21997
rect 14038 21994 14044 21996
rect 9397 21992 11346 21994
rect 9397 21936 9402 21992
rect 9458 21936 11242 21992
rect 11298 21936 11346 21992
rect 9397 21934 11346 21936
rect 9397 21931 9463 21934
rect 11237 21931 11346 21934
rect 11421 21992 14044 21994
rect 11421 21936 11426 21992
rect 11482 21936 14044 21992
rect 11421 21934 14044 21936
rect 11421 21931 11487 21934
rect 14038 21932 14044 21934
rect 14108 21932 14114 21996
rect 18321 21994 18387 21997
rect 14782 21992 18387 21994
rect 14782 21936 18326 21992
rect 18382 21936 18387 21992
rect 14782 21934 18387 21936
rect 11286 21858 11346 21931
rect 14782 21858 14842 21934
rect 18321 21931 18387 21934
rect 11286 21798 14842 21858
rect 16941 21858 17007 21861
rect 20437 21858 20503 21861
rect 16941 21856 20503 21858
rect 16941 21800 16946 21856
rect 17002 21800 20442 21856
rect 20498 21800 20503 21856
rect 16941 21798 20503 21800
rect 16941 21795 17007 21798
rect 20437 21795 20503 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 23473 21722 23539 21725
rect 17174 21720 23539 21722
rect 17174 21664 23478 21720
rect 23534 21664 23539 21720
rect 17174 21662 23539 21664
rect 0 21586 480 21616
rect 1577 21586 1643 21589
rect 0 21584 1643 21586
rect 0 21528 1582 21584
rect 1638 21528 1643 21584
rect 0 21526 1643 21528
rect 0 21496 480 21526
rect 1577 21523 1643 21526
rect 4889 21586 4955 21589
rect 11697 21586 11763 21589
rect 4889 21584 11763 21586
rect 4889 21528 4894 21584
rect 4950 21528 11702 21584
rect 11758 21528 11763 21584
rect 4889 21526 11763 21528
rect 4889 21523 4955 21526
rect 11697 21523 11763 21526
rect 13721 21586 13787 21589
rect 15377 21586 15443 21589
rect 16665 21586 16731 21589
rect 13721 21584 16731 21586
rect 13721 21528 13726 21584
rect 13782 21528 15382 21584
rect 15438 21528 16670 21584
rect 16726 21528 16731 21584
rect 13721 21526 16731 21528
rect 13721 21523 13787 21526
rect 15377 21523 15443 21526
rect 16665 21523 16731 21526
rect 8109 21450 8175 21453
rect 17174 21450 17234 21662
rect 23473 21659 23539 21662
rect 24025 21586 24091 21589
rect 27520 21586 28000 21616
rect 24025 21584 28000 21586
rect 24025 21528 24030 21584
rect 24086 21528 28000 21584
rect 24025 21526 28000 21528
rect 24025 21523 24091 21526
rect 27520 21496 28000 21526
rect 25405 21450 25471 21453
rect 8109 21448 17234 21450
rect 8109 21392 8114 21448
rect 8170 21392 17234 21448
rect 8109 21390 17234 21392
rect 17358 21448 25471 21450
rect 17358 21392 25410 21448
rect 25466 21392 25471 21448
rect 17358 21390 25471 21392
rect 8109 21387 8175 21390
rect 7005 21314 7071 21317
rect 10041 21314 10107 21317
rect 7005 21312 10107 21314
rect 7005 21256 7010 21312
rect 7066 21256 10046 21312
rect 10102 21256 10107 21312
rect 7005 21254 10107 21256
rect 7005 21251 7071 21254
rect 10041 21251 10107 21254
rect 11973 21314 12039 21317
rect 17358 21314 17418 21390
rect 25405 21387 25471 21390
rect 23473 21316 23539 21317
rect 11973 21312 17418 21314
rect 11973 21256 11978 21312
rect 12034 21256 17418 21312
rect 11973 21254 17418 21256
rect 11973 21251 12039 21254
rect 23422 21252 23428 21316
rect 23492 21314 23539 21316
rect 23492 21312 23584 21314
rect 23534 21256 23584 21312
rect 23492 21254 23584 21256
rect 23492 21252 23539 21254
rect 23473 21251 23539 21252
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 2405 21178 2471 21181
rect 4521 21178 4587 21181
rect 2405 21176 4587 21178
rect 2405 21120 2410 21176
rect 2466 21120 4526 21176
rect 4582 21120 4587 21176
rect 2405 21118 4587 21120
rect 2405 21115 2471 21118
rect 4521 21115 4587 21118
rect 6453 21178 6519 21181
rect 9673 21178 9739 21181
rect 6453 21176 9739 21178
rect 6453 21120 6458 21176
rect 6514 21120 9678 21176
rect 9734 21120 9739 21176
rect 6453 21118 9739 21120
rect 6453 21115 6519 21118
rect 9673 21115 9739 21118
rect 16389 21178 16455 21181
rect 17677 21178 17743 21181
rect 19149 21178 19215 21181
rect 16389 21176 19215 21178
rect 16389 21120 16394 21176
rect 16450 21120 17682 21176
rect 17738 21120 19154 21176
rect 19210 21120 19215 21176
rect 16389 21118 19215 21120
rect 16389 21115 16455 21118
rect 17677 21115 17743 21118
rect 19149 21115 19215 21118
rect 23841 21176 23907 21181
rect 23841 21120 23846 21176
rect 23902 21120 23907 21176
rect 23841 21115 23907 21120
rect 0 21042 480 21072
rect 3049 21042 3115 21045
rect 0 21040 3115 21042
rect 0 20984 3054 21040
rect 3110 20984 3115 21040
rect 0 20982 3115 20984
rect 0 20952 480 20982
rect 3049 20979 3115 20982
rect 11881 21042 11947 21045
rect 20713 21042 20779 21045
rect 11881 21040 20779 21042
rect 11881 20984 11886 21040
rect 11942 20984 20718 21040
rect 20774 20984 20779 21040
rect 11881 20982 20779 20984
rect 11881 20979 11947 20982
rect 20713 20979 20779 20982
rect 22185 21042 22251 21045
rect 23844 21042 23904 21115
rect 22185 21040 23904 21042
rect 22185 20984 22190 21040
rect 22246 20984 23904 21040
rect 22185 20982 23904 20984
rect 24209 21042 24275 21045
rect 27520 21042 28000 21072
rect 24209 21040 28000 21042
rect 24209 20984 24214 21040
rect 24270 20984 28000 21040
rect 24209 20982 28000 20984
rect 22185 20979 22251 20982
rect 24209 20979 24275 20982
rect 27520 20952 28000 20982
rect 14733 20906 14799 20909
rect 16113 20906 16179 20909
rect 18137 20906 18203 20909
rect 24577 20906 24643 20909
rect 14733 20904 18203 20906
rect 14733 20848 14738 20904
rect 14794 20848 16118 20904
rect 16174 20848 18142 20904
rect 18198 20848 18203 20904
rect 14733 20846 18203 20848
rect 14733 20843 14799 20846
rect 16113 20843 16179 20846
rect 18137 20843 18203 20846
rect 24120 20904 24643 20906
rect 24120 20848 24582 20904
rect 24638 20848 24643 20904
rect 24120 20846 24643 20848
rect 15377 20770 15443 20773
rect 17493 20770 17559 20773
rect 15377 20768 17559 20770
rect 15377 20712 15382 20768
rect 15438 20712 17498 20768
rect 17554 20712 17559 20768
rect 15377 20710 17559 20712
rect 15377 20707 15443 20710
rect 17493 20707 17559 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 10869 20634 10935 20637
rect 12433 20634 12499 20637
rect 24120 20634 24180 20846
rect 24577 20843 24643 20846
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 10869 20632 12499 20634
rect 10869 20576 10874 20632
rect 10930 20576 12438 20632
rect 12494 20576 12499 20632
rect 10869 20574 12499 20576
rect 10869 20571 10935 20574
rect 12433 20571 12499 20574
rect 15334 20574 24180 20634
rect 3969 20498 4035 20501
rect 5165 20498 5231 20501
rect 6729 20498 6795 20501
rect 3969 20496 6795 20498
rect 3969 20440 3974 20496
rect 4030 20440 5170 20496
rect 5226 20440 6734 20496
rect 6790 20440 6795 20496
rect 3969 20438 6795 20440
rect 3969 20435 4035 20438
rect 5165 20435 5231 20438
rect 6729 20435 6795 20438
rect 10961 20498 11027 20501
rect 12709 20498 12775 20501
rect 10961 20496 12775 20498
rect 10961 20440 10966 20496
rect 11022 20440 12714 20496
rect 12770 20440 12775 20496
rect 10961 20438 12775 20440
rect 10961 20435 11027 20438
rect 12709 20435 12775 20438
rect 12985 20498 13051 20501
rect 15334 20498 15394 20574
rect 12985 20496 15394 20498
rect 12985 20440 12990 20496
rect 13046 20440 15394 20496
rect 12985 20438 15394 20440
rect 18229 20498 18295 20501
rect 23565 20498 23631 20501
rect 18229 20496 23631 20498
rect 18229 20440 18234 20496
rect 18290 20440 23570 20496
rect 23626 20440 23631 20496
rect 18229 20438 23631 20440
rect 12985 20435 13051 20438
rect 18229 20435 18295 20438
rect 23565 20435 23631 20438
rect 0 20362 480 20392
rect 1393 20362 1459 20365
rect 0 20360 1459 20362
rect 0 20304 1398 20360
rect 1454 20304 1459 20360
rect 0 20302 1459 20304
rect 0 20272 480 20302
rect 1393 20299 1459 20302
rect 6821 20362 6887 20365
rect 13261 20362 13327 20365
rect 23565 20362 23631 20365
rect 6821 20360 13186 20362
rect 6821 20304 6826 20360
rect 6882 20304 13186 20360
rect 6821 20302 13186 20304
rect 6821 20299 6887 20302
rect 13126 20226 13186 20302
rect 13261 20360 23631 20362
rect 13261 20304 13266 20360
rect 13322 20304 23570 20360
rect 23626 20304 23631 20360
rect 13261 20302 23631 20304
rect 13261 20299 13327 20302
rect 23565 20299 23631 20302
rect 23749 20362 23815 20365
rect 27520 20362 28000 20392
rect 23749 20360 28000 20362
rect 23749 20304 23754 20360
rect 23810 20304 28000 20360
rect 23749 20302 28000 20304
rect 23749 20299 23815 20302
rect 27520 20272 28000 20302
rect 18873 20226 18939 20229
rect 13126 20224 18939 20226
rect 13126 20168 18878 20224
rect 18934 20168 18939 20224
rect 13126 20166 18939 20168
rect 18873 20163 18939 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 1669 20090 1735 20093
rect 7649 20090 7715 20093
rect 1669 20088 7715 20090
rect 1669 20032 1674 20088
rect 1730 20032 7654 20088
rect 7710 20032 7715 20088
rect 1669 20030 7715 20032
rect 1669 20027 1735 20030
rect 7649 20027 7715 20030
rect 18321 19954 18387 19957
rect 25221 19954 25287 19957
rect 18321 19952 25287 19954
rect 18321 19896 18326 19952
rect 18382 19896 25226 19952
rect 25282 19896 25287 19952
rect 18321 19894 25287 19896
rect 18321 19891 18387 19894
rect 25221 19891 25287 19894
rect 0 19818 480 19848
rect 3969 19818 4035 19821
rect 0 19816 4035 19818
rect 0 19760 3974 19816
rect 4030 19760 4035 19816
rect 0 19758 4035 19760
rect 0 19728 480 19758
rect 3969 19755 4035 19758
rect 9489 19818 9555 19821
rect 12341 19818 12407 19821
rect 9489 19816 12407 19818
rect 9489 19760 9494 19816
rect 9550 19760 12346 19816
rect 12402 19760 12407 19816
rect 9489 19758 12407 19760
rect 9489 19755 9555 19758
rect 12341 19755 12407 19758
rect 21265 19818 21331 19821
rect 27520 19818 28000 19848
rect 21265 19816 28000 19818
rect 21265 19760 21270 19816
rect 21326 19760 28000 19816
rect 21265 19758 28000 19760
rect 21265 19755 21331 19758
rect 27520 19728 28000 19758
rect 9213 19682 9279 19685
rect 14089 19682 14155 19685
rect 9213 19680 14155 19682
rect 9213 19624 9218 19680
rect 9274 19624 14094 19680
rect 14150 19624 14155 19680
rect 9213 19622 14155 19624
rect 9213 19619 9279 19622
rect 14089 19619 14155 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 9622 19484 9628 19548
rect 9692 19546 9698 19548
rect 16665 19546 16731 19549
rect 17125 19546 17191 19549
rect 21817 19546 21883 19549
rect 9692 19486 12266 19546
rect 9692 19484 9698 19486
rect 7373 19412 7439 19413
rect 7373 19410 7420 19412
rect 7328 19408 7420 19410
rect 7328 19352 7378 19408
rect 7328 19350 7420 19352
rect 7373 19348 7420 19350
rect 7484 19348 7490 19412
rect 7557 19410 7623 19413
rect 12065 19410 12131 19413
rect 7557 19408 12131 19410
rect 7557 19352 7562 19408
rect 7618 19352 12070 19408
rect 12126 19352 12131 19408
rect 7557 19350 12131 19352
rect 12206 19410 12266 19486
rect 16665 19544 21883 19546
rect 16665 19488 16670 19544
rect 16726 19488 17130 19544
rect 17186 19488 21822 19544
rect 21878 19488 21883 19544
rect 16665 19486 21883 19488
rect 16665 19483 16731 19486
rect 17125 19483 17191 19486
rect 21817 19483 21883 19486
rect 16389 19410 16455 19413
rect 12206 19408 16455 19410
rect 12206 19352 16394 19408
rect 16450 19352 16455 19408
rect 12206 19350 16455 19352
rect 7373 19347 7439 19348
rect 7557 19347 7623 19350
rect 12065 19347 12131 19350
rect 16389 19347 16455 19350
rect 19149 19410 19215 19413
rect 21725 19410 21791 19413
rect 22461 19410 22527 19413
rect 24669 19410 24735 19413
rect 19149 19408 24735 19410
rect 19149 19352 19154 19408
rect 19210 19352 21730 19408
rect 21786 19352 22466 19408
rect 22522 19352 24674 19408
rect 24730 19352 24735 19408
rect 19149 19350 24735 19352
rect 19149 19347 19215 19350
rect 21725 19347 21791 19350
rect 22461 19347 22527 19350
rect 24669 19347 24735 19350
rect 2589 19274 2655 19277
rect 5993 19274 6059 19277
rect 2589 19272 6059 19274
rect 2589 19216 2594 19272
rect 2650 19216 5998 19272
rect 6054 19216 6059 19272
rect 2589 19214 6059 19216
rect 2589 19211 2655 19214
rect 5993 19211 6059 19214
rect 6269 19274 6335 19277
rect 17677 19274 17743 19277
rect 6269 19272 17743 19274
rect 6269 19216 6274 19272
rect 6330 19216 17682 19272
rect 17738 19216 17743 19272
rect 6269 19214 17743 19216
rect 6269 19211 6335 19214
rect 17677 19211 17743 19214
rect 17861 19274 17927 19277
rect 19609 19274 19675 19277
rect 17861 19272 19675 19274
rect 17861 19216 17866 19272
rect 17922 19216 19614 19272
rect 19670 19216 19675 19272
rect 17861 19214 19675 19216
rect 17861 19211 17927 19214
rect 19609 19211 19675 19214
rect 24894 19212 24900 19276
rect 24964 19274 24970 19276
rect 25221 19274 25287 19277
rect 24964 19272 25287 19274
rect 24964 19216 25226 19272
rect 25282 19216 25287 19272
rect 24964 19214 25287 19216
rect 24964 19212 24970 19214
rect 25221 19211 25287 19214
rect 0 19138 480 19168
rect 3693 19138 3759 19141
rect 0 19136 3759 19138
rect 0 19080 3698 19136
rect 3754 19080 3759 19136
rect 0 19078 3759 19080
rect 0 19048 480 19078
rect 3693 19075 3759 19078
rect 4797 19138 4863 19141
rect 9673 19138 9739 19141
rect 4797 19136 9739 19138
rect 4797 19080 4802 19136
rect 4858 19080 9678 19136
rect 9734 19080 9739 19136
rect 4797 19078 9739 19080
rect 4797 19075 4863 19078
rect 9673 19075 9739 19078
rect 13169 19138 13235 19141
rect 15745 19138 15811 19141
rect 13169 19136 15811 19138
rect 13169 19080 13174 19136
rect 13230 19080 15750 19136
rect 15806 19080 15811 19136
rect 13169 19078 15811 19080
rect 13169 19075 13235 19078
rect 15745 19075 15811 19078
rect 20529 19138 20595 19141
rect 22553 19138 22619 19141
rect 20529 19136 22619 19138
rect 20529 19080 20534 19136
rect 20590 19080 22558 19136
rect 22614 19080 22619 19136
rect 20529 19078 22619 19080
rect 20529 19075 20595 19078
rect 22553 19075 22619 19078
rect 23974 19076 23980 19140
rect 24044 19138 24050 19140
rect 24301 19138 24367 19141
rect 24044 19136 24367 19138
rect 24044 19080 24306 19136
rect 24362 19080 24367 19136
rect 24044 19078 24367 19080
rect 24044 19076 24050 19078
rect 24301 19075 24367 19078
rect 25773 19138 25839 19141
rect 27520 19138 28000 19168
rect 25773 19136 28000 19138
rect 25773 19080 25778 19136
rect 25834 19080 28000 19136
rect 25773 19078 28000 19080
rect 25773 19075 25839 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19078
rect 19610 19007 19930 19008
rect 2497 19002 2563 19005
rect 5257 19002 5323 19005
rect 2497 19000 5323 19002
rect 2497 18944 2502 19000
rect 2558 18944 5262 19000
rect 5318 18944 5323 19000
rect 2497 18942 5323 18944
rect 2497 18939 2563 18942
rect 5257 18939 5323 18942
rect 8477 19002 8543 19005
rect 22001 19002 22067 19005
rect 22921 19002 22987 19005
rect 25129 19002 25195 19005
rect 8477 19000 9552 19002
rect 8477 18944 8482 19000
rect 8538 18968 9552 19000
rect 22001 19000 25195 19002
rect 8538 18944 9644 18968
rect 8477 18942 9644 18944
rect 8477 18939 8543 18942
rect 9492 18908 9644 18942
rect 22001 18944 22006 19000
rect 22062 18944 22926 19000
rect 22982 18944 25134 19000
rect 25190 18944 25195 19000
rect 22001 18942 25195 18944
rect 22001 18939 22067 18942
rect 22921 18939 22987 18942
rect 25129 18939 25195 18942
rect 9584 18866 9644 18908
rect 14089 18866 14155 18869
rect 9584 18864 14155 18866
rect 9584 18808 14094 18864
rect 14150 18808 14155 18864
rect 9584 18806 14155 18808
rect 14089 18803 14155 18806
rect 16849 18866 16915 18869
rect 21633 18866 21699 18869
rect 16849 18864 21699 18866
rect 16849 18808 16854 18864
rect 16910 18808 21638 18864
rect 21694 18808 21699 18864
rect 16849 18806 21699 18808
rect 16849 18803 16915 18806
rect 21633 18803 21699 18806
rect 23841 18866 23907 18869
rect 25129 18866 25195 18869
rect 23841 18864 25195 18866
rect 23841 18808 23846 18864
rect 23902 18808 25134 18864
rect 25190 18808 25195 18864
rect 23841 18806 25195 18808
rect 23841 18803 23907 18806
rect 25129 18803 25195 18806
rect 8017 18730 8083 18733
rect 8385 18730 8451 18733
rect 8017 18728 8451 18730
rect 8017 18672 8022 18728
rect 8078 18672 8390 18728
rect 8446 18672 8451 18728
rect 8017 18670 8451 18672
rect 8017 18667 8083 18670
rect 8385 18667 8451 18670
rect 18413 18730 18479 18733
rect 21173 18730 21239 18733
rect 24577 18730 24643 18733
rect 25497 18730 25563 18733
rect 18413 18728 21239 18730
rect 18413 18672 18418 18728
rect 18474 18672 21178 18728
rect 21234 18672 21239 18728
rect 18413 18670 21239 18672
rect 18413 18667 18479 18670
rect 21173 18667 21239 18670
rect 24120 18728 25563 18730
rect 24120 18672 24582 18728
rect 24638 18672 25502 18728
rect 25558 18672 25563 18728
rect 24120 18670 25563 18672
rect 0 18594 480 18624
rect 3785 18594 3851 18597
rect 0 18592 3851 18594
rect 0 18536 3790 18592
rect 3846 18536 3851 18592
rect 0 18534 3851 18536
rect 0 18504 480 18534
rect 3785 18531 3851 18534
rect 15561 18594 15627 18597
rect 24120 18594 24180 18670
rect 24577 18667 24643 18670
rect 25497 18667 25563 18670
rect 27520 18594 28000 18624
rect 15561 18592 24180 18594
rect 15561 18536 15566 18592
rect 15622 18536 24180 18592
rect 15561 18534 24180 18536
rect 24672 18534 28000 18594
rect 15561 18531 15627 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 9489 18458 9555 18461
rect 11053 18458 11119 18461
rect 11421 18458 11487 18461
rect 9489 18456 11487 18458
rect 9489 18400 9494 18456
rect 9550 18400 11058 18456
rect 11114 18400 11426 18456
rect 11482 18400 11487 18456
rect 9489 18398 11487 18400
rect 9489 18395 9555 18398
rect 11053 18395 11119 18398
rect 11421 18395 11487 18398
rect 9397 18322 9463 18325
rect 10685 18322 10751 18325
rect 9397 18320 10751 18322
rect 9397 18264 9402 18320
rect 9458 18264 10690 18320
rect 10746 18264 10751 18320
rect 9397 18262 10751 18264
rect 9397 18259 9463 18262
rect 10685 18259 10751 18262
rect 11237 18322 11303 18325
rect 16389 18322 16455 18325
rect 23473 18322 23539 18325
rect 11237 18320 11530 18322
rect 11237 18264 11242 18320
rect 11298 18264 11530 18320
rect 11237 18262 11530 18264
rect 11237 18259 11303 18262
rect 8109 18186 8175 18189
rect 11237 18186 11303 18189
rect 8109 18184 11303 18186
rect 8109 18128 8114 18184
rect 8170 18128 11242 18184
rect 11298 18128 11303 18184
rect 8109 18126 11303 18128
rect 11470 18186 11530 18262
rect 16389 18320 23539 18322
rect 16389 18264 16394 18320
rect 16450 18264 23478 18320
rect 23534 18264 23539 18320
rect 16389 18262 23539 18264
rect 16389 18259 16455 18262
rect 23473 18259 23539 18262
rect 23749 18322 23815 18325
rect 24672 18322 24732 18534
rect 27520 18504 28000 18534
rect 23749 18320 24732 18322
rect 23749 18264 23754 18320
rect 23810 18264 24732 18320
rect 23749 18262 24732 18264
rect 23749 18259 23815 18262
rect 17769 18186 17835 18189
rect 11470 18184 17835 18186
rect 11470 18128 17774 18184
rect 17830 18128 17835 18184
rect 11470 18126 17835 18128
rect 8109 18123 8175 18126
rect 11237 18123 11303 18126
rect 17769 18123 17835 18126
rect 22737 18186 22803 18189
rect 23841 18186 23907 18189
rect 22737 18184 23907 18186
rect 22737 18128 22742 18184
rect 22798 18128 23846 18184
rect 23902 18128 23907 18184
rect 22737 18126 23907 18128
rect 22737 18123 22803 18126
rect 23841 18123 23907 18126
rect 3509 18050 3575 18053
rect 10041 18050 10107 18053
rect 3509 18048 10107 18050
rect 3509 17992 3514 18048
rect 3570 17992 10046 18048
rect 10102 17992 10107 18048
rect 3509 17990 10107 17992
rect 3509 17987 3575 17990
rect 10041 17987 10107 17990
rect 10277 17984 10597 17985
rect 0 17914 480 17944
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 3233 17914 3299 17917
rect 0 17912 3299 17914
rect 0 17856 3238 17912
rect 3294 17856 3299 17912
rect 0 17854 3299 17856
rect 0 17824 480 17854
rect 3233 17851 3299 17854
rect 3969 17914 4035 17917
rect 6729 17914 6795 17917
rect 3969 17912 6795 17914
rect 3969 17856 3974 17912
rect 4030 17856 6734 17912
rect 6790 17856 6795 17912
rect 3969 17854 6795 17856
rect 3969 17851 4035 17854
rect 6729 17851 6795 17854
rect 6913 17914 6979 17917
rect 9949 17914 10015 17917
rect 6913 17912 10015 17914
rect 6913 17856 6918 17912
rect 6974 17856 9954 17912
rect 10010 17856 10015 17912
rect 6913 17854 10015 17856
rect 6913 17851 6979 17854
rect 9949 17851 10015 17854
rect 10685 17914 10751 17917
rect 15285 17914 15351 17917
rect 10685 17912 15351 17914
rect 10685 17856 10690 17912
rect 10746 17856 15290 17912
rect 15346 17856 15351 17912
rect 10685 17854 15351 17856
rect 10685 17851 10751 17854
rect 15285 17851 15351 17854
rect 23473 17914 23539 17917
rect 27520 17914 28000 17944
rect 23473 17912 28000 17914
rect 23473 17856 23478 17912
rect 23534 17856 28000 17912
rect 23473 17854 28000 17856
rect 23473 17851 23539 17854
rect 27520 17824 28000 17854
rect 8017 17778 8083 17781
rect 15745 17778 15811 17781
rect 8017 17776 15811 17778
rect 8017 17720 8022 17776
rect 8078 17720 15750 17776
rect 15806 17720 15811 17776
rect 8017 17718 15811 17720
rect 8017 17715 8083 17718
rect 15745 17715 15811 17718
rect 16481 17778 16547 17781
rect 16481 17776 16682 17778
rect 16481 17720 16486 17776
rect 16542 17720 16682 17776
rect 16481 17718 16682 17720
rect 16481 17715 16547 17718
rect 9857 17642 9923 17645
rect 4846 17640 9923 17642
rect 4846 17584 9862 17640
rect 9918 17584 9923 17640
rect 4846 17582 9923 17584
rect 0 17370 480 17400
rect 4846 17370 4906 17582
rect 9857 17579 9923 17582
rect 10961 17642 11027 17645
rect 13629 17642 13695 17645
rect 10961 17640 13695 17642
rect 10961 17584 10966 17640
rect 11022 17584 13634 17640
rect 13690 17584 13695 17640
rect 10961 17582 13695 17584
rect 10961 17579 11027 17582
rect 13629 17579 13695 17582
rect 14457 17642 14523 17645
rect 16481 17642 16547 17645
rect 14457 17640 16547 17642
rect 14457 17584 14462 17640
rect 14518 17584 16486 17640
rect 16542 17584 16547 17640
rect 14457 17582 16547 17584
rect 16622 17642 16682 17718
rect 20161 17642 20227 17645
rect 16622 17640 20227 17642
rect 16622 17584 20166 17640
rect 20222 17584 20227 17640
rect 16622 17582 20227 17584
rect 14457 17579 14523 17582
rect 16481 17579 16547 17582
rect 20161 17579 20227 17582
rect 8569 17506 8635 17509
rect 14549 17506 14615 17509
rect 8569 17504 14615 17506
rect 8569 17448 8574 17504
rect 8630 17448 14554 17504
rect 14610 17448 14615 17504
rect 8569 17446 14615 17448
rect 8569 17443 8635 17446
rect 14549 17443 14615 17446
rect 16297 17506 16363 17509
rect 20621 17506 20687 17509
rect 16297 17504 20687 17506
rect 16297 17448 16302 17504
rect 16358 17448 20626 17504
rect 20682 17448 20687 17504
rect 16297 17446 20687 17448
rect 16297 17443 16363 17446
rect 20621 17443 20687 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 0 17310 4906 17370
rect 9949 17370 10015 17373
rect 10910 17370 10916 17372
rect 9949 17368 10916 17370
rect 9949 17312 9954 17368
rect 10010 17312 10916 17368
rect 9949 17310 10916 17312
rect 0 17280 480 17310
rect 9949 17307 10015 17310
rect 10910 17308 10916 17310
rect 10980 17308 10986 17372
rect 17493 17370 17559 17373
rect 18597 17370 18663 17373
rect 19425 17370 19491 17373
rect 17493 17368 19491 17370
rect 17493 17312 17498 17368
rect 17554 17312 18602 17368
rect 18658 17312 19430 17368
rect 19486 17312 19491 17368
rect 17493 17310 19491 17312
rect 17493 17307 17559 17310
rect 18597 17307 18663 17310
rect 19425 17307 19491 17310
rect 24761 17370 24827 17373
rect 27520 17370 28000 17400
rect 24761 17368 28000 17370
rect 24761 17312 24766 17368
rect 24822 17312 28000 17368
rect 24761 17310 28000 17312
rect 24761 17307 24827 17310
rect 27520 17280 28000 17310
rect 1761 17234 1827 17237
rect 6729 17234 6795 17237
rect 1761 17232 6795 17234
rect 1761 17176 1766 17232
rect 1822 17176 6734 17232
rect 6790 17176 6795 17232
rect 1761 17174 6795 17176
rect 1761 17171 1827 17174
rect 6729 17171 6795 17174
rect 9581 17234 9647 17237
rect 15929 17234 15995 17237
rect 9581 17232 15995 17234
rect 9581 17176 9586 17232
rect 9642 17176 15934 17232
rect 15990 17176 15995 17232
rect 9581 17174 15995 17176
rect 9581 17171 9647 17174
rect 15929 17171 15995 17174
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 4521 16826 4587 16829
rect 7557 16826 7623 16829
rect 4521 16824 7623 16826
rect 4521 16768 4526 16824
rect 4582 16768 7562 16824
rect 7618 16768 7623 16824
rect 4521 16766 7623 16768
rect 4521 16763 4587 16766
rect 7557 16763 7623 16766
rect 11421 16826 11487 16829
rect 13997 16826 14063 16829
rect 11421 16824 14063 16826
rect 11421 16768 11426 16824
rect 11482 16768 14002 16824
rect 14058 16768 14063 16824
rect 11421 16766 14063 16768
rect 11421 16763 11487 16766
rect 13997 16763 14063 16766
rect 22185 16826 22251 16829
rect 23749 16826 23815 16829
rect 22185 16824 23815 16826
rect 22185 16768 22190 16824
rect 22246 16768 23754 16824
rect 23810 16768 23815 16824
rect 22185 16766 23815 16768
rect 22185 16763 22251 16766
rect 23749 16763 23815 16766
rect 0 16690 480 16720
rect 6729 16690 6795 16693
rect 0 16688 6795 16690
rect 0 16632 6734 16688
rect 6790 16632 6795 16688
rect 0 16630 6795 16632
rect 0 16600 480 16630
rect 6729 16627 6795 16630
rect 7097 16690 7163 16693
rect 9673 16690 9739 16693
rect 7097 16688 9739 16690
rect 7097 16632 7102 16688
rect 7158 16632 9678 16688
rect 9734 16632 9739 16688
rect 7097 16630 9739 16632
rect 7097 16627 7163 16630
rect 9673 16627 9739 16630
rect 18873 16690 18939 16693
rect 22461 16690 22527 16693
rect 18873 16688 22527 16690
rect 18873 16632 18878 16688
rect 18934 16632 22466 16688
rect 22522 16632 22527 16688
rect 18873 16630 22527 16632
rect 18873 16627 18939 16630
rect 22461 16627 22527 16630
rect 26049 16690 26115 16693
rect 27520 16690 28000 16720
rect 26049 16688 28000 16690
rect 26049 16632 26054 16688
rect 26110 16632 28000 16688
rect 26049 16630 28000 16632
rect 26049 16627 26115 16630
rect 27520 16600 28000 16630
rect 6637 16554 6703 16557
rect 13721 16554 13787 16557
rect 19333 16554 19399 16557
rect 6637 16552 13787 16554
rect 6637 16496 6642 16552
rect 6698 16496 13726 16552
rect 13782 16496 13787 16552
rect 6637 16494 13787 16496
rect 6637 16491 6703 16494
rect 13721 16491 13787 16494
rect 14782 16552 19399 16554
rect 14782 16496 19338 16552
rect 19394 16496 19399 16552
rect 14782 16494 19399 16496
rect 6913 16418 6979 16421
rect 14782 16418 14842 16494
rect 19333 16491 19399 16494
rect 20069 16554 20135 16557
rect 21633 16554 21699 16557
rect 24761 16554 24827 16557
rect 20069 16552 20178 16554
rect 20069 16496 20074 16552
rect 20130 16496 20178 16552
rect 20069 16491 20178 16496
rect 21633 16552 24827 16554
rect 21633 16496 21638 16552
rect 21694 16496 24766 16552
rect 24822 16496 24827 16552
rect 21633 16494 24827 16496
rect 21633 16491 21699 16494
rect 24761 16491 24827 16494
rect 20118 16421 20178 16491
rect 6913 16416 14842 16418
rect 6913 16360 6918 16416
rect 6974 16360 14842 16416
rect 6913 16358 14842 16360
rect 16205 16418 16271 16421
rect 19977 16418 20043 16421
rect 16205 16416 20043 16418
rect 16205 16360 16210 16416
rect 16266 16360 19982 16416
rect 20038 16360 20043 16416
rect 16205 16358 20043 16360
rect 20118 16416 20227 16421
rect 20118 16360 20166 16416
rect 20222 16360 20227 16416
rect 20118 16358 20227 16360
rect 6913 16355 6979 16358
rect 16205 16355 16271 16358
rect 19977 16355 20043 16358
rect 20161 16355 20227 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 10961 16282 11027 16285
rect 12525 16282 12591 16285
rect 10961 16280 12591 16282
rect 10961 16224 10966 16280
rect 11022 16224 12530 16280
rect 12586 16224 12591 16280
rect 10961 16222 12591 16224
rect 10961 16219 11027 16222
rect 12525 16219 12591 16222
rect 0 16146 480 16176
rect 1577 16146 1643 16149
rect 0 16144 1643 16146
rect 0 16088 1582 16144
rect 1638 16088 1643 16144
rect 0 16086 1643 16088
rect 0 16056 480 16086
rect 1577 16083 1643 16086
rect 3785 16146 3851 16149
rect 7005 16146 7071 16149
rect 3785 16144 7071 16146
rect 3785 16088 3790 16144
rect 3846 16088 7010 16144
rect 7066 16088 7071 16144
rect 3785 16086 7071 16088
rect 3785 16083 3851 16086
rect 7005 16083 7071 16086
rect 7189 16146 7255 16149
rect 13445 16146 13511 16149
rect 7189 16144 13511 16146
rect 7189 16088 7194 16144
rect 7250 16088 13450 16144
rect 13506 16088 13511 16144
rect 7189 16086 13511 16088
rect 7189 16083 7255 16086
rect 13445 16083 13511 16086
rect 13629 16146 13695 16149
rect 24209 16146 24275 16149
rect 27520 16146 28000 16176
rect 13629 16144 23674 16146
rect 13629 16088 13634 16144
rect 13690 16088 23674 16144
rect 13629 16086 23674 16088
rect 13629 16083 13695 16086
rect 11697 16010 11763 16013
rect 21449 16010 21515 16013
rect 22737 16010 22803 16013
rect 11697 16008 21515 16010
rect 11697 15952 11702 16008
rect 11758 15952 21454 16008
rect 21510 15952 21515 16008
rect 11697 15950 21515 15952
rect 11697 15947 11763 15950
rect 21449 15947 21515 15950
rect 21590 16008 22803 16010
rect 21590 15952 22742 16008
rect 22798 15952 22803 16008
rect 21590 15950 22803 15952
rect 23614 16010 23674 16086
rect 24209 16144 28000 16146
rect 24209 16088 24214 16144
rect 24270 16088 28000 16144
rect 24209 16086 28000 16088
rect 24209 16083 24275 16086
rect 27520 16056 28000 16086
rect 24025 16010 24091 16013
rect 24710 16010 24716 16012
rect 23614 16008 24716 16010
rect 23614 15952 24030 16008
rect 24086 15952 24716 16008
rect 23614 15950 24716 15952
rect 197 15874 263 15877
rect 6453 15874 6519 15877
rect 197 15872 6519 15874
rect 197 15816 202 15872
rect 258 15816 6458 15872
rect 6514 15816 6519 15872
rect 197 15814 6519 15816
rect 197 15811 263 15814
rect 6453 15811 6519 15814
rect 13721 15874 13787 15877
rect 18781 15874 18847 15877
rect 13721 15872 18847 15874
rect 13721 15816 13726 15872
rect 13782 15816 18786 15872
rect 18842 15816 18847 15872
rect 13721 15814 18847 15816
rect 13721 15811 13787 15814
rect 18781 15811 18847 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 5441 15738 5507 15741
rect 7649 15738 7715 15741
rect 5441 15736 7715 15738
rect 5441 15680 5446 15736
rect 5502 15680 7654 15736
rect 7710 15680 7715 15736
rect 5441 15678 7715 15680
rect 5441 15675 5507 15678
rect 7649 15675 7715 15678
rect 10777 15738 10843 15741
rect 13445 15738 13511 15741
rect 10777 15736 13511 15738
rect 10777 15680 10782 15736
rect 10838 15680 13450 15736
rect 13506 15680 13511 15736
rect 10777 15678 13511 15680
rect 10777 15675 10843 15678
rect 13445 15675 13511 15678
rect 1761 15602 1827 15605
rect 3601 15602 3667 15605
rect 7465 15602 7531 15605
rect 1761 15600 7531 15602
rect 1761 15544 1766 15600
rect 1822 15544 3606 15600
rect 3662 15544 7470 15600
rect 7526 15544 7531 15600
rect 1761 15542 7531 15544
rect 1761 15539 1827 15542
rect 3601 15539 3667 15542
rect 7465 15539 7531 15542
rect 12985 15602 13051 15605
rect 13445 15602 13511 15605
rect 20069 15602 20135 15605
rect 21449 15602 21515 15605
rect 12985 15600 19994 15602
rect 12985 15544 12990 15600
rect 13046 15544 13450 15600
rect 13506 15544 19994 15600
rect 12985 15542 19994 15544
rect 12985 15539 13051 15542
rect 13445 15539 13511 15542
rect 0 15466 480 15496
rect 1485 15466 1551 15469
rect 0 15464 1551 15466
rect 0 15408 1490 15464
rect 1546 15408 1551 15464
rect 0 15406 1551 15408
rect 19934 15466 19994 15542
rect 20069 15600 21515 15602
rect 20069 15544 20074 15600
rect 20130 15544 21454 15600
rect 21510 15544 21515 15600
rect 20069 15542 21515 15544
rect 20069 15539 20135 15542
rect 21449 15539 21515 15542
rect 21590 15466 21650 15950
rect 22737 15947 22803 15950
rect 24025 15947 24091 15950
rect 24710 15948 24716 15950
rect 24780 15948 24786 16012
rect 22001 15738 22067 15741
rect 23473 15738 23539 15741
rect 22001 15736 23539 15738
rect 22001 15680 22006 15736
rect 22062 15680 23478 15736
rect 23534 15680 23539 15736
rect 22001 15678 23539 15680
rect 22001 15675 22067 15678
rect 23473 15675 23539 15678
rect 21909 15602 21975 15605
rect 24577 15602 24643 15605
rect 21909 15600 24643 15602
rect 21909 15544 21914 15600
rect 21970 15544 24582 15600
rect 24638 15544 24643 15600
rect 21909 15542 24643 15544
rect 21909 15539 21975 15542
rect 24577 15539 24643 15542
rect 19934 15406 21650 15466
rect 24025 15466 24091 15469
rect 27520 15466 28000 15496
rect 24025 15464 28000 15466
rect 24025 15408 24030 15464
rect 24086 15408 28000 15464
rect 24025 15406 28000 15408
rect 0 15376 480 15406
rect 1485 15403 1551 15406
rect 24025 15403 24091 15406
rect 27520 15376 28000 15406
rect 16481 15330 16547 15333
rect 18045 15330 18111 15333
rect 16481 15328 18111 15330
rect 16481 15272 16486 15328
rect 16542 15272 18050 15328
rect 18106 15272 18111 15328
rect 16481 15270 18111 15272
rect 16481 15267 16547 15270
rect 18045 15267 18111 15270
rect 19149 15330 19215 15333
rect 23238 15330 23244 15332
rect 19149 15328 23244 15330
rect 19149 15272 19154 15328
rect 19210 15272 23244 15328
rect 19149 15270 23244 15272
rect 19149 15267 19215 15270
rect 23238 15268 23244 15270
rect 23308 15268 23314 15332
rect 26509 15330 26575 15333
rect 24672 15328 26575 15330
rect 24672 15272 26514 15328
rect 26570 15272 26575 15328
rect 24672 15270 26575 15272
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 14273 15194 14339 15197
rect 6134 15192 14339 15194
rect 6134 15136 14278 15192
rect 14334 15136 14339 15192
rect 6134 15134 14339 15136
rect 4061 15058 4127 15061
rect 6134 15058 6194 15134
rect 14273 15131 14339 15134
rect 21725 15194 21791 15197
rect 23381 15194 23447 15197
rect 21725 15192 23447 15194
rect 21725 15136 21730 15192
rect 21786 15136 23386 15192
rect 23442 15136 23447 15192
rect 21725 15134 23447 15136
rect 21725 15131 21791 15134
rect 23381 15131 23447 15134
rect 4061 15056 6194 15058
rect 4061 15000 4066 15056
rect 4122 15000 6194 15056
rect 4061 14998 6194 15000
rect 7373 15058 7439 15061
rect 10041 15058 10107 15061
rect 7373 15056 10107 15058
rect 7373 15000 7378 15056
rect 7434 15000 10046 15056
rect 10102 15000 10107 15056
rect 7373 14998 10107 15000
rect 4061 14995 4127 14998
rect 7373 14995 7439 14998
rect 10041 14995 10107 14998
rect 12433 15058 12499 15061
rect 23381 15058 23447 15061
rect 24672 15058 24732 15270
rect 26509 15267 26575 15270
rect 12433 15056 20684 15058
rect 12433 15000 12438 15056
rect 12494 15000 20684 15056
rect 12433 14998 20684 15000
rect 12433 14995 12499 14998
rect 0 14922 480 14952
rect 3693 14922 3759 14925
rect 5809 14922 5875 14925
rect 0 14862 2744 14922
rect 0 14832 480 14862
rect 2684 14786 2744 14862
rect 3693 14920 5875 14922
rect 3693 14864 3698 14920
rect 3754 14864 5814 14920
rect 5870 14864 5875 14920
rect 3693 14862 5875 14864
rect 3693 14859 3759 14862
rect 5809 14859 5875 14862
rect 7465 14922 7531 14925
rect 10501 14922 10567 14925
rect 7465 14920 10567 14922
rect 7465 14864 7470 14920
rect 7526 14864 10506 14920
rect 10562 14864 10567 14920
rect 7465 14862 10567 14864
rect 7465 14859 7531 14862
rect 10501 14859 10567 14862
rect 5901 14786 5967 14789
rect 2684 14784 5967 14786
rect 2684 14728 5906 14784
rect 5962 14728 5967 14784
rect 2684 14726 5967 14728
rect 20624 14786 20684 14998
rect 23381 15056 24732 15058
rect 23381 15000 23386 15056
rect 23442 15000 24732 15056
rect 23381 14998 24732 15000
rect 23381 14995 23447 14998
rect 23422 14860 23428 14924
rect 23492 14922 23498 14924
rect 27520 14922 28000 14952
rect 23492 14862 28000 14922
rect 23492 14860 23498 14862
rect 27520 14832 28000 14862
rect 20805 14786 20871 14789
rect 25589 14786 25655 14789
rect 20624 14784 25655 14786
rect 20624 14728 20810 14784
rect 20866 14728 25594 14784
rect 25650 14728 25655 14784
rect 20624 14726 25655 14728
rect 5901 14723 5967 14726
rect 20805 14723 20871 14726
rect 25589 14723 25655 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 0 14378 480 14408
rect 4061 14378 4127 14381
rect 0 14376 4127 14378
rect 0 14320 4066 14376
rect 4122 14320 4127 14376
rect 0 14318 4127 14320
rect 0 14288 480 14318
rect 4061 14315 4127 14318
rect 7741 14378 7807 14381
rect 17401 14378 17467 14381
rect 19517 14378 19583 14381
rect 19701 14378 19767 14381
rect 7741 14376 17234 14378
rect 7741 14320 7746 14376
rect 7802 14320 17234 14376
rect 7741 14318 17234 14320
rect 7741 14315 7807 14318
rect 17174 14242 17234 14318
rect 17401 14376 19767 14378
rect 17401 14320 17406 14376
rect 17462 14320 19522 14376
rect 19578 14320 19706 14376
rect 19762 14320 19767 14376
rect 17401 14318 19767 14320
rect 17401 14315 17467 14318
rect 19517 14315 19583 14318
rect 19701 14315 19767 14318
rect 22553 14378 22619 14381
rect 27520 14378 28000 14408
rect 22553 14376 28000 14378
rect 22553 14320 22558 14376
rect 22614 14320 28000 14376
rect 22553 14318 28000 14320
rect 22553 14315 22619 14318
rect 27520 14288 28000 14318
rect 20069 14242 20135 14245
rect 17174 14240 20135 14242
rect 17174 14184 20074 14240
rect 20130 14184 20135 14240
rect 17174 14182 20135 14184
rect 20069 14179 20135 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 16389 14106 16455 14109
rect 18413 14106 18479 14109
rect 16389 14104 18479 14106
rect 16389 14048 16394 14104
rect 16450 14048 18418 14104
rect 18474 14048 18479 14104
rect 16389 14046 18479 14048
rect 16389 14043 16455 14046
rect 18413 14043 18479 14046
rect 7281 13970 7347 13973
rect 10869 13970 10935 13973
rect 16021 13970 16087 13973
rect 7281 13968 8402 13970
rect 7281 13912 7286 13968
rect 7342 13912 8402 13968
rect 7281 13910 8402 13912
rect 7281 13907 7347 13910
rect 4981 13834 5047 13837
rect 8201 13834 8267 13837
rect 4981 13832 8267 13834
rect 4981 13776 4986 13832
rect 5042 13776 8206 13832
rect 8262 13776 8267 13832
rect 4981 13774 8267 13776
rect 8342 13834 8402 13910
rect 10869 13968 16087 13970
rect 10869 13912 10874 13968
rect 10930 13912 16026 13968
rect 16082 13912 16087 13968
rect 10869 13910 16087 13912
rect 10869 13907 10935 13910
rect 16021 13907 16087 13910
rect 15653 13834 15719 13837
rect 8342 13832 15719 13834
rect 8342 13776 15658 13832
rect 15714 13776 15719 13832
rect 8342 13774 15719 13776
rect 4981 13771 5047 13774
rect 8201 13771 8267 13774
rect 15653 13771 15719 13774
rect 21817 13834 21883 13837
rect 24117 13834 24183 13837
rect 21817 13832 24183 13834
rect 21817 13776 21822 13832
rect 21878 13776 24122 13832
rect 24178 13776 24183 13832
rect 21817 13774 24183 13776
rect 21817 13771 21883 13774
rect 24117 13771 24183 13774
rect 0 13698 480 13728
rect 3785 13698 3851 13701
rect 5073 13698 5139 13701
rect 5533 13698 5599 13701
rect 0 13638 3618 13698
rect 0 13608 480 13638
rect 3558 13562 3618 13638
rect 3785 13696 5599 13698
rect 3785 13640 3790 13696
rect 3846 13640 5078 13696
rect 5134 13640 5538 13696
rect 5594 13640 5599 13696
rect 3785 13638 5599 13640
rect 3785 13635 3851 13638
rect 5073 13635 5139 13638
rect 5533 13635 5599 13638
rect 5809 13698 5875 13701
rect 9305 13698 9371 13701
rect 9581 13698 9647 13701
rect 5809 13696 9647 13698
rect 5809 13640 5814 13696
rect 5870 13640 9310 13696
rect 9366 13640 9586 13696
rect 9642 13640 9647 13696
rect 5809 13638 9647 13640
rect 5809 13635 5875 13638
rect 9305 13635 9371 13638
rect 9581 13635 9647 13638
rect 13997 13698 14063 13701
rect 17861 13698 17927 13701
rect 13997 13696 17927 13698
rect 13997 13640 14002 13696
rect 14058 13640 17866 13696
rect 17922 13640 17927 13696
rect 13997 13638 17927 13640
rect 13997 13635 14063 13638
rect 17861 13635 17927 13638
rect 20437 13698 20503 13701
rect 27520 13698 28000 13728
rect 20437 13696 28000 13698
rect 20437 13640 20442 13696
rect 20498 13640 28000 13696
rect 20437 13638 28000 13640
rect 20437 13635 20503 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 27520 13608 28000 13638
rect 19610 13567 19930 13568
rect 6913 13562 6979 13565
rect 3558 13560 6979 13562
rect 3558 13504 6918 13560
rect 6974 13504 6979 13560
rect 3558 13502 6979 13504
rect 6913 13499 6979 13502
rect 14549 13562 14615 13565
rect 17033 13562 17099 13565
rect 19333 13562 19399 13565
rect 14549 13560 19399 13562
rect 14549 13504 14554 13560
rect 14610 13504 17038 13560
rect 17094 13504 19338 13560
rect 19394 13504 19399 13560
rect 14549 13502 19399 13504
rect 14549 13499 14615 13502
rect 17033 13499 17099 13502
rect 19333 13499 19399 13502
rect 17585 13426 17651 13429
rect 21081 13426 21147 13429
rect 17585 13424 21147 13426
rect 17585 13368 17590 13424
rect 17646 13368 21086 13424
rect 21142 13368 21147 13424
rect 17585 13366 21147 13368
rect 17585 13363 17651 13366
rect 21081 13363 21147 13366
rect 21357 13426 21423 13429
rect 23565 13426 23631 13429
rect 21357 13424 23631 13426
rect 21357 13368 21362 13424
rect 21418 13368 23570 13424
rect 23626 13368 23631 13424
rect 21357 13366 23631 13368
rect 21357 13363 21423 13366
rect 23565 13363 23631 13366
rect 23749 13426 23815 13429
rect 23749 13424 24962 13426
rect 23749 13368 23754 13424
rect 23810 13368 24962 13424
rect 23749 13366 24962 13368
rect 23749 13363 23815 13366
rect 14181 13290 14247 13293
rect 24669 13290 24735 13293
rect 14181 13288 24735 13290
rect 14181 13232 14186 13288
rect 14242 13232 24674 13288
rect 24730 13232 24735 13288
rect 14181 13230 24735 13232
rect 14181 13227 14247 13230
rect 24669 13227 24735 13230
rect 0 13154 480 13184
rect 2865 13154 2931 13157
rect 0 13152 2931 13154
rect 0 13096 2870 13152
rect 2926 13096 2931 13152
rect 0 13094 2931 13096
rect 0 13064 480 13094
rect 2865 13091 2931 13094
rect 15929 13154 15995 13157
rect 18321 13154 18387 13157
rect 19701 13154 19767 13157
rect 15929 13152 18387 13154
rect 15929 13096 15934 13152
rect 15990 13096 18326 13152
rect 18382 13096 18387 13152
rect 15929 13094 18387 13096
rect 15929 13091 15995 13094
rect 18321 13091 18387 13094
rect 18508 13152 19767 13154
rect 18508 13096 19706 13152
rect 19762 13096 19767 13152
rect 18508 13094 19767 13096
rect 24902 13154 24962 13366
rect 27520 13154 28000 13184
rect 24902 13094 28000 13154
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 9581 13018 9647 13021
rect 13997 13018 14063 13021
rect 9581 13016 14063 13018
rect 9581 12960 9586 13016
rect 9642 12960 14002 13016
rect 14058 12960 14063 13016
rect 9581 12958 14063 12960
rect 9581 12955 9647 12958
rect 13997 12955 14063 12958
rect 6453 12882 6519 12885
rect 13997 12882 14063 12885
rect 18508 12882 18568 13094
rect 19701 13091 19767 13094
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 27520 13064 28000 13094
rect 24277 13023 24597 13024
rect 19149 13018 19215 13021
rect 20345 13018 20411 13021
rect 23289 13020 23355 13021
rect 23238 13018 23244 13020
rect 19149 13016 20411 13018
rect 19149 12960 19154 13016
rect 19210 12960 20350 13016
rect 20406 12960 20411 13016
rect 19149 12958 20411 12960
rect 23198 12958 23244 13018
rect 23308 13016 23355 13020
rect 24025 13018 24091 13021
rect 23350 12960 23355 13016
rect 19149 12955 19215 12958
rect 20345 12955 20411 12958
rect 23238 12956 23244 12958
rect 23308 12956 23355 12960
rect 23289 12955 23355 12956
rect 23798 13016 24091 13018
rect 23798 12960 24030 13016
rect 24086 12960 24091 13016
rect 23798 12958 24091 12960
rect 6453 12880 18568 12882
rect 6453 12824 6458 12880
rect 6514 12824 14002 12880
rect 14058 12824 18568 12880
rect 6453 12822 18568 12824
rect 18689 12882 18755 12885
rect 20989 12882 21055 12885
rect 18689 12880 21055 12882
rect 18689 12824 18694 12880
rect 18750 12824 20994 12880
rect 21050 12824 21055 12880
rect 18689 12822 21055 12824
rect 6453 12819 6519 12822
rect 13997 12819 14063 12822
rect 18689 12819 18755 12822
rect 20989 12819 21055 12822
rect 10777 12746 10843 12749
rect 23798 12746 23858 12958
rect 24025 12955 24091 12958
rect 24117 12882 24183 12885
rect 24117 12880 24226 12882
rect 24117 12824 24122 12880
rect 24178 12824 24226 12880
rect 24117 12819 24226 12824
rect 10777 12744 23858 12746
rect 10777 12688 10782 12744
rect 10838 12688 23858 12744
rect 10777 12686 23858 12688
rect 24166 12746 24226 12819
rect 24577 12746 24643 12749
rect 24166 12744 24643 12746
rect 24166 12688 24582 12744
rect 24638 12688 24643 12744
rect 24166 12686 24643 12688
rect 10777 12683 10843 12686
rect 24577 12683 24643 12686
rect 3693 12610 3759 12613
rect 6085 12610 6151 12613
rect 15009 12610 15075 12613
rect 3693 12608 6151 12610
rect 3693 12552 3698 12608
rect 3754 12552 6090 12608
rect 6146 12552 6151 12608
rect 3693 12550 6151 12552
rect 3693 12547 3759 12550
rect 6085 12547 6151 12550
rect 10734 12608 15075 12610
rect 10734 12552 15014 12608
rect 15070 12552 15075 12608
rect 10734 12550 15075 12552
rect 10277 12544 10597 12545
rect 0 12474 480 12504
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 0 12414 10058 12474
rect 0 12384 480 12414
rect 9998 12338 10058 12414
rect 10734 12338 10794 12550
rect 15009 12547 15075 12550
rect 15285 12610 15351 12613
rect 16481 12610 16547 12613
rect 15285 12608 16547 12610
rect 15285 12552 15290 12608
rect 15346 12552 16486 12608
rect 16542 12552 16547 12608
rect 15285 12550 16547 12552
rect 15285 12547 15351 12550
rect 16481 12547 16547 12550
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 14365 12474 14431 12477
rect 16481 12474 16547 12477
rect 14365 12472 16547 12474
rect 14365 12416 14370 12472
rect 14426 12416 16486 12472
rect 16542 12416 16547 12472
rect 14365 12414 16547 12416
rect 14365 12411 14431 12414
rect 16481 12411 16547 12414
rect 20345 12474 20411 12477
rect 27520 12474 28000 12504
rect 20345 12472 28000 12474
rect 20345 12416 20350 12472
rect 20406 12416 28000 12472
rect 20345 12414 28000 12416
rect 20345 12411 20411 12414
rect 27520 12384 28000 12414
rect 9998 12278 10794 12338
rect 14089 12338 14155 12341
rect 15745 12338 15811 12341
rect 17309 12338 17375 12341
rect 22553 12338 22619 12341
rect 14089 12336 16498 12338
rect 14089 12280 14094 12336
rect 14150 12280 15750 12336
rect 15806 12280 16498 12336
rect 14089 12278 16498 12280
rect 14089 12275 14155 12278
rect 15745 12275 15811 12278
rect 12065 12202 12131 12205
rect 2868 12200 12131 12202
rect 2868 12144 12070 12200
rect 12126 12144 12131 12200
rect 2868 12142 12131 12144
rect 2868 12066 2928 12142
rect 12065 12139 12131 12142
rect 13077 12202 13143 12205
rect 16205 12202 16271 12205
rect 13077 12200 16271 12202
rect 13077 12144 13082 12200
rect 13138 12144 16210 12200
rect 16266 12144 16271 12200
rect 13077 12142 16271 12144
rect 13077 12139 13143 12142
rect 16205 12139 16271 12142
rect 2684 12006 2928 12066
rect 16205 12066 16271 12069
rect 16438 12066 16498 12278
rect 17309 12336 22619 12338
rect 17309 12280 17314 12336
rect 17370 12280 22558 12336
rect 22614 12280 22619 12336
rect 17309 12278 22619 12280
rect 17309 12275 17375 12278
rect 22553 12275 22619 12278
rect 24669 12338 24735 12341
rect 25681 12338 25747 12341
rect 24669 12336 25747 12338
rect 24669 12280 24674 12336
rect 24730 12280 25686 12336
rect 25742 12280 25747 12336
rect 24669 12278 25747 12280
rect 24669 12275 24735 12278
rect 25681 12275 25747 12278
rect 20529 12202 20595 12205
rect 20529 12200 24962 12202
rect 20529 12144 20534 12200
rect 20590 12144 24962 12200
rect 20529 12142 24962 12144
rect 20529 12139 20595 12142
rect 21633 12066 21699 12069
rect 16205 12064 16498 12066
rect 16205 12008 16210 12064
rect 16266 12008 16498 12064
rect 16205 12006 16498 12008
rect 16622 12064 21699 12066
rect 16622 12008 21638 12064
rect 21694 12008 21699 12064
rect 16622 12006 21699 12008
rect 0 11930 480 11960
rect 2684 11930 2744 12006
rect 16205 12003 16271 12006
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 16622 11930 16682 12006
rect 21633 12003 21699 12006
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 0 11870 2744 11930
rect 15334 11870 16682 11930
rect 18781 11930 18847 11933
rect 23197 11930 23263 11933
rect 18781 11928 23263 11930
rect 18781 11872 18786 11928
rect 18842 11872 23202 11928
rect 23258 11872 23263 11928
rect 18781 11870 23263 11872
rect 24902 11930 24962 12142
rect 27520 11930 28000 11960
rect 24902 11870 28000 11930
rect 0 11840 480 11870
rect 14365 11794 14431 11797
rect 15334 11794 15394 11870
rect 18781 11867 18847 11870
rect 23197 11867 23263 11870
rect 27520 11840 28000 11870
rect 14365 11792 15394 11794
rect 14365 11736 14370 11792
rect 14426 11736 15394 11792
rect 14365 11734 15394 11736
rect 16021 11794 16087 11797
rect 25497 11794 25563 11797
rect 16021 11792 25563 11794
rect 16021 11736 16026 11792
rect 16082 11736 25502 11792
rect 25558 11736 25563 11792
rect 16021 11734 25563 11736
rect 14365 11731 14431 11734
rect 16021 11731 16087 11734
rect 25497 11731 25563 11734
rect 3969 11658 4035 11661
rect 13813 11658 13879 11661
rect 3969 11656 13879 11658
rect 3969 11600 3974 11656
rect 4030 11600 13818 11656
rect 13874 11600 13879 11656
rect 3969 11598 13879 11600
rect 3969 11595 4035 11598
rect 13813 11595 13879 11598
rect 15561 11658 15627 11661
rect 21449 11658 21515 11661
rect 15561 11656 21515 11658
rect 15561 11600 15566 11656
rect 15622 11600 21454 11656
rect 21510 11600 21515 11656
rect 15561 11598 21515 11600
rect 15561 11595 15627 11598
rect 21449 11595 21515 11598
rect 21633 11658 21699 11661
rect 25037 11658 25103 11661
rect 21633 11656 25103 11658
rect 21633 11600 21638 11656
rect 21694 11600 25042 11656
rect 25098 11600 25103 11656
rect 21633 11598 25103 11600
rect 21633 11595 21699 11598
rect 25037 11595 25103 11598
rect 23197 11522 23263 11525
rect 23565 11522 23631 11525
rect 23197 11520 23631 11522
rect 23197 11464 23202 11520
rect 23258 11464 23570 11520
rect 23626 11464 23631 11520
rect 23197 11462 23631 11464
rect 23197 11459 23263 11462
rect 23565 11459 23631 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 4705 11386 4771 11389
rect 7833 11386 7899 11389
rect 4705 11384 7899 11386
rect 4705 11328 4710 11384
rect 4766 11328 7838 11384
rect 7894 11328 7899 11384
rect 4705 11326 7899 11328
rect 4705 11323 4771 11326
rect 7833 11323 7899 11326
rect 14089 11386 14155 11389
rect 19425 11386 19491 11389
rect 14089 11384 19491 11386
rect 14089 11328 14094 11384
rect 14150 11328 19430 11384
rect 19486 11328 19491 11384
rect 14089 11326 19491 11328
rect 14089 11323 14155 11326
rect 19425 11323 19491 11326
rect 0 11250 480 11280
rect 11053 11250 11119 11253
rect 0 11248 11119 11250
rect 0 11192 11058 11248
rect 11114 11192 11119 11248
rect 0 11190 11119 11192
rect 0 11160 480 11190
rect 11053 11187 11119 11190
rect 24577 11250 24643 11253
rect 24710 11250 24716 11252
rect 24577 11248 24716 11250
rect 24577 11192 24582 11248
rect 24638 11192 24716 11248
rect 24577 11190 24716 11192
rect 24577 11187 24643 11190
rect 24710 11188 24716 11190
rect 24780 11188 24786 11252
rect 25589 11250 25655 11253
rect 27520 11250 28000 11280
rect 25589 11248 28000 11250
rect 25589 11192 25594 11248
rect 25650 11192 28000 11248
rect 25589 11190 28000 11192
rect 25589 11187 25655 11190
rect 27520 11160 28000 11190
rect 4521 11114 4587 11117
rect 5993 11114 6059 11117
rect 19333 11114 19399 11117
rect 23749 11114 23815 11117
rect 4521 11112 23815 11114
rect 4521 11056 4526 11112
rect 4582 11056 5998 11112
rect 6054 11056 19338 11112
rect 19394 11056 23754 11112
rect 23810 11056 23815 11112
rect 4521 11054 23815 11056
rect 4521 11051 4587 11054
rect 5993 11051 6059 11054
rect 19333 11051 19399 11054
rect 23749 11051 23815 11054
rect 23982 11054 24778 11114
rect 23982 10978 24042 11054
rect 17174 10918 24042 10978
rect 24718 10978 24778 11054
rect 25221 10978 25287 10981
rect 24718 10976 25287 10978
rect 24718 10920 25226 10976
rect 25282 10920 25287 10976
rect 24718 10918 25287 10920
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 12433 10842 12499 10845
rect 12617 10842 12683 10845
rect 13169 10842 13235 10845
rect 12433 10840 13235 10842
rect 12433 10784 12438 10840
rect 12494 10784 12622 10840
rect 12678 10784 13174 10840
rect 13230 10784 13235 10840
rect 12433 10782 13235 10784
rect 12433 10779 12499 10782
rect 12617 10779 12683 10782
rect 13169 10779 13235 10782
rect 0 10706 480 10736
rect 17174 10706 17234 10918
rect 25221 10915 25287 10918
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 23933 10842 23999 10845
rect 0 10646 17234 10706
rect 17358 10840 23999 10842
rect 17358 10784 23938 10840
rect 23994 10784 23999 10840
rect 17358 10782 23999 10784
rect 0 10616 480 10646
rect 12433 10570 12499 10573
rect 17358 10570 17418 10782
rect 23933 10779 23999 10782
rect 24577 10706 24643 10709
rect 27520 10706 28000 10736
rect 12433 10568 17418 10570
rect 12433 10512 12438 10568
rect 12494 10512 17418 10568
rect 12433 10510 17418 10512
rect 17496 10704 24643 10706
rect 17496 10648 24582 10704
rect 24638 10648 24643 10704
rect 17496 10646 24643 10648
rect 12433 10507 12499 10510
rect 17496 10434 17556 10646
rect 24577 10643 24643 10646
rect 24718 10646 28000 10706
rect 23473 10570 23539 10573
rect 24718 10570 24778 10646
rect 27520 10616 28000 10646
rect 23473 10568 24778 10570
rect 23473 10512 23478 10568
rect 23534 10512 24778 10568
rect 23473 10510 24778 10512
rect 23473 10507 23539 10510
rect 16806 10374 17556 10434
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 3693 10162 3759 10165
rect 13721 10162 13787 10165
rect 16806 10162 16866 10374
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 23790 10162 23796 10164
rect 3693 10160 16866 10162
rect 3693 10104 3698 10160
rect 3754 10104 13726 10160
rect 13782 10104 16866 10160
rect 3693 10102 16866 10104
rect 17174 10102 23796 10162
rect 3693 10099 3759 10102
rect 13721 10099 13787 10102
rect 0 10026 480 10056
rect 1301 10026 1367 10029
rect 0 10024 1367 10026
rect 0 9968 1306 10024
rect 1362 9968 1367 10024
rect 0 9966 1367 9968
rect 0 9936 480 9966
rect 1301 9963 1367 9966
rect 6177 10026 6243 10029
rect 17174 10026 17234 10102
rect 23790 10100 23796 10102
rect 23860 10100 23866 10164
rect 6177 10024 17234 10026
rect 6177 9968 6182 10024
rect 6238 9968 17234 10024
rect 6177 9966 17234 9968
rect 21541 10026 21607 10029
rect 27520 10026 28000 10056
rect 21541 10024 28000 10026
rect 21541 9968 21546 10024
rect 21602 9968 28000 10024
rect 21541 9966 28000 9968
rect 6177 9963 6243 9966
rect 21541 9963 21607 9966
rect 27520 9936 28000 9966
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 9673 9754 9739 9757
rect 12065 9754 12131 9757
rect 9673 9752 12131 9754
rect 9673 9696 9678 9752
rect 9734 9696 12070 9752
rect 12126 9696 12131 9752
rect 9673 9694 12131 9696
rect 9673 9691 9739 9694
rect 12065 9691 12131 9694
rect 12801 9618 12867 9621
rect 1350 9616 12867 9618
rect 1350 9560 12806 9616
rect 12862 9560 12867 9616
rect 1350 9558 12867 9560
rect 0 9482 480 9512
rect 1350 9482 1410 9558
rect 12801 9555 12867 9558
rect 14825 9618 14891 9621
rect 17769 9618 17835 9621
rect 14825 9616 17835 9618
rect 14825 9560 14830 9616
rect 14886 9560 17774 9616
rect 17830 9560 17835 9616
rect 14825 9558 17835 9560
rect 14825 9555 14891 9558
rect 17769 9555 17835 9558
rect 26233 9618 26299 9621
rect 26509 9618 26575 9621
rect 26233 9616 26575 9618
rect 26233 9560 26238 9616
rect 26294 9560 26514 9616
rect 26570 9560 26575 9616
rect 26233 9558 26575 9560
rect 26233 9555 26299 9558
rect 26509 9555 26575 9558
rect 0 9422 1410 9482
rect 1577 9482 1643 9485
rect 23606 9482 23612 9484
rect 1577 9480 23612 9482
rect 1577 9424 1582 9480
rect 1638 9424 23612 9480
rect 1577 9422 23612 9424
rect 0 9392 480 9422
rect 1577 9419 1643 9422
rect 23606 9420 23612 9422
rect 23676 9420 23682 9484
rect 23974 9420 23980 9484
rect 24044 9482 24050 9484
rect 27520 9482 28000 9512
rect 24044 9422 28000 9482
rect 24044 9420 24050 9422
rect 27520 9392 28000 9422
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 3877 9074 3943 9077
rect 13905 9074 13971 9077
rect 3877 9072 13971 9074
rect 3877 9016 3882 9072
rect 3938 9016 13910 9072
rect 13966 9016 13971 9072
rect 3877 9014 13971 9016
rect 3877 9011 3943 9014
rect 13905 9011 13971 9014
rect 22277 9074 22343 9077
rect 22277 9072 24962 9074
rect 22277 9016 22282 9072
rect 22338 9016 24962 9072
rect 22277 9014 24962 9016
rect 22277 9011 22343 9014
rect 13629 8938 13695 8941
rect 2454 8936 13695 8938
rect 2454 8880 13634 8936
rect 13690 8880 13695 8936
rect 2454 8878 13695 8880
rect 0 8802 480 8832
rect 2454 8802 2514 8878
rect 13629 8875 13695 8878
rect 16021 8938 16087 8941
rect 24669 8938 24735 8941
rect 16021 8936 24735 8938
rect 16021 8880 16026 8936
rect 16082 8880 24674 8936
rect 24730 8880 24735 8936
rect 16021 8878 24735 8880
rect 16021 8875 16087 8878
rect 24669 8875 24735 8878
rect 0 8742 2514 8802
rect 24902 8802 24962 9014
rect 27520 8802 28000 8832
rect 24902 8742 28000 8802
rect 0 8712 480 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 27520 8712 28000 8742
rect 24277 8671 24597 8672
rect 19149 8530 19215 8533
rect 19149 8528 24778 8530
rect 19149 8472 19154 8528
rect 19210 8472 24778 8528
rect 19149 8470 24778 8472
rect 19149 8467 19215 8470
rect 17953 8394 18019 8397
rect 23657 8394 23723 8397
rect 17953 8392 23723 8394
rect 17953 8336 17958 8392
rect 18014 8336 23662 8392
rect 23718 8336 23723 8392
rect 17953 8334 23723 8336
rect 17953 8331 18019 8334
rect 23657 8331 23723 8334
rect 0 8258 480 8288
rect 4061 8258 4127 8261
rect 0 8256 4127 8258
rect 0 8200 4066 8256
rect 4122 8200 4127 8256
rect 0 8198 4127 8200
rect 24718 8258 24778 8470
rect 27520 8258 28000 8288
rect 24718 8198 28000 8258
rect 0 8168 480 8198
rect 4061 8195 4127 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 27520 8168 28000 8198
rect 19610 8127 19930 8128
rect 14549 7850 14615 7853
rect 3190 7848 14615 7850
rect 3190 7792 14554 7848
rect 14610 7792 14615 7848
rect 3190 7790 14615 7792
rect 3190 7714 3250 7790
rect 14549 7787 14615 7790
rect 16205 7850 16271 7853
rect 23657 7850 23723 7853
rect 16205 7848 23723 7850
rect 16205 7792 16210 7848
rect 16266 7792 23662 7848
rect 23718 7792 23723 7848
rect 16205 7790 23723 7792
rect 16205 7787 16271 7790
rect 23657 7787 23723 7790
rect 2684 7654 3250 7714
rect 0 7578 480 7608
rect 2684 7578 2744 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 0 7518 2744 7578
rect 24761 7578 24827 7581
rect 27520 7578 28000 7608
rect 24761 7576 28000 7578
rect 24761 7520 24766 7576
rect 24822 7520 28000 7576
rect 24761 7518 28000 7520
rect 0 7488 480 7518
rect 24761 7515 24827 7518
rect 27520 7488 28000 7518
rect 4061 7442 4127 7445
rect 17953 7442 18019 7445
rect 4061 7440 18019 7442
rect 4061 7384 4066 7440
rect 4122 7384 17958 7440
rect 18014 7384 18019 7440
rect 4061 7382 18019 7384
rect 4061 7379 4127 7382
rect 17953 7379 18019 7382
rect 10277 7104 10597 7105
rect 0 7034 480 7064
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 3877 7034 3943 7037
rect 0 7032 3943 7034
rect 0 6976 3882 7032
rect 3938 6976 3943 7032
rect 0 6974 3943 6976
rect 0 6944 480 6974
rect 3877 6971 3943 6974
rect 23565 7034 23631 7037
rect 27520 7034 28000 7064
rect 23565 7032 28000 7034
rect 23565 6976 23570 7032
rect 23626 6976 28000 7032
rect 23565 6974 28000 6976
rect 23565 6971 23631 6974
rect 27520 6944 28000 6974
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 0 6354 480 6384
rect 3693 6354 3759 6357
rect 0 6352 3759 6354
rect 0 6296 3698 6352
rect 3754 6296 3759 6352
rect 0 6294 3759 6296
rect 0 6264 480 6294
rect 3693 6291 3759 6294
rect 23749 6354 23815 6357
rect 27520 6354 28000 6384
rect 23749 6352 28000 6354
rect 23749 6296 23754 6352
rect 23810 6296 28000 6352
rect 23749 6294 28000 6296
rect 23749 6291 23815 6294
rect 27520 6264 28000 6294
rect 23473 6082 23539 6085
rect 23473 6080 26250 6082
rect 23473 6024 23478 6080
rect 23534 6024 26250 6080
rect 23473 6022 26250 6024
rect 23473 6019 23539 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 0 5810 480 5840
rect 24025 5810 24091 5813
rect 0 5808 24091 5810
rect 0 5752 24030 5808
rect 24086 5752 24091 5808
rect 0 5750 24091 5752
rect 26190 5810 26250 6022
rect 27520 5810 28000 5840
rect 26190 5750 28000 5810
rect 0 5720 480 5750
rect 24025 5747 24091 5750
rect 27520 5720 28000 5750
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 0 5130 480 5160
rect 3969 5130 4035 5133
rect 0 5128 4035 5130
rect 0 5072 3974 5128
rect 4030 5072 4035 5128
rect 0 5070 4035 5072
rect 0 5040 480 5070
rect 3969 5067 4035 5070
rect 13537 5130 13603 5133
rect 23473 5130 23539 5133
rect 13537 5128 23539 5130
rect 13537 5072 13542 5128
rect 13598 5072 23478 5128
rect 23534 5072 23539 5128
rect 13537 5070 23539 5072
rect 13537 5067 13603 5070
rect 23473 5067 23539 5070
rect 24669 5130 24735 5133
rect 27520 5130 28000 5160
rect 24669 5128 28000 5130
rect 24669 5072 24674 5128
rect 24730 5072 28000 5128
rect 24669 5070 28000 5072
rect 24669 5067 24735 5070
rect 27520 5040 28000 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 0 4586 480 4616
rect 565 4586 631 4589
rect 0 4584 631 4586
rect 0 4528 570 4584
rect 626 4528 631 4584
rect 0 4526 631 4528
rect 0 4496 480 4526
rect 565 4523 631 4526
rect 17033 4586 17099 4589
rect 27520 4586 28000 4616
rect 17033 4584 28000 4586
rect 17033 4528 17038 4584
rect 17094 4528 28000 4584
rect 17033 4526 28000 4528
rect 17033 4523 17099 4526
rect 27520 4496 28000 4526
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 17953 4212 18019 4215
rect 17910 4210 18019 4212
rect 8201 4178 8267 4181
rect 17910 4178 17958 4210
rect 8201 4176 17958 4178
rect 8201 4120 8206 4176
rect 8262 4154 17958 4176
rect 18014 4154 18019 4210
rect 8262 4149 18019 4154
rect 8262 4120 17970 4149
rect 8201 4118 17970 4120
rect 8201 4115 8267 4118
rect 2773 4042 2839 4045
rect 9673 4042 9739 4045
rect 2773 4040 9739 4042
rect 2773 3984 2778 4040
rect 2834 3984 9678 4040
rect 9734 3984 9739 4040
rect 2773 3982 9739 3984
rect 2773 3979 2839 3982
rect 9673 3979 9739 3982
rect 0 3906 480 3936
rect 24577 3906 24643 3909
rect 27520 3906 28000 3936
rect 0 3846 4906 3906
rect 0 3816 480 3846
rect 4846 3498 4906 3846
rect 24577 3904 28000 3906
rect 24577 3848 24582 3904
rect 24638 3848 28000 3904
rect 24577 3846 28000 3848
rect 24577 3843 24643 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 27520 3816 28000 3846
rect 19610 3775 19930 3776
rect 14181 3770 14247 3773
rect 14181 3768 15762 3770
rect 14181 3712 14186 3768
rect 14242 3712 15762 3768
rect 14181 3710 15762 3712
rect 14181 3707 14247 3710
rect 9121 3634 9187 3637
rect 13905 3634 13971 3637
rect 9121 3632 13971 3634
rect 9121 3576 9126 3632
rect 9182 3576 13910 3632
rect 13966 3576 13971 3632
rect 9121 3574 13971 3576
rect 9121 3571 9187 3574
rect 13905 3571 13971 3574
rect 15561 3498 15627 3501
rect 4846 3496 15627 3498
rect 4846 3440 15566 3496
rect 15622 3440 15627 3496
rect 4846 3438 15627 3440
rect 15702 3498 15762 3710
rect 15702 3438 24962 3498
rect 15561 3435 15627 3438
rect 0 3362 480 3392
rect 24902 3362 24962 3438
rect 27520 3362 28000 3392
rect 0 3302 1226 3362
rect 24902 3302 28000 3362
rect 0 3272 480 3302
rect 1166 3226 1226 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 27520 3272 28000 3302
rect 24277 3231 24597 3232
rect 1945 3226 2011 3229
rect 1166 3224 2011 3226
rect 1166 3168 1950 3224
rect 2006 3168 2011 3224
rect 1166 3166 2011 3168
rect 1945 3163 2011 3166
rect 8293 2954 8359 2957
rect 12433 2954 12499 2957
rect 8293 2952 12499 2954
rect 8293 2896 8298 2952
rect 8354 2896 12438 2952
rect 12494 2896 12499 2952
rect 8293 2894 12499 2896
rect 8293 2891 8359 2894
rect 12433 2891 12499 2894
rect 19517 2954 19583 2957
rect 25129 2954 25195 2957
rect 19517 2952 25195 2954
rect 19517 2896 19522 2952
rect 19578 2896 25134 2952
rect 25190 2896 25195 2952
rect 19517 2894 25195 2896
rect 19517 2891 19583 2894
rect 25129 2891 25195 2894
rect 3141 2818 3207 2821
rect 1580 2816 3207 2818
rect 1580 2760 3146 2816
rect 3202 2760 3207 2816
rect 1580 2758 3207 2760
rect 0 2682 480 2712
rect 1580 2682 1640 2758
rect 3141 2755 3207 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 0 2622 1640 2682
rect 23657 2682 23723 2685
rect 27520 2682 28000 2712
rect 23657 2680 28000 2682
rect 23657 2624 23662 2680
rect 23718 2624 28000 2680
rect 23657 2622 28000 2624
rect 0 2592 480 2622
rect 23657 2619 23723 2622
rect 27520 2592 28000 2622
rect 23473 2410 23539 2413
rect 23473 2408 27538 2410
rect 23473 2352 23478 2408
rect 23534 2352 27538 2408
rect 23473 2350 27538 2352
rect 23473 2347 23539 2350
rect 5610 2208 5930 2209
rect 0 2138 480 2168
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 27478 2168 27538 2350
rect 3325 2138 3391 2141
rect 0 2136 3391 2138
rect 0 2080 3330 2136
rect 3386 2080 3391 2136
rect 0 2078 3391 2080
rect 27478 2078 28000 2168
rect 0 2048 480 2078
rect 3325 2075 3391 2078
rect 27520 2048 28000 2078
rect 0 1458 480 1488
rect 3693 1458 3759 1461
rect 0 1456 3759 1458
rect 0 1400 3698 1456
rect 3754 1400 3759 1456
rect 0 1398 3759 1400
rect 0 1368 480 1398
rect 3693 1395 3759 1398
rect 23933 1458 23999 1461
rect 27520 1458 28000 1488
rect 23933 1456 28000 1458
rect 23933 1400 23938 1456
rect 23994 1400 28000 1456
rect 23933 1398 28000 1400
rect 23933 1395 23999 1398
rect 27520 1368 28000 1398
rect 0 914 480 944
rect 933 914 999 917
rect 0 912 999 914
rect 0 856 938 912
rect 994 856 999 912
rect 0 854 999 856
rect 0 824 480 854
rect 933 851 999 854
rect 20345 914 20411 917
rect 27520 914 28000 944
rect 20345 912 28000 914
rect 20345 856 20350 912
rect 20406 856 28000 912
rect 20345 854 28000 856
rect 20345 851 20411 854
rect 27520 824 28000 854
rect 0 370 480 400
rect 1301 370 1367 373
rect 27520 370 28000 400
rect 0 368 1367 370
rect 0 312 1306 368
rect 1362 312 1367 368
rect 0 310 1367 312
rect 0 280 480 310
rect 1301 307 1367 310
rect 27478 280 28000 370
rect 13169 234 13235 237
rect 27478 234 27538 280
rect 13169 232 27538 234
rect 13169 176 13174 232
rect 13230 176 27538 232
rect 13169 174 27538 176
rect 13169 171 13235 174
rect 13445 98 13511 101
rect 20345 98 20411 101
rect 13445 96 20411 98
rect 13445 40 13450 96
rect 13506 40 20350 96
rect 20406 40 20411 96
rect 13445 38 20411 40
rect 13445 35 13511 38
rect 20345 35 20411 38
<< via3 >>
rect 9996 26012 10060 26076
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 8892 24712 8956 24716
rect 8892 24656 8906 24712
rect 8906 24656 8956 24712
rect 8892 24652 8956 24656
rect 21036 24652 21100 24716
rect 23612 24788 23676 24852
rect 23796 24652 23860 24716
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 9444 23428 9508 23492
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 14044 23292 14108 23356
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 5028 22748 5092 22812
rect 9996 22672 10060 22676
rect 9996 22616 10010 22672
rect 10010 22616 10060 22672
rect 9996 22612 10060 22616
rect 19012 22748 19076 22812
rect 7420 22340 7484 22404
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 14044 21932 14108 21996
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 23428 21312 23492 21316
rect 23428 21256 23478 21312
rect 23478 21256 23492 21312
rect 23428 21252 23492 21256
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 9628 19484 9692 19548
rect 7420 19408 7484 19412
rect 7420 19352 7434 19408
rect 7434 19352 7484 19408
rect 7420 19348 7484 19352
rect 24900 19212 24964 19276
rect 23980 19076 24044 19140
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10916 17308 10980 17372
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 24716 15948 24780 16012
rect 23244 15268 23308 15332
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 23428 14860 23492 14924
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 23244 13016 23308 13020
rect 23244 12960 23294 13016
rect 23294 12960 23308 13016
rect 23244 12956 23308 12960
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 24716 11188 24780 11252
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 23796 10100 23860 10164
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 23612 9420 23676 9484
rect 23980 9420 24044 9484
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 9995 26076 10061 26077
rect 9995 26012 9996 26076
rect 10060 26012 10061 26076
rect 9995 26011 10061 26012
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 8891 24652 8892 24702
rect 8956 24652 8957 24702
rect 8891 24651 8957 24652
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 9443 23492 9509 23493
rect 9443 23428 9444 23492
rect 9508 23428 9509 23492
rect 9443 23427 9509 23428
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 7419 22404 7485 22405
rect 7419 22340 7420 22404
rect 7484 22340 7485 22404
rect 7419 22339 7485 22340
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 7422 19413 7482 22339
rect 7419 19412 7485 19413
rect 7419 19348 7420 19412
rect 7484 19348 7485 19412
rect 9446 19410 9506 23427
rect 9998 22677 10058 26011
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 9995 22676 10061 22677
rect 9995 22612 9996 22676
rect 10060 22612 10061 22676
rect 9995 22611 10061 22612
rect 10277 22336 10597 23360
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14043 23356 14109 23357
rect 14043 23292 14044 23356
rect 14108 23292 14109 23356
rect 14043 23291 14109 23292
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 14046 21997 14106 23291
rect 14944 22880 15264 23904
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 23611 24852 23677 24853
rect 23611 24788 23612 24852
rect 23676 24788 23677 24852
rect 23611 24787 23677 24788
rect 21035 24652 21036 24702
rect 21100 24652 21101 24702
rect 21035 24651 21101 24652
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14043 21996 14109 21997
rect 14043 21932 14044 21996
rect 14108 21932 14109 21996
rect 14043 21931 14109 21932
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 9627 19548 9693 19549
rect 9627 19484 9628 19548
rect 9692 19484 9693 19548
rect 9627 19483 9693 19484
rect 9630 19410 9690 19483
rect 9446 19350 9690 19410
rect 7419 19347 7485 19348
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 23427 21316 23493 21317
rect 23427 21252 23428 21316
rect 23492 21252 23493 21316
rect 23427 21251 23493 21252
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 23243 15332 23309 15333
rect 23243 15268 23244 15332
rect 23308 15268 23309 15332
rect 23243 15267 23309 15268
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 23246 13021 23306 15267
rect 23430 14925 23490 21251
rect 23427 14924 23493 14925
rect 23427 14860 23428 14924
rect 23492 14860 23493 14924
rect 23427 14859 23493 14860
rect 23243 13020 23309 13021
rect 23243 12956 23244 13020
rect 23308 12956 23309 13020
rect 23243 12955 23309 12956
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 23614 9485 23674 24787
rect 23795 24716 23861 24717
rect 23795 24652 23796 24716
rect 23860 24652 23861 24716
rect 23795 24651 23861 24652
rect 23798 10165 23858 24651
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 23979 19140 24045 19141
rect 23979 19076 23980 19140
rect 24044 19076 24045 19140
rect 23979 19075 24045 19076
rect 23795 10164 23861 10165
rect 23795 10100 23796 10164
rect 23860 10100 23861 10164
rect 23795 10099 23861 10100
rect 23982 9485 24042 19075
rect 24277 18528 24597 19552
rect 24899 19276 24965 19277
rect 24899 19212 24900 19276
rect 24964 19212 24965 19276
rect 24899 19211 24965 19212
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24902 17458 24962 19211
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24715 16012 24781 16013
rect 24715 15948 24716 16012
rect 24780 15948 24781 16012
rect 24715 15947 24781 15948
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24718 11253 24778 15947
rect 24715 11252 24781 11253
rect 24715 11188 24716 11252
rect 24780 11188 24781 11252
rect 24715 11187 24781 11188
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 23611 9484 23677 9485
rect 23611 9420 23612 9484
rect 23676 9420 23677 9484
rect 23611 9419 23677 9420
rect 23979 9484 24045 9485
rect 23979 9420 23980 9484
rect 24044 9420 24045 9484
rect 23979 9419 24045 9420
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 8806 24716 9042 24938
rect 8806 24702 8892 24716
rect 8892 24702 8956 24716
rect 8956 24702 9042 24716
rect 4942 22812 5178 22898
rect 4942 22748 5028 22812
rect 5028 22748 5092 22812
rect 5092 22748 5178 22812
rect 4942 22662 5178 22748
rect 20950 24716 21186 24938
rect 20950 24702 21036 24716
rect 21036 24702 21100 24716
rect 21100 24702 21186 24716
rect 18926 22812 19162 22898
rect 18926 22748 19012 22812
rect 19012 22748 19076 22812
rect 19076 22748 19162 22812
rect 18926 22662 19162 22748
rect 10830 17372 11066 17458
rect 10830 17308 10916 17372
rect 10916 17308 10980 17372
rect 10980 17308 11066 17372
rect 10830 17222 11066 17308
rect 24814 17222 25050 17458
<< metal5 >>
rect 8764 24938 21228 24980
rect 8764 24702 8806 24938
rect 9042 24702 20950 24938
rect 21186 24702 21228 24938
rect 8764 24660 21228 24702
rect 4900 22898 19204 22940
rect 4900 22662 4942 22898
rect 5178 22662 18926 22898
rect 19162 22662 19204 22898
rect 4900 22620 19204 22662
rect 10788 17458 25092 17500
rect 10788 17222 10830 17458
rect 11066 17222 24814 17458
rect 25050 17222 25092 17458
rect 10788 17180 25092 17222
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1604681595
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1604681595
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__D tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604681595
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_144
timestamp 1604681595
transform 1 0 14352 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1604681595
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_152
timestamp 1604681595
transform 1 0 15088 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1604681595
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1604681595
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604681595
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1604681595
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1604681595
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1604681595
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1604681595
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1604681595
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _057_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1604681595
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1604681595
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1604681595
transform 1 0 25116 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__A
timestamp 1604681595
transform 1 0 25668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1604681595
transform 1 0 24380 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_265
timestamp 1604681595
transform 1 0 25484 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_269
timestamp 1604681595
transform 1 0 25852 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1604681595
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604681595
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1604681595
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1604681595
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1604681595
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1604681595
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1604681595
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1604681595
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1604681595
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1604681595
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1604681595
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1604681595
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604681595
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1604681595
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1604681595
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1604681595
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1604681595
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1604681595
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 24104 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1604681595
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_249
timestamp 1604681595
transform 1 0 24012 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_252
timestamp 1604681595
transform 1 0 24288 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_256
timestamp 1604681595
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_260
timestamp 1604681595
transform 1 0 25024 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_272
timestamp 1604681595
transform 1 0 26128 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_276
timestamp 1604681595
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1604681595
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1604681595
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1604681595
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1604681595
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1604681595
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1604681595
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 24104 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_239
timestamp 1604681595
transform 1 0 23092 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_247
timestamp 1604681595
transform 1 0 23828 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_259
timestamp 1604681595
transform 1 0 24932 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_271
timestamp 1604681595
transform 1 0 26036 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604681595
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1604681595
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1604681595
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1604681595
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1604681595
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1604681595
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1604681595
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604681595
transform 1 0 24012 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_251
timestamp 1604681595
transform 1 0 24196 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_263
timestamp 1604681595
transform 1 0 25300 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_275
timestamp 1604681595
transform 1 0 26404 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1604681595
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1604681595
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1604681595
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1604681595
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1604681595
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1604681595
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1604681595
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1604681595
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1604681595
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1604681595
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1604681595
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1604681595
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1604681595
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 24012 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_239
timestamp 1604681595
transform 1 0 23092 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_247
timestamp 1604681595
transform 1 0 23828 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1604681595
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1604681595
transform 1 0 24380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_265
timestamp 1604681595
transform 1 0 25484 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604681595
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1604681595
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_273
timestamp 1604681595
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1604681595
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1604681595
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1604681595
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1604681595
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1604681595
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1604681595
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1604681595
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1604681595
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604681595
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1604681595
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1604681595
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1604681595
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_110
timestamp 1604681595
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1604681595
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1604681595
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1604681595
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1604681595
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1604681595
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_220
timestamp 1604681595
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1604681595
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1604681595
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1604681595
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1604681595
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1604681595
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1604681595
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1604681595
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1604681595
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1604681595
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1604681595
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1604681595
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1604681595
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1604681595
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1604681595
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1604681595
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_98
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_110
timestamp 1604681595
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1604681595
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1604681595
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1604681595
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1604681595
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_249
timestamp 1604681595
transform 1 0 24012 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604681595
transform 1 0 24196 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_253
timestamp 1604681595
transform 1 0 24380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_265
timestamp 1604681595
transform 1 0 25484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604681595
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_7
timestamp 1604681595
transform 1 0 1748 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_19
timestamp 1604681595
transform 1 0 2852 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1604681595
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1604681595
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1604681595
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1604681595
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1604681595
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_143
timestamp 1604681595
transform 1 0 14260 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1604681595
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1604681595
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1604681595
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1604681595
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604681595
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1604681595
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1604681595
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_7
timestamp 1604681595
transform 1 0 1748 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604681595
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_19
timestamp 1604681595
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_12
timestamp 1604681595
transform 1 0 2208 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_11
timestamp 1604681595
transform 1 0 2116 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 2484 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_17
timestamp 1604681595
transform 1 0 2668 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_29
timestamp 1604681595
transform 1 0 3772 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_41
timestamp 1604681595
transform 1 0 4876 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_23
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_53
timestamp 1604681595
transform 1 0 5980 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1604681595
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1604681595
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1604681595
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1604681595
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1604681595
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_110
timestamp 1604681595
transform 1 0 11224 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_117
timestamp 1604681595
transform 1 0 11868 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1604681595
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12604 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 12052 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12236 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1604681595
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_134
timestamp 1604681595
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_130
timestamp 1604681595
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_131
timestamp 1604681595
transform 1 0 13156 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_127
timestamp 1604681595
transform 1 0 12788 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12972 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_143
timestamp 1604681595
transform 1 0 14260 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_138
timestamp 1604681595
transform 1 0 13800 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13616 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 13892 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 14076 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1604681595
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_148
timestamp 1604681595
transform 1 0 14720 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1604681595
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_150
timestamp 1604681595
transform 1 0 14904 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14904 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14536 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_160
timestamp 1604681595
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_163
timestamp 1604681595
transform 1 0 16100 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_164
timestamp 1604681595
transform 1 0 16192 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_176
timestamp 1604681595
transform 1 0 17296 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1604681595
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_175
timestamp 1604681595
transform 1 0 17204 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_187
timestamp 1604681595
transform 1 0 18308 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1604681595
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_199
timestamp 1604681595
transform 1 0 19412 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_220
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_211
timestamp 1604681595
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_232
timestamp 1604681595
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1604681595
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 24564 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604681595
transform 1 0 24564 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_253
timestamp 1604681595
transform 1 0 24380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1604681595
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1604681595
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_251
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_259
timestamp 1604681595
transform 1 0 24932 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_271
timestamp 1604681595
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 2392 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 2024 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 1656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_8
timestamp 1604681595
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_12
timestamp 1604681595
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_23
timestamp 1604681595
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1604681595
transform 1 0 3588 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_31
timestamp 1604681595
transform 1 0 3956 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_34
timestamp 1604681595
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_38
timestamp 1604681595
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_42
timestamp 1604681595
transform 1 0 4968 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_54
timestamp 1604681595
transform 1 0 6072 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1604681595
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1604681595
transform 1 0 12512 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12052 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_110
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_114
timestamp 1604681595
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_117
timestamp 1604681595
transform 1 0 11868 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1604681595
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 13524 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_133
timestamp 1604681595
transform 1 0 13340 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_137
timestamp 1604681595
transform 1 0 13708 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_141
timestamp 1604681595
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_145
timestamp 1604681595
transform 1 0 14444 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14536 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_155
timestamp 1604681595
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_159
timestamp 1604681595
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_163
timestamp 1604681595
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_167
timestamp 1604681595
transform 1 0 16468 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_171
timestamp 1604681595
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1604681595
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_220
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604681595
transform 1 0 23828 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_232
timestamp 1604681595
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_249
timestamp 1604681595
transform 1 0 24012 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 24564 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604681595
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604681595
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_259
timestamp 1604681595
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_263
timestamp 1604681595
transform 1 0 25300 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_275
timestamp 1604681595
transform 1 0 26404 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1604681595
transform 1 0 2024 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1604681595
transform 1 0 1748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_19
timestamp 1604681595
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_41
timestamp 1604681595
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 5428 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_45
timestamp 1604681595
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_49
timestamp 1604681595
transform 1 0 5612 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_61
timestamp 1604681595
transform 1 0 6716 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_73
timestamp 1604681595
transform 1 0 7820 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_85
timestamp 1604681595
transform 1 0 8924 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1604681595
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12052 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_107
timestamp 1604681595
transform 1 0 10948 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_111
timestamp 1604681595
transform 1 0 11316 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_128
timestamp 1604681595
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_132
timestamp 1604681595
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_145
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 14904 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_149
timestamp 1604681595
transform 1 0 14812 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1604681595
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1604681595
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _055_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 16836 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_167
timestamp 1604681595
transform 1 0 16468 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_174
timestamp 1604681595
transform 1 0 17112 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_186
timestamp 1604681595
transform 1 0 18216 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_198
timestamp 1604681595
transform 1 0 19320 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1604681595
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_227
timestamp 1604681595
transform 1 0 21988 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1604681595
transform 1 0 22356 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 23460 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24012 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604681595
transform 1 0 22816 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_234
timestamp 1604681595
transform 1 0 22632 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_238
timestamp 1604681595
transform 1 0 23000 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_242
timestamp 1604681595
transform 1 0 23368 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_247
timestamp 1604681595
transform 1 0 23828 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 24564 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_251
timestamp 1604681595
transform 1 0 24196 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_259
timestamp 1604681595
transform 1 0 24932 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_271
timestamp 1604681595
transform 1 0 26036 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 1656 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_8
timestamp 1604681595
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_12
timestamp 1604681595
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 3956 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 3772 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_23
timestamp 1604681595
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1604681595
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_40
timestamp 1604681595
transform 1 0 4784 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 5520 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_45
timestamp 1604681595
transform 1 0 5244 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1604681595
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 8556 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_67
timestamp 1604681595
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_71
timestamp 1604681595
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_75
timestamp 1604681595
transform 1 0 8004 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_84
timestamp 1604681595
transform 1 0 8832 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_96
timestamp 1604681595
transform 1 0 9936 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_101
timestamp 1604681595
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1604681595
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604681595
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_132
timestamp 1604681595
transform 1 0 13248 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_137
timestamp 1604681595
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_141
timestamp 1604681595
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_145
timestamp 1604681595
transform 1 0 14444 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 14904 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_159
timestamp 1604681595
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_163
timestamp 1604681595
transform 1 0 16100 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_170
timestamp 1604681595
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1604681595
transform 1 0 16468 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_174
timestamp 1604681595
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_178
timestamp 1604681595
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_182
timestamp 1604681595
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17664 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1604681595
transform 1 0 19596 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 18676 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_188
timestamp 1604681595
transform 1 0 18400 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1604681595
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_197
timestamp 1604681595
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_204
timestamp 1604681595
transform 1 0 19872 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 21436 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604681595
transform 1 0 21896 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_216
timestamp 1604681595
transform 1 0 20976 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_220
timestamp 1604681595
transform 1 0 21344 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_224
timestamp 1604681595
transform 1 0 21712 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_228
timestamp 1604681595
transform 1 0 22080 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 22448 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23920 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604681595
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1604681595
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1604681595
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 25484 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_257
timestamp 1604681595
transform 1 0 24748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_261
timestamp 1604681595
transform 1 0 25116 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604681595
transform 1 0 26036 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_273
timestamp 1604681595
transform 1 0 26220 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2024 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1604681595
transform 1 0 1748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_19
timestamp 1604681595
transform 1 0 2852 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 3036 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_36
timestamp 1604681595
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 4232 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_40
timestamp 1604681595
transform 1 0 4784 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5060 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6072 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 6440 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_52
timestamp 1604681595
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_56
timestamp 1604681595
transform 1 0 6256 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_60
timestamp 1604681595
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7084 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8096 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8464 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_64
timestamp 1604681595
transform 1 0 6992 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_74
timestamp 1604681595
transform 1 0 7912 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_78
timestamp 1604681595
transform 1 0 8280 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_82
timestamp 1604681595
transform 1 0 8648 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 10028 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_100
timestamp 1604681595
transform 1 0 10304 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_104
timestamp 1604681595
transform 1 0 10672 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11040 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_107
timestamp 1604681595
transform 1 0 10948 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13524 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 13340 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_127
timestamp 1604681595
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_131
timestamp 1604681595
transform 1 0 13156 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_144
timestamp 1604681595
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 14904 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_148
timestamp 1604681595
transform 1 0 14720 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1604681595
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16836 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 18216 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17848 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1604681595
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_180
timestamp 1604681595
transform 1 0 17664 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_184
timestamp 1604681595
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18676 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19780 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20148 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_188
timestamp 1604681595
transform 1 0 18400 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_200
timestamp 1604681595
transform 1 0 19504 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_205
timestamp 1604681595
transform 1 0 19964 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 21436 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_209
timestamp 1604681595
transform 1 0 20332 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1604681595
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_225
timestamp 1604681595
transform 1 0 21804 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 22540 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23644 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 23460 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_237
timestamp 1604681595
transform 1 0 22908 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_264
timestamp 1604681595
transform 1 0 25392 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_272
timestamp 1604681595
transform 1 0 26128 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_6
timestamp 1604681595
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1748 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_10
timestamp 1604681595
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_16
timestamp 1604681595
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1604681595
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_20
timestamp 1604681595
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 3128 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 3312 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_38
timestamp 1604681595
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_40
timestamp 1604681595
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_37
timestamp 1604681595
transform 1 0 4508 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_33
timestamp 1604681595
transform 1 0 4140 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 4784 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_46
timestamp 1604681595
transform 1 0 5336 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_42
timestamp 1604681595
transform 1 0 4968 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 5520 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_81
timestamp 1604681595
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_67
timestamp 1604681595
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_71
timestamp 1604681595
transform 1 0 7636 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_85
timestamp 1604681595
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9292 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_88
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_92
timestamp 1604681595
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1604681595
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_97
timestamp 1604681595
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 9752 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 9936 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 10212 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_122
timestamp 1604681595
transform 1 0 12328 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_118
timestamp 1604681595
transform 1 0 11960 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_125
timestamp 1604681595
transform 1 0 12604 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 14352 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12696 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_19_132
timestamp 1604681595
transform 1 0 13248 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14720 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_163
timestamp 1604681595
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_146
timestamp 1604681595
transform 1 0 14536 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_150
timestamp 1604681595
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_173
timestamp 1604681595
transform 1 0 17020 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_174
timestamp 1604681595
transform 1 0 17112 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_167
timestamp 1604681595
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1604681595
transform 1 0 16836 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17480 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1604681595
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_177
timestamp 1604681595
transform 1 0 17388 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_180
timestamp 1604681595
transform 1 0 17664 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17848 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1604681595
transform 1 0 18216 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18032 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1604681595
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_193
timestamp 1604681595
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_195
timestamp 1604681595
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_204
timestamp 1604681595
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_199
timestamp 1604681595
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19780 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 19596 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_208
timestamp 1604681595
transform 1 0 20240 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_212
timestamp 1604681595
transform 1 0 20608 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_218
timestamp 1604681595
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604681595
transform 1 0 20976 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 20976 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_220
timestamp 1604681595
transform 1 0 21344 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 21528 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 21344 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_224
timestamp 1604681595
transform 1 0 21712 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_224
timestamp 1604681595
transform 1 0 21712 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604681595
transform 1 0 21896 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604681595
transform 1 0 22080 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 22080 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_236
timestamp 1604681595
transform 1 0 22816 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_232
timestamp 1604681595
transform 1 0 22448 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1604681595
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_230
timestamp 1604681595
transform 1 0 22264 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 22632 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604681595
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 22448 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_247
timestamp 1604681595
transform 1 0 23828 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_244
timestamp 1604681595
transform 1 0 23552 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_240
timestamp 1604681595
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 23644 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24104 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23828 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 25392 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24840 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_266
timestamp 1604681595
transform 1 0 25576 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_256
timestamp 1604681595
transform 1 0 24656 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_260
timestamp 1604681595
transform 1 0 25024 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_267
timestamp 1604681595
transform 1 0 25668 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_274
timestamp 1604681595
transform 1 0 26312 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 2392 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_9
timestamp 1604681595
transform 1 0 1932 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 4876 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4692 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_33
timestamp 1604681595
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_37
timestamp 1604681595
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8740 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604681595
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1604681595
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_75
timestamp 1604681595
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_79
timestamp 1604681595
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_102
timestamp 1604681595
transform 1 0 10488 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_110
timestamp 1604681595
transform 1 0 11224 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_106
timestamp 1604681595
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 11316 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 13984 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_136
timestamp 1604681595
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 14996 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_149
timestamp 1604681595
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_153
timestamp 1604681595
transform 1 0 15180 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_158
timestamp 1604681595
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_162
timestamp 1604681595
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1604681595
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_179
timestamp 1604681595
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_203
timestamp 1604681595
transform 1 0 19780 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_208
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_2_
timestamp 1604681595
transform 1 0 20976 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 20792 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 20424 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 21988 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_212
timestamp 1604681595
transform 1 0 20608 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1604681595
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_229
timestamp 1604681595
transform 1 0 22172 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 22540 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 22356 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_236
timestamp 1604681595
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604681595
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604681595
transform 1 0 25576 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1604681595
transform 1 0 25392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_268
timestamp 1604681595
transform 1 0 25760 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_276
timestamp 1604681595
transform 1 0 26496 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1472 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_41
timestamp 1604681595
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 5612 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 5428 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_45
timestamp 1604681595
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 8096 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7912 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_68
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_72
timestamp 1604681595
transform 1 0 7728 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_80
timestamp 1604681595
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1604681595
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12144 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 11960 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 11592 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_112
timestamp 1604681595
transform 1 0 11408 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_116
timestamp 1604681595
transform 1 0 11776 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13156 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 13524 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_129
timestamp 1604681595
transform 1 0 12972 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_133
timestamp 1604681595
transform 1 0 13340 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_137
timestamp 1604681595
transform 1 0 13708 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 15732 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 15548 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1604681595
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_162
timestamp 1604681595
transform 1 0 16008 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18308 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16744 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_168
timestamp 1604681595
transform 1 0 16560 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_179
timestamp 1604681595
transform 1 0 17572 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_183
timestamp 1604681595
transform 1 0 17940 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_186
timestamp 1604681595
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1604681595
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_3_
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 21896 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_210
timestamp 1604681595
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_224
timestamp 1604681595
transform 1 0 21712 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_228
timestamp 1604681595
transform 1 0 22080 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24012 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_1_
timestamp 1604681595
transform 1 0 22448 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23644 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604681595
transform 1 0 22264 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_241
timestamp 1604681595
transform 1 0 23276 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_247
timestamp 1604681595
transform 1 0 23828 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 25300 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24748 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604681595
transform 1 0 25116 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_255
timestamp 1604681595
transform 1 0 24564 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_259
timestamp 1604681595
transform 1 0 24932 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_267
timestamp 1604681595
transform 1 0 25668 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 1564 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_14
timestamp 1604681595
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_18
timestamp 1604681595
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3128 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_23_41
timestamp 1604681595
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_45
timestamp 1604681595
transform 1 0 5244 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 5060 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5428 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 5612 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7820 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604681595
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_65
timestamp 1604681595
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_69
timestamp 1604681595
transform 1 0 7452 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_92
timestamp 1604681595
transform 1 0 9568 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_96
timestamp 1604681595
transform 1 0 9936 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_99
timestamp 1604681595
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_112
timestamp 1604681595
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_116
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 14168 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_132
timestamp 1604681595
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_136
timestamp 1604681595
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_140
timestamp 1604681595
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_144
timestamp 1604681595
transform 1 0 14352 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 14812 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 14628 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 17664 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16744 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_168
timestamp 1604681595
transform 1 0 16560 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_172
timestamp 1604681595
transform 1 0 16928 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_176
timestamp 1604681595
transform 1 0 17296 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_179
timestamp 1604681595
transform 1 0 17572 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 19780 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19596 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_193
timestamp 1604681595
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_197
timestamp 1604681595
transform 1 0 19228 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604681595
transform 1 0 22080 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1604681595
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_226
timestamp 1604681595
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 22264 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_234
timestamp 1604681595
transform 1 0 22632 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1604681595
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 25208 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604681595
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_254
timestamp 1604681595
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_258
timestamp 1604681595
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_266
timestamp 1604681595
transform 1 0 25576 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_270
timestamp 1604681595
transform 1 0 25944 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_276
timestamp 1604681595
transform 1 0 26496 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 1748 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_16
timestamp 1604681595
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_20
timestamp 1604681595
transform 1 0 2944 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_24
timestamp 1604681595
transform 1 0 3312 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3128 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_28
timestamp 1604681595
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3496 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_35
timestamp 1604681595
transform 1 0 4324 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_39
timestamp 1604681595
transform 1 0 4692 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 4508 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 6624 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 5060 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6440 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6072 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_52
timestamp 1604681595
transform 1 0 5888 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_56
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7912 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_64
timestamp 1604681595
transform 1 0 6992 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_70
timestamp 1604681595
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_83
timestamp 1604681595
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 10304 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9936 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_87
timestamp 1604681595
transform 1 0 9108 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_98
timestamp 1604681595
transform 1 0 10120 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_121
timestamp 1604681595
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_125
timestamp 1604681595
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13984 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1604681595
transform 1 0 13800 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_142
timestamp 1604681595
transform 1 0 14168 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15732 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 14904 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 15456 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 14536 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_148
timestamp 1604681595
transform 1 0 14720 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1604681595
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_158
timestamp 1604681595
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18216 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17664 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_178
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_182
timestamp 1604681595
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20148 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_205
timestamp 1604681595
transform 1 0 19964 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21988 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_209
timestamp 1604681595
transform 1 0 20332 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_224
timestamp 1604681595
transform 1 0 21712 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_229
timestamp 1604681595
transform 1 0 22172 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 22448 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23552 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 23000 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_236
timestamp 1604681595
transform 1 0 22816 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_240
timestamp 1604681595
transform 1 0 23184 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 25116 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 24564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 24932 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1604681595
transform 1 0 24380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_257
timestamp 1604681595
transform 1 0 24748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_265
timestamp 1604681595
transform 1 0 25484 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_273
timestamp 1604681595
transform 1 0 26220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2668 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_9
timestamp 1604681595
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_13
timestamp 1604681595
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3680 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_26
timestamp 1604681595
transform 1 0 3496 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_30
timestamp 1604681595
transform 1 0 3864 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_34
timestamp 1604681595
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_38
timestamp 1604681595
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4968 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_51
timestamp 1604681595
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_55
timestamp 1604681595
transform 1 0 6164 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8004 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7544 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_66
timestamp 1604681595
transform 1 0 7176 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_72
timestamp 1604681595
transform 1 0 7728 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604681595
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_94
timestamp 1604681595
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_102
timestamp 1604681595
transform 1 0 10488 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14352 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_142
timestamp 1604681595
transform 1 0 14168 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 14904 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 15916 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_146
timestamp 1604681595
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_159
timestamp 1604681595
transform 1 0 15732 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_163
timestamp 1604681595
transform 1 0 16100 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16652 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_167
timestamp 1604681595
transform 1 0 16468 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1604681595
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_179
timestamp 1604681595
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19872 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_193
timestamp 1604681595
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_197
timestamp 1604681595
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_201
timestamp 1604681595
transform 1 0 19596 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 21712 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21528 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 21160 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_213
timestamp 1604681595
transform 1 0 20700 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_217
timestamp 1604681595
transform 1 0 21068 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_220
timestamp 1604681595
transform 1 0 21344 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1604681595
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1604681595
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_264
timestamp 1604681595
transform 1 0 25392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_268
timestamp 1604681595
transform 1 0 25760 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_276
timestamp 1604681595
transform 1 0 26496 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1656 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_19
timestamp 1604681595
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1932 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_28
timestamp 1604681595
transform 1 0 3680 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_34
timestamp 1604681595
transform 1 0 4232 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_35
timestamp 1604681595
transform 1 0 4324 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_39
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_39
timestamp 1604681595
transform 1 0 4692 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 4508 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 4876 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5060 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_3_
timestamp 1604681595
transform 1 0 5060 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_62
timestamp 1604681595
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_52
timestamp 1604681595
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_56
timestamp 1604681595
transform 1 0 6256 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_68
timestamp 1604681595
transform 1 0 7360 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_66
timestamp 1604681595
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7544 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_73
timestamp 1604681595
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_83
timestamp 1604681595
transform 1 0 8740 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_79
timestamp 1604681595
transform 1 0 8372 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 8556 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 8188 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_26_87
timestamp 1604681595
transform 1 0 9108 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8924 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_100
timestamp 1604681595
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_96
timestamp 1604681595
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_102
timestamp 1604681595
transform 1 0 10488 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_97
timestamp 1604681595
transform 1 0 10028 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10304 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10488 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10672 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10672 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 11132 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_106
timestamp 1604681595
transform 1 0 10856 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_113
timestamp 1604681595
transform 1 0 11500 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_118
timestamp 1604681595
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_132
timestamp 1604681595
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_132
timestamp 1604681595
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_128
timestamp 1604681595
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 13064 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_136
timestamp 1604681595
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_145
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 13984 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_26_149
timestamp 1604681595
transform 1 0 14812 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 14628 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_163
timestamp 1604681595
transform 1 0 16100 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_159
timestamp 1604681595
transform 1 0 15732 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1604681595
transform 1 0 16100 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16284 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 15916 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16468 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16836 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_169
timestamp 1604681595
transform 1 0 16652 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17204 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_173
timestamp 1604681595
transform 1 0 17020 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_173
timestamp 1604681595
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_177
timestamp 1604681595
transform 1 0 17388 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16468 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 17388 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_186
timestamp 1604681595
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_26_190
timestamp 1604681595
transform 1 0 18584 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 18768 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18952 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_27_207
timestamp 1604681595
transform 1 0 20148 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_203
timestamp 1604681595
transform 1 0 19780 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_207
timestamp 1604681595
transform 1 0 20148 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_203
timestamp 1604681595
transform 1 0 19780 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19964 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 19964 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_211
timestamp 1604681595
transform 1 0 20516 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 21068 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20424 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_223
timestamp 1604681595
transform 1 0 21620 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_219
timestamp 1604681595
transform 1 0 21252 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21436 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 21712 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 20608 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_236
timestamp 1604681595
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_231
timestamp 1604681595
transform 1 0 22356 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 22632 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_240
timestamp 1604681595
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_247
timestamp 1604681595
transform 1 0 23828 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_243
timestamp 1604681595
transform 1 0 23460 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 24012 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23644 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 23736 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25668 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25208 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_260
timestamp 1604681595
transform 1 0 25024 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_264
timestamp 1604681595
transform 1 0 25392 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_265
timestamp 1604681595
transform 1 0 25484 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_269
timestamp 1604681595
transform 1 0 25852 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 26036 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_272
timestamp 1604681595
transform 1 0 26128 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_273
timestamp 1604681595
transform 1 0 26220 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 1748 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 2760 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_16
timestamp 1604681595
transform 1 0 2576 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_20
timestamp 1604681595
transform 1 0 2944 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3128 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3496 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_24
timestamp 1604681595
transform 1 0 3312 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_28
timestamp 1604681595
transform 1 0 3680 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 6532 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 5980 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6348 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_51
timestamp 1604681595
transform 1 0 5796 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_55
timestamp 1604681595
transform 1 0 6164 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_63
timestamp 1604681595
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_67
timestamp 1604681595
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_71
timestamp 1604681595
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10396 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_88
timestamp 1604681595
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_99
timestamp 1604681595
transform 1 0 10212 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_103
timestamp 1604681595
transform 1 0 10580 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10948 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13432 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12880 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_126
timestamp 1604681595
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_130
timestamp 1604681595
transform 1 0 13064 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_143
timestamp 1604681595
transform 1 0 14260 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_147
timestamp 1604681595
transform 1 0 14628 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_163
timestamp 1604681595
transform 1 0 16100 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 17020 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16836 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 16468 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_169
timestamp 1604681595
transform 1 0 16652 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 18952 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19320 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_192
timestamp 1604681595
transform 1 0 18768 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_196
timestamp 1604681595
transform 1 0 19136 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_206
timestamp 1604681595
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_210
timestamp 1604681595
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23368 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22816 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 23184 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_234
timestamp 1604681595
transform 1 0 22632 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_238
timestamp 1604681595
transform 1 0 23000 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24932 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 24380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 24748 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_251
timestamp 1604681595
transform 1 0 24196 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_255
timestamp 1604681595
transform 1 0 24564 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_265
timestamp 1604681595
transform 1 0 25484 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_273
timestamp 1604681595
transform 1 0 26220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 2116 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_7
timestamp 1604681595
transform 1 0 1748 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4692 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_30
timestamp 1604681595
transform 1 0 3864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_35
timestamp 1604681595
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5704 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6072 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_48
timestamp 1604681595
transform 1 0 5520 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_52
timestamp 1604681595
transform 1 0 5888 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_56
timestamp 1604681595
transform 1 0 6256 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8280 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_68
timestamp 1604681595
transform 1 0 7360 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_73
timestamp 1604681595
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_77
timestamp 1604681595
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_97
timestamp 1604681595
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_101
timestamp 1604681595
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604681595
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14352 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_142
timestamp 1604681595
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 14904 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_146
timestamp 1604681595
transform 1 0 14536 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_169
timestamp 1604681595
transform 1 0 16652 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_174
timestamp 1604681595
transform 1 0 17112 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_179
timestamp 1604681595
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19872 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19688 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_193
timestamp 1604681595
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_197
timestamp 1604681595
transform 1 0 19228 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_201
timestamp 1604681595
transform 1 0 19596 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21436 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21252 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_213
timestamp 1604681595
transform 1 0 20700 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_217
timestamp 1604681595
transform 1 0 21068 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604681595
transform 1 0 22540 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_230
timestamp 1604681595
transform 1 0 22264 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_235
timestamp 1604681595
transform 1 0 22724 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_240
timestamp 1604681595
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_264
timestamp 1604681595
transform 1 0 25392 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_276
timestamp 1604681595
transform 1 0 26496 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1604681595
transform 1 0 2024 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 1840 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp 1604681595
transform 1 0 1748 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_19
timestamp 1604681595
transform 1 0 2852 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_23
timestamp 1604681595
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3036 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_36
timestamp 1604681595
transform 1 0 4416 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 4232 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4692 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6624 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_58
timestamp 1604681595
transform 1 0 6440 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_62
timestamp 1604681595
transform 1 0 6808 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_67
timestamp 1604681595
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_71
timestamp 1604681595
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10304 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10120 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 9292 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_84
timestamp 1604681595
transform 1 0 8832 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_88
timestamp 1604681595
transform 1 0 9200 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1604681595
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_97
timestamp 1604681595
transform 1 0 10028 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_119
timestamp 1604681595
transform 1 0 12052 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_125
timestamp 1604681595
transform 1 0 12604 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12788 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 14076 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1604681595
transform 1 0 13616 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_140
timestamp 1604681595
transform 1 0 13984 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_143
timestamp 1604681595
transform 1 0 14260 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 16284 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_147
timestamp 1604681595
transform 1 0 14628 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_163
timestamp 1604681595
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16928 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18032 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16652 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_167
timestamp 1604681595
transform 1 0 16468 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_171
timestamp 1604681595
transform 1 0 16836 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_181
timestamp 1604681595
transform 1 0 17756 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_186
timestamp 1604681595
transform 1 0 18216 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18492 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 20056 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19872 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19504 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_198
timestamp 1604681595
transform 1 0 19320 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_202
timestamp 1604681595
transform 1 0 19688 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 21896 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_209
timestamp 1604681595
transform 1 0 20332 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_224
timestamp 1604681595
transform 1 0 21712 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_228
timestamp 1604681595
transform 1 0 22080 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 22540 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23644 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22264 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 23092 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 23460 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_232
timestamp 1604681595
transform 1 0 22448 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_237
timestamp 1604681595
transform 1 0 22908 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_241
timestamp 1604681595
transform 1 0 23276 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 25576 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_264
timestamp 1604681595
transform 1 0 25392 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_268
timestamp 1604681595
transform 1 0 25760 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_274
timestamp 1604681595
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1840 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 1656 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_17
timestamp 1604681595
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4232 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4048 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_21
timestamp 1604681595
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_25
timestamp 1604681595
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_29
timestamp 1604681595
transform 1 0 3772 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_53
timestamp 1604681595
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604681595
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8556 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_71
timestamp 1604681595
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_75
timestamp 1604681595
transform 1 0 8004 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9936 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_90
timestamp 1604681595
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_94
timestamp 1604681595
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_107
timestamp 1604681595
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_111
timestamp 1604681595
transform 1 0 11316 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_115
timestamp 1604681595
transform 1 0 11684 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604681595
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12880 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 14444 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 12696 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 14260 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_137
timestamp 1604681595
transform 1 0 13708 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_141
timestamp 1604681595
transform 1 0 14076 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 16008 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15456 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 15824 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_154
timestamp 1604681595
transform 1 0 15272 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_158
timestamp 1604681595
transform 1 0 15640 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_171
timestamp 1604681595
transform 1 0 16836 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_175
timestamp 1604681595
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_179
timestamp 1604681595
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19596 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_193
timestamp 1604681595
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_197
timestamp 1604681595
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_207
timestamp 1604681595
transform 1 0 20148 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 21068 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_211
timestamp 1604681595
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_236
timestamp 1604681595
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_240
timestamp 1604681595
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 25208 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 24656 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 25024 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_254
timestamp 1604681595
transform 1 0 24472 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_258
timestamp 1604681595
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_266
timestamp 1604681595
transform 1 0 25576 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_270
timestamp 1604681595
transform 1 0 25944 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 26128 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_274
timestamp 1604681595
transform 1 0 26312 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1604681595
transform 1 0 1840 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 1656 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2852 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_17
timestamp 1604681595
transform 1 0 2668 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4600 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4232 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_21
timestamp 1604681595
transform 1 0 3036 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_25
timestamp 1604681595
transform 1 0 3404 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_36
timestamp 1604681595
transform 1 0 4416 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6532 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_57
timestamp 1604681595
transform 1 0 6348 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_61
timestamp 1604681595
transform 1 0 6716 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7084 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8096 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8556 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6900 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_74
timestamp 1604681595
transform 1 0 7912 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_78
timestamp 1604681595
transform 1 0 8280 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_83
timestamp 1604681595
transform 1 0 8740 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 10212 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 9292 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8924 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10028 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_87
timestamp 1604681595
transform 1 0 9108 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_118
timestamp 1604681595
transform 1 0 11960 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_122
timestamp 1604681595
transform 1 0 12328 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_125
timestamp 1604681595
transform 1 0 12604 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12696 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 13708 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_135
timestamp 1604681595
transform 1 0 13524 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_139
timestamp 1604681595
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_143
timestamp 1604681595
transform 1 0 14260 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 14904 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 16284 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_147
timestamp 1604681595
transform 1 0 14628 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_163
timestamp 1604681595
transform 1 0 16100 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18308 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16836 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16652 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 17572 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_167
timestamp 1604681595
transform 1 0 16468 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_177
timestamp 1604681595
transform 1 0 17388 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_181
timestamp 1604681595
transform 1 0 17756 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_186
timestamp 1604681595
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_206
timestamp 1604681595
transform 1 0 20056 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 21896 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 21620 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_210
timestamp 1604681595
transform 1 0 20424 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_218
timestamp 1604681595
transform 1 0 21160 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_222
timestamp 1604681595
transform 1 0 21528 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_225
timestamp 1604681595
transform 1 0 21804 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23828 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_245
timestamp 1604681595
transform 1 0 23644 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_249
timestamp 1604681595
transform 1 0 24012 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24380 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 24196 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604681595
transform 1 0 25392 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_262
timestamp 1604681595
transform 1 0 25208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_266
timestamp 1604681595
transform 1 0 25576 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_274
timestamp 1604681595
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2024 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 1840 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_8
timestamp 1604681595
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_7
timestamp 1604681595
transform 1 0 1748 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2024 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_19
timestamp 1604681595
transform 1 0 2852 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 2208 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_23
timestamp 1604681595
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3036 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_35
timestamp 1604681595
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_31
timestamp 1604681595
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4140 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4508 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_41
timestamp 1604681595
transform 1 0 4876 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_49
timestamp 1604681595
transform 1 0 5612 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_45
timestamp 1604681595
transform 1 0 5244 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_48
timestamp 1604681595
transform 1 0 5520 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5796 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 5428 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5060 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5704 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_53
timestamp 1604681595
transform 1 0 5980 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_52
timestamp 1604681595
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6072 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 6256 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6072 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_72
timestamp 1604681595
transform 1 0 7728 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_63
timestamp 1604681595
transform 1 0 6900 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_69
timestamp 1604681595
transform 1 0 7452 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_65
timestamp 1604681595
transform 1 0 7084 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7176 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 7268 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7544 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 7820 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_88
timestamp 1604681595
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_84
timestamp 1604681595
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_92
timestamp 1604681595
transform 1 0 9568 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604681595
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_97
timestamp 1604681595
transform 1 0 10028 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_99
timestamp 1604681595
transform 1 0 10212 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_96
timestamp 1604681595
transform 1 0 9936 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10028 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9844 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10396 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10580 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10212 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_33_116
timestamp 1604681595
transform 1 0 11776 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_112
timestamp 1604681595
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_122
timestamp 1604681595
transform 1 0 12328 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_118
timestamp 1604681595
transform 1 0 11960 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_125
timestamp 1604681595
transform 1 0 12604 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_135
timestamp 1604681595
transform 1 0 13524 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_133
timestamp 1604681595
transform 1 0 13340 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_129
timestamp 1604681595
transform 1 0 12972 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 13524 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 13156 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12696 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_143
timestamp 1604681595
transform 1 0 14260 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_139
timestamp 1604681595
transform 1 0 13892 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13708 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13708 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_34_151
timestamp 1604681595
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_147
timestamp 1604681595
transform 1 0 14628 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_156
timestamp 1604681595
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 14812 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_160
timestamp 1604681595
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16008 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16192 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_34_177
timestamp 1604681595
transform 1 0 17388 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_173
timestamp 1604681595
transform 1 0 17020 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_177
timestamp 1604681595
transform 1 0 17388 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_173
timestamp 1604681595
transform 1 0 17020 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17204 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17572 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 17756 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_33_192
timestamp 1604681595
transform 1 0 18768 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_188
timestamp 1604681595
transform 1 0 18400 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18952 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604681595
transform 1 0 18584 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_208
timestamp 1604681595
transform 1 0 20240 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_204
timestamp 1604681595
transform 1 0 19872 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_200
timestamp 1604681595
transform 1 0 19504 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20056 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1604681595
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1604681595
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21068 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 20424 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_225
timestamp 1604681595
transform 1 0 21804 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_221
timestamp 1604681595
transform 1 0 21436 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_219
timestamp 1604681595
transform 1 0 21252 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 21620 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 21436 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_3_
timestamp 1604681595
transform 1 0 21620 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 22172 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_238
timestamp 1604681595
transform 1 0 23000 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_236
timestamp 1604681595
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_232
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22632 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_242
timestamp 1604681595
transform 1 0 23368 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_240
timestamp 1604681595
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23552 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23184 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23736 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 25208 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604681595
transform 1 0 25760 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 24656 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25024 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_254
timestamp 1604681595
transform 1 0 24472 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_258
timestamp 1604681595
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_266
timestamp 1604681595
transform 1 0 25576 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_270
timestamp 1604681595
transform 1 0 25944 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_265
timestamp 1604681595
transform 1 0 25484 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_274
timestamp 1604681595
transform 1 0 26312 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_273
timestamp 1604681595
transform 1 0 26220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 2300 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_9
timestamp 1604681595
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4876 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4232 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_32
timestamp 1604681595
transform 1 0 4048 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_36
timestamp 1604681595
transform 1 0 4416 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_40
timestamp 1604681595
transform 1 0 4784 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5060 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_52
timestamp 1604681595
transform 1 0 5888 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1604681595
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7544 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A
timestamp 1604681595
transform 1 0 7360 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_66
timestamp 1604681595
transform 1 0 7176 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10488 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10028 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_89
timestamp 1604681595
transform 1 0 9292 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_95
timestamp 1604681595
transform 1 0 9844 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_99
timestamp 1604681595
transform 1 0 10212 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_111
timestamp 1604681595
transform 1 0 11316 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_115
timestamp 1604681595
transform 1 0 11684 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 14352 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 14168 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 13800 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_132
timestamp 1604681595
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_136
timestamp 1604681595
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_140
timestamp 1604681595
transform 1 0 13984 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16284 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_163
timestamp 1604681595
transform 1 0 16100 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604681595
transform 1 0 16836 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1604681595
transform 1 0 16652 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_167
timestamp 1604681595
transform 1 0 16468 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_175
timestamp 1604681595
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_179
timestamp 1604681595
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19044 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 20240 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19412 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19780 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_193
timestamp 1604681595
transform 1 0 18860 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_197
timestamp 1604681595
transform 1 0 19228 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_201
timestamp 1604681595
transform 1 0 19596 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_205
timestamp 1604681595
transform 1 0 19964 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_1_
timestamp 1604681595
transform 1 0 20424 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21804 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 21436 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_219
timestamp 1604681595
transform 1 0 21252 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_223
timestamp 1604681595
transform 1 0 21620 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1604681595
transform 1 0 22816 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1604681595
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 24656 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25024 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_254
timestamp 1604681595
transform 1 0 24472 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_258
timestamp 1604681595
transform 1 0 24840 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_268
timestamp 1604681595
transform 1 0 25760 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 26312 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_272
timestamp 1604681595
transform 1 0 26128 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_276
timestamp 1604681595
transform 1 0 26496 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 2208 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 1840 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_6
timestamp 1604681595
transform 1 0 1656 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_10
timestamp 1604681595
transform 1 0 2024 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_23
timestamp 1604681595
transform 1 0 3220 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1604681595
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6532 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5980 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 6348 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_51
timestamp 1604681595
transform 1 0 5796 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_55
timestamp 1604681595
transform 1 0 6164 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1604681595
transform 1 0 8096 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7544 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7912 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8648 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_68
timestamp 1604681595
transform 1 0 7360 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_72
timestamp 1604681595
transform 1 0 7728 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_80
timestamp 1604681595
transform 1 0 8464 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_84
timestamp 1604681595
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_88
timestamp 1604681595
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_102
timestamp 1604681595
transform 1 0 10488 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 11224 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12328 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12144 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_106
timestamp 1604681595
transform 1 0 10856 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_114
timestamp 1604681595
transform 1 0 11592 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_118
timestamp 1604681595
transform 1 0 11960 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13432 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_131
timestamp 1604681595
transform 1 0 13156 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_136
timestamp 1604681595
transform 1 0 13616 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_145
timestamp 1604681595
transform 1 0 14444 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15732 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14904 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 15456 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_149
timestamp 1604681595
transform 1 0 14812 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_152
timestamp 1604681595
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_154
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_158
timestamp 1604681595
transform 1 0 15640 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18216 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18032 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17664 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_178
timestamp 1604681595
transform 1 0 17480 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_182
timestamp 1604681595
transform 1 0 17848 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 19780 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19320 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_195
timestamp 1604681595
transform 1 0 19044 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_200
timestamp 1604681595
transform 1 0 19504 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_206
timestamp 1604681595
transform 1 0 20056 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20424 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_212
timestamp 1604681595
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23736 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22816 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 23184 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 23552 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_234
timestamp 1604681595
transform 1 0 22632 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_238
timestamp 1604681595
transform 1 0 23000 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_242
timestamp 1604681595
transform 1 0 23368 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_265
timestamp 1604681595
transform 1 0 25484 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_273
timestamp 1604681595
transform 1 0 26220 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2116 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2484 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_9
timestamp 1604681595
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_13
timestamp 1604681595
transform 1 0 2300 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_17
timestamp 1604681595
transform 1 0 2668 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 3588 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3404 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4600 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 3036 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_23
timestamp 1604681595
transform 1 0 3220 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_36
timestamp 1604681595
transform 1 0 4416 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_40
timestamp 1604681595
transform 1 0 4784 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_53
timestamp 1604681595
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1604681595
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6900 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_37_82
timestamp 1604681595
transform 1 0 8648 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9476 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9108 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10672 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_86
timestamp 1604681595
transform 1 0 9016 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_89
timestamp 1604681595
transform 1 0 9292 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_102
timestamp 1604681595
transform 1 0 10488 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604681595
transform 1 0 11224 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11040 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1604681595
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_106
timestamp 1604681595
transform 1 0 10856 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_114
timestamp 1604681595
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_118
timestamp 1604681595
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14352 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_142
timestamp 1604681595
transform 1 0 14168 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14904 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14720 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 15916 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 16284 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_146
timestamp 1604681595
transform 1 0 14536 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_159
timestamp 1604681595
transform 1 0 15732 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_163
timestamp 1604681595
transform 1 0 16100 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16652 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_167
timestamp 1604681595
transform 1 0 16468 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_175
timestamp 1604681595
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_179
timestamp 1604681595
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 19320 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19136 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18768 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_190
timestamp 1604681595
transform 1 0 18584 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_194
timestamp 1604681595
transform 1 0 18952 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21804 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21436 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_217
timestamp 1604681595
transform 1 0 21068 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_223
timestamp 1604681595
transform 1 0 21620 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_236
timestamp 1604681595
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_240
timestamp 1604681595
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25576 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 25944 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_264
timestamp 1604681595
transform 1 0 25392 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_268
timestamp 1604681595
transform 1 0 25760 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26312 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_272
timestamp 1604681595
transform 1 0 26128 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_276
timestamp 1604681595
transform 1 0 26496 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1748 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604681595
transform 1 0 1564 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604681595
transform 1 0 2852 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_13
timestamp 1604681595
transform 1 0 2300 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4508 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 4876 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1604681595
transform 1 0 3036 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1604681595
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_35
timestamp 1604681595
transform 1 0 4324 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_39
timestamp 1604681595
transform 1 0 4692 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5060 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_38_62
timestamp 1604681595
transform 1 0 6808 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7544 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6992 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7360 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8556 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_66
timestamp 1604681595
transform 1 0 7176 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_79
timestamp 1604681595
transform 1 0 8372 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_83
timestamp 1604681595
transform 1 0 8740 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10396 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604681595
transform 1 0 8924 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_87
timestamp 1604681595
transform 1 0 9108 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_99
timestamp 1604681595
transform 1 0 10212 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_103
timestamp 1604681595
transform 1 0 10580 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10948 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13432 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 12880 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14444 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_126
timestamp 1604681595
transform 1 0 12696 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_130
timestamp 1604681595
transform 1 0 13064 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_143
timestamp 1604681595
transform 1 0 14260 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14904 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_147
timestamp 1604681595
transform 1 0 14628 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_152
timestamp 1604681595
transform 1 0 15088 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17940 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17756 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17204 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_173
timestamp 1604681595
transform 1 0 17020 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_177
timestamp 1604681595
transform 1 0 17388 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18952 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_189
timestamp 1604681595
transform 1 0 18492 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_193
timestamp 1604681595
transform 1 0 18860 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_196
timestamp 1604681595
transform 1 0 19136 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_206
timestamp 1604681595
transform 1 0 20056 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_215
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_213
timestamp 1604681595
transform 1 0 20700 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_210
timestamp 1604681595
transform 1 0 20424 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20516 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21068 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_223
timestamp 1604681595
transform 1 0 21620 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_219
timestamp 1604681595
transform 1 0 21252 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21436 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 21804 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 23736 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 24104 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_244
timestamp 1604681595
transform 1 0 23552 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_248
timestamp 1604681595
transform 1 0 23920 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24288 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25300 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_261
timestamp 1604681595
transform 1 0 25116 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_265
timestamp 1604681595
transform 1 0 25484 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_273
timestamp 1604681595
transform 1 0 26220 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_7
timestamp 1604681595
transform 1 0 1748 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1932 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_11
timestamp 1604681595
transform 1 0 2116 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_17
timestamp 1604681595
transform 1 0 2668 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_11
timestamp 1604681595
transform 1 0 2116 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 2852 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_19
timestamp 1604681595
transform 1 0 2852 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_30
timestamp 1604681595
transform 1 0 3864 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_27
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_23
timestamp 1604681595
transform 1 0 3220 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3680 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_40
timestamp 1604681595
transform 1 0 4784 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_36
timestamp 1604681595
transform 1 0 4416 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_34
timestamp 1604681595
transform 1 0 4232 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4600 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1604681595
transform 1 0 4048 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4416 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_48
timestamp 1604681595
transform 1 0 5520 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_49
timestamp 1604681595
transform 1 0 5612 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_45
timestamp 1604681595
transform 1 0 5244 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 5428 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 5796 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1604681595
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_53
timestamp 1604681595
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 5796 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 8464 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8372 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7728 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8188 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_71
timestamp 1604681595
transform 1 0 7636 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_75
timestamp 1604681595
transform 1 0 8004 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_70
timestamp 1604681595
transform 1 0 7544 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_74
timestamp 1604681595
transform 1 0 7912 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_84
timestamp 1604681595
transform 1 0 8832 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_92
timestamp 1604681595
transform 1 0 9568 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_88
timestamp 1604681595
transform 1 0 9200 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9660 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_102
timestamp 1604681595
transform 1 0 10488 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_99
timestamp 1604681595
transform 1 0 10212 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_95
timestamp 1604681595
transform 1 0 9844 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10028 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10396 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_110
timestamp 1604681595
transform 1 0 11224 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_106
timestamp 1604681595
transform 1 0 10856 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_114
timestamp 1604681595
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1604681595
transform 1 0 11224 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11040 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11592 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11408 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_125
timestamp 1604681595
transform 1 0 12604 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1604681595
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11776 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1604681595
transform 1 0 13340 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 12788 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1604681595
transform 1 0 13156 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_142
timestamp 1604681595
transform 1 0 14168 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_129
timestamp 1604681595
transform 1 0 12972 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_142
timestamp 1604681595
transform 1 0 14168 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 14720 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_146
timestamp 1604681595
transform 1 0 14536 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_150
timestamp 1604681595
transform 1 0 14904 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_146
timestamp 1604681595
transform 1 0 14536 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_149
timestamp 1604681595
transform 1 0 14812 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 15088 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1604681595
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_154
timestamp 1604681595
transform 1 0 15272 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15364 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_162
timestamp 1604681595
transform 1 0 16008 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_158
timestamp 1604681595
transform 1 0 15640 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_164
timestamp 1604681595
transform 1 0 16192 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16192 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15824 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_166
timestamp 1604681595
transform 1 0 16376 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16376 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_175
timestamp 1604681595
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_168
timestamp 1604681595
transform 1 0 16560 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16744 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 16928 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_186
timestamp 1604681595
transform 1 0 18216 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_179
timestamp 1604681595
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 16468 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_40_190
timestamp 1604681595
transform 1 0 18584 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18768 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18400 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18952 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_40_207
timestamp 1604681595
transform 1 0 20148 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_203
timestamp 1604681595
transform 1 0 19780 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_207
timestamp 1604681595
transform 1 0 20148 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_203
timestamp 1604681595
transform 1 0 19780 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19964 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19964 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_213
timestamp 1604681595
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20516 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 20332 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20516 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_228
timestamp 1604681595
transform 1 0 22080 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_224
timestamp 1604681595
transform 1 0 21712 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_224
timestamp 1604681595
transform 1 0 21712 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_220
timestamp 1604681595
transform 1 0 21344 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 21896 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 22080 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21528 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_236
timestamp 1604681595
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 22264 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22264 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l3_in_0_
timestamp 1604681595
transform 1 0 22448 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_40_247
timestamp 1604681595
transform 1 0 23828 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_241
timestamp 1604681595
transform 1 0 23276 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_240
timestamp 1604681595
transform 1 0 23184 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23644 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 24564 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 25208 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604681595
transform 1 0 24656 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604681595
transform 1 0 25760 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_254
timestamp 1604681595
transform 1 0 24472 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_258
timestamp 1604681595
transform 1 0 24840 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_266
timestamp 1604681595
transform 1 0 25576 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_270
timestamp 1604681595
transform 1 0 25944 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_259
timestamp 1604681595
transform 1 0 24932 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_276
timestamp 1604681595
transform 1 0 26496 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1604681595
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1604681595
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604681595
transform 1 0 2300 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_7
timestamp 1604681595
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_11
timestamp 1604681595
transform 1 0 2116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_19
timestamp 1604681595
transform 1 0 2852 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1604681595
transform 1 0 4692 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1604681595
transform 1 0 3036 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1604681595
transform 1 0 4140 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1604681595
transform 1 0 4508 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1604681595
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_23
timestamp 1604681595
transform 1 0 3220 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_31
timestamp 1604681595
transform 1 0 3956 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_35
timestamp 1604681595
transform 1 0 4324 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_43
timestamp 1604681595
transform 1 0 5060 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1604681595
transform 1 0 5244 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_47
timestamp 1604681595
transform 1 0 5428 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5796 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_53
timestamp 1604681595
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1604681595
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8464 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6900 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 8280 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_72
timestamp 1604681595
transform 1 0 7728 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_76
timestamp 1604681595
transform 1 0 8096 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604681595
transform 1 0 10028 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9476 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604681595
transform 1 0 10488 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_89
timestamp 1604681595
transform 1 0 9292 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_93
timestamp 1604681595
transform 1 0 9660 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_100
timestamp 1604681595
transform 1 0 10304 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_104
timestamp 1604681595
transform 1 0 10672 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604681595
transform 1 0 12512 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604681595
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10856 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_114
timestamp 1604681595
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1604681595
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13616 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 13432 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13064 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_128
timestamp 1604681595
transform 1 0 12880 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_132
timestamp 1604681595
transform 1 0 13248 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_145
timestamp 1604681595
transform 1 0 14444 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15180 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 14996 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16192 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14628 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_149
timestamp 1604681595
transform 1 0 14812 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_162
timestamp 1604681595
transform 1 0 16008 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1604681595
transform 1 0 16376 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_175
timestamp 1604681595
transform 1 0 17204 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_170
timestamp 1604681595
transform 1 0 16744 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16560 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1604681595
transform 1 0 16836 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_184
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_179
timestamp 1604681595
transform 1 0 17572 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18216 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19780 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19596 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19228 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_195
timestamp 1604681595
transform 1 0 19044 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_199
timestamp 1604681595
transform 1 0 19412 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21344 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604681595
transform 1 0 20792 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21160 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_212
timestamp 1604681595
transform 1 0 20608 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_216
timestamp 1604681595
transform 1 0 20976 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_229
timestamp 1604681595
transform 1 0 22172 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22356 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_233
timestamp 1604681595
transform 1 0 22540 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_241
timestamp 1604681595
transform 1 0 23276 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 24564 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604681595
transform 1 0 25116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604681595
transform 1 0 24380 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_259
timestamp 1604681595
transform 1 0 24932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_263
timestamp 1604681595
transform 1 0 25300 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_275
timestamp 1604681595
transform 1 0 26404 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_7
timestamp 1604681595
transform 1 0 1748 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_19
timestamp 1604681595
transform 1 0 2852 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1604681595
transform 1 0 4692 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_36
timestamp 1604681595
transform 1 0 4416 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_41
timestamp 1604681595
transform 1 0 4876 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6624 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_48
timestamp 1604681595
transform 1 0 5520 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604681595
transform 1 0 8648 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7084 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 8464 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_74
timestamp 1604681595
transform 1 0 7912 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604681595
transform 1 0 10304 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 1604681595
transform 1 0 8924 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_94
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_104
timestamp 1604681595
transform 1 0 10672 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 11408 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_116
timestamp 1604681595
transform 1 0 11776 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604681595
transform 1 0 14260 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 13616 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13984 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_134
timestamp 1604681595
transform 1 0 13432 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1604681595
transform 1 0 13800 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_142
timestamp 1604681595
transform 1 0 14168 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15548 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_147
timestamp 1604681595
transform 1 0 14628 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_151
timestamp 1604681595
transform 1 0 14996 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_156
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_166
timestamp 1604681595
transform 1 0 16376 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_170
timestamp 1604681595
transform 1 0 16744 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 16560 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1604681595
transform 1 0 16928 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604681595
transform 1 0 17112 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_182
timestamp 1604681595
transform 1 0 17848 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_178
timestamp 1604681595
transform 1 0 17480 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17664 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18032 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 19964 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19780 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19320 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_196
timestamp 1604681595
transform 1 0 19136 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_200
timestamp 1604681595
transform 1 0 19504 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 21896 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21344 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21712 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_209
timestamp 1604681595
transform 1 0 20332 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_222
timestamp 1604681595
transform 1 0 21528 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_232
timestamp 1604681595
transform 1 0 22448 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_244
timestamp 1604681595
transform 1 0 23552 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 24564 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_259
timestamp 1604681595
transform 1 0 24932 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_271
timestamp 1604681595
transform 1 0 26036 0 -1 25568
box -38 -48 590 592
<< labels >>
rlabel metal2 s 19522 0 19578 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 27066 27520 27122 28000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 25134 0 25190 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 27618 27520 27674 28000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 8298 0 8354 480 6 ccff_head
port 4 nsew default input
rlabel metal2 s 13910 0 13966 480 6 ccff_tail
port 5 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_in[0]
port 6 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[10]
port 7 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_left_in[11]
port 8 nsew default input
rlabel metal3 s 0 11160 480 11280 6 chanx_left_in[12]
port 9 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[13]
port 10 nsew default input
rlabel metal3 s 0 12384 480 12504 6 chanx_left_in[14]
port 11 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_in[15]
port 12 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_in[16]
port 13 nsew default input
rlabel metal3 s 0 14288 480 14408 6 chanx_left_in[17]
port 14 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_left_in[18]
port 15 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[19]
port 16 nsew default input
rlabel metal3 s 0 4496 480 4616 6 chanx_left_in[1]
port 17 nsew default input
rlabel metal3 s 0 5040 480 5160 6 chanx_left_in[2]
port 18 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[3]
port 19 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_left_in[4]
port 20 nsew default input
rlabel metal3 s 0 6944 480 7064 6 chanx_left_in[5]
port 21 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[6]
port 22 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[7]
port 23 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[8]
port 24 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[9]
port 25 nsew default input
rlabel metal3 s 0 16056 480 16176 6 chanx_left_out[0]
port 26 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 chanx_left_out[10]
port 27 nsew default tristate
rlabel metal3 s 0 22720 480 22840 6 chanx_left_out[11]
port 28 nsew default tristate
rlabel metal3 s 0 23400 480 23520 6 chanx_left_out[12]
port 29 nsew default tristate
rlabel metal3 s 0 23944 480 24064 6 chanx_left_out[13]
port 30 nsew default tristate
rlabel metal3 s 0 24624 480 24744 6 chanx_left_out[14]
port 31 nsew default tristate
rlabel metal3 s 0 25168 480 25288 6 chanx_left_out[15]
port 32 nsew default tristate
rlabel metal3 s 0 25848 480 25968 6 chanx_left_out[16]
port 33 nsew default tristate
rlabel metal3 s 0 26392 480 26512 6 chanx_left_out[17]
port 34 nsew default tristate
rlabel metal3 s 0 27072 480 27192 6 chanx_left_out[18]
port 35 nsew default tristate
rlabel metal3 s 0 27616 480 27736 6 chanx_left_out[19]
port 36 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[1]
port 37 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[2]
port 38 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[3]
port 39 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 chanx_left_out[4]
port 40 nsew default tristate
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[5]
port 41 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[6]
port 42 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[7]
port 43 nsew default tristate
rlabel metal3 s 0 20952 480 21072 6 chanx_left_out[8]
port 44 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[9]
port 45 nsew default tristate
rlabel metal3 s 27520 3816 28000 3936 6 chanx_right_in[0]
port 46 nsew default input
rlabel metal3 s 27520 9936 28000 10056 6 chanx_right_in[10]
port 47 nsew default input
rlabel metal3 s 27520 10616 28000 10736 6 chanx_right_in[11]
port 48 nsew default input
rlabel metal3 s 27520 11160 28000 11280 6 chanx_right_in[12]
port 49 nsew default input
rlabel metal3 s 27520 11840 28000 11960 6 chanx_right_in[13]
port 50 nsew default input
rlabel metal3 s 27520 12384 28000 12504 6 chanx_right_in[14]
port 51 nsew default input
rlabel metal3 s 27520 13064 28000 13184 6 chanx_right_in[15]
port 52 nsew default input
rlabel metal3 s 27520 13608 28000 13728 6 chanx_right_in[16]
port 53 nsew default input
rlabel metal3 s 27520 14288 28000 14408 6 chanx_right_in[17]
port 54 nsew default input
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_in[18]
port 55 nsew default input
rlabel metal3 s 27520 15376 28000 15496 6 chanx_right_in[19]
port 56 nsew default input
rlabel metal3 s 27520 4496 28000 4616 6 chanx_right_in[1]
port 57 nsew default input
rlabel metal3 s 27520 5040 28000 5160 6 chanx_right_in[2]
port 58 nsew default input
rlabel metal3 s 27520 5720 28000 5840 6 chanx_right_in[3]
port 59 nsew default input
rlabel metal3 s 27520 6264 28000 6384 6 chanx_right_in[4]
port 60 nsew default input
rlabel metal3 s 27520 6944 28000 7064 6 chanx_right_in[5]
port 61 nsew default input
rlabel metal3 s 27520 7488 28000 7608 6 chanx_right_in[6]
port 62 nsew default input
rlabel metal3 s 27520 8168 28000 8288 6 chanx_right_in[7]
port 63 nsew default input
rlabel metal3 s 27520 8712 28000 8832 6 chanx_right_in[8]
port 64 nsew default input
rlabel metal3 s 27520 9392 28000 9512 6 chanx_right_in[9]
port 65 nsew default input
rlabel metal3 s 27520 16056 28000 16176 6 chanx_right_out[0]
port 66 nsew default tristate
rlabel metal3 s 27520 22176 28000 22296 6 chanx_right_out[10]
port 67 nsew default tristate
rlabel metal3 s 27520 22720 28000 22840 6 chanx_right_out[11]
port 68 nsew default tristate
rlabel metal3 s 27520 23400 28000 23520 6 chanx_right_out[12]
port 69 nsew default tristate
rlabel metal3 s 27520 23944 28000 24064 6 chanx_right_out[13]
port 70 nsew default tristate
rlabel metal3 s 27520 24624 28000 24744 6 chanx_right_out[14]
port 71 nsew default tristate
rlabel metal3 s 27520 25168 28000 25288 6 chanx_right_out[15]
port 72 nsew default tristate
rlabel metal3 s 27520 25848 28000 25968 6 chanx_right_out[16]
port 73 nsew default tristate
rlabel metal3 s 27520 26392 28000 26512 6 chanx_right_out[17]
port 74 nsew default tristate
rlabel metal3 s 27520 27072 28000 27192 6 chanx_right_out[18]
port 75 nsew default tristate
rlabel metal3 s 27520 27616 28000 27736 6 chanx_right_out[19]
port 76 nsew default tristate
rlabel metal3 s 27520 16600 28000 16720 6 chanx_right_out[1]
port 77 nsew default tristate
rlabel metal3 s 27520 17280 28000 17400 6 chanx_right_out[2]
port 78 nsew default tristate
rlabel metal3 s 27520 17824 28000 17944 6 chanx_right_out[3]
port 79 nsew default tristate
rlabel metal3 s 27520 18504 28000 18624 6 chanx_right_out[4]
port 80 nsew default tristate
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_out[5]
port 81 nsew default tristate
rlabel metal3 s 27520 19728 28000 19848 6 chanx_right_out[6]
port 82 nsew default tristate
rlabel metal3 s 27520 20272 28000 20392 6 chanx_right_out[7]
port 83 nsew default tristate
rlabel metal3 s 27520 20952 28000 21072 6 chanx_right_out[8]
port 84 nsew default tristate
rlabel metal3 s 27520 21496 28000 21616 6 chanx_right_out[9]
port 85 nsew default tristate
rlabel metal2 s 4710 27520 4766 28000 6 chany_top_in[0]
port 86 nsew default input
rlabel metal2 s 10322 27520 10378 28000 6 chany_top_in[10]
port 87 nsew default input
rlabel metal2 s 10874 27520 10930 28000 6 chany_top_in[11]
port 88 nsew default input
rlabel metal2 s 11426 27520 11482 28000 6 chany_top_in[12]
port 89 nsew default input
rlabel metal2 s 11978 27520 12034 28000 6 chany_top_in[13]
port 90 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 chany_top_in[14]
port 91 nsew default input
rlabel metal2 s 13082 27520 13138 28000 6 chany_top_in[15]
port 92 nsew default input
rlabel metal2 s 13634 27520 13690 28000 6 chany_top_in[16]
port 93 nsew default input
rlabel metal2 s 14278 27520 14334 28000 6 chany_top_in[17]
port 94 nsew default input
rlabel metal2 s 14830 27520 14886 28000 6 chany_top_in[18]
port 95 nsew default input
rlabel metal2 s 15382 27520 15438 28000 6 chany_top_in[19]
port 96 nsew default input
rlabel metal2 s 5262 27520 5318 28000 6 chany_top_in[1]
port 97 nsew default input
rlabel metal2 s 5814 27520 5870 28000 6 chany_top_in[2]
port 98 nsew default input
rlabel metal2 s 6366 27520 6422 28000 6 chany_top_in[3]
port 99 nsew default input
rlabel metal2 s 6918 27520 6974 28000 6 chany_top_in[4]
port 100 nsew default input
rlabel metal2 s 7562 27520 7618 28000 6 chany_top_in[5]
port 101 nsew default input
rlabel metal2 s 8114 27520 8170 28000 6 chany_top_in[6]
port 102 nsew default input
rlabel metal2 s 8666 27520 8722 28000 6 chany_top_in[7]
port 103 nsew default input
rlabel metal2 s 9218 27520 9274 28000 6 chany_top_in[8]
port 104 nsew default input
rlabel metal2 s 9770 27520 9826 28000 6 chany_top_in[9]
port 105 nsew default input
rlabel metal2 s 15934 27520 15990 28000 6 chany_top_out[0]
port 106 nsew default tristate
rlabel metal2 s 21546 27520 21602 28000 6 chany_top_out[10]
port 107 nsew default tristate
rlabel metal2 s 22098 27520 22154 28000 6 chany_top_out[11]
port 108 nsew default tristate
rlabel metal2 s 22650 27520 22706 28000 6 chany_top_out[12]
port 109 nsew default tristate
rlabel metal2 s 23202 27520 23258 28000 6 chany_top_out[13]
port 110 nsew default tristate
rlabel metal2 s 23754 27520 23810 28000 6 chany_top_out[14]
port 111 nsew default tristate
rlabel metal2 s 24306 27520 24362 28000 6 chany_top_out[15]
port 112 nsew default tristate
rlabel metal2 s 24858 27520 24914 28000 6 chany_top_out[16]
port 113 nsew default tristate
rlabel metal2 s 25410 27520 25466 28000 6 chany_top_out[17]
port 114 nsew default tristate
rlabel metal2 s 25962 27520 26018 28000 6 chany_top_out[18]
port 115 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[19]
port 116 nsew default tristate
rlabel metal2 s 16486 27520 16542 28000 6 chany_top_out[1]
port 117 nsew default tristate
rlabel metal2 s 17038 27520 17094 28000 6 chany_top_out[2]
port 118 nsew default tristate
rlabel metal2 s 17590 27520 17646 28000 6 chany_top_out[3]
port 119 nsew default tristate
rlabel metal2 s 18142 27520 18198 28000 6 chany_top_out[4]
port 120 nsew default tristate
rlabel metal2 s 18694 27520 18750 28000 6 chany_top_out[5]
port 121 nsew default tristate
rlabel metal2 s 19246 27520 19302 28000 6 chany_top_out[6]
port 122 nsew default tristate
rlabel metal2 s 19798 27520 19854 28000 6 chany_top_out[7]
port 123 nsew default tristate
rlabel metal2 s 20350 27520 20406 28000 6 chany_top_out[8]
port 124 nsew default tristate
rlabel metal2 s 20902 27520 20958 28000 6 chany_top_out[9]
port 125 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 left_bottom_grid_pin_11_
port 126 nsew default input
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_1_
port 127 nsew default input
rlabel metal3 s 0 824 480 944 6 left_bottom_grid_pin_3_
port 128 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_5_
port 129 nsew default input
rlabel metal3 s 0 2048 480 2168 6 left_bottom_grid_pin_7_
port 130 nsew default input
rlabel metal3 s 0 2592 480 2712 6 left_bottom_grid_pin_9_
port 131 nsew default input
rlabel metal2 s 2778 0 2834 480 6 prog_clk
port 132 nsew default input
rlabel metal3 s 27520 3272 28000 3392 6 right_bottom_grid_pin_11_
port 133 nsew default input
rlabel metal3 s 27520 280 28000 400 6 right_bottom_grid_pin_1_
port 134 nsew default input
rlabel metal3 s 27520 824 28000 944 6 right_bottom_grid_pin_3_
port 135 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 right_bottom_grid_pin_5_
port 136 nsew default input
rlabel metal3 s 27520 2048 28000 2168 6 right_bottom_grid_pin_7_
port 137 nsew default input
rlabel metal3 s 27520 2592 28000 2712 6 right_bottom_grid_pin_9_
port 138 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_42_
port 139 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_43_
port 140 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_44_
port 141 nsew default input
rlabel metal2 s 1950 27520 2006 28000 6 top_left_grid_pin_45_
port 142 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 top_left_grid_pin_46_
port 143 nsew default input
rlabel metal2 s 3054 27520 3110 28000 6 top_left_grid_pin_47_
port 144 nsew default input
rlabel metal2 s 3606 27520 3662 28000 6 top_left_grid_pin_48_
port 145 nsew default input
rlabel metal2 s 4158 27520 4214 28000 6 top_left_grid_pin_49_
port 146 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 147 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 148 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
